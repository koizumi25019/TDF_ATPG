module s1423 (G0, G1, G2, G3, G4
    , G5, G6, G7, G8, G9
    , G10, G11, G12, G13, G14
    , G15, G16, CLK
    , G726, G729, G702, G727, G701BF
    ) ;

input   G0, G1, G2, G3, G4
    , G5, G6, G7, G8, G9
    , G10, G11, G12, G13, G14
    , G15, G16, CLK ;

output  G726, G729, G702, G727, G701BF
     ;

INV     gate0  (.A(II1260), .Z(G726) ) ;
INV     gate1  (.A(II1267), .Z(G729) ) ;
AND2    gate2  (.A(G703), .B(G645), .Z(G702) ) ;
AND2    gate3  (.A(G476), .B(G645), .Z(G727) ) ;
INV     gate4  (.A(II1211), .Z(G701BF) ) ;
INV     gate5  (.A(II1), .Z(G332BF) ) ;
DFF     gate6  (.D(G332BF), .CP(CLK), .Q(G22) ) ;
INV     gate7  (.A(II12), .Z(G328BF) ) ;
DFF     gate8  (.D(G328BF), .CP(CLK), .Q(G23) ) ;
AND2    gate9  (.A(G106), .B(G108), .Z(G109) ) ;
DFF     gate10  (.D(G109), .CP(CLK), .Q(G24) ) ;
AND2    gate11  (.A(G114), .B(G112), .Z(G113) ) ;
DFF     gate12  (.D(G113), .CP(CLK), .Q(G25) ) ;
AND2    gate13  (.A(G119), .B(G117), .Z(G118) ) ;
DFF     gate14  (.D(G118), .CP(CLK), .Q(G26) ) ;
AND2    gate15  (.A(G122), .B(G124), .Z(G125) ) ;
DFF     gate16  (.D(G125), .CP(CLK), .Q(G27) ) ;
AND2    gate17  (.A(G130), .B(G128), .Z(G129) ) ;
DFF     gate18  (.D(G129), .CP(CLK), .Q(G28) ) ;
AND2    gate19  (.A(G137), .B(G139), .Z(G140) ) ;
DFF     gate20  (.D(G140), .CP(CLK), .Q(G29) ) ;
AND2    gate21  (.A(G145), .B(G143), .Z(G144) ) ;
DFF     gate22  (.D(G144), .CP(CLK), .Q(G30) ) ;
AND2    gate23  (.A(G150), .B(G148), .Z(G149) ) ;
DFF     gate24  (.D(G149), .CP(CLK), .Q(G31) ) ;
AND2    gate25  (.A(G155), .B(G153), .Z(G154) ) ;
DFF     gate26  (.D(G154), .CP(CLK), .Q(G32) ) ;
AND2    gate27  (.A(G160), .B(G158), .Z(G159) ) ;
DFF     gate28  (.D(G159), .CP(CLK), .Q(G33) ) ;
AND2    gate29  (.A(G163), .B(G165), .Z(G166) ) ;
DFF     gate30  (.D(G166), .CP(CLK), .Q(G34) ) ;
AND2    gate31  (.A(G176), .B(G174), .Z(G175) ) ;
DFF     gate32  (.D(G175), .CP(CLK), .Q(G35) ) ;
AND2    gate33  (.A(G186), .B(G188), .Z(G189) ) ;
DFF     gate34  (.D(G189), .CP(CLK), .Q(G36) ) ;
AND2    gate35  (.A(G194), .B(G192), .Z(G193) ) ;
DFF     gate36  (.D(G193), .CP(CLK), .Q(G37) ) ;
AND2    gate37  (.A(G199), .B(G197), .Z(G198) ) ;
DFF     gate38  (.D(G198), .CP(CLK), .Q(G38) ) ;
AND2    gate39  (.A(G205), .B(G207), .Z(G208) ) ;
DFF     gate40  (.D(G208), .CP(CLK), .Q(G39) ) ;
AND2    gate41  (.A(G211), .B(G213), .Z(G214) ) ;
DFF     gate42  (.D(G214), .CP(CLK), .Q(G40) ) ;
AND2    gate43  (.A(G219), .B(G217), .Z(G218) ) ;
DFF     gate44  (.D(G218), .CP(CLK), .Q(G41) ) ;
AND2    gate45  (.A(G238), .B(G236), .Z(G237) ) ;
DFF     gate46  (.D(G237), .CP(CLK), .Q(G42) ) ;
AND2    gate47  (.A(G243), .B(G241), .Z(G242) ) ;
DFF     gate48  (.D(G242), .CP(CLK), .Q(G43) ) ;
AND2    gate49  (.A(G248), .B(G246), .Z(G247) ) ;
DFF     gate50  (.D(G247), .CP(CLK), .Q(G44) ) ;
AND2    gate51  (.A(G253), .B(G251), .Z(G252) ) ;
DFF     gate52  (.D(G252), .CP(CLK), .Q(G45) ) ;
AND2    gate53  (.A(G256), .B(G258), .Z(G260) ) ;
DFF     gate54  (.D(G260), .CP(CLK), .Q(G46) ) ;
AND2    gate55  (.A(G304), .B(G302), .Z(G303) ) ;
DFF     gate56  (.D(G303), .CP(CLK), .Q(G47) ) ;
AND2    gate57  (.A(G310), .B(G308), .Z(G309) ) ;
DFF     gate58  (.D(G309), .CP(CLK), .Q(G48) ) ;
AND2    gate59  (.A(G316), .B(G314), .Z(G315) ) ;
DFF     gate60  (.D(G315), .CP(CLK), .Q(G49) ) ;
AND2    gate61  (.A(G322), .B(G320), .Z(G321) ) ;
DFF     gate62  (.D(G321), .CP(CLK), .Q(G50) ) ;
AND2    gate63  (.A(G361), .B(G359), .Z(G360) ) ;
DFF     gate64  (.D(G360), .CP(CLK), .Q(G51) ) ;
AND2    gate65  (.A(G366), .B(G364), .Z(G365) ) ;
DFF     gate66  (.D(G365), .CP(CLK), .Q(G52) ) ;
AND2    gate67  (.A(G369), .B(G371), .Z(G373) ) ;
DFF     gate68  (.D(G373), .CP(CLK), .Q(G53) ) ;
AND2    gate69  (.A(G380), .B(G378), .Z(G379) ) ;
DFF     gate70  (.D(G379), .CP(CLK), .Q(G54) ) ;
AND2    gate71  (.A(G385), .B(G383), .Z(G384) ) ;
DFF     gate72  (.D(G384), .CP(CLK), .Q(G55) ) ;
AND2    gate73  (.A(G388), .B(G390), .Z(G392) ) ;
DFF     gate74  (.D(G392), .CP(CLK), .Q(G56) ) ;
AND2    gate75  (.A(G398), .B(G396), .Z(G397) ) ;
DFF     gate76  (.D(G397), .CP(CLK), .Q(G57) ) ;
AND2    gate77  (.A(G401), .B(G403), .Z(G405) ) ;
DFF     gate78  (.D(G405), .CP(CLK), .Q(G58) ) ;
AND2    gate79  (.A(G409), .B(G407), .Z(G408) ) ;
DFF     gate80  (.D(G408), .CP(CLK), .Q(G59) ) ;
AND2    gate81  (.A(G417), .B(G415), .Z(G416) ) ;
DFF     gate82  (.D(G416), .CP(CLK), .Q(G60) ) ;
AND2    gate83  (.A(G420), .B(G422), .Z(G424) ) ;
DFF     gate84  (.D(G424), .CP(CLK), .Q(G61) ) ;
AND2    gate85  (.A(G428), .B(G426), .Z(G427) ) ;
DFF     gate86  (.D(G427), .CP(CLK), .Q(G62) ) ;
AND2    gate87  (.A(G439), .B(G437), .Z(G438) ) ;
DFF     gate88  (.D(G438), .CP(CLK), .Q(G63) ) ;
AND2    gate89  (.A(G442), .B(G440), .Z(G441) ) ;
DFF     gate90  (.D(G441), .CP(CLK), .Q(G64) ) ;
AND2    gate91  (.A(G448), .B(G446), .Z(G447) ) ;
DFF     gate92  (.D(G447), .CP(CLK), .Q(G65) ) ;
AND2    gate93  (.A(G452), .B(G450), .Z(G451) ) ;
DFF     gate94  (.D(G451), .CP(CLK), .Q(G66) ) ;
AND2    gate95  (.A(G460), .B(G458), .Z(G459) ) ;
DFF     gate96  (.D(G459), .CP(CLK), .Q(G67) ) ;
AND2    gate97  (.A(G465), .B(G463), .Z(G464) ) ;
DFF     gate98  (.D(G464), .CP(CLK), .Q(G68) ) ;
AND2    gate99  (.A(G470), .B(G468), .Z(G469) ) ;
DFF     gate100  (.D(G469), .CP(CLK), .Q(G69) ) ;
AND2    gate101  (.A(G473), .B(G475), .Z(G477) ) ;
DFF     gate102  (.D(G477), .CP(CLK), .Q(G70) ) ;
AND2    gate103  (.A(G492), .B(G493), .Z(G494) ) ;
DFF     gate104  (.D(G494), .CP(CLK), .Q(G71) ) ;
AND2    gate105  (.A(G496), .B(G497), .Z(G498) ) ;
DFF     gate106  (.D(G498), .CP(CLK), .Q(G72) ) ;
AND2    gate107  (.A(G501), .B(G502), .Z(G503) ) ;
DFF     gate108  (.D(G503), .CP(CLK), .Q(G73) ) ;
AND2    gate109  (.A(G527), .B(G525), .Z(G526) ) ;
DFF     gate110  (.D(G526), .CP(CLK), .Q(G74) ) ;
AND2    gate111  (.A(G532), .B(G530), .Z(G531) ) ;
DFF     gate112  (.D(G531), .CP(CLK), .Q(G75) ) ;
AND2    gate113  (.A(G537), .B(G535), .Z(G536) ) ;
DFF     gate114  (.D(G536), .CP(CLK), .Q(G76) ) ;
AND2    gate115  (.A(G542), .B(G540), .Z(G541) ) ;
DFF     gate116  (.D(G541), .CP(CLK), .Q(G77) ) ;
AND2    gate117  (.A(G545), .B(G547), .Z(G548) ) ;
DFF     gate118  (.D(G548), .CP(CLK), .Q(G78) ) ;
AND2    gate119  (.A(G563), .B(G564), .Z(G565) ) ;
DFF     gate120  (.D(G565), .CP(CLK), .Q(G79) ) ;
AND2    gate121  (.A(G567), .B(G568), .Z(G569) ) ;
DFF     gate122  (.D(G569), .CP(CLK), .Q(G80) ) ;
AND2    gate123  (.A(G571), .B(G572), .Z(G573) ) ;
DFF     gate124  (.D(G573), .CP(CLK), .Q(G81) ) ;
AND2    gate125  (.A(G575), .B(G576), .Z(G577) ) ;
DFF     gate126  (.D(G577), .CP(CLK), .Q(G82) ) ;
AND2    gate127  (.A(G591), .B(G588), .Z(G590) ) ;
DFF     gate128  (.D(G590), .CP(CLK), .Q(G83) ) ;
AND2    gate129  (.A(G606), .B(G607), .Z(G608) ) ;
DFF     gate130  (.D(G608), .CP(CLK), .Q(G84) ) ;
AND2    gate131  (.A(G611), .B(G612), .Z(G613) ) ;
DFF     gate132  (.D(G613), .CP(CLK), .Q(G85) ) ;
AND2    gate133  (.A(G659), .B(G656), .Z(G657) ) ;
DFF     gate134  (.D(G657), .CP(CLK), .Q(G86) ) ;
AND2    gate135  (.A(G664), .B(G662), .Z(G663) ) ;
DFF     gate136  (.D(G663), .CP(CLK), .Q(G87) ) ;
AND2    gate137  (.A(G670), .B(G668), .Z(G669) ) ;
DFF     gate138  (.D(G669), .CP(CLK), .Q(G88) ) ;
AND2    gate139  (.A(G676), .B(G674), .Z(G675) ) ;
DFF     gate140  (.D(G675), .CP(CLK), .Q(G89) ) ;
OR2     gate141  (.A(G681), .B(G699), .Z(G682) ) ;
DFF     gate142  (.D(G682), .CP(CLK), .Q(G90) ) ;
OR2     gate143  (.A(G686), .B(G699), .Z(G687) ) ;
DFF     gate144  (.D(G687), .CP(CLK), .Q(G91) ) ;
OR2     gate145  (.A(G692), .B(G699), .Z(G693) ) ;
DFF     gate146  (.D(G693), .CP(CLK), .Q(G92) ) ;
AND2    gate147  (.A(G230), .B(G704), .Z(G705) ) ;
DFF     gate148  (.D(G705), .CP(CLK), .Q(G93) ) ;
AND2    gate149  (.A(G708), .B(G706), .Z(G707) ) ;
DFF     gate150  (.D(G707), .CP(CLK), .Q(G94) ) ;
AND2    gate151  (.A(G599), .B(G711), .Z(G713) ) ;
DFF     gate152  (.D(G713), .CP(CLK), .Q(G95) ) ;
NAND2   gate153  (.A(G334), .B(G331), .Z(G332) ) ;
INV     gate154  (.A(G332), .Z(II1) ) ;
NOR2    gate155  (.A(G329), .B(G327), .Z(G328) ) ;
INV     gate156  (.A(G328), .Z(II12) ) ;
INV     gate157  (.A(G14), .Z(G712) ) ;
INV     gate158  (.A(G712), .Z(G108) ) ;
INV     gate159  (.A(G24), .Z(G111) ) ;
INV     gate160  (.A(G712), .Z(G112) ) ;
INV     gate161  (.A(G712), .Z(G117) ) ;
INV     gate162  (.A(G712), .Z(G124) ) ;
INV     gate163  (.A(G27), .Z(G127) ) ;
INV     gate164  (.A(G712), .Z(G128) ) ;
INV     gate165  (.A(G712), .Z(G139) ) ;
INV     gate166  (.A(G29), .Z(G142) ) ;
INV     gate167  (.A(G712), .Z(G143) ) ;
INV     gate168  (.A(G712), .Z(G148) ) ;
INV     gate169  (.A(G712), .Z(G153) ) ;
INV     gate170  (.A(G712), .Z(G158) ) ;
INV     gate171  (.A(G712), .Z(G165) ) ;
INV     gate172  (.A(G712), .Z(G174) ) ;
INV     gate173  (.A(G35), .Z(G176) ) ;
INV     gate174  (.A(G34), .Z(G178) ) ;
INV     gate175  (.A(G92), .Z(G180) ) ;
INV     gate176  (.A(G180), .Z(G179) ) ;
INV     gate177  (.A(G712), .Z(G188) ) ;
INV     gate178  (.A(G36), .Z(G191) ) ;
INV     gate179  (.A(G712), .Z(G192) ) ;
INV     gate180  (.A(G712), .Z(G197) ) ;
INV     gate181  (.A(G38), .Z(G204) ) ;
INV     gate182  (.A(G712), .Z(G207) ) ;
INV     gate183  (.A(G39), .Z(G210) ) ;
INV     gate184  (.A(G712), .Z(G213) ) ;
INV     gate185  (.A(G40), .Z(G216) ) ;
INV     gate186  (.A(G712), .Z(G217) ) ;
AND2    gate187  (.A(G624), .B(G625), .Z(G259) ) ;
INV     gate188  (.A(G259), .Z(G236) ) ;
INV     gate189  (.A(G259), .Z(G241) ) ;
INV     gate190  (.A(G259), .Z(G246) ) ;
INV     gate191  (.A(G259), .Z(G251) ) ;
INV     gate192  (.A(G259), .Z(G258) ) ;
NAND2   gate193  (.A(G289), .B(G290), .Z(G297) ) ;
INV     gate194  (.A(G297), .Z(G296) ) ;
INV     gate195  (.A(G712), .Z(G302) ) ;
OR2     gate196  (.A(G377), .B(G348), .Z(G324) ) ;
INV     gate197  (.A(G324), .Z(G305) ) ;
INV     gate198  (.A(G712), .Z(G308) ) ;
INV     gate199  (.A(G324), .Z(G311) ) ;
INV     gate200  (.A(G712), .Z(G314) ) ;
INV     gate201  (.A(G324), .Z(G317) ) ;
INV     gate202  (.A(G712), .Z(G320) ) ;
INV     gate203  (.A(G324), .Z(G323) ) ;
OR2     gate204  (.A(G457), .B(G645), .Z(G355) ) ;
INV     gate205  (.A(G355), .Z(G336) ) ;
INV     gate206  (.A(G355), .Z(G339) ) ;
INV     gate207  (.A(G91), .Z(G348) ) ;
INV     gate208  (.A(G348), .Z(G343) ) ;
INV     gate209  (.A(G348), .Z(G347) ) ;
INV     gate210  (.A(G90), .Z(G645) ) ;
INV     gate211  (.A(G645), .Z(G351) ) ;
INV     gate212  (.A(G355), .Z(G354) ) ;
OR2     gate213  (.A(G712), .B(G358), .Z(G372) ) ;
INV     gate214  (.A(G372), .Z(G359) ) ;
INV     gate215  (.A(G372), .Z(G364) ) ;
INV     gate216  (.A(G372), .Z(G371) ) ;
OR2     gate217  (.A(G712), .B(G377), .Z(G391) ) ;
INV     gate218  (.A(G391), .Z(G378) ) ;
INV     gate219  (.A(G391), .Z(G383) ) ;
INV     gate220  (.A(G391), .Z(G390) ) ;
OR2     gate221  (.A(G712), .B(G413), .Z(G404) ) ;
INV     gate222  (.A(G404), .Z(G396) ) ;
INV     gate223  (.A(G404), .Z(G403) ) ;
INV     gate224  (.A(G712), .Z(G407) ) ;
OR2     gate225  (.A(G712), .B(G432), .Z(G423) ) ;
INV     gate226  (.A(G423), .Z(G415) ) ;
INV     gate227  (.A(G423), .Z(G422) ) ;
INV     gate228  (.A(G712), .Z(G426) ) ;
INV     gate229  (.A(G712), .Z(G437) ) ;
INV     gate230  (.A(G712), .Z(G440) ) ;
INV     gate231  (.A(G65), .Z(G445) ) ;
INV     gate232  (.A(G712), .Z(G446) ) ;
INV     gate233  (.A(G66), .Z(G449) ) ;
INV     gate234  (.A(G712), .Z(G450) ) ;
OR2     gate235  (.A(G83), .B(G524), .Z(G456) ) ;
INV     gate236  (.A(G456), .Z(G455) ) ;
NAND2   gate237  (.A(G486), .B(G616), .Z(G476) ) ;
INV     gate238  (.A(G476), .Z(G458) ) ;
INV     gate239  (.A(G476), .Z(G463) ) ;
INV     gate240  (.A(G476), .Z(G468) ) ;
INV     gate241  (.A(G476), .Z(G475) ) ;
INV     gate242  (.A(G712), .Z(G486) ) ;
OR2     gate243  (.A(G654), .B(G712), .Z(G500) ) ;
INV     gate244  (.A(G500), .Z(G491) ) ;
INV     gate245  (.A(G500), .Z(G495) ) ;
INV     gate246  (.A(G500), .Z(G499) ) ;
INV     gate247  (.A(G63), .Z(G511) ) ;
INV     gate248  (.A(G511), .Z(G504) ) ;
INV     gate249  (.A(G511), .Z(G507) ) ;
INV     gate250  (.A(G511), .Z(G510) ) ;
AND2    gate251  (.A(G627), .B(G628), .Z(G589) ) ;
INV     gate252  (.A(G589), .Z(G525) ) ;
INV     gate253  (.A(G589), .Z(G530) ) ;
INV     gate254  (.A(G589), .Z(G535) ) ;
INV     gate255  (.A(G589), .Z(G540) ) ;
INV     gate256  (.A(G589), .Z(G547) ) ;
OR2     gate257  (.A(G655), .B(G712), .Z(G610) ) ;
INV     gate258  (.A(G610), .Z(G562) ) ;
INV     gate259  (.A(G610), .Z(G566) ) ;
INV     gate260  (.A(G610), .Z(G570) ) ;
INV     gate261  (.A(G610), .Z(G574) ) ;
INV     gate262  (.A(G589), .Z(G588) ) ;
NOR2    gate263  (.A(G435), .B(G524), .Z(G593) ) ;
INV     gate264  (.A(G593), .Z(G595) ) ;
NAND2   gate265  (.A(G602), .B(G603), .Z(G597) ) ;
INV     gate266  (.A(G597), .Z(G596) ) ;
AND2    gate267  (.A(G621), .B(G622), .Z(G601) ) ;
INV     gate268  (.A(G601), .Z(G600) ) ;
INV     gate269  (.A(G610), .Z(G605) ) ;
INV     gate270  (.A(G610), .Z(G609) ) ;
INV     gate271  (.A(G64), .Z(G614) ) ;
NAND4   gate272  (.A(G482), .B(G483), .C(G484), .D(G485), .Z(G616) ) ;
INV     gate273  (.A(G616), .Z(G615) ) ;
INV     gate274  (.A(G645), .Z(G617) ) ;
INV     gate275  (.A(G645), .Z(G620) ) ;
INV     gate276  (.A(G645), .Z(G623) ) ;
INV     gate277  (.A(G645), .Z(G626) ) ;
INV     gate278  (.A(G645), .Z(G629) ) ;
INV     gate279  (.A(G645), .Z(G632) ) ;
INV     gate280  (.A(G645), .Z(G635) ) ;
INV     gate281  (.A(G645), .Z(G638) ) ;
INV     gate282  (.A(G645), .Z(G641) ) ;
INV     gate283  (.A(G645), .Z(G644) ) ;
INV     gate284  (.A(G712), .Z(G656) ) ;
INV     gate285  (.A(II1162), .Z(G659) ) ;
INV     gate286  (.A(G659), .Z(G658) ) ;
INV     gate287  (.A(G13), .Z(II1162) ) ;
INV     gate288  (.A(G94), .Z(G661) ) ;
INV     gate289  (.A(G712), .Z(G662) ) ;
INV     gate290  (.A(II1183), .Z(G678) ) ;
INV     gate291  (.A(G678), .Z(G665) ) ;
INV     gate292  (.A(G712), .Z(G668) ) ;
INV     gate293  (.A(G678), .Z(G671) ) ;
INV     gate294  (.A(G712), .Z(G674) ) ;
INV     gate295  (.A(G678), .Z(G677) ) ;
INV     gate296  (.A(G11), .Z(II1183) ) ;
INV     gate297  (.A(II1203), .Z(G696) ) ;
INV     gate298  (.A(G696), .Z(G685) ) ;
INV     gate299  (.A(G696), .Z(G689) ) ;
INV     gate300  (.A(G696), .Z(G695) ) ;
INV     gate301  (.A(G10), .Z(II1203) ) ;
INV     gate302  (.A(G15), .Z(G701) ) ;
INV     gate303  (.A(G701), .Z(II1211) ) ;
INV     gate304  (.A(G712), .Z(G704) ) ;
INV     gate305  (.A(G712), .Z(G706) ) ;
INV     gate306  (.A(G712), .Z(G711) ) ;
INV     gate307  (.A(G701), .Z(G714) ) ;
INV     gate308  (.A(G6), .Z(II1227) ) ;
INV     gate309  (.A(II1227), .Z(G715) ) ;
INV     gate310  (.A(G7), .Z(II1230) ) ;
INV     gate311  (.A(II1230), .Z(G716) ) ;
INV     gate312  (.A(G8), .Z(II1233) ) ;
INV     gate313  (.A(II1233), .Z(G717) ) ;
INV     gate314  (.A(G9), .Z(II1236) ) ;
INV     gate315  (.A(II1236), .Z(G718) ) ;
INV     gate316  (.A(G12), .Z(II1239) ) ;
INV     gate317  (.A(II1239), .Z(G719) ) ;
INV     gate318  (.A(G0), .Z(II1242) ) ;
INV     gate319  (.A(II1242), .Z(G720) ) ;
INV     gate320  (.A(G1), .Z(II1245) ) ;
INV     gate321  (.A(II1245), .Z(G721) ) ;
INV     gate322  (.A(G2), .Z(II1248) ) ;
INV     gate323  (.A(II1248), .Z(G722) ) ;
INV     gate324  (.A(G3), .Z(II1251) ) ;
INV     gate325  (.A(II1251), .Z(G723) ) ;
INV     gate326  (.A(G4), .Z(II1254) ) ;
INV     gate327  (.A(II1254), .Z(G724) ) ;
INV     gate328  (.A(G5), .Z(II1257) ) ;
INV     gate329  (.A(II1257), .Z(G725) ) ;
INV     gate330  (.A(G93), .Z(II1260) ) ;
INV     gate331  (.A(G16), .Z(II1264) ) ;
INV     gate332  (.A(II1264), .Z(G728) ) ;
INV     gate333  (.A(G95), .Z(II1267) ) ;
OR2     gate334  (.A(G96), .B(G645), .Z(G630) ) ;
OR2     gate335  (.A(G720), .B(G629), .Z(G631) ) ;
AND2    gate336  (.A(G630), .B(G631), .Z(G101) ) ;
OR2     gate337  (.A(G97), .B(G645), .Z(G633) ) ;
OR2     gate338  (.A(G721), .B(G632), .Z(G634) ) ;
AND2    gate339  (.A(G633), .B(G634), .Z(G102) ) ;
OR2     gate340  (.A(G98), .B(G645), .Z(G636) ) ;
OR2     gate341  (.A(G722), .B(G635), .Z(G637) ) ;
AND2    gate342  (.A(G636), .B(G637), .Z(G103) ) ;
OR2     gate343  (.A(G99), .B(G645), .Z(G639) ) ;
OR2     gate344  (.A(G723), .B(G638), .Z(G640) ) ;
AND2    gate345  (.A(G639), .B(G640), .Z(G104) ) ;
OR2     gate346  (.A(G100), .B(G645), .Z(G642) ) ;
OR2     gate347  (.A(G724), .B(G641), .Z(G643) ) ;
AND2    gate348  (.A(G642), .B(G643), .Z(G105) ) ;
NAND2   gate349  (.A(G107), .B(G110), .Z(G106) ) ;
NOR2    gate350  (.A(G115), .B(G116), .Z(G114) ) ;
AND2    gate351  (.A(G700), .B(G111), .Z(G133) ) ;
AND2    gate352  (.A(G133), .B(G25), .Z(G116) ) ;
NOR2    gate353  (.A(G120), .B(G121), .Z(G119) ) ;
AND2    gate354  (.A(G133), .B(G25), .Z(G134) ) ;
AND2    gate355  (.A(G134), .B(G26), .Z(G121) ) ;
NAND2   gate356  (.A(G123), .B(G126), .Z(G122) ) ;
NOR2    gate357  (.A(G131), .B(G132), .Z(G130) ) ;
AND2    gate358  (.A(G135), .B(G127), .Z(G136) ) ;
AND2    gate359  (.A(G136), .B(G28), .Z(G132) ) ;
NAND2   gate360  (.A(G282), .B(G283), .Z(G700) ) ;
AND2    gate361  (.A(G134), .B(G26), .Z(G135) ) ;
NAND2   gate362  (.A(G138), .B(G141), .Z(G137) ) ;
NOR2    gate363  (.A(G146), .B(G147), .Z(G145) ) ;
AND2    gate364  (.A(G177), .B(G142), .Z(G168) ) ;
AND2    gate365  (.A(G168), .B(G30), .Z(G147) ) ;
NOR2    gate366  (.A(G151), .B(G152), .Z(G150) ) ;
AND2    gate367  (.A(G168), .B(G30), .Z(G169) ) ;
AND2    gate368  (.A(G169), .B(G31), .Z(G152) ) ;
NOR2    gate369  (.A(G156), .B(G157), .Z(G155) ) ;
AND2    gate370  (.A(G169), .B(G31), .Z(G170) ) ;
AND2    gate371  (.A(G170), .B(G32), .Z(G157) ) ;
NOR2    gate372  (.A(G161), .B(G162), .Z(G160) ) ;
AND2    gate373  (.A(G170), .B(G32), .Z(G171) ) ;
AND2    gate374  (.A(G171), .B(G33), .Z(G162) ) ;
NAND2   gate375  (.A(G164), .B(G167), .Z(G163) ) ;
OR2     gate376  (.A(G180), .B(G226), .Z(G177) ) ;
AND2    gate377  (.A(G171), .B(G33), .Z(G172) ) ;
AND2    gate378  (.A(G172), .B(G34), .Z(G173) ) ;
OR2     gate379  (.A(G178), .B(G180), .Z(G181) ) ;
OR2     gate380  (.A(G35), .B(G179), .Z(G182) ) ;
AND2    gate381  (.A(G181), .B(G182), .Z(G185) ) ;
NAND2   gate382  (.A(G187), .B(G190), .Z(G186) ) ;
NOR2    gate383  (.A(G195), .B(G196), .Z(G194) ) ;
AND2    gate384  (.A(G522), .B(G191), .Z(G202) ) ;
AND2    gate385  (.A(G202), .B(G37), .Z(G196) ) ;
NOR2    gate386  (.A(G200), .B(G201), .Z(G199) ) ;
AND2    gate387  (.A(G202), .B(G37), .Z(G203) ) ;
AND2    gate388  (.A(G203), .B(G38), .Z(G201) ) ;
OR2     gate389  (.A(G348), .B(G228), .Z(G522) ) ;
NAND2   gate390  (.A(G206), .B(G209), .Z(G205) ) ;
NAND2   gate391  (.A(G212), .B(G215), .Z(G211) ) ;
NOR2    gate392  (.A(G220), .B(G221), .Z(G219) ) ;
AND2    gate393  (.A(G222), .B(G216), .Z(G223) ) ;
AND2    gate394  (.A(G223), .B(G41), .Z(G221) ) ;
OR2     gate395  (.A(G180), .B(G227), .Z(G183) ) ;
AND2    gate396  (.A(G183), .B(G210), .Z(G222) ) ;
AND2    gate397  (.A(G203), .B(G38), .Z(G224) ) ;
AND2    gate398  (.A(G204), .B(G203), .Z(G225) ) ;
AND2    gate399  (.A(G136), .B(G28), .Z(G226) ) ;
AND2    gate400  (.A(G172), .B(G178), .Z(G227) ) ;
AND2    gate401  (.A(G223), .B(G41), .Z(G228) ) ;
AND2    gate402  (.A(G358), .B(G61), .Z(G432) ) ;
AND2    gate403  (.A(G432), .B(G62), .Z(G229) ) ;
NOR2    gate404  (.A(G239), .B(G240), .Z(G238) ) ;
NOR2    gate405  (.A(G301), .B(G328), .Z(G299) ) ;
AND2    gate406  (.A(G299), .B(G42), .Z(G240) ) ;
NOR2    gate407  (.A(G244), .B(G245), .Z(G243) ) ;
AND2    gate408  (.A(G299), .B(G42), .Z(G262) ) ;
AND2    gate409  (.A(G262), .B(G43), .Z(G245) ) ;
NOR2    gate410  (.A(G249), .B(G250), .Z(G248) ) ;
AND2    gate411  (.A(G262), .B(G43), .Z(G263) ) ;
AND2    gate412  (.A(G263), .B(G44), .Z(G250) ) ;
NOR2    gate413  (.A(G254), .B(G255), .Z(G253) ) ;
AND2    gate414  (.A(G263), .B(G44), .Z(G264) ) ;
AND2    gate415  (.A(G264), .B(G45), .Z(G255) ) ;
OR2     gate416  (.A(G476), .B(G645), .Z(G624) ) ;
OR2     gate417  (.A(G716), .B(G623), .Z(G625) ) ;
NOR2    gate418  (.A(G257), .B(G261), .Z(G256) ) ;
AND2    gate419  (.A(G264), .B(G45), .Z(G265) ) ;
AND2    gate420  (.A(G265), .B(G46), .Z(G261) ) ;
OR2     gate421  (.A(G101), .B(G42), .Z(G275) ) ;
NAND2   gate422  (.A(G286), .B(G291), .Z(G266) ) ;
AND2    gate423  (.A(G275), .B(G266), .Z(G271) ) ;
OR2     gate424  (.A(G102), .B(G43), .Z(G276) ) ;
OR2     gate425  (.A(G267), .B(G271), .Z(G277) ) ;
AND2    gate426  (.A(G276), .B(G277), .Z(G272) ) ;
OR2     gate427  (.A(G103), .B(G44), .Z(G278) ) ;
OR2     gate428  (.A(G268), .B(G272), .Z(G279) ) ;
AND2    gate429  (.A(G278), .B(G279), .Z(G273) ) ;
OR2     gate430  (.A(G104), .B(G45), .Z(G280) ) ;
OR2     gate431  (.A(G269), .B(G273), .Z(G281) ) ;
AND2    gate432  (.A(G280), .B(G281), .Z(G274) ) ;
AND2    gate433  (.A(G306), .B(G307), .Z(G304) ) ;
OR2     gate434  (.A(G47), .B(G324), .Z(G306) ) ;
OR2     gate435  (.A(G719), .B(G305), .Z(G307) ) ;
AND2    gate436  (.A(G312), .B(G313), .Z(G310) ) ;
OR2     gate437  (.A(G48), .B(G324), .Z(G312) ) ;
OR2     gate438  (.A(G47), .B(G311), .Z(G313) ) ;
AND2    gate439  (.A(G318), .B(G319), .Z(G316) ) ;
OR2     gate440  (.A(G49), .B(G324), .Z(G318) ) ;
OR2     gate441  (.A(G48), .B(G317), .Z(G319) ) ;
AND2    gate442  (.A(G325), .B(G326), .Z(G322) ) ;
OR2     gate443  (.A(G50), .B(G324), .Z(G325) ) ;
OR2     gate444  (.A(G49), .B(G323), .Z(G326) ) ;
NAND2   gate445  (.A(G333), .B(G22), .Z(G331) ) ;
AND2    gate446  (.A(G331), .B(G714), .Z(G329) ) ;
AND2    gate447  (.A(G332), .B(G714), .Z(G330) ) ;
OR2     gate448  (.A(G224), .B(G355), .Z(G337) ) ;
OR2     gate449  (.A(G183), .B(G336), .Z(G338) ) ;
AND2    gate450  (.A(G337), .B(G338), .Z(G335) ) ;
OR2     gate451  (.A(G229), .B(G348), .Z(G344) ) ;
OR2     gate452  (.A(G414), .B(G343), .Z(G345) ) ;
AND2    gate453  (.A(G344), .B(G345), .Z(G342) ) ;
OR2     gate454  (.A(G62), .B(G348), .Z(G349) ) ;
OR2     gate455  (.A(G59), .B(G347), .Z(G350) ) ;
AND2    gate456  (.A(G349), .B(G350), .Z(G346) ) ;
OR2     gate457  (.A(G348), .B(G414), .Z(G523) ) ;
AND2    gate458  (.A(G523), .B(G53), .Z(G358) ) ;
NOR2    gate459  (.A(G362), .B(G363), .Z(G361) ) ;
AND2    gate460  (.A(G523), .B(G51), .Z(G363) ) ;
NOR2    gate461  (.A(G367), .B(G368), .Z(G366) ) ;
AND2    gate462  (.A(G523), .B(G51), .Z(G375) ) ;
AND2    gate463  (.A(G375), .B(G52), .Z(G368) ) ;
NOR2    gate464  (.A(G370), .B(G374), .Z(G369) ) ;
AND2    gate465  (.A(G375), .B(G52), .Z(G376) ) ;
AND2    gate466  (.A(G376), .B(G53), .Z(G374) ) ;
AND3    gate467  (.A(G183), .B(G54), .C(G56), .Z(G377) ) ;
NOR2    gate468  (.A(G381), .B(G382), .Z(G380) ) ;
AND2    gate469  (.A(G183), .B(G54), .Z(G382) ) ;
NOR2    gate470  (.A(G386), .B(G387), .Z(G385) ) ;
AND2    gate471  (.A(G183), .B(G54), .Z(G394) ) ;
AND2    gate472  (.A(G394), .B(G55), .Z(G387) ) ;
NOR2    gate473  (.A(G389), .B(G393), .Z(G388) ) ;
AND2    gate474  (.A(G394), .B(G55), .Z(G395) ) ;
AND2    gate475  (.A(G395), .B(G56), .Z(G393) ) ;
NOR2    gate476  (.A(G399), .B(G400), .Z(G398) ) ;
AND2    gate477  (.A(G335), .B(G57), .Z(G400) ) ;
NOR2    gate478  (.A(G402), .B(G406), .Z(G401) ) ;
AND2    gate479  (.A(G335), .B(G57), .Z(G412) ) ;
AND2    gate480  (.A(G412), .B(G58), .Z(G406) ) ;
NOR2    gate481  (.A(G410), .B(G411), .Z(G409) ) ;
AND2    gate482  (.A(G335), .B(G58), .Z(G413) ) ;
AND2    gate483  (.A(G413), .B(G59), .Z(G411) ) ;
AND2    gate484  (.A(G413), .B(G59), .Z(G414) ) ;
NOR2    gate485  (.A(G418), .B(G419), .Z(G417) ) ;
AND2    gate486  (.A(G358), .B(G60), .Z(G419) ) ;
NOR2    gate487  (.A(G421), .B(G425), .Z(G420) ) ;
AND2    gate488  (.A(G358), .B(G60), .Z(G431) ) ;
AND2    gate489  (.A(G431), .B(G61), .Z(G425) ) ;
NOR2    gate490  (.A(G429), .B(G430), .Z(G428) ) ;
AND2    gate491  (.A(G432), .B(G62), .Z(G430) ) ;
OR2     gate492  (.A(G225), .B(G355), .Z(G356) ) ;
OR2     gate493  (.A(G184), .B(G354), .Z(G357) ) ;
AND2    gate494  (.A(G356), .B(G357), .Z(G433) ) ;
OR2     gate495  (.A(G38), .B(G355), .Z(G340) ) ;
OR2     gate496  (.A(G185), .B(G339), .Z(G341) ) ;
AND2    gate497  (.A(G340), .B(G341), .Z(G435) ) ;
OR2     gate498  (.A(G346), .B(G645), .Z(G352) ) ;
OR2     gate499  (.A(G35), .B(G351), .Z(G353) ) ;
AND2    gate500  (.A(G352), .B(G353), .Z(G436) ) ;
OR2     gate501  (.A(G435), .B(G63), .Z(G439) ) ;
NOR2    gate502  (.A(G443), .B(G444), .Z(G442) ) ;
AND2    gate503  (.A(G615), .B(G511), .Z(G443) ) ;
OR2     gate504  (.A(G615), .B(G65), .Z(G448) ) ;
NOR2    gate505  (.A(G453), .B(G454), .Z(G452) ) ;
AND2    gate506  (.A(G615), .B(G445), .Z(G453) ) ;
AND3    gate507  (.A(G455), .B(G449), .C(G728), .Z(G457) ) ;
NOR2    gate508  (.A(G461), .B(G462), .Z(G460) ) ;
OR2     gate509  (.A(G342), .B(G645), .Z(G434) ) ;
AND2    gate510  (.A(G434), .B(G67), .Z(G462) ) ;
NOR2    gate511  (.A(G466), .B(G467), .Z(G465) ) ;
AND2    gate512  (.A(G434), .B(G67), .Z(G479) ) ;
AND2    gate513  (.A(G479), .B(G68), .Z(G467) ) ;
NOR2    gate514  (.A(G471), .B(G472), .Z(G470) ) ;
AND2    gate515  (.A(G479), .B(G68), .Z(G480) ) ;
AND2    gate516  (.A(G480), .B(G69), .Z(G472) ) ;
NOR2    gate517  (.A(G474), .B(G478), .Z(G473) ) ;
AND2    gate518  (.A(G480), .B(G69), .Z(G481) ) ;
AND2    gate519  (.A(G481), .B(G70), .Z(G478) ) ;
OR2     gate520  (.A(G723), .B(G511), .Z(G505) ) ;
OR2     gate521  (.A(G720), .B(G504), .Z(G506) ) ;
AND2    gate522  (.A(G505), .B(G506), .Z(G488) ) ;
OR2     gate523  (.A(G724), .B(G511), .Z(G508) ) ;
OR2     gate524  (.A(G721), .B(G507), .Z(G509) ) ;
AND2    gate525  (.A(G508), .B(G509), .Z(G489) ) ;
OR2     gate526  (.A(G725), .B(G511), .Z(G512) ) ;
OR2     gate527  (.A(G722), .B(G510), .Z(G513) ) ;
AND2    gate528  (.A(G512), .B(G513), .Z(G490) ) ;
OR2     gate529  (.A(G71), .B(G500), .Z(G492) ) ;
OR2     gate530  (.A(G488), .B(G491), .Z(G493) ) ;
OR2     gate531  (.A(G72), .B(G500), .Z(G496) ) ;
OR2     gate532  (.A(G489), .B(G495), .Z(G497) ) ;
OR2     gate533  (.A(G73), .B(G500), .Z(G501) ) ;
OR2     gate534  (.A(G490), .B(G499), .Z(G502) ) ;
NOR2    gate535  (.A(G528), .B(G529), .Z(G527) ) ;
AND2    gate536  (.A(G433), .B(G524), .Z(G604) ) ;
AND2    gate537  (.A(G604), .B(G74), .Z(G529) ) ;
NOR2    gate538  (.A(G533), .B(G534), .Z(G532) ) ;
AND2    gate539  (.A(G604), .B(G74), .Z(G550) ) ;
AND2    gate540  (.A(G550), .B(G75), .Z(G534) ) ;
NOR2    gate541  (.A(G538), .B(G539), .Z(G537) ) ;
AND2    gate542  (.A(G550), .B(G75), .Z(G551) ) ;
AND2    gate543  (.A(G551), .B(G76), .Z(G539) ) ;
NOR2    gate544  (.A(G543), .B(G544), .Z(G542) ) ;
AND2    gate545  (.A(G551), .B(G76), .Z(G552) ) ;
AND2    gate546  (.A(G552), .B(G77), .Z(G544) ) ;
NOR2    gate547  (.A(G546), .B(G549), .Z(G545) ) ;
AND2    gate548  (.A(G552), .B(G77), .Z(G553) ) ;
AND2    gate549  (.A(G553), .B(G78), .Z(G549) ) ;
OR2     gate550  (.A(G79), .B(G610), .Z(G563) ) ;
OR2     gate551  (.A(G715), .B(G562), .Z(G564) ) ;
OR2     gate552  (.A(G80), .B(G610), .Z(G567) ) ;
OR2     gate553  (.A(G716), .B(G566), .Z(G568) ) ;
OR2     gate554  (.A(G81), .B(G610), .Z(G571) ) ;
OR2     gate555  (.A(G717), .B(G570), .Z(G572) ) ;
OR2     gate556  (.A(G82), .B(G610), .Z(G575) ) ;
OR2     gate557  (.A(G718), .B(G574), .Z(G576) ) ;
OR2     gate558  (.A(G476), .B(G645), .Z(G627) ) ;
OR2     gate559  (.A(G718), .B(G626), .Z(G628) ) ;
OR2     gate560  (.A(G592), .B(G604), .Z(G591) ) ;
OR2     gate561  (.A(G83), .B(G593), .Z(G594) ) ;
AND2    gate562  (.A(G594), .B(G595), .Z(G592) ) ;
OR2     gate563  (.A(G614), .B(G645), .Z(G621) ) ;
OR2     gate564  (.A(G717), .B(G620), .Z(G622) ) ;
OR2     gate565  (.A(G554), .B(G555), .Z(G524) ) ;
OR2     gate566  (.A(G84), .B(G610), .Z(G606) ) ;
OR2     gate567  (.A(G696), .B(G605), .Z(G607) ) ;
OR2     gate568  (.A(G85), .B(G610), .Z(G611) ) ;
OR2     gate569  (.A(G678), .B(G609), .Z(G612) ) ;
OR2     gate570  (.A(G456), .B(G645), .Z(G646) ) ;
OR2     gate571  (.A(G725), .B(G644), .Z(G647) ) ;
AND2    gate572  (.A(G646), .B(G647), .Z(G648) ) ;
OR2     gate573  (.A(G457), .B(G645), .Z(G618) ) ;
OR2     gate574  (.A(G715), .B(G617), .Z(G619) ) ;
AND2    gate575  (.A(G618), .B(G619), .Z(G649) ) ;
AND2    gate576  (.A(G226), .B(G661), .Z(G650) ) ;
AND2    gate577  (.A(G227), .B(G87), .Z(G651) ) ;
AND2    gate578  (.A(G228), .B(G88), .Z(G652) ) ;
AND2    gate579  (.A(G229), .B(G89), .Z(G653) ) ;
AND2    gate580  (.A(G90), .B(G476), .Z(G654) ) ;
AND2    gate581  (.A(G91), .B(G476), .Z(G655) ) ;
AND2    gate582  (.A(G666), .B(G667), .Z(G664) ) ;
OR2     gate583  (.A(G87), .B(G678), .Z(G666) ) ;
OR2     gate584  (.A(G661), .B(G665), .Z(G667) ) ;
AND2    gate585  (.A(G672), .B(G673), .Z(G670) ) ;
OR2     gate586  (.A(G88), .B(G678), .Z(G672) ) ;
OR2     gate587  (.A(G87), .B(G671), .Z(G673) ) ;
AND2    gate588  (.A(G679), .B(G680), .Z(G676) ) ;
OR2     gate589  (.A(G89), .B(G678), .Z(G679) ) ;
OR2     gate590  (.A(G88), .B(G677), .Z(G680) ) ;
OR2     gate591  (.A(G645), .B(G696), .Z(G684) ) ;
AND2    gate592  (.A(G684), .B(G685), .Z(G683) ) ;
OR2     gate593  (.A(G348), .B(G696), .Z(G690) ) ;
OR2     gate594  (.A(G645), .B(G689), .Z(G691) ) ;
AND2    gate595  (.A(G690), .B(G691), .Z(G688) ) ;
OR2     gate596  (.A(G180), .B(G696), .Z(G697) ) ;
OR2     gate597  (.A(G348), .B(G695), .Z(G698) ) ;
AND2    gate598  (.A(G697), .B(G698), .Z(G694) ) ;
NOR4    gate599  (.A(G650), .B(G651), .C(G652), .D(G653), .Z(G703) ) ;
NAND2   gate600  (.A(G234), .B(G235), .Z(G230) ) ;
NOR2    gate601  (.A(G709), .B(G710), .Z(G708) ) ;
AND2    gate602  (.A(G678), .B(G89), .Z(G709) ) ;
NOR2    gate603  (.A(G598), .B(G597), .Z(G599) ) ;
OR2     gate604  (.A(G700), .B(G111), .Z(G110) ) ;
OR2     gate605  (.A(G135), .B(G127), .Z(G126) ) ;
OR2     gate606  (.A(G177), .B(G142), .Z(G141) ) ;
OR2     gate607  (.A(G172), .B(G178), .Z(G167) ) ;
OR2     gate608  (.A(G180), .B(G173), .Z(G184) ) ;
OR2     gate609  (.A(G522), .B(G191), .Z(G190) ) ;
OR2     gate610  (.A(G183), .B(G210), .Z(G209) ) ;
OR2     gate611  (.A(G222), .B(G216), .Z(G215) ) ;
NAND3   gate612  (.A(G700), .B(G232), .C(G231), .Z(G233) ) ;
OR2     gate613  (.A(G649), .B(G233), .Z(G235) ) ;
NAND2   gate614  (.A(G287), .B(G292), .Z(G267) ) ;
NAND2   gate615  (.A(G288), .B(G293), .Z(G268) ) ;
NAND2   gate616  (.A(G284), .B(G294), .Z(G269) ) ;
OR2     gate617  (.A(G105), .B(G46), .Z(G282) ) ;
NAND2   gate618  (.A(G285), .B(G295), .Z(G270) ) ;
OR2     gate619  (.A(G270), .B(G274), .Z(G283) ) ;
OR2     gate620  (.A(G42), .B(G101), .Z(G291) ) ;
OR2     gate621  (.A(G43), .B(G102), .Z(G292) ) ;
OR2     gate622  (.A(G44), .B(G103), .Z(G293) ) ;
OR2     gate623  (.A(G45), .B(G104), .Z(G294) ) ;
OR2     gate624  (.A(G46), .B(G105), .Z(G295) ) ;
OR4     gate625  (.A(G50), .B(G49), .C(G48), .D(G47), .Z(G300) ) ;
OR2     gate626  (.A(G300), .B(G714), .Z(G333) ) ;
NAND4   gate627  (.A(G50), .B(G49), .C(G48), .D(G47), .Z(G301) ) ;
OR2     gate628  (.A(G301), .B(G714), .Z(G334) ) ;
OR2     gate629  (.A(G71), .B(G67), .Z(G518) ) ;
OR2     gate630  (.A(G72), .B(G68), .Z(G519) ) ;
OR2     gate631  (.A(G73), .B(G69), .Z(G520) ) ;
NOR3    gate632  (.A(G71), .B(G72), .C(G73), .Z(G487) ) ;
OR2     gate633  (.A(G487), .B(G70), .Z(G521) ) ;
NAND3   gate634  (.A(G556), .B(G557), .C(G558), .Z(G554) ) ;
NAND2   gate635  (.A(G559), .B(G560), .Z(G555) ) ;
OR2     gate636  (.A(G79), .B(G74), .Z(G583) ) ;
OR2     gate637  (.A(G80), .B(G75), .Z(G584) ) ;
OR2     gate638  (.A(G81), .B(G76), .Z(G585) ) ;
OR2     gate639  (.A(G82), .B(G77), .Z(G586) ) ;
NOR4    gate640  (.A(G79), .B(G80), .C(G81), .D(G82), .Z(G561) ) ;
OR2     gate641  (.A(G561), .B(G78), .Z(G587) ) ;
OR2     gate642  (.A(G85), .B(G601), .Z(G602) ) ;
OR2     gate643  (.A(G600), .B(G84), .Z(G603) ) ;
NAND2   gate644  (.A(G74), .B(G596), .Z(G96) ) ;
NAND2   gate645  (.A(G75), .B(G596), .Z(G97) ) ;
NAND2   gate646  (.A(G76), .B(G596), .Z(G98) ) ;
NAND2   gate647  (.A(G77), .B(G596), .Z(G99) ) ;
NAND2   gate648  (.A(G78), .B(G596), .Z(G100) ) ;
NOR2    gate649  (.A(G683), .B(G660), .Z(G681) ) ;
OR2     gate650  (.A(G658), .B(G712), .Z(G699) ) ;
NOR2    gate651  (.A(G688), .B(G660), .Z(G686) ) ;
NOR2    gate652  (.A(G694), .B(G660), .Z(G692) ) ;
NAND2   gate653  (.A(G700), .B(G111), .Z(G107) ) ;
NAND2   gate654  (.A(G135), .B(G127), .Z(G123) ) ;
NAND2   gate655  (.A(G177), .B(G142), .Z(G138) ) ;
NAND2   gate656  (.A(G172), .B(G178), .Z(G164) ) ;
NAND2   gate657  (.A(G522), .B(G191), .Z(G187) ) ;
NAND2   gate658  (.A(G183), .B(G210), .Z(G206) ) ;
NAND2   gate659  (.A(G222), .B(G216), .Z(G212) ) ;
NAND2   gate660  (.A(G649), .B(G436), .Z(G234) ) ;
NAND2   gate661  (.A(G435), .B(G648), .Z(G231) ) ;
NAND2   gate662  (.A(G297), .B(G700), .Z(G298) ) ;
NAND3   gate663  (.A(G296), .B(G298), .C(G435), .Z(G232) ) ;
NAND2   gate664  (.A(G42), .B(G101), .Z(G286) ) ;
NAND2   gate665  (.A(G43), .B(G102), .Z(G287) ) ;
NAND2   gate666  (.A(G44), .B(G103), .Z(G288) ) ;
NAND2   gate667  (.A(G45), .B(G104), .Z(G284) ) ;
NAND2   gate668  (.A(G46), .B(G105), .Z(G285) ) ;
NOR3    gate669  (.A(G270), .B(G269), .C(G268), .Z(G289) ) ;
NOR2    gate670  (.A(G267), .B(G266), .Z(G290) ) ;
NAND2   gate671  (.A(G71), .B(G67), .Z(G514) ) ;
NAND2   gate672  (.A(G514), .B(G518), .Z(G482) ) ;
NAND2   gate673  (.A(G72), .B(G68), .Z(G515) ) ;
NAND2   gate674  (.A(G515), .B(G519), .Z(G483) ) ;
NAND2   gate675  (.A(G73), .B(G69), .Z(G516) ) ;
NAND2   gate676  (.A(G516), .B(G520), .Z(G484) ) ;
NAND2   gate677  (.A(G487), .B(G70), .Z(G517) ) ;
NAND2   gate678  (.A(G517), .B(G521), .Z(G485) ) ;
NAND2   gate679  (.A(G578), .B(G583), .Z(G556) ) ;
NAND2   gate680  (.A(G579), .B(G584), .Z(G557) ) ;
NAND2   gate681  (.A(G580), .B(G585), .Z(G558) ) ;
NAND2   gate682  (.A(G581), .B(G586), .Z(G559) ) ;
NAND2   gate683  (.A(G582), .B(G587), .Z(G560) ) ;
NAND2   gate684  (.A(G79), .B(G74), .Z(G578) ) ;
NAND2   gate685  (.A(G80), .B(G75), .Z(G579) ) ;
NAND2   gate686  (.A(G81), .B(G76), .Z(G580) ) ;
NAND2   gate687  (.A(G82), .B(G77), .Z(G581) ) ;
NAND2   gate688  (.A(G561), .B(G78), .Z(G582) ) ;
NAND2   gate689  (.A(G435), .B(G83), .Z(G598) ) ;
NOR2    gate690  (.A(G133), .B(G25), .Z(G115) ) ;
NOR2    gate691  (.A(G134), .B(G26), .Z(G120) ) ;
NOR2    gate692  (.A(G136), .B(G28), .Z(G131) ) ;
NOR2    gate693  (.A(G168), .B(G30), .Z(G146) ) ;
NOR2    gate694  (.A(G169), .B(G31), .Z(G151) ) ;
NOR2    gate695  (.A(G170), .B(G32), .Z(G156) ) ;
NOR2    gate696  (.A(G171), .B(G33), .Z(G161) ) ;
NOR2    gate697  (.A(G202), .B(G37), .Z(G195) ) ;
NOR2    gate698  (.A(G203), .B(G38), .Z(G200) ) ;
NOR2    gate699  (.A(G223), .B(G41), .Z(G220) ) ;
NOR2    gate700  (.A(G299), .B(G42), .Z(G239) ) ;
NOR2    gate701  (.A(G262), .B(G43), .Z(G244) ) ;
NOR2    gate702  (.A(G263), .B(G44), .Z(G249) ) ;
NOR2    gate703  (.A(G264), .B(G45), .Z(G254) ) ;
NOR2    gate704  (.A(G265), .B(G46), .Z(G257) ) ;
NOR2    gate705  (.A(G330), .B(G23), .Z(G327) ) ;
NOR2    gate706  (.A(G523), .B(G51), .Z(G362) ) ;
NOR2    gate707  (.A(G375), .B(G52), .Z(G367) ) ;
NOR2    gate708  (.A(G376), .B(G53), .Z(G370) ) ;
NOR2    gate709  (.A(G183), .B(G54), .Z(G381) ) ;
NOR2    gate710  (.A(G394), .B(G55), .Z(G386) ) ;
NOR2    gate711  (.A(G395), .B(G56), .Z(G389) ) ;
NOR2    gate712  (.A(G335), .B(G57), .Z(G399) ) ;
NOR2    gate713  (.A(G412), .B(G58), .Z(G402) ) ;
NOR2    gate714  (.A(G413), .B(G59), .Z(G410) ) ;
NOR2    gate715  (.A(G358), .B(G60), .Z(G418) ) ;
NOR2    gate716  (.A(G431), .B(G61), .Z(G421) ) ;
NOR2    gate717  (.A(G432), .B(G62), .Z(G429) ) ;
NOR2    gate718  (.A(G615), .B(G64), .Z(G444) ) ;
NOR2    gate719  (.A(G615), .B(G66), .Z(G454) ) ;
NOR2    gate720  (.A(G434), .B(G67), .Z(G461) ) ;
NOR2    gate721  (.A(G479), .B(G68), .Z(G466) ) ;
NOR2    gate722  (.A(G480), .B(G69), .Z(G471) ) ;
NOR2    gate723  (.A(G481), .B(G70), .Z(G474) ) ;
NOR2    gate724  (.A(G604), .B(G74), .Z(G528) ) ;
NOR2    gate725  (.A(G550), .B(G75), .Z(G533) ) ;
NOR2    gate726  (.A(G551), .B(G76), .Z(G538) ) ;
NOR2    gate727  (.A(G552), .B(G77), .Z(G543) ) ;
NOR2    gate728  (.A(G553), .B(G78), .Z(G546) ) ;
NOR2    gate729  (.A(G658), .B(G86), .Z(G660) ) ;
NOR2    gate730  (.A(G678), .B(G94), .Z(G710) ) ;

endmodule
