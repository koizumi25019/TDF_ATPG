module s13207 (g43, g49, g633, g634, g635
    , g645, g647, g648, g690, g694
    , g698, g702, g722, g723, g751
    , g752, g753, g754, g755, g756
    , g757, g781, g941, g962, g1000
    , g1008, g1016, g1080, g1234, g1553
    , g1554, CLK
    , g206, g291, g372, g453, g534
    , g594, g785, g1006, g1015, g1017
    , g1246, g1724, g1783, g1798, g1804
    , g1810, g1817, g1824, g1829, g1870
    , g1871, g1894, g1911, g1944, g2662
    , g2844, g2888, g3077, g3096, g3130
    , g3159, g3191, g3829, g3859, g3860
    , g4267, g4316, g4370, g4371, g4372
    , g4373, g4655, g4657, g4660, g4661
    , g4663, g4664, g5143, g5164, g5571
    , g5669, g5678, g5682, g5684, g5687
    , g5729, g6207, g6212, g6223, g6236
    , g6269, g6425, g6648, g6653, g6675
    , g6849, g6850, g6895, g6909, g7048
    , g7063, g7103, g7283, g7284, g7285
    , g7286, g7287, g7288, g7289, g7290
    , g7291, g7292, g7293, g7294, g7295
    , g7298, g7423, g7424, g7425, g7474
    , g7504, g7505, g7506, g7507, g7508
    , g7514, g7729, g7730, g7731, g7732
    , g8216, g8217, g8218, g8219, g8234
    , g8661, g8663, g8872, g8958, g9128
    , g9132, g9204, g9280, g9297, g9299
    , g9305, g9308, g9310, g9312, g9314
    , g9378) ;

input   g43, g49, g633, g634, g635
    , g645, g647, g648, g690, g694
    , g698, g702, g722, g723, g751
    , g752, g753, g754, g755, g756
    , g757, g781, g941, g962, g1000
    , g1008, g1016, g1080, g1234, g1553
    , g1554, CLK ;

output  g206, g291, g372, g453, g534
    , g594, g785, g1006, g1015, g1017
    , g1246, g1724, g1783, g1798, g1804
    , g1810, g1817, g1824, g1829, g1870
    , g1871, g1894, g1911, g1944, g2662
    , g2844, g2888, g3077, g3096, g3130
    , g3159, g3191, g3829, g3859, g3860
    , g4267, g4316, g4370, g4371, g4372
    , g4373, g4655, g4657, g4660, g4661
    , g4663, g4664, g5143, g5164, g5571
    , g5669, g5678, g5682, g5684, g5687
    , g5729, g6207, g6212, g6223, g6236
    , g6269, g6425, g6648, g6653, g6675
    , g6849, g6850, g6895, g6909, g7048
    , g7063, g7103, g7283, g7284, g7285
    , g7286, g7287, g7288, g7289, g7290
    , g7291, g7292, g7293, g7294, g7295
    , g7298, g7423, g7424, g7425, g7474
    , g7504, g7505, g7506, g7507, g7508
    , g7514, g7729, g7730, g7731, g7732
    , g8216, g8217, g8218, g8219, g8234
    , g8661, g8663, g8872, g8958, g9128
    , g9132, g9204, g9280, g9297, g9299
    , g9305, g9308, g9310, g9312, g9314
    , g9378 ;

INV     gate0  (.A(II5353), .Z(g206) ) ;
INV     gate1  (.A(II5356), .Z(g291) ) ;
INV     gate2  (.A(II5359), .Z(g372) ) ;
INV     gate3  (.A(II5362), .Z(g453) ) ;
INV     gate4  (.A(II5365), .Z(g534) ) ;
INV     gate5  (.A(II5368), .Z(g594) ) ;
INV     gate6  (.A(II5407), .Z(g785) ) ;
INV     gate7  (.A(II5410), .Z(g1006) ) ;
INV     gate8  (.A(II5416), .Z(g1015) ) ;
INV     gate9  (.A(II5419), .Z(g1017) ) ;
INV     gate10  (.A(II5425), .Z(g1246) ) ;
INV     gate11  (.A(II5568), .Z(g1724) ) ;
INV     gate12  (.A(II5633), .Z(g1783) ) ;
INV     gate13  (.A(II5654), .Z(g1798) ) ;
INV     gate14  (.A(II5664), .Z(g1804) ) ;
INV     gate15  (.A(II5676), .Z(g1810) ) ;
INV     gate16  (.A(II5689), .Z(g1817) ) ;
INV     gate17  (.A(II5706), .Z(g1824) ) ;
INV     gate18  (.A(II5715), .Z(g1829) ) ;
INV     gate19  (.A(II5751), .Z(g1870) ) ;
INV     gate20  (.A(II5754), .Z(g1871) ) ;
INV     gate21  (.A(II5772), .Z(g1894) ) ;
INV     gate22  (.A(II5789), .Z(g1911) ) ;
INV     gate23  (.A(II5817), .Z(g1944) ) ;
INV     gate24  (.A(II6457), .Z(g2662) ) ;
INV     gate25  (.A(II6574), .Z(g2844) ) ;
INV     gate26  (.A(II6608), .Z(g2888) ) ;
INV     gate27  (.A(II6805), .Z(g3077) ) ;
INV     gate28  (.A(II6834), .Z(g3096) ) ;
INV     gate29  (.A(II6849), .Z(g3130) ) ;
INV     gate30  (.A(II6856), .Z(g3159) ) ;
INV     gate31  (.A(II6868), .Z(g3191) ) ;
INV     gate32  (.A(II7290), .Z(g3829) ) ;
INV     gate33  (.A(II7380), .Z(g3859) ) ;
INV     gate34  (.A(II7383), .Z(g3860) ) ;
INV     gate35  (.A(II8205), .Z(g4267) ) ;
INV     gate36  (.A(II8291), .Z(g4316) ) ;
INV     gate37  (.A(II8351), .Z(g4370) ) ;
INV     gate38  (.A(II8354), .Z(g4371) ) ;
INV     gate39  (.A(II8357), .Z(g4372) ) ;
INV     gate40  (.A(II8360), .Z(g4373) ) ;
INV     gate41  (.A(II8880), .Z(g4655) ) ;
INV     gate42  (.A(II8886), .Z(g4657) ) ;
INV     gate43  (.A(II8895), .Z(g4660) ) ;
INV     gate44  (.A(II8898), .Z(g4661) ) ;
INV     gate45  (.A(II8904), .Z(g4663) ) ;
INV     gate46  (.A(II8907), .Z(g4664) ) ;
INV     gate47  (.A(II9555), .Z(g5143) ) ;
INV     gate48  (.A(II9618), .Z(g5164) ) ;
INV     gate49  (.A(II10032), .Z(g5571) ) ;
INV     gate50  (.A(II10154), .Z(g5669) ) ;
INV     gate51  (.A(II10169), .Z(g5678) ) ;
INV     gate52  (.A(II10177), .Z(g5682) ) ;
INV     gate53  (.A(II10183), .Z(g5684) ) ;
INV     gate54  (.A(II10190), .Z(g5687) ) ;
INV     gate55  (.A(g5144), .Z(g5729) ) ;
INV     gate56  (.A(II10962), .Z(g6207) ) ;
INV     gate57  (.A(II10973), .Z(g6212) ) ;
INV     gate58  (.A(II11008), .Z(g6223) ) ;
INV     gate59  (.A(II11037), .Z(g6236) ) ;
INV     gate60  (.A(II11090), .Z(g6269) ) ;
INV     gate61  (.A(II11556), .Z(g6425) ) ;
INV     gate62  (.A(II11926), .Z(g6648) ) ;
INV     gate63  (.A(II11939), .Z(g6653) ) ;
INV     gate64  (.A(II11981), .Z(g6675) ) ;
INV     gate65  (.A(II12418), .Z(g6849) ) ;
INV     gate66  (.A(II12421), .Z(g6850) ) ;
INV     gate67  (.A(II12558), .Z(g6895) ) ;
INV     gate68  (.A(II12592), .Z(g6909) ) ;
INV     gate69  (.A(II12810), .Z(g7048) ) ;
INV     gate70  (.A(II12826), .Z(g7063) ) ;
INV     gate71  (.A(II12897), .Z(g7103) ) ;
INV     gate72  (.A(II13281), .Z(g7283) ) ;
INV     gate73  (.A(II13284), .Z(g7284) ) ;
INV     gate74  (.A(II13287), .Z(g7285) ) ;
INV     gate75  (.A(II13290), .Z(g7286) ) ;
INV     gate76  (.A(II13293), .Z(g7287) ) ;
INV     gate77  (.A(II13296), .Z(g7288) ) ;
INV     gate78  (.A(II13299), .Z(g7289) ) ;
INV     gate79  (.A(II13302), .Z(g7290) ) ;
INV     gate80  (.A(II13305), .Z(g7291) ) ;
INV     gate81  (.A(II13308), .Z(g7292) ) ;
INV     gate82  (.A(II13311), .Z(g7293) ) ;
INV     gate83  (.A(II13314), .Z(g7294) ) ;
INV     gate84  (.A(II13317), .Z(g7295) ) ;
INV     gate85  (.A(II13326), .Z(g7298) ) ;
INV     gate86  (.A(II13544), .Z(g7423) ) ;
INV     gate87  (.A(II13547), .Z(g7424) ) ;
INV     gate88  (.A(II13550), .Z(g7425) ) ;
INV     gate89  (.A(II13628), .Z(g7474) ) ;
INV     gate90  (.A(II13692), .Z(g7504) ) ;
INV     gate91  (.A(II13695), .Z(g7505) ) ;
INV     gate92  (.A(II13698), .Z(g7506) ) ;
INV     gate93  (.A(II13701), .Z(g7507) ) ;
INV     gate94  (.A(II13704), .Z(g7508) ) ;
INV     gate95  (.A(II13722), .Z(g7514) ) ;
INV     gate96  (.A(II14058), .Z(g7729) ) ;
INV     gate97  (.A(II14061), .Z(g7730) ) ;
INV     gate98  (.A(II14064), .Z(g7731) ) ;
INV     gate99  (.A(II14067), .Z(g7732) ) ;
INV     gate100  (.A(II14427), .Z(g8216) ) ;
INV     gate101  (.A(II14430), .Z(g8217) ) ;
INV     gate102  (.A(II14433), .Z(g8218) ) ;
INV     gate103  (.A(II14436), .Z(g8219) ) ;
INV     gate104  (.A(II14489), .Z(g8234) ) ;
INV     gate105  (.A(II14777), .Z(g8661) ) ;
INV     gate106  (.A(II14783), .Z(g8663) ) ;
INV     gate107  (.A(II15202), .Z(g8872) ) ;
INV     gate108  (.A(II15388), .Z(g8958) ) ;
INV     gate109  (.A(II15762), .Z(g9128) ) ;
INV     gate110  (.A(II15770), .Z(g9132) ) ;
INV     gate111  (.A(II15894), .Z(g9204) ) ;
INV     gate112  (.A(II16006), .Z(g9280) ) ;
INV     gate113  (.A(II16017), .Z(g9297) ) ;
INV     gate114  (.A(II16023), .Z(g9299) ) ;
INV     gate115  (.A(II16033), .Z(g9305) ) ;
INV     gate116  (.A(II16040), .Z(g9308) ) ;
INV     gate117  (.A(II16046), .Z(g9310) ) ;
INV     gate118  (.A(II16052), .Z(g9312) ) ;
INV     gate119  (.A(II16058), .Z(g9314) ) ;
INV     gate120  (.A(II16158), .Z(g9378) ) ;
INV     gate121  (.A(II11233), .Z(g6302) ) ;
DFF     gate122  (.D(g6302), .CP(CLK), .Q(g31) ) ;
INV     gate123  (.A(II11230), .Z(g6301) ) ;
DFF     gate124  (.D(g6301), .CP(CLK), .Q(g30) ) ;
INV     gate125  (.A(II11227), .Z(g6300) ) ;
DFF     gate126  (.D(g6300), .CP(CLK), .Q(g29) ) ;
INV     gate127  (.A(II11221), .Z(g6298) ) ;
DFF     gate128  (.D(g6298), .CP(CLK), .Q(g28) ) ;
INV     gate129  (.A(II11218), .Z(g6297) ) ;
DFF     gate130  (.D(g6297), .CP(CLK), .Q(g27) ) ;
INV     gate131  (.A(II11215), .Z(g6296) ) ;
DFF     gate132  (.D(g6296), .CP(CLK), .Q(g26) ) ;
INV     gate133  (.A(II11212), .Z(g6295) ) ;
DFF     gate134  (.D(g6295), .CP(CLK), .Q(g25) ) ;
INV     gate135  (.A(II11209), .Z(g6294) ) ;
DFF     gate136  (.D(g6294), .CP(CLK), .Q(g24) ) ;
INV     gate137  (.A(II11206), .Z(g6293) ) ;
DFF     gate138  (.D(g6293), .CP(CLK), .Q(g23) ) ;
INV     gate139  (.A(II11203), .Z(g6292) ) ;
DFF     gate140  (.D(g6292), .CP(CLK), .Q(g22) ) ;
INV     gate141  (.A(II14780), .Z(g8662) ) ;
DFF     gate142  (.D(g8662), .CP(CLK), .Q(g12) ) ;
INV     gate143  (.A(II11197), .Z(g6290) ) ;
DFF     gate144  (.D(g6290), .CP(CLK), .Q(g11) ) ;
INV     gate145  (.A(II11191), .Z(g6288) ) ;
DFF     gate146  (.D(g6288), .CP(CLK), .Q(g9) ) ;
INV     gate147  (.A(II16154), .Z(g9376) ) ;
DFF     gate148  (.D(g9376), .CP(CLK), .Q(g8) ) ;
INV     gate149  (.A(II16151), .Z(g9375) ) ;
DFF     gate150  (.D(g9375), .CP(CLK), .Q(g7) ) ;
INV     gate151  (.A(II16148), .Z(g9374) ) ;
DFF     gate152  (.D(g9374), .CP(CLK), .Q(g6) ) ;
INV     gate153  (.A(II16145), .Z(g9373) ) ;
DFF     gate154  (.D(g9373), .CP(CLK), .Q(g5) ) ;
INV     gate155  (.A(II16142), .Z(g9372) ) ;
DFF     gate156  (.D(g9372), .CP(CLK), .Q(g4) ) ;
INV     gate157  (.A(II16119), .Z(g9361) ) ;
DFF     gate158  (.D(g9361), .CP(CLK), .Q(g2) ) ;
INV     gate159  (.A(II16116), .Z(g9360) ) ;
DFF     gate160  (.D(g9360), .CP(CLK), .Q(g3) ) ;
INV     gate161  (.A(II16122), .Z(g9362) ) ;
DFF     gate162  (.D(g9362), .CP(CLK), .Q(g48) ) ;
INV     gate163  (.A(II11224), .Z(g6299) ) ;
DFF     gate164  (.D(g6299), .CP(CLK), .Q(g21) ) ;
INV     gate165  (.A(II11200), .Z(g6291) ) ;
DFF     gate166  (.D(g6291), .CP(CLK), .Q(g10) ) ;
INV     gate167  (.A(II11194), .Z(g6289) ) ;
DFF     gate168  (.D(g6289), .CP(CLK), .Q(g1) ) ;
INV     gate169  (.A(II16183), .Z(g9389) ) ;
DFF     gate170  (.D(g9389), .CP(CLK), .Q(g47) ) ;
INV     gate171  (.A(II15379), .Z(g8955) ) ;
DFF     gate172  (.D(g8955), .CP(CLK), .Q(g46) ) ;
INV     gate173  (.A(II11251), .Z(g6308) ) ;
DFF     gate174  (.D(g6308), .CP(CLK), .Q(g45) ) ;
INV     gate175  (.A(II11248), .Z(g6307) ) ;
DFF     gate176  (.D(g6307), .CP(CLK), .Q(g44) ) ;
INV     gate177  (.A(II11245), .Z(g6306) ) ;
DFF     gate178  (.D(g6306), .CP(CLK), .Q(g42) ) ;
INV     gate179  (.A(II11242), .Z(g6305) ) ;
DFF     gate180  (.D(g6305), .CP(CLK), .Q(g41) ) ;
INV     gate181  (.A(II11239), .Z(g6304) ) ;
DFF     gate182  (.D(g6304), .CP(CLK), .Q(g37) ) ;
INV     gate183  (.A(II11236), .Z(g6303) ) ;
DFF     gate184  (.D(g6303), .CP(CLK), .Q(g32) ) ;
INV     gate185  (.A(II9645), .Z(g5173) ) ;
DFF     gate186  (.D(g5173), .CP(CLK), .Q(g1207) ) ;
INV     gate187  (.A(II9648), .Z(g5174) ) ;
DFF     gate188  (.D(g5174), .CP(CLK), .Q(g1211) ) ;
INV     gate189  (.A(II10265), .Z(g5736) ) ;
DFF     gate190  (.D(g5736), .CP(CLK), .Q(g1214) ) ;
INV     gate191  (.A(II11458), .Z(g6377) ) ;
DFF     gate192  (.D(g6377), .CP(CLK), .Q(g1217) ) ;
INV     gate193  (.A(II11461), .Z(g6378) ) ;
DFF     gate194  (.D(g6378), .CP(CLK), .Q(g1220) ) ;
INV     gate195  (.A(II11464), .Z(g6379) ) ;
DFF     gate196  (.D(g6379), .CP(CLK), .Q(g1223) ) ;
INV     gate197  (.A(II12442), .Z(g6857) ) ;
DFF     gate198  (.D(g6857), .CP(CLK), .Q(g1224) ) ;
INV     gate199  (.A(II12445), .Z(g6858) ) ;
DFF     gate200  (.D(g6858), .CP(CLK), .Q(g1225) ) ;
INV     gate201  (.A(II12448), .Z(g6859) ) ;
DFF     gate202  (.D(g6859), .CP(CLK), .Q(g1226) ) ;
INV     gate203  (.A(II12912), .Z(g7108) ) ;
DFF     gate204  (.D(g7108), .CP(CLK), .Q(g1227) ) ;
INV     gate205  (.A(II12915), .Z(g7109) ) ;
DFF     gate206  (.D(g7109), .CP(CLK), .Q(g1228) ) ;
INV     gate207  (.A(II12918), .Z(g7110) ) ;
DFF     gate208  (.D(g7110), .CP(CLK), .Q(g1229) ) ;
INV     gate209  (.A(II13332), .Z(g7300) ) ;
DFF     gate210  (.D(g7300), .CP(CLK), .Q(g1230) ) ;
INV     gate211  (.A(II5422), .Z(g1235) ) ;
DFF     gate212  (.D(g1235), .CP(CLK), .Q(g1240) ) ;
DFF     gate213  (.D(g1240), .CP(CLK), .Q(g1236) ) ;
DFF     gate214  (.D(g1236), .CP(CLK), .Q(g1231) ) ;
INV     gate215  (.A(g1655), .Z(g2659) ) ;
DFF     gate216  (.D(g2659), .CP(CLK), .Q(g1244) ) ;
DFF     gate217  (.D(g1244), .CP(CLK), .Q(g1245) ) ;
INV     gate218  (.A(II6451), .Z(g2660) ) ;
DFF     gate219  (.D(g2660), .CP(CLK), .Q(g1243) ) ;
INV     gate220  (.A(II11476), .Z(g6383) ) ;
DFF     gate221  (.D(g6383), .CP(CLK), .Q(g1272) ) ;
INV     gate222  (.A(II11479), .Z(g6384) ) ;
DFF     gate223  (.D(g6384), .CP(CLK), .Q(g1276) ) ;
INV     gate224  (.A(II12924), .Z(g7112) ) ;
DFF     gate225  (.D(g7112), .CP(CLK), .Q(g1280) ) ;
INV     gate226  (.A(II13335), .Z(g7301) ) ;
DFF     gate227  (.D(g7301), .CP(CLK), .Q(g1284) ) ;
INV     gate228  (.A(II13761), .Z(g7527) ) ;
DFF     gate229  (.D(g7527), .CP(CLK), .Q(g1288) ) ;
INV     gate230  (.A(II13338), .Z(g7302) ) ;
DFF     gate231  (.D(g7302), .CP(CLK), .Q(g1292) ) ;
INV     gate232  (.A(II13341), .Z(g7303) ) ;
DFF     gate233  (.D(g7303), .CP(CLK), .Q(g1300) ) ;
INV     gate234  (.A(II13344), .Z(g7304) ) ;
DFF     gate235  (.D(g7304), .CP(CLK), .Q(g1296) ) ;
INV     gate236  (.A(II10280), .Z(g5741) ) ;
DFF     gate237  (.D(g5741), .CP(CLK), .Q(g1253) ) ;
INV     gate238  (.A(II11482), .Z(g6385) ) ;
DFF     gate239  (.D(g6385), .CP(CLK), .Q(g1308) ) ;
DFF     gate240  (.D(g1308), .CP(CLK), .Q(g1309) ) ;
DFF     gate241  (.D(g1309), .CP(CLK), .Q(g1310) ) ;
DFF     gate242  (.D(g1310), .CP(CLK), .Q(g1311) ) ;
DFF     gate243  (.D(g1311), .CP(CLK), .Q(g1312) ) ;
DFF     gate244  (.D(g1312), .CP(CLK), .Q(g1304) ) ;
INV     gate245  (.A(II7377), .Z(g3858) ) ;
DFF     gate246  (.D(g3858), .CP(CLK), .Q(g1307) ) ;
INV     gate247  (.A(II12457), .Z(g6862) ) ;
DFF     gate248  (.D(g6862), .CP(CLK), .Q(g1330) ) ;
INV     gate249  (.A(II12460), .Z(g6863) ) ;
DFF     gate250  (.D(g6863), .CP(CLK), .Q(g1333) ) ;
INV     gate251  (.A(II12463), .Z(g6864) ) ;
DFF     gate252  (.D(g6864), .CP(CLK), .Q(g1336) ) ;
INV     gate253  (.A(II12466), .Z(g6865) ) ;
DFF     gate254  (.D(g6865), .CP(CLK), .Q(g1339) ) ;
INV     gate255  (.A(II12945), .Z(g7119) ) ;
DFF     gate256  (.D(g7119), .CP(CLK), .Q(g1342) ) ;
INV     gate257  (.A(II13764), .Z(g7528) ) ;
DFF     gate258  (.D(g7528), .CP(CLK), .Q(g1345) ) ;
INV     gate259  (.A(II13767), .Z(g7529) ) ;
DFF     gate260  (.D(g7529), .CP(CLK), .Q(g1348) ) ;
INV     gate261  (.A(II13770), .Z(g7530) ) ;
DFF     gate262  (.D(g7530), .CP(CLK), .Q(g1351) ) ;
INV     gate263  (.A(II14175), .Z(g7768) ) ;
DFF     gate264  (.D(g7768), .CP(CLK), .Q(g1354) ) ;
INV     gate265  (.A(II14819), .Z(g8675) ) ;
DFF     gate266  (.D(g8675), .CP(CLK), .Q(g1357) ) ;
INV     gate267  (.A(II14822), .Z(g8676) ) ;
DFF     gate268  (.D(g8676), .CP(CLK), .Q(g1360) ) ;
INV     gate269  (.A(II14825), .Z(g8677) ) ;
DFF     gate270  (.D(g8677), .CP(CLK), .Q(g1190) ) ;
INV     gate271  (.A(II11446), .Z(g6373) ) ;
DFF     gate272  (.D(g6373), .CP(CLK), .Q(g1191) ) ;
DFF     gate273  (.D(g1191), .CP(CLK), .Q(g1192) ) ;
DFF     gate274  (.D(g1192), .CP(CLK), .Q(g1193) ) ;
DFF     gate275  (.D(g1193), .CP(CLK), .Q(g1194) ) ;
INV     gate276  (.A(II11449), .Z(g6374) ) ;
DFF     gate277  (.D(g6374), .CP(CLK), .Q(g1195) ) ;
DFF     gate278  (.D(g1195), .CP(CLK), .Q(g1196) ) ;
DFF     gate279  (.D(g1196), .CP(CLK), .Q(g1197) ) ;
DFF     gate280  (.D(g1197), .CP(CLK), .Q(g1198) ) ;
INV     gate281  (.A(II11452), .Z(g6375) ) ;
DFF     gate282  (.D(g6375), .CP(CLK), .Q(g1199) ) ;
DFF     gate283  (.D(g1199), .CP(CLK), .Q(g1200) ) ;
DFF     gate284  (.D(g1200), .CP(CLK), .Q(g1201) ) ;
DFF     gate285  (.D(g1201), .CP(CLK), .Q(g1202) ) ;
INV     gate286  (.A(II11455), .Z(g6376) ) ;
DFF     gate287  (.D(g6376), .CP(CLK), .Q(g1203) ) ;
DFF     gate288  (.D(g1203), .CP(CLK), .Q(g1204) ) ;
DFF     gate289  (.D(g1204), .CP(CLK), .Q(g1205) ) ;
DFF     gate290  (.D(g1205), .CP(CLK), .Q(g1206) ) ;
INV     gate291  (.A(II6454), .Z(g2661) ) ;
DFF     gate292  (.D(g2661), .CP(CLK), .Q(g1252) ) ;
INV     gate293  (.A(II12921), .Z(g7111) ) ;
DFF     gate294  (.D(g7111), .CP(CLK), .Q(g1250) ) ;
INV     gate295  (.A(II12451), .Z(g6860) ) ;
DFF     gate296  (.D(g6860), .CP(CLK), .Q(g1251) ) ;
INV     gate297  (.A(II11467), .Z(g6380) ) ;
DFF     gate298  (.D(g6380), .CP(CLK), .Q(g1247) ) ;
INV     gate299  (.A(II11470), .Z(g6381) ) ;
DFF     gate300  (.D(g6381), .CP(CLK), .Q(g1254) ) ;
INV     gate301  (.A(II10274), .Z(g5739) ) ;
DFF     gate302  (.D(g5739), .CP(CLK), .Q(g1266) ) ;
INV     gate303  (.A(II11473), .Z(g6382) ) ;
DFF     gate304  (.D(g6382), .CP(CLK), .Q(g1260) ) ;
INV     gate305  (.A(II10271), .Z(g5738) ) ;
DFF     gate306  (.D(g5738), .CP(CLK), .Q(g1257) ) ;
INV     gate307  (.A(II10268), .Z(g5737) ) ;
DFF     gate308  (.D(g5737), .CP(CLK), .Q(g1263) ) ;
INV     gate309  (.A(II8883), .Z(g4656) ) ;
DFF     gate310  (.D(g4656), .CP(CLK), .Q(g1267) ) ;
INV     gate311  (.A(II9651), .Z(g5175) ) ;
DFF     gate312  (.D(g5175), .CP(CLK), .Q(g1268) ) ;
INV     gate313  (.A(II10277), .Z(g5740) ) ;
DFF     gate314  (.D(g5740), .CP(CLK), .Q(g1269) ) ;
INV     gate315  (.A(II9654), .Z(g5176) ) ;
DFF     gate316  (.D(g5176), .CP(CLK), .Q(g1271) ) ;
DFF     gate317  (.D(g1271), .CP(CLK), .Q(g1270) ) ;
DFF     gate318  (.D(g1270), .CP(CLK), .Q(g172) ) ;
INV     gate319  (.A(II10283), .Z(g5742) ) ;
DFF     gate320  (.D(g5742), .CP(CLK), .Q(g1313) ) ;
INV     gate321  (.A(II10286), .Z(g5743) ) ;
DFF     gate322  (.D(g5743), .CP(CLK), .Q(g1317) ) ;
INV     gate323  (.A(II12454), .Z(g6861) ) ;
DFF     gate324  (.D(g6861), .CP(CLK), .Q(g1318) ) ;
INV     gate325  (.A(II12927), .Z(g7113) ) ;
DFF     gate326  (.D(g7113), .CP(CLK), .Q(g1319) ) ;
INV     gate327  (.A(II12930), .Z(g7114) ) ;
DFF     gate328  (.D(g7114), .CP(CLK), .Q(g1320) ) ;
INV     gate329  (.A(II12933), .Z(g7115) ) ;
DFF     gate330  (.D(g7115), .CP(CLK), .Q(g1321) ) ;
INV     gate331  (.A(II12936), .Z(g7116) ) ;
DFF     gate332  (.D(g7116), .CP(CLK), .Q(g1322) ) ;
INV     gate333  (.A(II12939), .Z(g7117) ) ;
DFF     gate334  (.D(g7117), .CP(CLK), .Q(g1323) ) ;
INV     gate335  (.A(II12942), .Z(g7118) ) ;
DFF     gate336  (.D(g7118), .CP(CLK), .Q(g1324) ) ;
INV     gate337  (.A(II13347), .Z(g7305) ) ;
DFF     gate338  (.D(g7305), .CP(CLK), .Q(g1325) ) ;
INV     gate339  (.A(II13350), .Z(g7306) ) ;
DFF     gate340  (.D(g7306), .CP(CLK), .Q(g1326) ) ;
INV     gate341  (.A(II13353), .Z(g7307) ) ;
DFF     gate342  (.D(g7307), .CP(CLK), .Q(g1327) ) ;
INV     gate343  (.A(II13359), .Z(g7309) ) ;
DFF     gate344  (.D(g7309), .CP(CLK), .Q(g1328) ) ;
INV     gate345  (.A(II13356), .Z(g7308) ) ;
DFF     gate346  (.D(g7308), .CP(CLK), .Q(g13) ) ;
INV     gate347  (.A(II6460), .Z(g2663) ) ;
DFF     gate348  (.D(g2663), .CP(CLK), .Q(g1329) ) ;
INV     gate349  (.A(II11485), .Z(g6386) ) ;
DFF     gate350  (.D(g6386), .CP(CLK), .Q(g20) ) ;
INV     gate351  (.A(II12469), .Z(g6866) ) ;
DFF     gate352  (.D(g6866), .CP(CLK), .Q(g1366) ) ;
INV     gate353  (.A(II12505), .Z(g6878) ) ;
DFF     gate354  (.D(g6878), .CP(CLK), .Q(g1364) ) ;
INV     gate355  (.A(II12499), .Z(g6876) ) ;
DFF     gate356  (.D(g6876), .CP(CLK), .Q(g1370) ) ;
INV     gate357  (.A(II12493), .Z(g6874) ) ;
DFF     gate358  (.D(g6874), .CP(CLK), .Q(g1368) ) ;
INV     gate359  (.A(II12487), .Z(g6872) ) ;
DFF     gate360  (.D(g6872), .CP(CLK), .Q(g1374) ) ;
INV     gate361  (.A(II12481), .Z(g6870) ) ;
DFF     gate362  (.D(g6870), .CP(CLK), .Q(g1372) ) ;
INV     gate363  (.A(II12478), .Z(g6869) ) ;
DFF     gate364  (.D(g6869), .CP(CLK), .Q(g1375) ) ;
INV     gate365  (.A(II12472), .Z(g6867) ) ;
DFF     gate366  (.D(g6867), .CP(CLK), .Q(g1365) ) ;
INV     gate367  (.A(II12502), .Z(g6877) ) ;
DFF     gate368  (.D(g6877), .CP(CLK), .Q(g1363) ) ;
INV     gate369  (.A(II12496), .Z(g6875) ) ;
DFF     gate370  (.D(g6875), .CP(CLK), .Q(g1369) ) ;
INV     gate371  (.A(II12490), .Z(g6873) ) ;
DFF     gate372  (.D(g6873), .CP(CLK), .Q(g1367) ) ;
INV     gate373  (.A(II12484), .Z(g6871) ) ;
DFF     gate374  (.D(g6871), .CP(CLK), .Q(g1373) ) ;
INV     gate375  (.A(II12475), .Z(g6868) ) ;
DFF     gate376  (.D(g6868), .CP(CLK), .Q(g1371) ) ;
INV     gate377  (.A(II8889), .Z(g4658) ) ;
DFF     gate378  (.D(g4658), .CP(CLK), .Q(g1389) ) ;
INV     gate379  (.A(II12508), .Z(g6879) ) ;
DFF     gate380  (.D(g6879), .CP(CLK), .Q(g1379) ) ;
INV     gate381  (.A(II12544), .Z(g6891) ) ;
DFF     gate382  (.D(g6891), .CP(CLK), .Q(g1377) ) ;
INV     gate383  (.A(II12538), .Z(g6889) ) ;
DFF     gate384  (.D(g6889), .CP(CLK), .Q(g1383) ) ;
INV     gate385  (.A(II12532), .Z(g6887) ) ;
DFF     gate386  (.D(g6887), .CP(CLK), .Q(g1381) ) ;
INV     gate387  (.A(II12526), .Z(g6885) ) ;
DFF     gate388  (.D(g6885), .CP(CLK), .Q(g1387) ) ;
INV     gate389  (.A(II12520), .Z(g6883) ) ;
DFF     gate390  (.D(g6883), .CP(CLK), .Q(g1385) ) ;
INV     gate391  (.A(II12517), .Z(g6882) ) ;
DFF     gate392  (.D(g6882), .CP(CLK), .Q(g1388) ) ;
INV     gate393  (.A(II12511), .Z(g6880) ) ;
DFF     gate394  (.D(g6880), .CP(CLK), .Q(g1378) ) ;
INV     gate395  (.A(II12541), .Z(g6890) ) ;
DFF     gate396  (.D(g6890), .CP(CLK), .Q(g1376) ) ;
INV     gate397  (.A(II12535), .Z(g6888) ) ;
DFF     gate398  (.D(g6888), .CP(CLK), .Q(g1382) ) ;
INV     gate399  (.A(II12529), .Z(g6886) ) ;
DFF     gate400  (.D(g6886), .CP(CLK), .Q(g1380) ) ;
INV     gate401  (.A(II12523), .Z(g6884) ) ;
DFF     gate402  (.D(g6884), .CP(CLK), .Q(g1386) ) ;
INV     gate403  (.A(II12514), .Z(g6881) ) ;
DFF     gate404  (.D(g6881), .CP(CLK), .Q(g1384) ) ;
INV     gate405  (.A(II8892), .Z(g4659) ) ;
DFF     gate406  (.D(g4659), .CP(CLK), .Q(g1390) ) ;
DFF     gate407  (.D(g1390), .CP(CLK), .Q(g1391) ) ;
INV     gate408  (.A(II11488), .Z(g6387) ) ;
DFF     gate409  (.D(g6387), .CP(CLK), .Q(g1392) ) ;
INV     gate410  (.A(II6463), .Z(g2664) ) ;
DFF     gate411  (.D(g2664), .CP(CLK), .Q(g1393) ) ;
DFF     gate412  (.D(g1393), .CP(CLK), .Q(g1395) ) ;
INV     gate413  (.A(II11491), .Z(g6388) ) ;
DFF     gate414  (.D(g6388), .CP(CLK), .Q(g1394) ) ;
INV     gate415  (.A(II8901), .Z(g4662) ) ;
DFF     gate416  (.D(g4662), .CP(CLK), .Q(g1396) ) ;
DFF     gate417  (.D(g1396), .CP(CLK), .Q(g1398) ) ;
INV     gate418  (.A(II11494), .Z(g6389) ) ;
DFF     gate419  (.D(g6389), .CP(CLK), .Q(g1397) ) ;
INV     gate420  (.A(II7386), .Z(g3861) ) ;
DFF     gate421  (.D(g3861), .CP(CLK), .Q(g1399) ) ;
DFF     gate422  (.D(g1399), .CP(CLK), .Q(g1401) ) ;
INV     gate423  (.A(II11497), .Z(g6390) ) ;
DFF     gate424  (.D(g6390), .CP(CLK), .Q(g1400) ) ;
INV     gate425  (.A(II11500), .Z(g6391) ) ;
DFF     gate426  (.D(g6391), .CP(CLK), .Q(g1402) ) ;
DFF     gate427  (.D(g1402), .CP(CLK), .Q(g1403) ) ;
DFF     gate428  (.D(g1403), .CP(CLK), .Q(g1404) ) ;
DFF     gate429  (.D(g1404), .CP(CLK), .Q(g16) ) ;
INV     gate430  (.A(II11503), .Z(g6392) ) ;
DFF     gate431  (.D(g6392), .CP(CLK), .Q(g1189) ) ;
INV     gate432  (.A(II10292), .Z(g5745) ) ;
DFF     gate433  (.D(g5745), .CP(CLK), .Q(g1412) ) ;
INV     gate434  (.A(II9666), .Z(g5180) ) ;
DFF     gate435  (.D(g5180), .CP(CLK), .Q(g1415) ) ;
INV     gate436  (.A(II9660), .Z(g5178) ) ;
DFF     gate437  (.D(g5178), .CP(CLK), .Q(g1409) ) ;
INV     gate438  (.A(II8910), .Z(g4665) ) ;
DFF     gate439  (.D(g4665), .CP(CLK), .Q(g1416) ) ;
INV     gate440  (.A(II9663), .Z(g5179) ) ;
DFF     gate441  (.D(g5179), .CP(CLK), .Q(g1421) ) ;
INV     gate442  (.A(II10289), .Z(g5744) ) ;
DFF     gate443  (.D(g5744), .CP(CLK), .Q(g1405) ) ;
INV     gate444  (.A(II9657), .Z(g5177) ) ;
DFF     gate445  (.D(g5177), .CP(CLK), .Q(g1408) ) ;
INV     gate446  (.A(II6468), .Z(g2671) ) ;
DFF     gate447  (.D(g2671), .CP(CLK), .Q(g1429) ) ;
INV     gate448  (.A(II6471), .Z(g2672) ) ;
DFF     gate449  (.D(g2672), .CP(CLK), .Q(g1428) ) ;
INV     gate450  (.A(II6474), .Z(g2673) ) ;
DFF     gate451  (.D(g2673), .CP(CLK), .Q(g1431) ) ;
INV     gate452  (.A(II8913), .Z(g4666) ) ;
DFF     gate453  (.D(g4666), .CP(CLK), .Q(g1430) ) ;
INV     gate454  (.A(II7389), .Z(g3862) ) ;
DFF     gate455  (.D(g3862), .CP(CLK), .Q(g1424) ) ;
INV     gate456  (.A(II11506), .Z(g6393) ) ;
DFF     gate457  (.D(g6393), .CP(CLK), .Q(g1524) ) ;
DFF     gate458  (.D(g1524), .CP(CLK), .Q(g1513) ) ;
INV     gate459  (.A(II14457), .Z(g8226) ) ;
DFF     gate460  (.D(g8226), .CP(CLK), .Q(g1486) ) ;
INV     gate461  (.A(II14178), .Z(g7769) ) ;
DFF     gate462  (.D(g7769), .CP(CLK), .Q(g1481) ) ;
INV     gate463  (.A(II14181), .Z(g7770) ) ;
DFF     gate464  (.D(g7770), .CP(CLK), .Q(g1489) ) ;
INV     gate465  (.A(II14184), .Z(g7771) ) ;
DFF     gate466  (.D(g7771), .CP(CLK), .Q(g1494) ) ;
INV     gate467  (.A(II14187), .Z(g7772) ) ;
DFF     gate468  (.D(g7772), .CP(CLK), .Q(g1499) ) ;
INV     gate469  (.A(II14190), .Z(g7773) ) ;
DFF     gate470  (.D(g7773), .CP(CLK), .Q(g1504) ) ;
INV     gate471  (.A(II14193), .Z(g7774) ) ;
DFF     gate472  (.D(g7774), .CP(CLK), .Q(g1509) ) ;
INV     gate473  (.A(II14196), .Z(g7775) ) ;
DFF     gate474  (.D(g7775), .CP(CLK), .Q(g1514) ) ;
INV     gate475  (.A(II14460), .Z(g8227) ) ;
DFF     gate476  (.D(g8227), .CP(CLK), .Q(g1519) ) ;
INV     gate477  (.A(II14828), .Z(g8678) ) ;
DFF     gate478  (.D(g8678), .CP(CLK), .Q(g1462) ) ;
INV     gate479  (.A(II15211), .Z(g8875) ) ;
DFF     gate480  (.D(g8875), .CP(CLK), .Q(g1467) ) ;
INV     gate481  (.A(II15394), .Z(g8960) ) ;
DFF     gate482  (.D(g8960), .CP(CLK), .Q(g1472) ) ;
INV     gate483  (.A(II15522), .Z(g9036) ) ;
DFF     gate484  (.D(g9036), .CP(CLK), .Q(g1477) ) ;
INV     gate485  (.A(II14463), .Z(g8228) ) ;
DFF     gate486  (.D(g8228), .CP(CLK), .Q(g727) ) ;
INV     gate487  (.A(II14214), .Z(g7781) ) ;
DFF     gate488  (.D(g7781), .CP(CLK), .Q(g1532) ) ;
INV     gate489  (.A(II14199), .Z(g7776) ) ;
DFF     gate490  (.D(g7776), .CP(CLK), .Q(g1528) ) ;
INV     gate491  (.A(II14202), .Z(g7777) ) ;
DFF     gate492  (.D(g7777), .CP(CLK), .Q(g1537) ) ;
INV     gate493  (.A(II14205), .Z(g7778) ) ;
DFF     gate494  (.D(g7778), .CP(CLK), .Q(g1541) ) ;
INV     gate495  (.A(II14208), .Z(g7779) ) ;
DFF     gate496  (.D(g7779), .CP(CLK), .Q(g1545) ) ;
INV     gate497  (.A(II14211), .Z(g7780) ) ;
DFF     gate498  (.D(g7780), .CP(CLK), .Q(g1549) ) ;
INV     gate499  (.A(II9669), .Z(g5181) ) ;
DFF     gate500  (.D(g5181), .CP(CLK), .Q(g1435) ) ;
INV     gate501  (.A(II9672), .Z(g5182) ) ;
DFF     gate502  (.D(g5182), .CP(CLK), .Q(g1439) ) ;
INV     gate503  (.A(II9675), .Z(g5183) ) ;
DFF     gate504  (.D(g5183), .CP(CLK), .Q(g1432) ) ;
INV     gate505  (.A(II8916), .Z(g4667) ) ;
DFF     gate506  (.D(g4667), .CP(CLK), .Q(g1443) ) ;
INV     gate507  (.A(II9678), .Z(g5184) ) ;
DFF     gate508  (.D(g5184), .CP(CLK), .Q(g33) ) ;
INV     gate509  (.A(II10295), .Z(g5746) ) ;
DFF     gate510  (.D(g5746), .CP(CLK), .Q(g38) ) ;
INV     gate511  (.A(II8922), .Z(g4669) ) ;
DFF     gate512  (.D(g4669), .CP(CLK), .Q(g1461) ) ;
INV     gate513  (.A(II9681), .Z(g5185) ) ;
DFF     gate514  (.D(g5185), .CP(CLK), .Q(g1444) ) ;
INV     gate515  (.A(II9684), .Z(g5186) ) ;
DFF     gate516  (.D(g5186), .CP(CLK), .Q(g1450) ) ;
INV     gate517  (.A(II9687), .Z(g5187) ) ;
DFF     gate518  (.D(g5187), .CP(CLK), .Q(g1454) ) ;
INV     gate519  (.A(II7392), .Z(g3863) ) ;
DFF     gate520  (.D(g3863), .CP(CLK), .Q(g1459) ) ;
INV     gate521  (.A(II8919), .Z(g4668) ) ;
DFF     gate522  (.D(g4668), .CP(CLK), .Q(g1460) ) ;
INV     gate523  (.A(II12900), .Z(g7104) ) ;
DFF     gate524  (.D(g7104), .CP(CLK), .Q(g979) ) ;
INV     gate525  (.A(II14448), .Z(g8223) ) ;
DFF     gate526  (.D(g8223), .CP(CLK), .Q(g966) ) ;
DFF     gate527  (.D(g966), .CP(CLK), .Q(g969) ) ;
INV     gate528  (.A(II14163), .Z(g7764) ) ;
DFF     gate529  (.D(g7764), .CP(CLK), .Q(g963) ) ;
DFF     gate530  (.D(g963), .CP(CLK), .Q(g970) ) ;
INV     gate531  (.A(II9639), .Z(g5171) ) ;
DFF     gate532  (.D(g5171), .CP(CLK), .Q(g971) ) ;
INV     gate533  (.A(II6443), .Z(g2653) ) ;
DFF     gate534  (.D(g2653), .CP(CLK), .Q(g972) ) ;
INV     gate535  (.A(II14810), .Z(g8672) ) ;
DFF     gate536  (.D(g8672), .CP(CLK), .Q(g973) ) ;
INV     gate537  (.A(II15178), .Z(g8864) ) ;
DFF     gate538  (.D(g8864), .CP(CLK), .Q(g976) ) ;
INV     gate539  (.A(II15773), .Z(g9133) ) ;
DFF     gate540  (.D(g9133), .CP(CLK), .Q(g984) ) ;
INV     gate541  (.A(II13725), .Z(g7515) ) ;
DFF     gate542  (.D(g7515), .CP(CLK), .Q(g985) ) ;
INV     gate543  (.A(II13728), .Z(g7516) ) ;
DFF     gate544  (.D(g7516), .CP(CLK), .Q(g990) ) ;
INV     gate545  (.A(II13731), .Z(g7517) ) ;
DFF     gate546  (.D(g7517), .CP(CLK), .Q(g995) ) ;
INV     gate547  (.A(II12903), .Z(g7105) ) ;
DFF     gate548  (.D(g7105), .CP(CLK), .Q(g1004) ) ;
DFF     gate549  (.D(g1004), .CP(CLK), .Q(g1005) ) ;
DFF     gate550  (.D(g1005), .CP(CLK), .Q(g998) ) ;
INV     gate551  (.A(II15181), .Z(g8865) ) ;
DFF     gate552  (.D(g8865), .CP(CLK), .Q(g999) ) ;
INV     gate553  (.A(II15187), .Z(g8867) ) ;
DFF     gate554  (.D(g8867), .CP(CLK), .Q(g1007) ) ;
INV     gate555  (.A(II12424), .Z(g6851) ) ;
DFF     gate556  (.D(g6851), .CP(CLK), .Q(g1012) ) ;
DFF     gate557  (.D(g1012), .CP(CLK), .Q(g1014) ) ;
DFF     gate558  (.D(g1014), .CP(CLK), .Q(g1013) ) ;
INV     gate559  (.A(II6446), .Z(g2654) ) ;
DFF     gate560  (.D(g2654), .CP(CLK), .Q(g1029) ) ;
INV     gate561  (.A(II15193), .Z(g8869) ) ;
DFF     gate562  (.D(g8869), .CP(CLK), .Q(g1018) ) ;
INV     gate563  (.A(II15196), .Z(g8870) ) ;
DFF     gate564  (.D(g8870), .CP(CLK), .Q(g1021) ) ;
INV     gate565  (.A(II15199), .Z(g8871) ) ;
DFF     gate566  (.D(g8871), .CP(CLK), .Q(g1025) ) ;
INV     gate567  (.A(II15516), .Z(g9034) ) ;
DFF     gate568  (.D(g9034), .CP(CLK), .Q(g1033) ) ;
INV     gate569  (.A(II15385), .Z(g8957) ) ;
DFF     gate570  (.D(g8957), .CP(CLK), .Q(g1034) ) ;
INV     gate571  (.A(II13734), .Z(g7518) ) ;
DFF     gate572  (.D(g7518), .CP(CLK), .Q(g1030) ) ;
INV     gate573  (.A(II12427), .Z(g6852) ) ;
DFF     gate574  (.D(g6852), .CP(CLK), .Q(g1081) ) ;
DFF     gate575  (.D(g1081), .CP(CLK), .Q(g1156) ) ;
DFF     gate576  (.D(g1156), .CP(CLK), .Q(g1157) ) ;
DFF     gate577  (.D(g1157), .CP(CLK), .Q(g1159) ) ;
DFF     gate578  (.D(g1159), .CP(CLK), .Q(g1158) ) ;
INV     gate579  (.A(II12906), .Z(g7106) ) ;
DFF     gate580  (.D(g7106), .CP(CLK), .Q(g1084) ) ;
INV     gate581  (.A(II5475), .Z(g1612) ) ;
DFF     gate582  (.D(g1612), .CP(CLK), .Q(g1146) ) ;
DFF     gate583  (.D(g1146), .CP(CLK), .Q(g1147) ) ;
DFF     gate584  (.D(g1147), .CP(CLK), .Q(g1148) ) ;
INV     gate585  (.A(II12430), .Z(g6853) ) ;
DFF     gate586  (.D(g6853), .CP(CLK), .Q(g1087) ) ;
INV     gate587  (.A(II12433), .Z(g6854) ) ;
DFF     gate588  (.D(g6854), .CP(CLK), .Q(g1098) ) ;
INV     gate589  (.A(II12436), .Z(g6855) ) ;
DFF     gate590  (.D(g6855), .CP(CLK), .Q(g1102) ) ;
INV     gate591  (.A(II12909), .Z(g7107) ) ;
DFF     gate592  (.D(g7107), .CP(CLK), .Q(g1106) ) ;
INV     gate593  (.A(II13329), .Z(g7299) ) ;
DFF     gate594  (.D(g7299), .CP(CLK), .Q(g1110) ) ;
INV     gate595  (.A(II13743), .Z(g7521) ) ;
DFF     gate596  (.D(g7521), .CP(CLK), .Q(g1114) ) ;
INV     gate597  (.A(II14169), .Z(g7766) ) ;
DFF     gate598  (.D(g7766), .CP(CLK), .Q(g1118) ) ;
INV     gate599  (.A(II14454), .Z(g8225) ) ;
DFF     gate600  (.D(g8225), .CP(CLK), .Q(g1122) ) ;
INV     gate601  (.A(II14816), .Z(g8674) ) ;
DFF     gate602  (.D(g8674), .CP(CLK), .Q(g1126) ) ;
INV     gate603  (.A(II15208), .Z(g8874) ) ;
DFF     gate604  (.D(g8874), .CP(CLK), .Q(g1142) ) ;
INV     gate605  (.A(II13758), .Z(g7526) ) ;
DFF     gate606  (.D(g7526), .CP(CLK), .Q(g1173) ) ;
DFF     gate607  (.D(g1173), .CP(CLK), .Q(g1170) ) ;
DFF     gate608  (.D(g1170), .CP(CLK), .Q(g1167) ) ;
DFF     gate609  (.D(g1167), .CP(CLK), .Q(g1166) ) ;
INV     gate610  (.A(II14172), .Z(g7767) ) ;
DFF     gate611  (.D(g7767), .CP(CLK), .Q(g1077) ) ;
INV     gate612  (.A(II12439), .Z(g6856) ) ;
DFF     gate613  (.D(g6856), .CP(CLK), .Q(g1153) ) ;
DFF     gate614  (.D(g1153), .CP(CLK), .Q(g1154) ) ;
DFF     gate615  (.D(g1154), .CP(CLK), .Q(g1155) ) ;
DFF     gate616  (.D(g1155), .CP(CLK), .Q(g1185) ) ;
DFF     gate617  (.D(g1185), .CP(CLK), .Q(g1097) ) ;
INV     gate618  (.A(II13740), .Z(g7520) ) ;
DFF     gate619  (.D(g7520), .CP(CLK), .Q(g1092) ) ;
INV     gate620  (.A(II13746), .Z(g7522) ) ;
DFF     gate621  (.D(g7522), .CP(CLK), .Q(g1130) ) ;
INV     gate622  (.A(II13749), .Z(g7523) ) ;
DFF     gate623  (.D(g7523), .CP(CLK), .Q(g1134) ) ;
INV     gate624  (.A(II13752), .Z(g7524) ) ;
DFF     gate625  (.D(g7524), .CP(CLK), .Q(g1138) ) ;
INV     gate626  (.A(II13755), .Z(g7525) ) ;
DFF     gate627  (.D(g7525), .CP(CLK), .Q(g1149) ) ;
INV     gate628  (.A(II13737), .Z(g7519) ) ;
DFF     gate629  (.D(g7519), .CP(CLK), .Q(g1037) ) ;
INV     gate630  (.A(II14166), .Z(g7765) ) ;
DFF     gate631  (.D(g7765), .CP(CLK), .Q(g1041) ) ;
INV     gate632  (.A(II14451), .Z(g8224) ) ;
DFF     gate633  (.D(g8224), .CP(CLK), .Q(g1045) ) ;
INV     gate634  (.A(II14813), .Z(g8673) ) ;
DFF     gate635  (.D(g8673), .CP(CLK), .Q(g1049) ) ;
INV     gate636  (.A(II15205), .Z(g8873) ) ;
DFF     gate637  (.D(g8873), .CP(CLK), .Q(g1053) ) ;
INV     gate638  (.A(II15391), .Z(g8959) ) ;
DFF     gate639  (.D(g8959), .CP(CLK), .Q(g1057) ) ;
INV     gate640  (.A(II15519), .Z(g9035) ) ;
DFF     gate641  (.D(g9035), .CP(CLK), .Q(g1061) ) ;
INV     gate642  (.A(II15741), .Z(g9117) ) ;
DFF     gate643  (.D(g9117), .CP(CLK), .Q(g1065) ) ;
INV     gate644  (.A(II15776), .Z(g9134) ) ;
DFF     gate645  (.D(g9134), .CP(CLK), .Q(g1069) ) ;
INV     gate646  (.A(II15791), .Z(g9145) ) ;
DFF     gate647  (.D(g9145), .CP(CLK), .Q(g1073) ) ;
INV     gate648  (.A(g1611), .Z(g2655) ) ;
DFF     gate649  (.D(g2655), .CP(CLK), .Q(g1163) ) ;
DFF     gate650  (.D(g1163), .CP(CLK), .Q(g1160) ) ;
DFF     gate651  (.D(g1160), .CP(CLK), .Q(g1182) ) ;
DFF     gate652  (.D(g1182), .CP(CLK), .Q(g1186) ) ;
DFF     gate653  (.D(g1186), .CP(CLK), .Q(g1179) ) ;
INV     gate654  (.A(II9642), .Z(g5172) ) ;
DFF     gate655  (.D(g5172), .CP(CLK), .Q(g1176) ) ;
INV     gate656  (.A(II12193), .Z(g6774) ) ;
DFF     gate657  (.D(g6774), .CP(CLK), .Q(g68) ) ;
INV     gate658  (.A(II12196), .Z(g6775) ) ;
DFF     gate659  (.D(g6775), .CP(CLK), .Q(g71) ) ;
INV     gate660  (.A(II12199), .Z(g6776) ) ;
DFF     gate661  (.D(g6776), .CP(CLK), .Q(g74) ) ;
INV     gate662  (.A(II12202), .Z(g6777) ) ;
DFF     gate663  (.D(g6777), .CP(CLK), .Q(g77) ) ;
INV     gate664  (.A(II12205), .Z(g6778) ) ;
DFF     gate665  (.D(g6778), .CP(CLK), .Q(g80) ) ;
INV     gate666  (.A(II12208), .Z(g6779) ) ;
DFF     gate667  (.D(g6779), .CP(CLK), .Q(g83) ) ;
INV     gate668  (.A(II12211), .Z(g6780) ) ;
DFF     gate669  (.D(g6780), .CP(CLK), .Q(g86) ) ;
INV     gate670  (.A(II12214), .Z(g6781) ) ;
DFF     gate671  (.D(g6781), .CP(CLK), .Q(g52) ) ;
INV     gate672  (.A(II14070), .Z(g7733) ) ;
DFF     gate673  (.D(g7733), .CP(CLK), .Q(g55) ) ;
INV     gate674  (.A(II13707), .Z(g7509) ) ;
DFF     gate675  (.D(g7509), .CP(CLK), .Q(g62) ) ;
INV     gate676  (.A(II14073), .Z(g7734) ) ;
DFF     gate677  (.D(g7734), .CP(CLK), .Q(g58) ) ;
INV     gate678  (.A(II8709), .Z(g4598) ) ;
DFF     gate679  (.D(g4598), .CP(CLK), .Q(g65) ) ;
INV     gate680  (.A(II7299), .Z(g3832) ) ;
DFF     gate681  (.D(g3832), .CP(CLK), .Q(g199) ) ;
DFF     gate682  (.D(g199), .CP(CLK), .Q(g200) ) ;
DFF     gate683  (.D(g200), .CP(CLK), .Q(g201) ) ;
DFF     gate684  (.D(g201), .CP(CLK), .Q(g190) ) ;
INV     gate685  (.A(II7296), .Z(g3831) ) ;
DFF     gate686  (.D(g3831), .CP(CLK), .Q(g195) ) ;
INV     gate687  (.A(II10250), .Z(g5731) ) ;
DFF     gate688  (.D(g5731), .CP(CLK), .Q(g196) ) ;
INV     gate689  (.A(II9603), .Z(g5159) ) ;
DFF     gate690  (.D(g5159), .CP(CLK), .Q(g179) ) ;
INV     gate691  (.A(II7293), .Z(g3830) ) ;
DFF     gate692  (.D(g3830), .CP(CLK), .Q(g186) ) ;
INV     gate693  (.A(II10247), .Z(g5730) ) ;
DFF     gate694  (.D(g5730), .CP(CLK), .Q(g187) ) ;
INV     gate695  (.A(II9600), .Z(g5158) ) ;
DFF     gate696  (.D(g5158), .CP(CLK), .Q(g180) ) ;
INV     gate697  (.A(II7308), .Z(g3835) ) ;
DFF     gate698  (.D(g3835), .CP(CLK), .Q(g205) ) ;
INV     gate699  (.A(II10253), .Z(g5732) ) ;
DFF     gate700  (.D(g5732), .CP(CLK), .Q(g202) ) ;
INV     gate701  (.A(II9606), .Z(g5160) ) ;
DFF     gate702  (.D(g5160), .CP(CLK), .Q(g181) ) ;
INV     gate703  (.A(II7305), .Z(g3834) ) ;
DFF     gate704  (.D(g3834), .CP(CLK), .Q(g210) ) ;
INV     gate705  (.A(II10256), .Z(g5733) ) ;
DFF     gate706  (.D(g5733), .CP(CLK), .Q(g207) ) ;
INV     gate707  (.A(II9609), .Z(g5161) ) ;
DFF     gate708  (.D(g5161), .CP(CLK), .Q(g182) ) ;
INV     gate709  (.A(II14076), .Z(g7735) ) ;
DFF     gate710  (.D(g7735), .CP(CLK), .Q(g146) ) ;
INV     gate711  (.A(II14079), .Z(g7736) ) ;
DFF     gate712  (.D(g7736), .CP(CLK), .Q(g173) ) ;
INV     gate713  (.A(II14085), .Z(g7738) ) ;
DFF     gate714  (.D(g7738), .CP(CLK), .Q(g150) ) ;
INV     gate715  (.A(II14082), .Z(g7737) ) ;
DFF     gate716  (.D(g7737), .CP(CLK), .Q(g174) ) ;
INV     gate717  (.A(II14088), .Z(g7739) ) ;
DFF     gate718  (.D(g7739), .CP(CLK), .Q(g154) ) ;
INV     gate719  (.A(II14091), .Z(g7740) ) ;
DFF     gate720  (.D(g7740), .CP(CLK), .Q(g158) ) ;
INV     gate721  (.A(II14094), .Z(g7741) ) ;
DFF     gate722  (.D(g7741), .CP(CLK), .Q(g162) ) ;
INV     gate723  (.A(II14097), .Z(g7742) ) ;
DFF     gate724  (.D(g7742), .CP(CLK), .Q(g168) ) ;
INV     gate725  (.A(II11254), .Z(g6309) ) ;
DFF     gate726  (.D(g6309), .CP(CLK), .Q(g183) ) ;
INV     gate727  (.A(II11257), .Z(g6310) ) ;
DFF     gate728  (.D(g6310), .CP(CLK), .Q(g184) ) ;
INV     gate729  (.A(II8712), .Z(g4599) ) ;
DFF     gate730  (.D(g4599), .CP(CLK), .Q(g185) ) ;
INV     gate731  (.A(II12253), .Z(g6794) ) ;
DFF     gate732  (.D(g6794), .CP(CLK), .Q(g92) ) ;
DFF     gate733  (.D(g92), .CP(CLK), .Q(g89) ) ;
INV     gate734  (.A(II9561), .Z(g5145) ) ;
DFF     gate735  (.D(g5145), .CP(CLK), .Q(g93) ) ;
INV     gate736  (.A(II12217), .Z(g6782) ) ;
DFF     gate737  (.D(g6782), .CP(CLK), .Q(g94) ) ;
DFF     gate738  (.D(g94), .CP(CLK), .Q(g95) ) ;
INV     gate739  (.A(II9564), .Z(g5146) ) ;
DFF     gate740  (.D(g5146), .CP(CLK), .Q(g98) ) ;
INV     gate741  (.A(II12220), .Z(g6783) ) ;
DFF     gate742  (.D(g6783), .CP(CLK), .Q(g99) ) ;
DFF     gate743  (.D(g99), .CP(CLK), .Q(g100) ) ;
INV     gate744  (.A(II9597), .Z(g5157) ) ;
DFF     gate745  (.D(g5157), .CP(CLK), .Q(g103) ) ;
INV     gate746  (.A(II12223), .Z(g6784) ) ;
DFF     gate747  (.D(g6784), .CP(CLK), .Q(g104) ) ;
DFF     gate748  (.D(g104), .CP(CLK), .Q(g105) ) ;
INV     gate749  (.A(II9567), .Z(g5147) ) ;
DFF     gate750  (.D(g5147), .CP(CLK), .Q(g108) ) ;
INV     gate751  (.A(II12226), .Z(g6785) ) ;
DFF     gate752  (.D(g6785), .CP(CLK), .Q(g109) ) ;
DFF     gate753  (.D(g109), .CP(CLK), .Q(g110) ) ;
INV     gate754  (.A(II9570), .Z(g5148) ) ;
DFF     gate755  (.D(g5148), .CP(CLK), .Q(g113) ) ;
INV     gate756  (.A(II12229), .Z(g6786) ) ;
DFF     gate757  (.D(g6786), .CP(CLK), .Q(g114) ) ;
INV     gate758  (.A(II9585), .Z(g5153) ) ;
DFF     gate759  (.D(g5153), .CP(CLK), .Q(g117) ) ;
INV     gate760  (.A(II12232), .Z(g6787) ) ;
DFF     gate761  (.D(g6787), .CP(CLK), .Q(g118) ) ;
INV     gate762  (.A(II9588), .Z(g5154) ) ;
DFF     gate763  (.D(g5154), .CP(CLK), .Q(g121) ) ;
INV     gate764  (.A(II12235), .Z(g6788) ) ;
DFF     gate765  (.D(g6788), .CP(CLK), .Q(g122) ) ;
INV     gate766  (.A(II9591), .Z(g5155) ) ;
DFF     gate767  (.D(g5155), .CP(CLK), .Q(g125) ) ;
INV     gate768  (.A(II12238), .Z(g6789) ) ;
DFF     gate769  (.D(g6789), .CP(CLK), .Q(g126) ) ;
INV     gate770  (.A(II9594), .Z(g5156) ) ;
DFF     gate771  (.D(g5156), .CP(CLK), .Q(g129) ) ;
INV     gate772  (.A(II12241), .Z(g6790) ) ;
DFF     gate773  (.D(g6790), .CP(CLK), .Q(g130) ) ;
INV     gate774  (.A(II9573), .Z(g5149) ) ;
DFF     gate775  (.D(g5149), .CP(CLK), .Q(g133) ) ;
INV     gate776  (.A(II12244), .Z(g6791) ) ;
DFF     gate777  (.D(g6791), .CP(CLK), .Q(g134) ) ;
INV     gate778  (.A(II9576), .Z(g5150) ) ;
DFF     gate779  (.D(g5150), .CP(CLK), .Q(g137) ) ;
INV     gate780  (.A(II12247), .Z(g6792) ) ;
DFF     gate781  (.D(g6792), .CP(CLK), .Q(g138) ) ;
INV     gate782  (.A(II9579), .Z(g5151) ) ;
DFF     gate783  (.D(g5151), .CP(CLK), .Q(g141) ) ;
INV     gate784  (.A(II12250), .Z(g6793) ) ;
DFF     gate785  (.D(g6793), .CP(CLK), .Q(g142) ) ;
INV     gate786  (.A(II9582), .Z(g5152) ) ;
DFF     gate787  (.D(g5152), .CP(CLK), .Q(g145) ) ;
INV     gate788  (.A(II7311), .Z(g3836) ) ;
DFF     gate789  (.D(g3836), .CP(CLK), .Q(g287) ) ;
DFF     gate790  (.D(g287), .CP(CLK), .Q(g290) ) ;
INV     gate791  (.A(II15651), .Z(g9087) ) ;
DFF     gate792  (.D(g9087), .CP(CLK), .Q(g255) ) ;
INV     gate793  (.A(II15654), .Z(g9088) ) ;
DFF     gate794  (.D(g9088), .CP(CLK), .Q(g258) ) ;
INV     gate795  (.A(II15657), .Z(g9089) ) ;
DFF     gate796  (.D(g9089), .CP(CLK), .Q(g261) ) ;
INV     gate797  (.A(II15660), .Z(g9090) ) ;
DFF     gate798  (.D(g9090), .CP(CLK), .Q(g264) ) ;
INV     gate799  (.A(II15663), .Z(g9091) ) ;
DFF     gate800  (.D(g9091), .CP(CLK), .Q(g267) ) ;
INV     gate801  (.A(II15666), .Z(g9092) ) ;
DFF     gate802  (.D(g9092), .CP(CLK), .Q(g270) ) ;
INV     gate803  (.A(II15645), .Z(g9085) ) ;
DFF     gate804  (.D(g9085), .CP(CLK), .Q(g281) ) ;
INV     gate805  (.A(II15648), .Z(g9086) ) ;
DFF     gate806  (.D(g9086), .CP(CLK), .Q(g284) ) ;
INV     gate807  (.A(II8715), .Z(g4600) ) ;
DFF     gate808  (.D(g4600), .CP(CLK), .Q(g211) ) ;
INV     gate809  (.A(II11260), .Z(g6311) ) ;
DFF     gate810  (.D(g6311), .CP(CLK), .Q(g216) ) ;
INV     gate811  (.A(II8718), .Z(g4601) ) ;
DFF     gate812  (.D(g4601), .CP(CLK), .Q(g212) ) ;
INV     gate813  (.A(II11263), .Z(g6312) ) ;
DFF     gate814  (.D(g6312), .CP(CLK), .Q(g219) ) ;
INV     gate815  (.A(II8721), .Z(g4602) ) ;
DFF     gate816  (.D(g4602), .CP(CLK), .Q(g213) ) ;
INV     gate817  (.A(II11266), .Z(g6313) ) ;
DFF     gate818  (.D(g6313), .CP(CLK), .Q(g222) ) ;
INV     gate819  (.A(II8724), .Z(g4603) ) ;
DFF     gate820  (.D(g4603), .CP(CLK), .Q(g214) ) ;
INV     gate821  (.A(II11269), .Z(g6314) ) ;
DFF     gate822  (.D(g6314), .CP(CLK), .Q(g225) ) ;
INV     gate823  (.A(II8727), .Z(g4604) ) ;
DFF     gate824  (.D(g4604), .CP(CLK), .Q(g215) ) ;
INV     gate825  (.A(II11272), .Z(g6315) ) ;
DFF     gate826  (.D(g6315), .CP(CLK), .Q(g228) ) ;
INV     gate827  (.A(II8730), .Z(g4605) ) ;
DFF     gate828  (.D(g4605), .CP(CLK), .Q(g231) ) ;
INV     gate829  (.A(II11275), .Z(g6316) ) ;
DFF     gate830  (.D(g6316), .CP(CLK), .Q(g237) ) ;
INV     gate831  (.A(II8733), .Z(g4606) ) ;
DFF     gate832  (.D(g4606), .CP(CLK), .Q(g232) ) ;
INV     gate833  (.A(II11278), .Z(g6317) ) ;
DFF     gate834  (.D(g6317), .CP(CLK), .Q(g240) ) ;
INV     gate835  (.A(II8736), .Z(g4607) ) ;
DFF     gate836  (.D(g4607), .CP(CLK), .Q(g233) ) ;
INV     gate837  (.A(II11281), .Z(g6318) ) ;
DFF     gate838  (.D(g6318), .CP(CLK), .Q(g243) ) ;
INV     gate839  (.A(II8739), .Z(g4608) ) ;
DFF     gate840  (.D(g4608), .CP(CLK), .Q(g234) ) ;
INV     gate841  (.A(II11284), .Z(g6319) ) ;
DFF     gate842  (.D(g6319), .CP(CLK), .Q(g246) ) ;
INV     gate843  (.A(II8742), .Z(g4609) ) ;
DFF     gate844  (.D(g4609), .CP(CLK), .Q(g235) ) ;
INV     gate845  (.A(II11287), .Z(g6320) ) ;
DFF     gate846  (.D(g6320), .CP(CLK), .Q(g249) ) ;
INV     gate847  (.A(II8745), .Z(g4610) ) ;
DFF     gate848  (.D(g4610), .CP(CLK), .Q(g236) ) ;
INV     gate849  (.A(II11290), .Z(g6321) ) ;
DFF     gate850  (.D(g6321), .CP(CLK), .Q(g252) ) ;
INV     gate851  (.A(II8748), .Z(g4611) ) ;
DFF     gate852  (.D(g4611), .CP(CLK), .Q(g273) ) ;
INV     gate853  (.A(II11293), .Z(g6322) ) ;
DFF     gate854  (.D(g6322), .CP(CLK), .Q(g275) ) ;
INV     gate855  (.A(II8751), .Z(g4612) ) ;
DFF     gate856  (.D(g4612), .CP(CLK), .Q(g274) ) ;
INV     gate857  (.A(II11296), .Z(g6323) ) ;
DFF     gate858  (.D(g6323), .CP(CLK), .Q(g278) ) ;
INV     gate859  (.A(II7317), .Z(g3838) ) ;
DFF     gate860  (.D(g3838), .CP(CLK), .Q(g368) ) ;
DFF     gate861  (.D(g368), .CP(CLK), .Q(g371) ) ;
INV     gate862  (.A(II15675), .Z(g9095) ) ;
DFF     gate863  (.D(g9095), .CP(CLK), .Q(g336) ) ;
INV     gate864  (.A(II15678), .Z(g9096) ) ;
DFF     gate865  (.D(g9096), .CP(CLK), .Q(g339) ) ;
INV     gate866  (.A(II15681), .Z(g9097) ) ;
DFF     gate867  (.D(g9097), .CP(CLK), .Q(g342) ) ;
INV     gate868  (.A(II15684), .Z(g9098) ) ;
DFF     gate869  (.D(g9098), .CP(CLK), .Q(g345) ) ;
INV     gate870  (.A(II15687), .Z(g9099) ) ;
DFF     gate871  (.D(g9099), .CP(CLK), .Q(g348) ) ;
INV     gate872  (.A(II15690), .Z(g9100) ) ;
DFF     gate873  (.D(g9100), .CP(CLK), .Q(g351) ) ;
INV     gate874  (.A(II15669), .Z(g9093) ) ;
DFF     gate875  (.D(g9093), .CP(CLK), .Q(g362) ) ;
INV     gate876  (.A(II15672), .Z(g9094) ) ;
DFF     gate877  (.D(g9094), .CP(CLK), .Q(g365) ) ;
INV     gate878  (.A(II8754), .Z(g4613) ) ;
DFF     gate879  (.D(g4613), .CP(CLK), .Q(g292) ) ;
INV     gate880  (.A(II11299), .Z(g6324) ) ;
DFF     gate881  (.D(g6324), .CP(CLK), .Q(g297) ) ;
INV     gate882  (.A(II8757), .Z(g4614) ) ;
DFF     gate883  (.D(g4614), .CP(CLK), .Q(g293) ) ;
INV     gate884  (.A(II11302), .Z(g6325) ) ;
DFF     gate885  (.D(g6325), .CP(CLK), .Q(g300) ) ;
INV     gate886  (.A(II8760), .Z(g4615) ) ;
DFF     gate887  (.D(g4615), .CP(CLK), .Q(g294) ) ;
INV     gate888  (.A(II11305), .Z(g6326) ) ;
DFF     gate889  (.D(g6326), .CP(CLK), .Q(g303) ) ;
INV     gate890  (.A(II8763), .Z(g4616) ) ;
DFF     gate891  (.D(g4616), .CP(CLK), .Q(g295) ) ;
INV     gate892  (.A(II11308), .Z(g6327) ) ;
DFF     gate893  (.D(g6327), .CP(CLK), .Q(g306) ) ;
INV     gate894  (.A(II8766), .Z(g4617) ) ;
DFF     gate895  (.D(g4617), .CP(CLK), .Q(g296) ) ;
INV     gate896  (.A(II11311), .Z(g6328) ) ;
DFF     gate897  (.D(g6328), .CP(CLK), .Q(g309) ) ;
INV     gate898  (.A(II8769), .Z(g4618) ) ;
DFF     gate899  (.D(g4618), .CP(CLK), .Q(g312) ) ;
INV     gate900  (.A(II11314), .Z(g6329) ) ;
DFF     gate901  (.D(g6329), .CP(CLK), .Q(g318) ) ;
INV     gate902  (.A(II8772), .Z(g4619) ) ;
DFF     gate903  (.D(g4619), .CP(CLK), .Q(g313) ) ;
INV     gate904  (.A(II11317), .Z(g6330) ) ;
DFF     gate905  (.D(g6330), .CP(CLK), .Q(g321) ) ;
INV     gate906  (.A(II8775), .Z(g4620) ) ;
DFF     gate907  (.D(g4620), .CP(CLK), .Q(g314) ) ;
INV     gate908  (.A(II11320), .Z(g6331) ) ;
DFF     gate909  (.D(g6331), .CP(CLK), .Q(g324) ) ;
INV     gate910  (.A(II8778), .Z(g4621) ) ;
DFF     gate911  (.D(g4621), .CP(CLK), .Q(g315) ) ;
INV     gate912  (.A(II11323), .Z(g6332) ) ;
DFF     gate913  (.D(g6332), .CP(CLK), .Q(g327) ) ;
INV     gate914  (.A(II8781), .Z(g4622) ) ;
DFF     gate915  (.D(g4622), .CP(CLK), .Q(g316) ) ;
INV     gate916  (.A(II11326), .Z(g6333) ) ;
DFF     gate917  (.D(g6333), .CP(CLK), .Q(g330) ) ;
INV     gate918  (.A(II8784), .Z(g4623) ) ;
DFF     gate919  (.D(g4623), .CP(CLK), .Q(g317) ) ;
INV     gate920  (.A(II11329), .Z(g6334) ) ;
DFF     gate921  (.D(g6334), .CP(CLK), .Q(g333) ) ;
INV     gate922  (.A(II8787), .Z(g4624) ) ;
DFF     gate923  (.D(g4624), .CP(CLK), .Q(g354) ) ;
INV     gate924  (.A(II11332), .Z(g6335) ) ;
DFF     gate925  (.D(g6335), .CP(CLK), .Q(g356) ) ;
INV     gate926  (.A(II8790), .Z(g4625) ) ;
DFF     gate927  (.D(g4625), .CP(CLK), .Q(g355) ) ;
INV     gate928  (.A(II11335), .Z(g6336) ) ;
DFF     gate929  (.D(g6336), .CP(CLK), .Q(g359) ) ;
INV     gate930  (.A(II7323), .Z(g3840) ) ;
DFF     gate931  (.D(g3840), .CP(CLK), .Q(g449) ) ;
DFF     gate932  (.D(g449), .CP(CLK), .Q(g452) ) ;
INV     gate933  (.A(II15699), .Z(g9103) ) ;
DFF     gate934  (.D(g9103), .CP(CLK), .Q(g417) ) ;
INV     gate935  (.A(II15702), .Z(g9104) ) ;
DFF     gate936  (.D(g9104), .CP(CLK), .Q(g420) ) ;
INV     gate937  (.A(II15705), .Z(g9105) ) ;
DFF     gate938  (.D(g9105), .CP(CLK), .Q(g423) ) ;
INV     gate939  (.A(II15708), .Z(g9106) ) ;
DFF     gate940  (.D(g9106), .CP(CLK), .Q(g426) ) ;
INV     gate941  (.A(II15711), .Z(g9107) ) ;
DFF     gate942  (.D(g9107), .CP(CLK), .Q(g429) ) ;
INV     gate943  (.A(II15714), .Z(g9108) ) ;
DFF     gate944  (.D(g9108), .CP(CLK), .Q(g432) ) ;
INV     gate945  (.A(II15693), .Z(g9101) ) ;
DFF     gate946  (.D(g9101), .CP(CLK), .Q(g443) ) ;
INV     gate947  (.A(II15696), .Z(g9102) ) ;
DFF     gate948  (.D(g9102), .CP(CLK), .Q(g446) ) ;
INV     gate949  (.A(II8793), .Z(g4626) ) ;
DFF     gate950  (.D(g4626), .CP(CLK), .Q(g373) ) ;
INV     gate951  (.A(II11338), .Z(g6337) ) ;
DFF     gate952  (.D(g6337), .CP(CLK), .Q(g378) ) ;
INV     gate953  (.A(II8796), .Z(g4627) ) ;
DFF     gate954  (.D(g4627), .CP(CLK), .Q(g374) ) ;
INV     gate955  (.A(II11341), .Z(g6338) ) ;
DFF     gate956  (.D(g6338), .CP(CLK), .Q(g381) ) ;
INV     gate957  (.A(II8799), .Z(g4628) ) ;
DFF     gate958  (.D(g4628), .CP(CLK), .Q(g375) ) ;
INV     gate959  (.A(II11344), .Z(g6339) ) ;
DFF     gate960  (.D(g6339), .CP(CLK), .Q(g384) ) ;
INV     gate961  (.A(II8802), .Z(g4629) ) ;
DFF     gate962  (.D(g4629), .CP(CLK), .Q(g376) ) ;
INV     gate963  (.A(II11347), .Z(g6340) ) ;
DFF     gate964  (.D(g6340), .CP(CLK), .Q(g387) ) ;
INV     gate965  (.A(II8805), .Z(g4630) ) ;
DFF     gate966  (.D(g4630), .CP(CLK), .Q(g377) ) ;
INV     gate967  (.A(II11350), .Z(g6341) ) ;
DFF     gate968  (.D(g6341), .CP(CLK), .Q(g390) ) ;
INV     gate969  (.A(II8808), .Z(g4631) ) ;
DFF     gate970  (.D(g4631), .CP(CLK), .Q(g393) ) ;
INV     gate971  (.A(II11353), .Z(g6342) ) ;
DFF     gate972  (.D(g6342), .CP(CLK), .Q(g399) ) ;
INV     gate973  (.A(II8811), .Z(g4632) ) ;
DFF     gate974  (.D(g4632), .CP(CLK), .Q(g394) ) ;
INV     gate975  (.A(II11356), .Z(g6343) ) ;
DFF     gate976  (.D(g6343), .CP(CLK), .Q(g402) ) ;
INV     gate977  (.A(II8814), .Z(g4633) ) ;
DFF     gate978  (.D(g4633), .CP(CLK), .Q(g395) ) ;
INV     gate979  (.A(II11359), .Z(g6344) ) ;
DFF     gate980  (.D(g6344), .CP(CLK), .Q(g405) ) ;
INV     gate981  (.A(II8817), .Z(g4634) ) ;
DFF     gate982  (.D(g4634), .CP(CLK), .Q(g396) ) ;
INV     gate983  (.A(II11362), .Z(g6345) ) ;
DFF     gate984  (.D(g6345), .CP(CLK), .Q(g408) ) ;
INV     gate985  (.A(II8820), .Z(g4635) ) ;
DFF     gate986  (.D(g4635), .CP(CLK), .Q(g397) ) ;
INV     gate987  (.A(II11365), .Z(g6346) ) ;
DFF     gate988  (.D(g6346), .CP(CLK), .Q(g411) ) ;
INV     gate989  (.A(II8823), .Z(g4636) ) ;
DFF     gate990  (.D(g4636), .CP(CLK), .Q(g398) ) ;
INV     gate991  (.A(II11368), .Z(g6347) ) ;
DFF     gate992  (.D(g6347), .CP(CLK), .Q(g414) ) ;
INV     gate993  (.A(II8826), .Z(g4637) ) ;
DFF     gate994  (.D(g4637), .CP(CLK), .Q(g435) ) ;
INV     gate995  (.A(II11371), .Z(g6348) ) ;
DFF     gate996  (.D(g6348), .CP(CLK), .Q(g437) ) ;
INV     gate997  (.A(II8829), .Z(g4638) ) ;
DFF     gate998  (.D(g4638), .CP(CLK), .Q(g436) ) ;
INV     gate999  (.A(II11374), .Z(g6349) ) ;
DFF     gate1000  (.D(g6349), .CP(CLK), .Q(g440) ) ;
INV     gate1001  (.A(II7329), .Z(g3842) ) ;
DFF     gate1002  (.D(g3842), .CP(CLK), .Q(g530) ) ;
DFF     gate1003  (.D(g530), .CP(CLK), .Q(g533) ) ;
INV     gate1004  (.A(II15723), .Z(g9111) ) ;
DFF     gate1005  (.D(g9111), .CP(CLK), .Q(g498) ) ;
INV     gate1006  (.A(II15726), .Z(g9112) ) ;
DFF     gate1007  (.D(g9112), .CP(CLK), .Q(g501) ) ;
INV     gate1008  (.A(II15729), .Z(g9113) ) ;
DFF     gate1009  (.D(g9113), .CP(CLK), .Q(g504) ) ;
INV     gate1010  (.A(II15732), .Z(g9114) ) ;
DFF     gate1011  (.D(g9114), .CP(CLK), .Q(g507) ) ;
INV     gate1012  (.A(II15735), .Z(g9115) ) ;
DFF     gate1013  (.D(g9115), .CP(CLK), .Q(g510) ) ;
INV     gate1014  (.A(II15738), .Z(g9116) ) ;
DFF     gate1015  (.D(g9116), .CP(CLK), .Q(g513) ) ;
INV     gate1016  (.A(II15717), .Z(g9109) ) ;
DFF     gate1017  (.D(g9109), .CP(CLK), .Q(g524) ) ;
INV     gate1018  (.A(II15720), .Z(g9110) ) ;
DFF     gate1019  (.D(g9110), .CP(CLK), .Q(g527) ) ;
INV     gate1020  (.A(II8832), .Z(g4639) ) ;
DFF     gate1021  (.D(g4639), .CP(CLK), .Q(g454) ) ;
INV     gate1022  (.A(II11377), .Z(g6350) ) ;
DFF     gate1023  (.D(g6350), .CP(CLK), .Q(g459) ) ;
INV     gate1024  (.A(II8835), .Z(g4640) ) ;
DFF     gate1025  (.D(g4640), .CP(CLK), .Q(g455) ) ;
INV     gate1026  (.A(II11380), .Z(g6351) ) ;
DFF     gate1027  (.D(g6351), .CP(CLK), .Q(g462) ) ;
INV     gate1028  (.A(II8838), .Z(g4641) ) ;
DFF     gate1029  (.D(g4641), .CP(CLK), .Q(g456) ) ;
INV     gate1030  (.A(II11383), .Z(g6352) ) ;
DFF     gate1031  (.D(g6352), .CP(CLK), .Q(g465) ) ;
INV     gate1032  (.A(II8841), .Z(g4642) ) ;
DFF     gate1033  (.D(g4642), .CP(CLK), .Q(g457) ) ;
INV     gate1034  (.A(II11386), .Z(g6353) ) ;
DFF     gate1035  (.D(g6353), .CP(CLK), .Q(g468) ) ;
INV     gate1036  (.A(II8844), .Z(g4643) ) ;
DFF     gate1037  (.D(g4643), .CP(CLK), .Q(g458) ) ;
INV     gate1038  (.A(II11389), .Z(g6354) ) ;
DFF     gate1039  (.D(g6354), .CP(CLK), .Q(g471) ) ;
INV     gate1040  (.A(II8847), .Z(g4644) ) ;
DFF     gate1041  (.D(g4644), .CP(CLK), .Q(g474) ) ;
INV     gate1042  (.A(II11392), .Z(g6355) ) ;
DFF     gate1043  (.D(g6355), .CP(CLK), .Q(g480) ) ;
INV     gate1044  (.A(II8850), .Z(g4645) ) ;
DFF     gate1045  (.D(g4645), .CP(CLK), .Q(g475) ) ;
INV     gate1046  (.A(II11395), .Z(g6356) ) ;
DFF     gate1047  (.D(g6356), .CP(CLK), .Q(g483) ) ;
INV     gate1048  (.A(II8853), .Z(g4646) ) ;
DFF     gate1049  (.D(g4646), .CP(CLK), .Q(g476) ) ;
INV     gate1050  (.A(II11398), .Z(g6357) ) ;
DFF     gate1051  (.D(g6357), .CP(CLK), .Q(g486) ) ;
INV     gate1052  (.A(II8856), .Z(g4647) ) ;
DFF     gate1053  (.D(g4647), .CP(CLK), .Q(g477) ) ;
INV     gate1054  (.A(II11401), .Z(g6358) ) ;
DFF     gate1055  (.D(g6358), .CP(CLK), .Q(g489) ) ;
INV     gate1056  (.A(II8859), .Z(g4648) ) ;
DFF     gate1057  (.D(g4648), .CP(CLK), .Q(g478) ) ;
INV     gate1058  (.A(II11404), .Z(g6359) ) ;
DFF     gate1059  (.D(g6359), .CP(CLK), .Q(g492) ) ;
INV     gate1060  (.A(II8862), .Z(g4649) ) ;
DFF     gate1061  (.D(g4649), .CP(CLK), .Q(g479) ) ;
INV     gate1062  (.A(II11407), .Z(g6360) ) ;
DFF     gate1063  (.D(g6360), .CP(CLK), .Q(g495) ) ;
INV     gate1064  (.A(II8865), .Z(g4650) ) ;
DFF     gate1065  (.D(g4650), .CP(CLK), .Q(g516) ) ;
INV     gate1066  (.A(II11410), .Z(g6361) ) ;
DFF     gate1067  (.D(g6361), .CP(CLK), .Q(g518) ) ;
INV     gate1068  (.A(II8868), .Z(g4651) ) ;
DFF     gate1069  (.D(g4651), .CP(CLK), .Q(g517) ) ;
INV     gate1070  (.A(II11413), .Z(g6362) ) ;
DFF     gate1071  (.D(g6362), .CP(CLK), .Q(g521) ) ;
INV     gate1072  (.A(II7335), .Z(g3844) ) ;
DFF     gate1073  (.D(g3844), .CP(CLK), .Q(g535) ) ;
INV     gate1074  (.A(II11416), .Z(g6363) ) ;
DFF     gate1075  (.D(g6363), .CP(CLK), .Q(g536) ) ;
INV     gate1076  (.A(II7338), .Z(g3845) ) ;
DFF     gate1077  (.D(g3845), .CP(CLK), .Q(g539) ) ;
INV     gate1078  (.A(II11419), .Z(g6364) ) ;
DFF     gate1079  (.D(g6364), .CP(CLK), .Q(g540) ) ;
INV     gate1080  (.A(II7341), .Z(g3846) ) ;
DFF     gate1081  (.D(g3846), .CP(CLK), .Q(g543) ) ;
INV     gate1082  (.A(II11422), .Z(g6365) ) ;
DFF     gate1083  (.D(g6365), .CP(CLK), .Q(g544) ) ;
INV     gate1084  (.A(II15492), .Z(g9026) ) ;
DFF     gate1085  (.D(g9026), .CP(CLK), .Q(g547) ) ;
INV     gate1086  (.A(II15495), .Z(g9027) ) ;
DFF     gate1087  (.D(g9027), .CP(CLK), .Q(g550) ) ;
INV     gate1088  (.A(II15498), .Z(g9028) ) ;
DFF     gate1089  (.D(g9028), .CP(CLK), .Q(g553) ) ;
INV     gate1090  (.A(II7344), .Z(g3847) ) ;
DFF     gate1091  (.D(g3847), .CP(CLK), .Q(g556) ) ;
INV     gate1092  (.A(II11425), .Z(g6366) ) ;
DFF     gate1093  (.D(g6366), .CP(CLK), .Q(g557) ) ;
INV     gate1094  (.A(II7347), .Z(g3848) ) ;
DFF     gate1095  (.D(g3848), .CP(CLK), .Q(g566) ) ;
INV     gate1096  (.A(II11428), .Z(g6367) ) ;
DFF     gate1097  (.D(g6367), .CP(CLK), .Q(g567) ) ;
INV     gate1098  (.A(II7353), .Z(g3850) ) ;
DFF     gate1099  (.D(g3850), .CP(CLK), .Q(g579) ) ;
INV     gate1100  (.A(II11431), .Z(g6368) ) ;
DFF     gate1101  (.D(g6368), .CP(CLK), .Q(g580) ) ;
INV     gate1102  (.A(II7356), .Z(g3851) ) ;
DFF     gate1103  (.D(g3851), .CP(CLK), .Q(g583) ) ;
INV     gate1104  (.A(II11434), .Z(g6369) ) ;
DFF     gate1105  (.D(g6369), .CP(CLK), .Q(g584) ) ;
INV     gate1106  (.A(II7359), .Z(g3852) ) ;
DFF     gate1107  (.D(g3852), .CP(CLK), .Q(g587) ) ;
INV     gate1108  (.A(II11437), .Z(g6370) ) ;
DFF     gate1109  (.D(g6370), .CP(CLK), .Q(g560) ) ;
INV     gate1110  (.A(II15501), .Z(g9029) ) ;
DFF     gate1111  (.D(g9029), .CP(CLK), .Q(g563) ) ;
INV     gate1112  (.A(II15504), .Z(g9030) ) ;
DFF     gate1113  (.D(g9030), .CP(CLK), .Q(g570) ) ;
INV     gate1114  (.A(II15507), .Z(g9031) ) ;
DFF     gate1115  (.D(g9031), .CP(CLK), .Q(g588) ) ;
INV     gate1116  (.A(II15510), .Z(g9032) ) ;
DFF     gate1117  (.D(g9032), .CP(CLK), .Q(g591) ) ;
INV     gate1118  (.A(II15513), .Z(g9033) ) ;
DFF     gate1119  (.D(g9033), .CP(CLK), .Q(g573) ) ;
INV     gate1120  (.A(II7350), .Z(g3849) ) ;
DFF     gate1121  (.D(g3849), .CP(CLK), .Q(g576) ) ;
DFF     gate1122  (.D(g576), .CP(CLK), .Q(g595) ) ;
INV     gate1123  (.A(II12256), .Z(g6795) ) ;
DFF     gate1124  (.D(g6795), .CP(CLK), .Q(g596) ) ;
INV     gate1125  (.A(II12259), .Z(g6796) ) ;
DFF     gate1126  (.D(g6796), .CP(CLK), .Q(g597) ) ;
INV     gate1127  (.A(II12262), .Z(g6797) ) ;
DFF     gate1128  (.D(g6797), .CP(CLK), .Q(g598) ) ;
INV     gate1129  (.A(II12265), .Z(g6798) ) ;
DFF     gate1130  (.D(g6798), .CP(CLK), .Q(g599) ) ;
INV     gate1131  (.A(II12292), .Z(g6807) ) ;
DFF     gate1132  (.D(g6807), .CP(CLK), .Q(g600) ) ;
INV     gate1133  (.A(II12268), .Z(g6799) ) ;
DFF     gate1134  (.D(g6799), .CP(CLK), .Q(g601) ) ;
INV     gate1135  (.A(II12271), .Z(g6800) ) ;
DFF     gate1136  (.D(g6800), .CP(CLK), .Q(g602) ) ;
INV     gate1137  (.A(II12274), .Z(g6801) ) ;
DFF     gate1138  (.D(g6801), .CP(CLK), .Q(g603) ) ;
INV     gate1139  (.A(II12277), .Z(g6802) ) ;
DFF     gate1140  (.D(g6802), .CP(CLK), .Q(g604) ) ;
INV     gate1141  (.A(II12280), .Z(g6803) ) ;
DFF     gate1142  (.D(g6803), .CP(CLK), .Q(g605) ) ;
INV     gate1143  (.A(II12283), .Z(g6804) ) ;
DFF     gate1144  (.D(g6804), .CP(CLK), .Q(g606) ) ;
INV     gate1145  (.A(II12286), .Z(g6805) ) ;
DFF     gate1146  (.D(g6805), .CP(CLK), .Q(g607) ) ;
INV     gate1147  (.A(II12289), .Z(g6806) ) ;
DFF     gate1148  (.D(g6806), .CP(CLK), .Q(g608) ) ;
INV     gate1149  (.A(II12295), .Z(g6808) ) ;
DFF     gate1150  (.D(g6808), .CP(CLK), .Q(g609) ) ;
INV     gate1151  (.A(II12298), .Z(g6809) ) ;
DFF     gate1152  (.D(g6809), .CP(CLK), .Q(g610) ) ;
INV     gate1153  (.A(II12301), .Z(g6810) ) ;
DFF     gate1154  (.D(g6810), .CP(CLK), .Q(g611) ) ;
INV     gate1155  (.A(II12304), .Z(g6811) ) ;
DFF     gate1156  (.D(g6811), .CP(CLK), .Q(g612) ) ;
INV     gate1157  (.A(II12331), .Z(g6820) ) ;
DFF     gate1158  (.D(g6820), .CP(CLK), .Q(g613) ) ;
INV     gate1159  (.A(II12307), .Z(g6812) ) ;
DFF     gate1160  (.D(g6812), .CP(CLK), .Q(g614) ) ;
INV     gate1161  (.A(II12310), .Z(g6813) ) ;
DFF     gate1162  (.D(g6813), .CP(CLK), .Q(g615) ) ;
INV     gate1163  (.A(II12313), .Z(g6814) ) ;
DFF     gate1164  (.D(g6814), .CP(CLK), .Q(g616) ) ;
INV     gate1165  (.A(II12316), .Z(g6815) ) ;
DFF     gate1166  (.D(g6815), .CP(CLK), .Q(g617) ) ;
INV     gate1167  (.A(II12319), .Z(g6816) ) ;
DFF     gate1168  (.D(g6816), .CP(CLK), .Q(g618) ) ;
INV     gate1169  (.A(II12322), .Z(g6817) ) ;
DFF     gate1170  (.D(g6817), .CP(CLK), .Q(g619) ) ;
INV     gate1171  (.A(II12325), .Z(g6818) ) ;
DFF     gate1172  (.D(g6818), .CP(CLK), .Q(g620) ) ;
INV     gate1173  (.A(II12328), .Z(g6819) ) ;
DFF     gate1174  (.D(g6819), .CP(CLK), .Q(g621) ) ;
INV     gate1175  (.A(II12334), .Z(g6821) ) ;
DFF     gate1176  (.D(g6821), .CP(CLK), .Q(g622) ) ;
INV     gate1177  (.A(II12337), .Z(g6822) ) ;
DFF     gate1178  (.D(g6822), .CP(CLK), .Q(g623) ) ;
INV     gate1179  (.A(II12364), .Z(g6831) ) ;
DFF     gate1180  (.D(g6831), .CP(CLK), .Q(g624) ) ;
INV     gate1181  (.A(II12340), .Z(g6823) ) ;
DFF     gate1182  (.D(g6823), .CP(CLK), .Q(g625) ) ;
INV     gate1183  (.A(II12343), .Z(g6824) ) ;
DFF     gate1184  (.D(g6824), .CP(CLK), .Q(g626) ) ;
INV     gate1185  (.A(II12346), .Z(g6825) ) ;
DFF     gate1186  (.D(g6825), .CP(CLK), .Q(g627) ) ;
INV     gate1187  (.A(II12349), .Z(g6826) ) ;
DFF     gate1188  (.D(g6826), .CP(CLK), .Q(g628) ) ;
INV     gate1189  (.A(II12352), .Z(g6827) ) ;
DFF     gate1190  (.D(g6827), .CP(CLK), .Q(g629) ) ;
INV     gate1191  (.A(II12355), .Z(g6828) ) ;
DFF     gate1192  (.D(g6828), .CP(CLK), .Q(g630) ) ;
INV     gate1193  (.A(II12358), .Z(g6829) ) ;
DFF     gate1194  (.D(g6829), .CP(CLK), .Q(g631) ) ;
INV     gate1195  (.A(II12361), .Z(g6830) ) ;
DFF     gate1196  (.D(g6830), .CP(CLK), .Q(g632) ) ;
INV     gate1197  (.A(II8871), .Z(g4652) ) ;
DFF     gate1198  (.D(g4652), .CP(CLK), .Q(g646) ) ;
DFF     gate1199  (.D(g646), .CP(CLK), .Q(g652) ) ;
INV     gate1200  (.A(II14100), .Z(g7743) ) ;
DFF     gate1201  (.D(g7743), .CP(CLK), .Q(g661) ) ;
INV     gate1202  (.A(II14103), .Z(g7744) ) ;
DFF     gate1203  (.D(g7744), .CP(CLK), .Q(g665) ) ;
INV     gate1204  (.A(II14106), .Z(g7745) ) ;
DFF     gate1205  (.D(g7745), .CP(CLK), .Q(g669) ) ;
INV     gate1206  (.A(II14109), .Z(g7746) ) ;
DFF     gate1207  (.D(g7746), .CP(CLK), .Q(g673) ) ;
INV     gate1208  (.A(II14112), .Z(g7747) ) ;
DFF     gate1209  (.D(g7747), .CP(CLK), .Q(g677) ) ;
INV     gate1210  (.A(II14115), .Z(g7748) ) ;
DFF     gate1211  (.D(g7748), .CP(CLK), .Q(g681) ) ;
INV     gate1212  (.A(II14118), .Z(g7749) ) ;
DFF     gate1213  (.D(g7749), .CP(CLK), .Q(g685) ) ;
INV     gate1214  (.A(II14121), .Z(g7750) ) ;
DFF     gate1215  (.D(g7750), .CP(CLK), .Q(g706) ) ;
INV     gate1216  (.A(II14124), .Z(g7751) ) ;
DFF     gate1217  (.D(g7751), .CP(CLK), .Q(g710) ) ;
INV     gate1218  (.A(II14127), .Z(g7752) ) ;
DFF     gate1219  (.D(g7752), .CP(CLK), .Q(g714) ) ;
INV     gate1220  (.A(II14130), .Z(g7753) ) ;
DFF     gate1221  (.D(g7753), .CP(CLK), .Q(g718) ) ;
INV     gate1222  (.A(II14136), .Z(g7755) ) ;
DFF     gate1223  (.D(g7755), .CP(CLK), .Q(g734) ) ;
INV     gate1224  (.A(II14133), .Z(g7754) ) ;
DFF     gate1225  (.D(g7754), .CP(CLK), .Q(g730) ) ;
INV     gate1226  (.A(II11440), .Z(g6371) ) ;
DFF     gate1227  (.D(g6371), .CP(CLK), .Q(g689) ) ;
INV     gate1228  (.A(II12391), .Z(g6840) ) ;
DFF     gate1229  (.D(g6840), .CP(CLK), .Q(g758) ) ;
INV     gate1230  (.A(II12367), .Z(g6832) ) ;
DFF     gate1231  (.D(g6832), .CP(CLK), .Q(g759) ) ;
INV     gate1232  (.A(II12370), .Z(g6833) ) ;
DFF     gate1233  (.D(g6833), .CP(CLK), .Q(g760) ) ;
INV     gate1234  (.A(II12373), .Z(g6834) ) ;
DFF     gate1235  (.D(g6834), .CP(CLK), .Q(g761) ) ;
INV     gate1236  (.A(II12376), .Z(g6835) ) ;
DFF     gate1237  (.D(g6835), .CP(CLK), .Q(g762) ) ;
INV     gate1238  (.A(II12379), .Z(g6836) ) ;
DFF     gate1239  (.D(g6836), .CP(CLK), .Q(g763) ) ;
INV     gate1240  (.A(II12382), .Z(g6837) ) ;
DFF     gate1241  (.D(g6837), .CP(CLK), .Q(g764) ) ;
INV     gate1242  (.A(II12385), .Z(g6838) ) ;
DFF     gate1243  (.D(g6838), .CP(CLK), .Q(g765) ) ;
INV     gate1244  (.A(II12388), .Z(g6839) ) ;
DFF     gate1245  (.D(g6839), .CP(CLK), .Q(g766) ) ;
INV     gate1246  (.A(II12394), .Z(g6841) ) ;
DFF     gate1247  (.D(g6841), .CP(CLK), .Q(g767) ) ;
INV     gate1248  (.A(II12397), .Z(g6842) ) ;
DFF     gate1249  (.D(g6842), .CP(CLK), .Q(g768) ) ;
INV     gate1250  (.A(II12400), .Z(g6843) ) ;
DFF     gate1251  (.D(g6843), .CP(CLK), .Q(g769) ) ;
INV     gate1252  (.A(II12403), .Z(g6844) ) ;
DFF     gate1253  (.D(g6844), .CP(CLK), .Q(g770) ) ;
INV     gate1254  (.A(II12406), .Z(g6845) ) ;
DFF     gate1255  (.D(g6845), .CP(CLK), .Q(g771) ) ;
INV     gate1256  (.A(II12409), .Z(g6846) ) ;
DFF     gate1257  (.D(g6846), .CP(CLK), .Q(g772) ) ;
INV     gate1258  (.A(II12412), .Z(g6847) ) ;
DFF     gate1259  (.D(g6847), .CP(CLK), .Q(g773) ) ;
INV     gate1260  (.A(II12415), .Z(g6848) ) ;
DFF     gate1261  (.D(g6848), .CP(CLK), .Q(g774) ) ;
INV     gate1262  (.A(II7365), .Z(g3854) ) ;
DFF     gate1263  (.D(g3854), .CP(CLK), .Q(g795) ) ;
INV     gate1264  (.A(II9612), .Z(g5162) ) ;
DFF     gate1265  (.D(g5162), .CP(CLK), .Q(g792) ) ;
INV     gate1266  (.A(II10259), .Z(g5734) ) ;
DFF     gate1267  (.D(g5734), .CP(CLK), .Q(g782) ) ;
INV     gate1268  (.A(II14139), .Z(g7756) ) ;
DFF     gate1269  (.D(g7756), .CP(CLK), .Q(g799) ) ;
INV     gate1270  (.A(II14142), .Z(g7757) ) ;
DFF     gate1271  (.D(g7757), .CP(CLK), .Q(g803) ) ;
INV     gate1272  (.A(II13710), .Z(g7510) ) ;
DFF     gate1273  (.D(g7510), .CP(CLK), .Q(g806) ) ;
INV     gate1274  (.A(II13713), .Z(g7511) ) ;
DFF     gate1275  (.D(g7511), .CP(CLK), .Q(g809) ) ;
INV     gate1276  (.A(II14145), .Z(g7758) ) ;
DFF     gate1277  (.D(g7758), .CP(CLK), .Q(g812) ) ;
INV     gate1278  (.A(II14148), .Z(g7759) ) ;
DFF     gate1279  (.D(g7759), .CP(CLK), .Q(g775) ) ;
INV     gate1280  (.A(II13320), .Z(g7296) ) ;
DFF     gate1281  (.D(g7296), .CP(CLK), .Q(g778) ) ;
INV     gate1282  (.A(II14151), .Z(g7760) ) ;
DFF     gate1283  (.D(g7760), .CP(CLK), .Q(g815) ) ;
INV     gate1284  (.A(II14154), .Z(g7761) ) ;
DFF     gate1285  (.D(g7761), .CP(CLK), .Q(g819) ) ;
INV     gate1286  (.A(II13716), .Z(g7512) ) ;
DFF     gate1287  (.D(g7512), .CP(CLK), .Q(g822) ) ;
INV     gate1288  (.A(II13719), .Z(g7513) ) ;
DFF     gate1289  (.D(g7513), .CP(CLK), .Q(g825) ) ;
INV     gate1290  (.A(II14157), .Z(g7762) ) ;
DFF     gate1291  (.D(g7762), .CP(CLK), .Q(g828) ) ;
INV     gate1292  (.A(II14160), .Z(g7763) ) ;
DFF     gate1293  (.D(g7763), .CP(CLK), .Q(g786) ) ;
INV     gate1294  (.A(II13323), .Z(g7297) ) ;
DFF     gate1295  (.D(g7297), .CP(CLK), .Q(g789) ) ;
INV     gate1296  (.A(II7374), .Z(g3857) ) ;
DFF     gate1297  (.D(g3857), .CP(CLK), .Q(g955) ) ;
INV     gate1298  (.A(II9633), .Z(g5169) ) ;
DFF     gate1299  (.D(g5169), .CP(CLK), .Q(g959) ) ;
INV     gate1300  (.A(II9636), .Z(g5170) ) ;
DFF     gate1301  (.D(g5170), .CP(CLK), .Q(g945) ) ;
INV     gate1302  (.A(II14786), .Z(g8664) ) ;
DFF     gate1303  (.D(g8664), .CP(CLK), .Q(g948) ) ;
INV     gate1304  (.A(II14789), .Z(g8665) ) ;
DFF     gate1305  (.D(g8665), .CP(CLK), .Q(g949) ) ;
INV     gate1306  (.A(II14792), .Z(g8666) ) ;
DFF     gate1307  (.D(g8666), .CP(CLK), .Q(g950) ) ;
INV     gate1308  (.A(II14795), .Z(g8667) ) ;
DFF     gate1309  (.D(g8667), .CP(CLK), .Q(g951) ) ;
INV     gate1310  (.A(II14798), .Z(g8668) ) ;
DFF     gate1311  (.D(g8668), .CP(CLK), .Q(g952) ) ;
INV     gate1312  (.A(II14801), .Z(g8669) ) ;
DFF     gate1313  (.D(g8669), .CP(CLK), .Q(g953) ) ;
INV     gate1314  (.A(II14804), .Z(g8670) ) ;
DFF     gate1315  (.D(g8670), .CP(CLK), .Q(g954) ) ;
INV     gate1316  (.A(II14807), .Z(g8671) ) ;
DFF     gate1317  (.D(g8671), .CP(CLK), .Q(g943) ) ;
INV     gate1318  (.A(II9630), .Z(g5168) ) ;
DFF     gate1319  (.D(g5168), .CP(CLK), .Q(g936) ) ;
INV     gate1320  (.A(II10262), .Z(g5735) ) ;
DFF     gate1321  (.D(g5735), .CP(CLK), .Q(g940) ) ;
INV     gate1322  (.A(II6440), .Z(g2652) ) ;
DFF     gate1323  (.D(g2652), .CP(CLK), .Q(g942) ) ;
INV     gate1324  (.A(II11443), .Z(g6372) ) ;
DFF     gate1325  (.D(g6372), .CP(CLK), .Q(g944) ) ;
INV     gate1326  (.A(II14439), .Z(g8220) ) ;
DFF     gate1327  (.D(g8220), .CP(CLK), .Q(g855) ) ;
INV     gate1328  (.A(II14442), .Z(g8221) ) ;
DFF     gate1329  (.D(g8221), .CP(CLK), .Q(g859) ) ;
INV     gate1330  (.A(II14445), .Z(g8222) ) ;
DFF     gate1331  (.D(g8222), .CP(CLK), .Q(g863) ) ;
INV     gate1332  (.A(II6437), .Z(g2651) ) ;
DFF     gate1333  (.D(g2651), .CP(CLK), .Q(g831) ) ;
INV     gate1334  (.A(II6434), .Z(g2650) ) ;
DFF     gate1335  (.D(g2650), .CP(CLK), .Q(g834) ) ;
INV     gate1336  (.A(II6431), .Z(g2649) ) ;
DFF     gate1337  (.D(g2649), .CP(CLK), .Q(g837) ) ;
INV     gate1338  (.A(II6428), .Z(g2648) ) ;
DFF     gate1339  (.D(g2648), .CP(CLK), .Q(g840) ) ;
INV     gate1340  (.A(II6425), .Z(g2647) ) ;
DFF     gate1341  (.D(g2647), .CP(CLK), .Q(g843) ) ;
INV     gate1342  (.A(II6422), .Z(g2646) ) ;
DFF     gate1343  (.D(g2646), .CP(CLK), .Q(g846) ) ;
INV     gate1344  (.A(II6419), .Z(g2645) ) ;
DFF     gate1345  (.D(g2645), .CP(CLK), .Q(g849) ) ;
INV     gate1346  (.A(II6416), .Z(g2644) ) ;
DFF     gate1347  (.D(g2644), .CP(CLK), .Q(g852) ) ;
INV     gate1348  (.A(II12894), .Z(g7102) ) ;
DFF     gate1349  (.D(g7102), .CP(CLK), .Q(g890) ) ;
DFF     gate1350  (.D(g890), .CP(CLK), .Q(g878) ) ;
DFF     gate1351  (.D(g878), .CP(CLK), .Q(g926) ) ;
INV     gate1352  (.A(II9621), .Z(g5165) ) ;
DFF     gate1353  (.D(g5165), .CP(CLK), .Q(g875) ) ;
INV     gate1354  (.A(II9615), .Z(g5163) ) ;
DFF     gate1355  (.D(g5163), .CP(CLK), .Q(g866) ) ;
INV     gate1356  (.A(II7371), .Z(g3856) ) ;
DFF     gate1357  (.D(g3856), .CP(CLK), .Q(g929) ) ;
INV     gate1358  (.A(II9624), .Z(g5166) ) ;
DFF     gate1359  (.D(g5166), .CP(CLK), .Q(g933) ) ;
INV     gate1360  (.A(II9627), .Z(g5167) ) ;
DFF     gate1361  (.D(g5167), .CP(CLK), .Q(g871) ) ;
INV     gate1362  (.A(II8877), .Z(g4654) ) ;
DFF     gate1363  (.D(g4654), .CP(CLK), .Q(g874) ) ;
INV     gate1364  (.A(II7368), .Z(g3855) ) ;
DFF     gate1365  (.D(g3855), .CP(CLK), .Q(g891) ) ;
DFF     gate1366  (.D(g891), .CP(CLK), .Q(g896) ) ;
DFF     gate1367  (.D(g896), .CP(CLK), .Q(g901) ) ;
DFF     gate1368  (.D(g901), .CP(CLK), .Q(g906) ) ;
DFF     gate1369  (.D(g906), .CP(CLK), .Q(g911) ) ;
DFF     gate1370  (.D(g911), .CP(CLK), .Q(g916) ) ;
DFF     gate1371  (.D(g916), .CP(CLK), .Q(g921) ) ;
DFF     gate1372  (.D(g921), .CP(CLK), .Q(g883) ) ;
INV     gate1373  (.A(II12885), .Z(g7099) ) ;
DFF     gate1374  (.D(g7099), .CP(CLK), .Q(g887) ) ;
INV     gate1375  (.A(II12888), .Z(g7100) ) ;
DFF     gate1376  (.D(g7100), .CP(CLK), .Q(g888) ) ;
INV     gate1377  (.A(II12891), .Z(g7101) ) ;
DFF     gate1378  (.D(g7101), .CP(CLK), .Q(g889) ) ;
INV     gate1379  (.A(II16176), .Z(g9386) ) ;
DFF     gate1380  (.D(g9386), .CP(CLK), .Q(g741) ) ;
INV     gate1381  (.A(II15382), .Z(g8956) ) ;
DFF     gate1382  (.D(g8956), .CP(CLK), .Q(g746) ) ;
INV     gate1383  (.A(II7302), .Z(g3833) ) ;
INV     gate1384  (.A(g3833), .Z(II5353) ) ;
INV     gate1385  (.A(II7314), .Z(g3837) ) ;
INV     gate1386  (.A(g3837), .Z(II5356) ) ;
INV     gate1387  (.A(II7320), .Z(g3839) ) ;
INV     gate1388  (.A(g3839), .Z(II5359) ) ;
INV     gate1389  (.A(II7326), .Z(g3841) ) ;
INV     gate1390  (.A(g3841), .Z(II5362) ) ;
INV     gate1391  (.A(II7332), .Z(g3843) ) ;
INV     gate1392  (.A(g3843), .Z(II5365) ) ;
INV     gate1393  (.A(II7362), .Z(g3853) ) ;
INV     gate1394  (.A(g3853), .Z(II5368) ) ;
INV     gate1395  (.A(g633), .Z(II5371) ) ;
INV     gate1396  (.A(II5371), .Z(g636) ) ;
INV     gate1397  (.A(g634), .Z(II5374) ) ;
INV     gate1398  (.A(II5374), .Z(g639) ) ;
INV     gate1399  (.A(g635), .Z(II5377) ) ;
INV     gate1400  (.A(II5377), .Z(g642) ) ;
INV     gate1401  (.A(g645), .Z(II5380) ) ;
INV     gate1402  (.A(II5380), .Z(g649) ) ;
INV     gate1403  (.A(g647), .Z(II5383) ) ;
INV     gate1404  (.A(II5383), .Z(g655) ) ;
INV     gate1405  (.A(g648), .Z(II5386) ) ;
INV     gate1406  (.A(II5386), .Z(g658) ) ;
INV     gate1407  (.A(g690), .Z(II5389) ) ;
INV     gate1408  (.A(II5389), .Z(g691) ) ;
INV     gate1409  (.A(g694), .Z(II5392) ) ;
INV     gate1410  (.A(II5392), .Z(g695) ) ;
INV     gate1411  (.A(g698), .Z(II5395) ) ;
INV     gate1412  (.A(II5395), .Z(g699) ) ;
INV     gate1413  (.A(g702), .Z(II5398) ) ;
INV     gate1414  (.A(II5398), .Z(g703) ) ;
INV     gate1415  (.A(g723), .Z(II5401) ) ;
INV     gate1416  (.A(II5401), .Z(g724) ) ;
INV     gate1417  (.A(g722), .Z(II5404) ) ;
INV     gate1418  (.A(II5404), .Z(g738) ) ;
INV     gate1419  (.A(II8874), .Z(g4653) ) ;
INV     gate1420  (.A(g4653), .Z(II5407) ) ;
INV     gate1421  (.A(II15184), .Z(g8866) ) ;
INV     gate1422  (.A(g8866), .Z(II5410) ) ;
INV     gate1423  (.A(g1016), .Z(II5413) ) ;
INV     gate1424  (.A(II5413), .Z(g1011) ) ;
INV     gate1425  (.A(II15190), .Z(g8868) ) ;
INV     gate1426  (.A(g8868), .Z(II5416) ) ;
INV     gate1427  (.A(II5471), .Z(g1603) ) ;
INV     gate1428  (.A(g1603), .Z(II5419) ) ;
INV     gate1429  (.A(g1234), .Z(II5422) ) ;
INV     gate1430  (.A(g1245), .Z(II5425) ) ;
INV     gate1431  (.A(g49), .Z(II5428) ) ;
INV     gate1432  (.A(II5428), .Z(g1555) ) ;
INV     gate1433  (.A(g65), .Z(g1556) ) ;
INV     gate1434  (.A(g1176), .Z(II5432) ) ;
INV     gate1435  (.A(II5432), .Z(g1557) ) ;
INV     gate1436  (.A(g1461), .Z(II5435) ) ;
INV     gate1437  (.A(II5435), .Z(g1558) ) ;
INV     gate1438  (.A(g636), .Z(g1562) ) ;
INV     gate1439  (.A(g639), .Z(g1563) ) ;
INV     gate1440  (.A(g642), .Z(g1564) ) ;
INV     gate1441  (.A(g649), .Z(g1565) ) ;
INV     gate1442  (.A(g652), .Z(g1566) ) ;
INV     gate1443  (.A(g655), .Z(g1567) ) ;
INV     gate1444  (.A(g658), .Z(g1568) ) ;
INV     gate1445  (.A(g661), .Z(g1569) ) ;
INV     gate1446  (.A(g665), .Z(g1570) ) ;
INV     gate1447  (.A(g669), .Z(g1571) ) ;
INV     gate1448  (.A(g673), .Z(g1572) ) ;
INV     gate1449  (.A(g677), .Z(g1573) ) ;
INV     gate1450  (.A(g681), .Z(g1574) ) ;
INV     gate1451  (.A(g685), .Z(g1575) ) ;
INV     gate1452  (.A(g691), .Z(g1576) ) ;
INV     gate1453  (.A(g695), .Z(g1577) ) ;
INV     gate1454  (.A(g699), .Z(g1578) ) ;
INV     gate1455  (.A(g703), .Z(g1579) ) ;
INV     gate1456  (.A(g706), .Z(g1580) ) ;
INV     gate1457  (.A(g710), .Z(g1581) ) ;
INV     gate1458  (.A(g714), .Z(g1582) ) ;
INV     gate1459  (.A(g718), .Z(g1583) ) ;
INV     gate1460  (.A(g738), .Z(g1584) ) ;
INV     gate1461  (.A(g724), .Z(g1585) ) ;
INV     gate1462  (.A(g730), .Z(g1586) ) ;
INV     gate1463  (.A(g734), .Z(g1587) ) ;
INV     gate1464  (.A(g741), .Z(g1588) ) ;
INV     gate1465  (.A(g746), .Z(g1589) ) ;
INV     gate1466  (.A(g926), .Z(II5466) ) ;
INV     gate1467  (.A(II5466), .Z(g1590) ) ;
INV     gate1468  (.A(g973), .Z(g1597) ) ;
INV     gate1469  (.A(g976), .Z(g1600) ) ;
INV     gate1470  (.A(g1029), .Z(II5471) ) ;
INV     gate1471  (.A(g1073), .Z(g1611) ) ;
INV     gate1472  (.A(g1084), .Z(II5475) ) ;
INV     gate1473  (.A(g1148), .Z(II5478) ) ;
INV     gate1474  (.A(II5478), .Z(g1616) ) ;
INV     gate1475  (.A(g1087), .Z(g1637) ) ;
INV     gate1476  (.A(g1092), .Z(g1638) ) ;
INV     gate1477  (.A(g1207), .Z(g1639) ) ;
INV     gate1478  (.A(g1211), .Z(g1643) ) ;
INV     gate1479  (.A(g1214), .Z(g1646) ) ;
INV     gate1480  (.A(g1217), .Z(g1649) ) ;
INV     gate1481  (.A(g1220), .Z(g1652) ) ;
INV     gate1482  (.A(g1231), .Z(g1655) ) ;
INV     gate1483  (.A(g1313), .Z(g1658) ) ;
INV     gate1484  (.A(g1405), .Z(g1661) ) ;
INV     gate1485  (.A(g1412), .Z(g1662) ) ;
INV     gate1486  (.A(g1416), .Z(g1663) ) ;
INV     gate1487  (.A(g1462), .Z(g1664) ) ;
INV     gate1488  (.A(g1467), .Z(g1665) ) ;
INV     gate1489  (.A(g1472), .Z(g1666) ) ;
INV     gate1490  (.A(g1481), .Z(g1667) ) ;
INV     gate1491  (.A(g1489), .Z(g1670) ) ;
INV     gate1492  (.A(g1494), .Z(g1671) ) ;
INV     gate1493  (.A(g1499), .Z(g1672) ) ;
INV     gate1494  (.A(g1504), .Z(g1673) ) ;
INV     gate1495  (.A(g1514), .Z(g1674) ) ;
INV     gate1496  (.A(g1519), .Z(g1675) ) ;
INV     gate1497  (.A(g727), .Z(g1676) ) ;
INV     gate1498  (.A(g1532), .Z(g1677) ) ;
INV     gate1499  (.A(g557), .Z(II5512) ) ;
INV     gate1500  (.A(II5512), .Z(g1679) ) ;
INV     gate1501  (.A(g567), .Z(II5515) ) ;
INV     gate1502  (.A(II5515), .Z(g1680) ) ;
INV     gate1503  (.A(g929), .Z(g1681) ) ;
INV     gate1504  (.A(g795), .Z(g1683) ) ;
INV     gate1505  (.A(g1), .Z(g1684) ) ;
INV     gate1506  (.A(g43), .Z(II5528) ) ;
INV     gate1507  (.A(II5528), .Z(g1685) ) ;
INV     gate1508  (.A(g866), .Z(II5531) ) ;
INV     gate1509  (.A(II5531), .Z(g1686) ) ;
INV     gate1510  (.A(g10), .Z(g1687) ) ;
INV     gate1511  (.A(g48), .Z(II5535) ) ;
INV     gate1512  (.A(II5535), .Z(g1688) ) ;
INV     gate1513  (.A(g855), .Z(g1689) ) ;
INV     gate1514  (.A(g21), .Z(g1694) ) ;
INV     gate1515  (.A(g778), .Z(g1695) ) ;
INV     gate1516  (.A(g1272), .Z(II5542) ) ;
INV     gate1517  (.A(II5542), .Z(g1698) ) ;
INV     gate1518  (.A(g1276), .Z(II5545) ) ;
INV     gate1519  (.A(II5545), .Z(g1701) ) ;
INV     gate1520  (.A(g1280), .Z(II5548) ) ;
INV     gate1521  (.A(II5548), .Z(g1704) ) ;
INV     gate1522  (.A(g955), .Z(g1707) ) ;
INV     gate1523  (.A(g1284), .Z(II5552) ) ;
INV     gate1524  (.A(II5552), .Z(g1708) ) ;
INV     gate1525  (.A(g1288), .Z(II5555) ) ;
INV     gate1526  (.A(II5555), .Z(g1711) ) ;
INV     gate1527  (.A(g1292), .Z(II5559) ) ;
INV     gate1528  (.A(II5559), .Z(g1715) ) ;
INV     gate1529  (.A(g1300), .Z(II5562) ) ;
INV     gate1530  (.A(II5562), .Z(g1718) ) ;
INV     gate1531  (.A(g1296), .Z(II5565) ) ;
INV     gate1532  (.A(II5565), .Z(g1721) ) ;
INV     gate1533  (.A(g1409), .Z(II5568) ) ;
INV     gate1534  (.A(g158), .Z(g1726) ) ;
INV     gate1535  (.A(g596), .Z(g1727) ) ;
INV     gate1536  (.A(g1439), .Z(g1732) ) ;
INV     gate1537  (.A(g172), .Z(II5577) ) ;
INV     gate1538  (.A(II5577), .Z(g1736) ) ;
INV     gate1539  (.A(g597), .Z(g1737) ) ;
INV     gate1540  (.A(g741), .Z(g1738) ) ;
INV     gate1541  (.A(g1486), .Z(g1742) ) ;
INV     gate1542  (.A(g598), .Z(g1743) ) ;
INV     gate1543  (.A(g600), .Z(g1744) ) ;
INV     gate1544  (.A(g746), .Z(g1745) ) ;
INV     gate1545  (.A(g290), .Z(g1746) ) ;
INV     gate1546  (.A(g599), .Z(g1747) ) ;
INV     gate1547  (.A(g601), .Z(g1748) ) ;
INV     gate1548  (.A(g371), .Z(g1749) ) ;
INV     gate1549  (.A(g602), .Z(g1750) ) ;
INV     gate1550  (.A(g452), .Z(g1751) ) ;
INV     gate1551  (.A(g603), .Z(g1752) ) ;
INV     gate1552  (.A(g533), .Z(g1756) ) ;
INV     gate1553  (.A(g604), .Z(g1757) ) ;
INV     gate1554  (.A(g1084), .Z(g1758) ) ;
INV     gate1555  (.A(g58), .Z(II5605) ) ;
INV     gate1556  (.A(II5605), .Z(g1760) ) ;
INV     gate1557  (.A(g605), .Z(g1768) ) ;
INV     gate1558  (.A(g16), .Z(II5609) ) ;
INV     gate1559  (.A(II5609), .Z(g1769) ) ;
INV     gate1560  (.A(g606), .Z(g1770) ) ;
INV     gate1561  (.A(g609), .Z(g1771) ) ;
INV     gate1562  (.A(g607), .Z(g1772) ) ;
INV     gate1563  (.A(g610), .Z(g1773) ) ;
INV     gate1564  (.A(g979), .Z(II5616) ) ;
INV     gate1565  (.A(II5616), .Z(g1774) ) ;
INV     gate1566  (.A(g608), .Z(g1776) ) ;
INV     gate1567  (.A(g611), .Z(g1777) ) ;
INV     gate1568  (.A(g613), .Z(g1778) ) ;
INV     gate1569  (.A(g612), .Z(g1779) ) ;
INV     gate1570  (.A(g614), .Z(g1780) ) ;
INV     gate1571  (.A(g622), .Z(g1781) ) ;
INV     gate1572  (.A(g624), .Z(g1782) ) ;
INV     gate1573  (.A(g891), .Z(II5633) ) ;
INV     gate1574  (.A(g891), .Z(II5636) ) ;
INV     gate1575  (.A(II5636), .Z(g1784) ) ;
INV     gate1576  (.A(g615), .Z(g1785) ) ;
INV     gate1577  (.A(g623), .Z(g1786) ) ;
INV     gate1578  (.A(g625), .Z(g1787) ) ;
INV     gate1579  (.A(g984), .Z(g1788) ) ;
INV     gate1580  (.A(g1034), .Z(g1789) ) ;
INV     gate1581  (.A(g616), .Z(g1792) ) ;
INV     gate1582  (.A(g626), .Z(g1793) ) ;
INV     gate1583  (.A(g883), .Z(II5646) ) ;
INV     gate1584  (.A(II5646), .Z(g1794) ) ;
INV     gate1585  (.A(g1389), .Z(II5649) ) ;
INV     gate1586  (.A(II5649), .Z(g1795) ) ;
INV     gate1587  (.A(g617), .Z(g1796) ) ;
INV     gate1588  (.A(g627), .Z(g1797) ) ;
INV     gate1589  (.A(g921), .Z(II5654) ) ;
INV     gate1590  (.A(g921), .Z(II5657) ) ;
INV     gate1591  (.A(II5657), .Z(g1799) ) ;
INV     gate1592  (.A(g1477), .Z(g1800) ) ;
INV     gate1593  (.A(g618), .Z(g1801) ) ;
INV     gate1594  (.A(g628), .Z(g1802) ) ;
INV     gate1595  (.A(g758), .Z(g1803) ) ;
INV     gate1596  (.A(g916), .Z(II5664) ) ;
INV     gate1597  (.A(g916), .Z(II5667) ) ;
INV     gate1598  (.A(II5667), .Z(g1805) ) ;
INV     gate1599  (.A(g941), .Z(II5670) ) ;
INV     gate1600  (.A(II5670), .Z(g1806) ) ;
INV     gate1601  (.A(g619), .Z(g1807) ) ;
INV     gate1602  (.A(g629), .Z(g1808) ) ;
INV     gate1603  (.A(g759), .Z(g1809) ) ;
INV     gate1604  (.A(g911), .Z(II5676) ) ;
INV     gate1605  (.A(g911), .Z(II5679) ) ;
INV     gate1606  (.A(II5679), .Z(g1811) ) ;
INV     gate1607  (.A(g168), .Z(II5682) ) ;
INV     gate1608  (.A(II5682), .Z(g1812) ) ;
INV     gate1609  (.A(g620), .Z(g1813) ) ;
INV     gate1610  (.A(g630), .Z(g1814) ) ;
INV     gate1611  (.A(g760), .Z(g1815) ) ;
INV     gate1612  (.A(g767), .Z(g1816) ) ;
INV     gate1613  (.A(g906), .Z(II5689) ) ;
INV     gate1614  (.A(g906), .Z(II5692) ) ;
INV     gate1615  (.A(II5692), .Z(g1818) ) ;
INV     gate1616  (.A(g621), .Z(g1820) ) ;
INV     gate1617  (.A(g631), .Z(g1821) ) ;
INV     gate1618  (.A(g761), .Z(g1822) ) ;
INV     gate1619  (.A(g768), .Z(g1823) ) ;
INV     gate1620  (.A(g901), .Z(II5706) ) ;
INV     gate1621  (.A(g901), .Z(II5709) ) ;
INV     gate1622  (.A(II5709), .Z(g1825) ) ;
INV     gate1623  (.A(g632), .Z(g1826) ) ;
INV     gate1624  (.A(g762), .Z(g1827) ) ;
INV     gate1625  (.A(g769), .Z(g1828) ) ;
INV     gate1626  (.A(g896), .Z(II5715) ) ;
INV     gate1627  (.A(g896), .Z(II5718) ) ;
INV     gate1628  (.A(II5718), .Z(g1830) ) ;
INV     gate1629  (.A(g689), .Z(g1831) ) ;
INV     gate1630  (.A(g763), .Z(g1832) ) ;
INV     gate1631  (.A(g770), .Z(g1833) ) ;
INV     gate1632  (.A(g1007), .Z(g1837) ) ;
INV     gate1633  (.A(g1450), .Z(g1838) ) ;
INV     gate1634  (.A(g764), .Z(g1842) ) ;
INV     gate1635  (.A(g771), .Z(g1843) ) ;
INV     gate1636  (.A(g765), .Z(g1847) ) ;
INV     gate1637  (.A(g772), .Z(g1848) ) ;
INV     gate1638  (.A(g859), .Z(II5732) ) ;
INV     gate1639  (.A(II5732), .Z(g1849) ) ;
INV     gate1640  (.A(g887), .Z(g1852) ) ;
INV     gate1641  (.A(g766), .Z(g1853) ) ;
INV     gate1642  (.A(g773), .Z(g1854) ) ;
INV     gate1643  (.A(g866), .Z(g1855) ) ;
INV     gate1644  (.A(g774), .Z(g1856) ) ;
INV     gate1645  (.A(g889), .Z(g1857) ) ;
INV     gate1646  (.A(g162), .Z(g1860) ) ;
INV     gate1647  (.A(g68), .Z(g1863) ) ;
INV     gate1648  (.A(g162), .Z(g1864) ) ;
INV     gate1649  (.A(g1013), .Z(g1865) ) ;
INV     gate1650  (.A(g71), .Z(g1866) ) ;
INV     gate1651  (.A(g878), .Z(g1867) ) ;
INV     gate1652  (.A(g1260), .Z(II5747) ) ;
INV     gate1653  (.A(II5747), .Z(g1868) ) ;
INV     gate1654  (.A(g74), .Z(g1869) ) ;
INV     gate1655  (.A(g963), .Z(II5751) ) ;
INV     gate1656  (.A(g966), .Z(II5754) ) ;
INV     gate1657  (.A(g77), .Z(g1876) ) ;
INV     gate1658  (.A(g595), .Z(g1877) ) ;
INV     gate1659  (.A(g80), .Z(g1878) ) ;
INV     gate1660  (.A(g1207), .Z(II5763) ) ;
INV     gate1661  (.A(II5763), .Z(g1879) ) ;
INV     gate1662  (.A(g1254), .Z(II5766) ) ;
INV     gate1663  (.A(II5766), .Z(g1886) ) ;
INV     gate1664  (.A(g83), .Z(g1887) ) ;
INV     gate1665  (.A(g781), .Z(g1888) ) ;
INV     gate1666  (.A(g1018), .Z(g1889) ) ;
INV     gate1667  (.A(g1240), .Z(II5772) ) ;
INV     gate1668  (.A(g1240), .Z(II5775) ) ;
INV     gate1669  (.A(II5775), .Z(g1895) ) ;
INV     gate1670  (.A(g86), .Z(g1896) ) ;
INV     gate1671  (.A(g789), .Z(g1897) ) ;
INV     gate1672  (.A(g979), .Z(II5781) ) ;
INV     gate1673  (.A(II5781), .Z(g1901) ) ;
INV     gate1674  (.A(g1021), .Z(g1904) ) ;
INV     gate1675  (.A(g52), .Z(g1907) ) ;
INV     gate1676  (.A(g812), .Z(g1908) ) ;
INV     gate1677  (.A(g998), .Z(g1909) ) ;
INV     gate1678  (.A(g1524), .Z(II5789) ) ;
INV     gate1679  (.A(g1524), .Z(g1912) ) ;
INV     gate1680  (.A(g775), .Z(g1916) ) ;
INV     gate1681  (.A(g1236), .Z(II5795) ) ;
INV     gate1682  (.A(II5795), .Z(g1917) ) ;
INV     gate1683  (.A(g822), .Z(g1918) ) ;
INV     gate1684  (.A(g1251), .Z(g1922) ) ;
INV     gate1685  (.A(g1424), .Z(II5801) ) ;
INV     gate1686  (.A(II5801), .Z(g1923) ) ;
INV     gate1687  (.A(g174), .Z(g1924) ) ;
INV     gate1688  (.A(g825), .Z(g1925) ) ;
INV     gate1689  (.A(g874), .Z(g1926) ) ;
INV     gate1690  (.A(g1224), .Z(g1929) ) ;
INV     gate1691  (.A(g1247), .Z(g1933) ) ;
INV     gate1692  (.A(g154), .Z(g1934) ) ;
INV     gate1693  (.A(g1280), .Z(g1935) ) ;
INV     gate1694  (.A(g1288), .Z(g1938) ) ;
INV     gate1695  (.A(g1243), .Z(II5812) ) ;
INV     gate1696  (.A(II5812), .Z(g1941) ) ;
INV     gate1697  (.A(g828), .Z(g1942) ) ;
INV     gate1698  (.A(g1025), .Z(g1943) ) ;
INV     gate1699  (.A(g1081), .Z(II5817) ) ;
INV     gate1700  (.A(g1081), .Z(g1945) ) ;
INV     gate1701  (.A(g1250), .Z(g1948) ) ;
INV     gate1702  (.A(g1292), .Z(g1949) ) ;
INV     gate1703  (.A(g1333), .Z(g1952) ) ;
INV     gate1704  (.A(g786), .Z(g1958) ) ;
INV     gate1705  (.A(g1252), .Z(g1959) ) ;
INV     gate1706  (.A(g1268), .Z(g1960) ) ;
INV     gate1707  (.A(g1345), .Z(g1961) ) ;
INV     gate1708  (.A(g1432), .Z(g1967) ) ;
INV     gate1709  (.A(g1194), .Z(II5831) ) ;
INV     gate1710  (.A(II5831), .Z(g1970) ) ;
INV     gate1711  (.A(g803), .Z(g1974) ) ;
INV     gate1712  (.A(g1253), .Z(g1975) ) ;
INV     gate1713  (.A(g1269), .Z(g1976) ) ;
INV     gate1714  (.A(g1357), .Z(g1977) ) ;
INV     gate1715  (.A(g1198), .Z(II5839) ) ;
INV     gate1716  (.A(II5839), .Z(g1983) ) ;
INV     gate1717  (.A(g68), .Z(II5842) ) ;
INV     gate1718  (.A(II5842), .Z(g1987) ) ;
INV     gate1719  (.A(g806), .Z(g2006) ) ;
INV     gate1720  (.A(g1223), .Z(g2007) ) ;
INV     gate1721  (.A(g1360), .Z(II5847) ) ;
INV     gate1722  (.A(II5847), .Z(g2011) ) ;
INV     gate1723  (.A(g33), .Z(g2015) ) ;
INV     gate1724  (.A(g1202), .Z(II5852) ) ;
INV     gate1725  (.A(II5852), .Z(g2016) ) ;
INV     gate1726  (.A(g71), .Z(II5855) ) ;
INV     gate1727  (.A(II5855), .Z(g2020) ) ;
INV     gate1728  (.A(g809), .Z(g2038) ) ;
INV     gate1729  (.A(g1228), .Z(g2039) ) ;
INV     gate1730  (.A(g1313), .Z(II5861) ) ;
INV     gate1731  (.A(II5861), .Z(g2044) ) ;
INV     gate1732  (.A(g1206), .Z(II5865) ) ;
INV     gate1733  (.A(II5865), .Z(g2052) ) ;
INV     gate1734  (.A(g74), .Z(II5868) ) ;
INV     gate1735  (.A(II5868), .Z(g2057) ) ;
INV     gate1736  (.A(g1254), .Z(g2073) ) ;
INV     gate1737  (.A(g77), .Z(II5872) ) ;
INV     gate1738  (.A(II5872), .Z(g2074) ) ;
INV     gate1739  (.A(g819), .Z(g2091) ) ;
INV     gate1740  (.A(g1225), .Z(g2092) ) ;
INV     gate1741  (.A(g1226), .Z(g2096) ) ;
INV     gate1742  (.A(g1227), .Z(g2100) ) ;
INV     gate1743  (.A(g1267), .Z(II5879) ) ;
INV     gate1744  (.A(II5879), .Z(g2104) ) ;
INV     gate1745  (.A(g1444), .Z(g2105) ) ;
INV     gate1746  (.A(g80), .Z(II5883) ) ;
INV     gate1747  (.A(II5883), .Z(g2106) ) ;
INV     gate1748  (.A(g1284), .Z(g2128) ) ;
INV     gate1749  (.A(g1300), .Z(g2131) ) ;
INV     gate1750  (.A(g1317), .Z(g2134) ) ;
INV     gate1751  (.A(g83), .Z(II5889) ) ;
INV     gate1752  (.A(II5889), .Z(g2137) ) ;
INV     gate1753  (.A(g1296), .Z(g2145) ) ;
INV     gate1754  (.A(g1304), .Z(g2148) ) ;
INV     gate1755  (.A(g86), .Z(II5894) ) ;
INV     gate1756  (.A(II5894), .Z(g2149) ) ;
INV     gate1757  (.A(g173), .Z(II5897) ) ;
INV     gate1758  (.A(II5897), .Z(g2157) ) ;
INV     gate1759  (.A(g1454), .Z(g2161) ) ;
INV     gate1760  (.A(g52), .Z(II5901) ) ;
INV     gate1761  (.A(II5901), .Z(g2162) ) ;
INV     gate1762  (.A(g1229), .Z(g2170) ) ;
INV     gate1763  (.A(g1319), .Z(g2174) ) ;
INV     gate1764  (.A(g1322), .Z(g2177) ) ;
INV     gate1765  (.A(g1318), .Z(g2180) ) ;
INV     gate1766  (.A(g196), .Z(II5908) ) ;
INV     gate1767  (.A(II5908), .Z(g2183) ) ;
INV     gate1768  (.A(g216), .Z(II5911) ) ;
INV     gate1769  (.A(II5911), .Z(g2184) ) ;
INV     gate1770  (.A(g1097), .Z(II5914) ) ;
INV     gate1771  (.A(II5914), .Z(g2185) ) ;
INV     gate1772  (.A(g1321), .Z(g2202) ) ;
INV     gate1773  (.A(g13), .Z(g2205) ) ;
INV     gate1774  (.A(g219), .Z(II5920) ) ;
INV     gate1775  (.A(II5920), .Z(g2207) ) ;
INV     gate1776  (.A(g252), .Z(II5923) ) ;
INV     gate1777  (.A(II5923), .Z(g2208) ) ;
INV     gate1778  (.A(g297), .Z(II5926) ) ;
INV     gate1779  (.A(II5926), .Z(g2209) ) ;
INV     gate1780  (.A(g1326), .Z(g2210) ) ;
INV     gate1781  (.A(g1416), .Z(g2215) ) ;
INV     gate1782  (.A(g1158), .Z(II5933) ) ;
INV     gate1783  (.A(II5933), .Z(g2216) ) ;
INV     gate1784  (.A(g222), .Z(II5936) ) ;
INV     gate1785  (.A(II5936), .Z(g2221) ) ;
INV     gate1786  (.A(g275), .Z(II5939) ) ;
INV     gate1787  (.A(II5939), .Z(g2222) ) ;
INV     gate1788  (.A(g300), .Z(II5942) ) ;
INV     gate1789  (.A(II5942), .Z(g2223) ) ;
INV     gate1790  (.A(g333), .Z(II5945) ) ;
INV     gate1791  (.A(II5945), .Z(g2224) ) ;
INV     gate1792  (.A(g378), .Z(II5948) ) ;
INV     gate1793  (.A(II5948), .Z(g2225) ) ;
INV     gate1794  (.A(g1320), .Z(g2226) ) ;
INV     gate1795  (.A(g89), .Z(II5954) ) ;
INV     gate1796  (.A(II5954), .Z(g2231) ) ;
INV     gate1797  (.A(g110), .Z(II5957) ) ;
INV     gate1798  (.A(II5957), .Z(g2232) ) ;
INV     gate1799  (.A(g187), .Z(II5960) ) ;
INV     gate1800  (.A(II5960), .Z(g2233) ) ;
INV     gate1801  (.A(g225), .Z(II5963) ) ;
INV     gate1802  (.A(II5963), .Z(g2234) ) ;
INV     gate1803  (.A(g278), .Z(II5966) ) ;
INV     gate1804  (.A(II5966), .Z(g2235) ) ;
INV     gate1805  (.A(g303), .Z(II5969) ) ;
INV     gate1806  (.A(II5969), .Z(g2236) ) ;
INV     gate1807  (.A(g356), .Z(II5972) ) ;
INV     gate1808  (.A(II5972), .Z(g2237) ) ;
INV     gate1809  (.A(g381), .Z(II5975) ) ;
INV     gate1810  (.A(II5975), .Z(g2238) ) ;
INV     gate1811  (.A(g414), .Z(II5978) ) ;
INV     gate1812  (.A(II5978), .Z(g2239) ) ;
INV     gate1813  (.A(g459), .Z(II5981) ) ;
INV     gate1814  (.A(II5981), .Z(g2240) ) ;
INV     gate1815  (.A(g540), .Z(II5984) ) ;
INV     gate1816  (.A(II5984), .Z(g2241) ) ;
INV     gate1817  (.A(g985), .Z(g2242) ) ;
INV     gate1818  (.A(g999), .Z(g2245) ) ;
INV     gate1819  (.A(g1460), .Z(II5989) ) ;
INV     gate1820  (.A(II5989), .Z(g2246) ) ;
INV     gate1821  (.A(g1323), .Z(g2253) ) ;
INV     gate1822  (.A(g1324), .Z(g2256) ) ;
INV     gate1823  (.A(g1325), .Z(g2259) ) ;
INV     gate1824  (.A(g1394), .Z(g2263) ) ;
INV     gate1825  (.A(g114), .Z(II5997) ) ;
INV     gate1826  (.A(II5997), .Z(g2264) ) ;
INV     gate1827  (.A(g202), .Z(II6000) ) ;
INV     gate1828  (.A(II6000), .Z(g2265) ) ;
INV     gate1829  (.A(g228), .Z(II6003) ) ;
INV     gate1830  (.A(II6003), .Z(g2266) ) ;
INV     gate1831  (.A(g306), .Z(II6006) ) ;
INV     gate1832  (.A(II6006), .Z(g2267) ) ;
INV     gate1833  (.A(g359), .Z(II6009) ) ;
INV     gate1834  (.A(II6009), .Z(g2268) ) ;
INV     gate1835  (.A(g384), .Z(II6012) ) ;
INV     gate1836  (.A(II6012), .Z(g2269) ) ;
INV     gate1837  (.A(g437), .Z(II6015) ) ;
INV     gate1838  (.A(II6015), .Z(g2270) ) ;
INV     gate1839  (.A(g462), .Z(II6018) ) ;
INV     gate1840  (.A(II6018), .Z(g2271) ) ;
INV     gate1841  (.A(g495), .Z(II6021) ) ;
INV     gate1842  (.A(II6021), .Z(g2272) ) ;
INV     gate1843  (.A(g544), .Z(II6024) ) ;
INV     gate1844  (.A(II6024), .Z(g2273) ) ;
INV     gate1845  (.A(g782), .Z(g2274) ) ;
INV     gate1846  (.A(g990), .Z(g2275) ) ;
INV     gate1847  (.A(g1207), .Z(II6029) ) ;
INV     gate1848  (.A(II6029), .Z(g2276) ) ;
INV     gate1849  (.A(g1400), .Z(g2282) ) ;
INV     gate1850  (.A(g3), .Z(II6033) ) ;
INV     gate1851  (.A(II6033), .Z(g2283) ) ;
INV     gate1852  (.A(g130), .Z(II6036) ) ;
INV     gate1853  (.A(II6036), .Z(g2284) ) ;
INV     gate1854  (.A(g207), .Z(II6039) ) ;
INV     gate1855  (.A(II6039), .Z(g2285) ) ;
INV     gate1856  (.A(g237), .Z(II6042) ) ;
INV     gate1857  (.A(II6042), .Z(g2286) ) ;
INV     gate1858  (.A(g309), .Z(II6045) ) ;
INV     gate1859  (.A(II6045), .Z(g2287) ) ;
INV     gate1860  (.A(g387), .Z(II6048) ) ;
INV     gate1861  (.A(II6048), .Z(g2288) ) ;
INV     gate1862  (.A(g440), .Z(II6051) ) ;
INV     gate1863  (.A(II6051), .Z(g2289) ) ;
INV     gate1864  (.A(g465), .Z(II6054) ) ;
INV     gate1865  (.A(II6054), .Z(g2290) ) ;
INV     gate1866  (.A(g518), .Z(II6057) ) ;
INV     gate1867  (.A(II6057), .Z(g2291) ) ;
INV     gate1868  (.A(g580), .Z(II6060) ) ;
INV     gate1869  (.A(II6060), .Z(g2292) ) ;
INV     gate1870  (.A(g888), .Z(g2293) ) ;
INV     gate1871  (.A(g995), .Z(g2295) ) ;
INV     gate1872  (.A(g1211), .Z(II6072) ) ;
INV     gate1873  (.A(II6072), .Z(g2298) ) ;
INV     gate1874  (.A(g2), .Z(II6075) ) ;
INV     gate1875  (.A(II6075), .Z(g2306) ) ;
INV     gate1876  (.A(g95), .Z(II6078) ) ;
INV     gate1877  (.A(II6078), .Z(g2307) ) ;
INV     gate1878  (.A(g118), .Z(II6081) ) ;
INV     gate1879  (.A(II6081), .Z(g2308) ) ;
INV     gate1880  (.A(g240), .Z(II6084) ) ;
INV     gate1881  (.A(II6084), .Z(g2309) ) ;
INV     gate1882  (.A(g318), .Z(II6087) ) ;
INV     gate1883  (.A(II6087), .Z(g2310) ) ;
INV     gate1884  (.A(g390), .Z(II6090) ) ;
INV     gate1885  (.A(II6090), .Z(g2311) ) ;
INV     gate1886  (.A(g468), .Z(II6093) ) ;
INV     gate1887  (.A(II6093), .Z(g2312) ) ;
INV     gate1888  (.A(g521), .Z(II6096) ) ;
INV     gate1889  (.A(II6096), .Z(g2313) ) ;
INV     gate1890  (.A(g584), .Z(II6099) ) ;
INV     gate1891  (.A(II6099), .Z(g2314) ) ;
INV     gate1892  (.A(g1214), .Z(II6109) ) ;
INV     gate1893  (.A(II6109), .Z(g2316) ) ;
INV     gate1894  (.A(g4), .Z(II6112) ) ;
INV     gate1895  (.A(II6112), .Z(g2323) ) ;
INV     gate1896  (.A(g134), .Z(II6115) ) ;
INV     gate1897  (.A(II6115), .Z(g2324) ) ;
INV     gate1898  (.A(g243), .Z(II6118) ) ;
INV     gate1899  (.A(II6118), .Z(g2325) ) ;
INV     gate1900  (.A(g321), .Z(II6121) ) ;
INV     gate1901  (.A(II6121), .Z(g2326) ) ;
INV     gate1902  (.A(g399), .Z(II6124) ) ;
INV     gate1903  (.A(II6124), .Z(g2327) ) ;
INV     gate1904  (.A(g471), .Z(II6127) ) ;
INV     gate1905  (.A(II6127), .Z(g2328) ) ;
INV     gate1906  (.A(g560), .Z(II6130) ) ;
INV     gate1907  (.A(II6130), .Z(g2329) ) ;
INV     gate1908  (.A(g933), .Z(g2331) ) ;
INV     gate1909  (.A(g926), .Z(g2332) ) ;
INV     gate1910  (.A(g1217), .Z(II6143) ) ;
INV     gate1911  (.A(II6143), .Z(g2334) ) ;
INV     gate1912  (.A(g1327), .Z(g2340) ) ;
INV     gate1913  (.A(g1392), .Z(g2343) ) ;
INV     gate1914  (.A(g5), .Z(II6148) ) ;
INV     gate1915  (.A(II6148), .Z(g2344) ) ;
INV     gate1916  (.A(g12), .Z(II6151) ) ;
INV     gate1917  (.A(II6151), .Z(g2345) ) ;
INV     gate1918  (.A(g122), .Z(II6154) ) ;
INV     gate1919  (.A(II6154), .Z(g2346) ) ;
INV     gate1920  (.A(g246), .Z(II6157) ) ;
INV     gate1921  (.A(II6157), .Z(g2347) ) ;
INV     gate1922  (.A(g324), .Z(II6160) ) ;
INV     gate1923  (.A(II6160), .Z(g2348) ) ;
INV     gate1924  (.A(g402), .Z(II6163) ) ;
INV     gate1925  (.A(II6163), .Z(g2349) ) ;
INV     gate1926  (.A(g480), .Z(II6166) ) ;
INV     gate1927  (.A(II6166), .Z(g2350) ) ;
INV     gate1928  (.A(g792), .Z(g2351) ) ;
INV     gate1929  (.A(g871), .Z(g2353) ) ;
INV     gate1930  (.A(g1220), .Z(II6178) ) ;
INV     gate1931  (.A(II6178), .Z(g2354) ) ;
INV     gate1932  (.A(g1397), .Z(g2359) ) ;
INV     gate1933  (.A(g1435), .Z(g2360) ) ;
INV     gate1934  (.A(g6), .Z(II6183) ) ;
INV     gate1935  (.A(II6183), .Z(g2361) ) ;
INV     gate1936  (.A(g138), .Z(II6186) ) ;
INV     gate1937  (.A(II6186), .Z(g2362) ) ;
INV     gate1938  (.A(g249), .Z(II6189) ) ;
INV     gate1939  (.A(II6189), .Z(g2363) ) ;
INV     gate1940  (.A(g327), .Z(II6192) ) ;
INV     gate1941  (.A(II6192), .Z(g2364) ) ;
INV     gate1942  (.A(g405), .Z(II6195) ) ;
INV     gate1943  (.A(II6195), .Z(g2365) ) ;
INV     gate1944  (.A(g483), .Z(II6198) ) ;
INV     gate1945  (.A(II6198), .Z(g2366) ) ;
INV     gate1946  (.A(g944), .Z(g2371) ) ;
INV     gate1947  (.A(g7), .Z(II6214) ) ;
INV     gate1948  (.A(II6214), .Z(g2372) ) ;
INV     gate1949  (.A(g105), .Z(II6217) ) ;
INV     gate1950  (.A(II6217), .Z(g2373) ) ;
INV     gate1951  (.A(g126), .Z(II6220) ) ;
INV     gate1952  (.A(II6220), .Z(g2374) ) ;
INV     gate1953  (.A(g330), .Z(II6223) ) ;
INV     gate1954  (.A(II6223), .Z(g2375) ) ;
INV     gate1955  (.A(g408), .Z(II6226) ) ;
INV     gate1956  (.A(II6226), .Z(g2376) ) ;
INV     gate1957  (.A(g486), .Z(II6229) ) ;
INV     gate1958  (.A(II6229), .Z(g2377) ) ;
INV     gate1959  (.A(g8), .Z(II6239) ) ;
INV     gate1960  (.A(II6239), .Z(g2379) ) ;
INV     gate1961  (.A(g1554), .Z(II6242) ) ;
INV     gate1962  (.A(II6242), .Z(g2380) ) ;
INV     gate1963  (.A(g142), .Z(II6245) ) ;
INV     gate1964  (.A(II6245), .Z(g2381) ) ;
INV     gate1965  (.A(g411), .Z(II6248) ) ;
INV     gate1966  (.A(II6248), .Z(g2382) ) ;
INV     gate1967  (.A(g489), .Z(II6251) ) ;
INV     gate1968  (.A(II6251), .Z(g2383) ) ;
INV     gate1969  (.A(g536), .Z(II6254) ) ;
INV     gate1970  (.A(II6254), .Z(g2384) ) ;
INV     gate1971  (.A(g1230), .Z(g2389) ) ;
INV     gate1972  (.A(g11), .Z(g2392) ) ;
INV     gate1973  (.A(g100), .Z(II6267) ) ;
INV     gate1974  (.A(II6267), .Z(g2393) ) ;
INV     gate1975  (.A(g492), .Z(II6270) ) ;
INV     gate1976  (.A(II6270), .Z(g2394) ) ;
INV     gate1977  (.A(g1033), .Z(g2396) ) ;
INV     gate1978  (.A(g1272), .Z(g2397) ) ;
INV     gate1979  (.A(g22), .Z(g2401) ) ;
INV     gate1980  (.A(g29), .Z(g2402) ) ;
INV     gate1981  (.A(g1176), .Z(g2403) ) ;
INV     gate1982  (.A(g1276), .Z(g2404) ) ;
INV     gate1983  (.A(g1307), .Z(II6286) ) ;
INV     gate1984  (.A(II6286), .Z(g2407) ) ;
INV     gate1985  (.A(g1329), .Z(g2424) ) ;
INV     gate1986  (.A(g23), .Z(g2452) ) ;
INV     gate1987  (.A(g46), .Z(II6291) ) ;
INV     gate1988  (.A(II6291), .Z(g2453) ) ;
INV     gate1989  (.A(g1330), .Z(II6294) ) ;
INV     gate1990  (.A(II6294), .Z(g2454) ) ;
INV     gate1991  (.A(g24), .Z(g2457) ) ;
INV     gate1992  (.A(g30), .Z(g2458) ) ;
INV     gate1993  (.A(g47), .Z(II6299) ) ;
INV     gate1994  (.A(II6299), .Z(g2459) ) ;
INV     gate1995  (.A(g1313), .Z(II6302) ) ;
INV     gate1996  (.A(II6302), .Z(g2460) ) ;
INV     gate1997  (.A(g1333), .Z(II6305) ) ;
INV     gate1998  (.A(II6305), .Z(g2467) ) ;
INV     gate1999  (.A(g42), .Z(g2470) ) ;
INV     gate2000  (.A(g1336), .Z(II6309) ) ;
INV     gate2001  (.A(II6309), .Z(g2471) ) ;
INV     gate2002  (.A(g25), .Z(g2477) ) ;
INV     gate2003  (.A(g31), .Z(g2478) ) ;
INV     gate2004  (.A(g32), .Z(g2479) ) ;
INV     gate2005  (.A(g44), .Z(g2480) ) ;
INV     gate2006  (.A(g1339), .Z(II6317) ) ;
INV     gate2007  (.A(II6317), .Z(g2481) ) ;
INV     gate2008  (.A(g45), .Z(g2484) ) ;
INV     gate2009  (.A(g62), .Z(g2485) ) ;
INV     gate2010  (.A(g959), .Z(g2486) ) ;
INV     gate2011  (.A(g1342), .Z(II6323) ) ;
INV     gate2012  (.A(II6323), .Z(g2487) ) ;
INV     gate2013  (.A(g1443), .Z(II6326) ) ;
INV     gate2014  (.A(II6326), .Z(g2490) ) ;
INV     gate2015  (.A(g9), .Z(g2494) ) ;
INV     gate2016  (.A(g26), .Z(g2495) ) ;
INV     gate2017  (.A(g942), .Z(g2496) ) ;
INV     gate2018  (.A(g945), .Z(g2497) ) ;
INV     gate2019  (.A(g1345), .Z(II6333) ) ;
INV     gate2020  (.A(II6333), .Z(g2498) ) ;
INV     gate2021  (.A(g27), .Z(g2501) ) ;
INV     gate2022  (.A(g1348), .Z(II6337) ) ;
INV     gate2023  (.A(II6337), .Z(g2502) ) ;
INV     gate2024  (.A(g28), .Z(g2505) ) ;
INV     gate2025  (.A(g1351), .Z(II6341) ) ;
INV     gate2026  (.A(II6341), .Z(g2506) ) ;
INV     gate2027  (.A(g37), .Z(g2509) ) ;
INV     gate2028  (.A(g58), .Z(g2510) ) ;
INV     gate2029  (.A(g1328), .Z(g2511) ) ;
INV     gate2030  (.A(g1330), .Z(g2514) ) ;
INV     gate2031  (.A(g1354), .Z(II6348) ) ;
INV     gate2032  (.A(II6348), .Z(g2517) ) ;
INV     gate2033  (.A(g41), .Z(g2520) ) ;
INV     gate2034  (.A(g1342), .Z(g2522) ) ;
INV     gate2035  (.A(g1357), .Z(II6354) ) ;
INV     gate2036  (.A(II6354), .Z(g2525) ) ;
INV     gate2037  (.A(g1260), .Z(g2528) ) ;
INV     gate2038  (.A(g13), .Z(II6358) ) ;
INV     gate2039  (.A(II6358), .Z(g2532) ) ;
INV     gate2040  (.A(g1336), .Z(g2533) ) ;
INV     gate2041  (.A(g1354), .Z(g2536) ) ;
INV     gate2042  (.A(g16), .Z(II6363) ) ;
INV     gate2043  (.A(II6363), .Z(g2539) ) ;
INV     gate2044  (.A(g1339), .Z(g2540) ) ;
INV     gate2045  (.A(g1348), .Z(g2543) ) ;
INV     gate2046  (.A(g20), .Z(II6368) ) ;
INV     gate2047  (.A(II6368), .Z(g2546) ) ;
INV     gate2048  (.A(g33), .Z(II6371) ) ;
INV     gate2049  (.A(II6371), .Z(g2547) ) ;
INV     gate2050  (.A(g1351), .Z(g2548) ) ;
INV     gate2051  (.A(g1360), .Z(g2551) ) ;
INV     gate2052  (.A(g38), .Z(II6376) ) ;
INV     gate2053  (.A(II6376), .Z(g2554) ) ;
INV     gate2054  (.A(g936), .Z(g2555) ) ;
INV     gate2055  (.A(g1190), .Z(g2556) ) ;
INV     gate2056  (.A(g940), .Z(g2557) ) ;
INV     gate2057  (.A(g1555), .Z(g2561) ) ;
INV     gate2058  (.A(g1652), .Z(g2562) ) ;
INV     gate2059  (.A(g1649), .Z(g2573) ) ;
INV     gate2060  (.A(g1646), .Z(g2584) ) ;
INV     gate2061  (.A(g1643), .Z(g2595) ) ;
INV     gate2062  (.A(g1639), .Z(g2605) ) ;
INV     gate2063  (.A(g1562), .Z(g2614) ) ;
INV     gate2064  (.A(g1563), .Z(g2615) ) ;
INV     gate2065  (.A(g1564), .Z(g2616) ) ;
INV     gate2066  (.A(g1565), .Z(g2617) ) ;
INV     gate2067  (.A(g1566), .Z(g2618) ) ;
INV     gate2068  (.A(g1567), .Z(g2621) ) ;
INV     gate2069  (.A(g1568), .Z(g2622) ) ;
INV     gate2070  (.A(g1585), .Z(g2623) ) ;
INV     gate2071  (.A(g1569), .Z(g2624) ) ;
INV     gate2072  (.A(g1570), .Z(g2625) ) ;
INV     gate2073  (.A(g1571), .Z(g2626) ) ;
INV     gate2074  (.A(g1572), .Z(g2627) ) ;
INV     gate2075  (.A(g1573), .Z(g2628) ) ;
INV     gate2076  (.A(g1574), .Z(g2629) ) ;
INV     gate2077  (.A(g1575), .Z(g2630) ) ;
INV     gate2078  (.A(g1586), .Z(g2631) ) ;
INV     gate2079  (.A(g1576), .Z(g2632) ) ;
INV     gate2080  (.A(g1577), .Z(g2633) ) ;
INV     gate2081  (.A(g1578), .Z(g2634) ) ;
INV     gate2082  (.A(g1579), .Z(g2635) ) ;
INV     gate2083  (.A(g1580), .Z(g2636) ) ;
INV     gate2084  (.A(g1581), .Z(g2637) ) ;
INV     gate2085  (.A(g1582), .Z(g2638) ) ;
INV     gate2086  (.A(g1583), .Z(g2639) ) ;
INV     gate2087  (.A(g1584), .Z(g2640) ) ;
INV     gate2088  (.A(g1587), .Z(g2641) ) ;
INV     gate2089  (.A(g1588), .Z(g2642) ) ;
INV     gate2090  (.A(g1589), .Z(g2643) ) ;
INV     gate2091  (.A(g1794), .Z(II6416) ) ;
INV     gate2092  (.A(g1799), .Z(II6419) ) ;
INV     gate2093  (.A(g1805), .Z(II6422) ) ;
INV     gate2094  (.A(g1811), .Z(II6425) ) ;
INV     gate2095  (.A(g1818), .Z(II6428) ) ;
INV     gate2096  (.A(g1825), .Z(II6431) ) ;
INV     gate2097  (.A(g1830), .Z(II6434) ) ;
INV     gate2098  (.A(g1784), .Z(II6437) ) ;
INV     gate2099  (.A(g1806), .Z(II6440) ) ;
INV     gate2100  (.A(g1774), .Z(II6443) ) ;
INV     gate2101  (.A(g1812), .Z(II6446) ) ;
INV     gate2102  (.A(g1895), .Z(II6451) ) ;
INV     gate2103  (.A(g1868), .Z(II6454) ) ;
INV     gate2104  (.A(g1886), .Z(II6457) ) ;
INV     gate2105  (.A(g2104), .Z(II6460) ) ;
INV     gate2106  (.A(g1769), .Z(II6463) ) ;
INV     gate2107  (.A(g1661), .Z(g2665) ) ;
INV     gate2108  (.A(g1662), .Z(g2668) ) ;
INV     gate2109  (.A(g1917), .Z(II6468) ) ;
INV     gate2110  (.A(g1923), .Z(II6471) ) ;
INV     gate2111  (.A(g1941), .Z(II6474) ) ;
INV     gate2112  (.A(g1675), .Z(g2674) ) ;
INV     gate2113  (.A(g1664), .Z(g2677) ) ;
INV     gate2114  (.A(g1665), .Z(g2680) ) ;
INV     gate2115  (.A(g1666), .Z(g2683) ) ;
INV     gate2116  (.A(g1667), .Z(g2686) ) ;
INV     gate2117  (.A(g1670), .Z(g2689) ) ;
INV     gate2118  (.A(g1671), .Z(g2692) ) ;
INV     gate2119  (.A(g1672), .Z(g2695) ) ;
INV     gate2120  (.A(g1673), .Z(g2698) ) ;
INV     gate2121  (.A(g1674), .Z(g2699) ) ;
INV     gate2122  (.A(g1744), .Z(g2700) ) ;
INV     gate2123  (.A(g1809), .Z(g2703) ) ;
INV     gate2124  (.A(g1821), .Z(g2706) ) ;
INV     gate2125  (.A(g1747), .Z(g2709) ) ;
INV     gate2126  (.A(g2039), .Z(g2712) ) ;
INV     gate2127  (.A(g1803), .Z(g2721) ) ;
INV     gate2128  (.A(g1814), .Z(g2724) ) ;
INV     gate2129  (.A(g2424), .Z(g2727) ) ;
INV     gate2130  (.A(g2256), .Z(g2728) ) ;
INV     gate2131  (.A(g2170), .Z(g2734) ) ;
INV     gate2132  (.A(g1808), .Z(g2743) ) ;
INV     gate2133  (.A(g2259), .Z(g2746) ) ;
INV     gate2134  (.A(g2389), .Z(g2752) ) ;
INV     gate2135  (.A(g1820), .Z(g2761) ) ;
INV     gate2136  (.A(g1802), .Z(g2764) ) ;
INV     gate2137  (.A(g1684), .Z(II6509) ) ;
INV     gate2138  (.A(II6509), .Z(g2767) ) ;
INV     gate2139  (.A(g2424), .Z(g2769) ) ;
INV     gate2140  (.A(g2210), .Z(g2770) ) ;
INV     gate2141  (.A(g1813), .Z(g2774) ) ;
INV     gate2142  (.A(g1797), .Z(g2777) ) ;
INV     gate2143  (.A(g1687), .Z(II6517) ) ;
INV     gate2144  (.A(II6517), .Z(g2780) ) ;
INV     gate2145  (.A(g1616), .Z(g2782) ) ;
INV     gate2146  (.A(g2340), .Z(g2784) ) ;
INV     gate2147  (.A(g1807), .Z(g2787) ) ;
INV     gate2148  (.A(g1793), .Z(g2790) ) ;
INV     gate2149  (.A(g1694), .Z(II6532) ) ;
INV     gate2150  (.A(II6532), .Z(g2793) ) ;
INV     gate2151  (.A(g2185), .Z(g2794) ) ;
INV     gate2152  (.A(g1801), .Z(g2795) ) ;
INV     gate2153  (.A(g1787), .Z(g2798) ) ;
INV     gate2154  (.A(g1796), .Z(g2804) ) ;
INV     gate2155  (.A(g1782), .Z(g2807) ) ;
INV     gate2156  (.A(g1922), .Z(g2810) ) ;
INV     gate2157  (.A(g1685), .Z(g2816) ) ;
INV     gate2158  (.A(g1849), .Z(g2817) ) ;
INV     gate2159  (.A(g1792), .Z(g2818) ) ;
INV     gate2160  (.A(g1786), .Z(g2821) ) ;
INV     gate2161  (.A(g1688), .Z(g2824) ) ;
INV     gate2162  (.A(g2246), .Z(II6553) ) ;
INV     gate2163  (.A(II6553), .Z(g2825) ) ;
INV     gate2164  (.A(g2183), .Z(g2826) ) ;
NOR2    gate2165  (.A(g1430), .B(g1431), .Z(g1980) ) ;
INV     gate2166  (.A(g1980), .Z(g2828) ) ;
INV     gate2167  (.A(g1785), .Z(g2829) ) ;
INV     gate2168  (.A(g2184), .Z(g2832) ) ;
INV     gate2169  (.A(g1715), .Z(II6561) ) ;
INV     gate2170  (.A(II6561), .Z(g2833) ) ;
INV     gate2171  (.A(g2073), .Z(II6564) ) ;
INV     gate2172  (.A(II6564), .Z(g2834) ) ;
INV     gate2173  (.A(g1780), .Z(g2837) ) ;
INV     gate2174  (.A(g2207), .Z(g2840) ) ;
INV     gate2175  (.A(g2208), .Z(g2841) ) ;
INV     gate2176  (.A(g2209), .Z(g2842) ) ;
INV     gate2177  (.A(g1711), .Z(II6571) ) ;
INV     gate2178  (.A(II6571), .Z(g2843) ) ;
INV     gate2179  (.A(g576), .Z(II6574) ) ;
INV     gate2180  (.A(g1603), .Z(II6578) ) ;
INV     gate2181  (.A(II6578), .Z(g2862) ) ;
INV     gate2182  (.A(g1778), .Z(g2863) ) ;
INV     gate2183  (.A(g2221), .Z(g2866) ) ;
INV     gate2184  (.A(g2222), .Z(g2867) ) ;
INV     gate2185  (.A(g2223), .Z(g2868) ) ;
INV     gate2186  (.A(g2224), .Z(g2869) ) ;
INV     gate2187  (.A(g2225), .Z(g2870) ) ;
INV     gate2188  (.A(g1708), .Z(II6587) ) ;
INV     gate2189  (.A(II6587), .Z(g2871) ) ;
INV     gate2190  (.A(g2467), .Z(II6590) ) ;
INV     gate2191  (.A(II6590), .Z(g2872) ) ;
INV     gate2192  (.A(g1779), .Z(g2873) ) ;
INV     gate2193  (.A(g2231), .Z(g2876) ) ;
INV     gate2194  (.A(g2232), .Z(g2877) ) ;
INV     gate2195  (.A(g2233), .Z(g2878) ) ;
INV     gate2196  (.A(g1970), .Z(II6597) ) ;
INV     gate2197  (.A(II6597), .Z(g2879) ) ;
INV     gate2198  (.A(g2234), .Z(g2880) ) ;
INV     gate2199  (.A(g2235), .Z(g2881) ) ;
INV     gate2200  (.A(g2236), .Z(g2882) ) ;
INV     gate2201  (.A(g2237), .Z(g2883) ) ;
INV     gate2202  (.A(g2238), .Z(g2884) ) ;
INV     gate2203  (.A(g2239), .Z(g2885) ) ;
INV     gate2204  (.A(g2240), .Z(g2886) ) ;
INV     gate2205  (.A(g2241), .Z(g2887) ) ;
INV     gate2206  (.A(g1612), .Z(II6608) ) ;
INV     gate2207  (.A(g2264), .Z(g2890) ) ;
INV     gate2208  (.A(g2265), .Z(g2891) ) ;
INV     gate2209  (.A(g2266), .Z(g2892) ) ;
INV     gate2210  (.A(g1983), .Z(II6615) ) ;
INV     gate2211  (.A(II6615), .Z(g2893) ) ;
INV     gate2212  (.A(g2267), .Z(g2894) ) ;
INV     gate2213  (.A(g2268), .Z(g2895) ) ;
INV     gate2214  (.A(g2269), .Z(g2896) ) ;
INV     gate2215  (.A(g2270), .Z(g2897) ) ;
INV     gate2216  (.A(g2271), .Z(g2898) ) ;
INV     gate2217  (.A(g2272), .Z(g2899) ) ;
INV     gate2218  (.A(g2273), .Z(g2900) ) ;
INV     gate2219  (.A(g2284), .Z(g2901) ) ;
INV     gate2220  (.A(g2285), .Z(g2902) ) ;
INV     gate2221  (.A(g2286), .Z(g2903) ) ;
INV     gate2222  (.A(g2287), .Z(g2904) ) ;
INV     gate2223  (.A(g2052), .Z(II6629) ) ;
INV     gate2224  (.A(II6629), .Z(g2905) ) ;
INV     gate2225  (.A(g2288), .Z(g2906) ) ;
INV     gate2226  (.A(g2289), .Z(g2907) ) ;
INV     gate2227  (.A(g2290), .Z(g2908) ) ;
INV     gate2228  (.A(g2291), .Z(g2909) ) ;
INV     gate2229  (.A(g1704), .Z(II6636) ) ;
INV     gate2230  (.A(II6636), .Z(g2910) ) ;
INV     gate2231  (.A(g2292), .Z(g2911) ) ;
INV     gate2232  (.A(g2307), .Z(g2913) ) ;
INV     gate2233  (.A(g2308), .Z(g2914) ) ;
INV     gate2234  (.A(g1970), .Z(II6643) ) ;
INV     gate2235  (.A(II6643), .Z(g2915) ) ;
INV     gate2236  (.A(g2246), .Z(II6646) ) ;
INV     gate2237  (.A(II6646), .Z(g2916) ) ;
INV     gate2238  (.A(g2309), .Z(g2917) ) ;
INV     gate2239  (.A(g2310), .Z(g2918) ) ;
INV     gate2240  (.A(g2311), .Z(g2919) ) ;
INV     gate2241  (.A(g2016), .Z(II6652) ) ;
INV     gate2242  (.A(II6652), .Z(g2920) ) ;
INV     gate2243  (.A(g2312), .Z(g2921) ) ;
INV     gate2244  (.A(g2313), .Z(g2922) ) ;
INV     gate2245  (.A(g1701), .Z(II6657) ) ;
INV     gate2246  (.A(II6657), .Z(g2923) ) ;
INV     gate2247  (.A(g2314), .Z(g2924) ) ;
INV     gate2248  (.A(g2324), .Z(g2925) ) ;
INV     gate2249  (.A(g2325), .Z(g2926) ) ;
INV     gate2250  (.A(g2246), .Z(II6663) ) ;
INV     gate2251  (.A(II6663), .Z(g2927) ) ;
INV     gate2252  (.A(g2326), .Z(g2928) ) ;
INV     gate2253  (.A(g2327), .Z(g2929) ) ;
INV     gate2254  (.A(g2328), .Z(g2930) ) ;
INV     gate2255  (.A(g1698), .Z(II6669) ) ;
INV     gate2256  (.A(II6669), .Z(g2931) ) ;
INV     gate2257  (.A(g2329), .Z(g2932) ) ;
INV     gate2258  (.A(g2246), .Z(II6673) ) ;
INV     gate2259  (.A(II6673), .Z(g2933) ) ;
INV     gate2260  (.A(g1603), .Z(II6676) ) ;
INV     gate2261  (.A(II6676), .Z(g2934) ) ;
INV     gate2262  (.A(g1558), .Z(II6680) ) ;
INV     gate2263  (.A(II6680), .Z(g2936) ) ;
INV     gate2264  (.A(g2346), .Z(g2937) ) ;
INV     gate2265  (.A(g2347), .Z(g2938) ) ;
INV     gate2266  (.A(g2348), .Z(g2939) ) ;
INV     gate2267  (.A(g2246), .Z(II6686) ) ;
INV     gate2268  (.A(II6686), .Z(g2940) ) ;
INV     gate2269  (.A(g2349), .Z(g2941) ) ;
INV     gate2270  (.A(g2350), .Z(g2942) ) ;
INV     gate2271  (.A(g2362), .Z(g2943) ) ;
INV     gate2272  (.A(g2363), .Z(g2944) ) ;
INV     gate2273  (.A(g2364), .Z(g2945) ) ;
INV     gate2274  (.A(g2365), .Z(g2946) ) ;
INV     gate2275  (.A(g2246), .Z(II6695) ) ;
INV     gate2276  (.A(II6695), .Z(g2947) ) ;
INV     gate2277  (.A(g2366), .Z(g2948) ) ;
INV     gate2278  (.A(g2373), .Z(g2953) ) ;
INV     gate2279  (.A(g2374), .Z(g2954) ) ;
INV     gate2280  (.A(g1983), .Z(II6703) ) ;
INV     gate2281  (.A(II6703), .Z(g2955) ) ;
INV     gate2282  (.A(g2375), .Z(g2956) ) ;
INV     gate2283  (.A(g2376), .Z(g2957) ) ;
INV     gate2284  (.A(g2377), .Z(g2958) ) ;
INV     gate2285  (.A(g1926), .Z(g2959) ) ;
INV     gate2286  (.A(g2381), .Z(g2960) ) ;
INV     gate2287  (.A(g1726), .Z(II6711) ) ;
INV     gate2288  (.A(II6711), .Z(g2961) ) ;
INV     gate2289  (.A(g2382), .Z(g2962) ) ;
INV     gate2290  (.A(g2383), .Z(g2963) ) ;
INV     gate2291  (.A(g1721), .Z(II6716) ) ;
INV     gate2292  (.A(II6716), .Z(g2964) ) ;
INV     gate2293  (.A(g2384), .Z(g2965) ) ;
INV     gate2294  (.A(g1856), .Z(g2966) ) ;
INV     gate2295  (.A(g2393), .Z(g2969) ) ;
INV     gate2296  (.A(g2394), .Z(g2970) ) ;
INV     gate2297  (.A(g2052), .Z(II6723) ) ;
INV     gate2298  (.A(II6723), .Z(g2971) ) ;
INV     gate2299  (.A(g1854), .Z(g2973) ) ;
INV     gate2300  (.A(g1959), .Z(II6728) ) ;
INV     gate2301  (.A(II6728), .Z(g2976) ) ;
INV     gate2302  (.A(g1848), .Z(g2982) ) ;
INV     gate2303  (.A(g1718), .Z(II6733) ) ;
INV     gate2304  (.A(II6733), .Z(g2985) ) ;
INV     gate2305  (.A(g1843), .Z(g2989) ) ;
INV     gate2306  (.A(g1833), .Z(g2992) ) ;
INV     gate2307  (.A(g1828), .Z(g2996) ) ;
INV     gate2308  (.A(g1823), .Z(g2999) ) ;
INV     gate2309  (.A(g1816), .Z(g3008) ) ;
OR2     gate2310  (.A(g1189), .B(g16), .Z(g1955) ) ;
INV     gate2311  (.A(g1955), .Z(II6764) ) ;
INV     gate2312  (.A(II6764), .Z(g3013) ) ;
INV     gate2313  (.A(g1933), .Z(II6767) ) ;
INV     gate2314  (.A(II6767), .Z(g3014) ) ;
INV     gate2315  (.A(g1590), .Z(II6770) ) ;
INV     gate2316  (.A(II6770), .Z(g3018) ) ;
INV     gate2317  (.A(g2007), .Z(g3019) ) ;
INV     gate2318  (.A(g1929), .Z(g3029) ) ;
INV     gate2319  (.A(g2092), .Z(g3038) ) ;
INV     gate2320  (.A(g1736), .Z(g3047) ) ;
INV     gate2321  (.A(g2052), .Z(II6784) ) ;
INV     gate2322  (.A(II6784), .Z(g3048) ) ;
INV     gate2323  (.A(g1681), .Z(II6788) ) ;
INV     gate2324  (.A(II6788), .Z(g3050) ) ;
INV     gate2325  (.A(g1967), .Z(II6791) ) ;
INV     gate2326  (.A(II6791), .Z(g3051) ) ;
INV     gate2327  (.A(g2096), .Z(g3052) ) ;
INV     gate2328  (.A(g1683), .Z(II6795) ) ;
INV     gate2329  (.A(II6795), .Z(g3061) ) ;
INV     gate2330  (.A(g2100), .Z(g3062) ) ;
INV     gate2331  (.A(g1948), .Z(g3071) ) ;
INV     gate2332  (.A(g2016), .Z(II6800) ) ;
INV     gate2333  (.A(II6800), .Z(g3074) ) ;
INV     gate2334  (.A(g2216), .Z(g3075) ) ;
INV     gate2335  (.A(g1831), .Z(g3076) ) ;
INV     gate2336  (.A(g1603), .Z(II6805) ) ;
INV     gate2337  (.A(g1603), .Z(g3078) ) ;
INV     gate2338  (.A(g1603), .Z(g3079) ) ;
INV     gate2339  (.A(g1679), .Z(g3080) ) ;
INV     gate2340  (.A(g1680), .Z(g3082) ) ;
INV     gate2341  (.A(g1707), .Z(II6820) ) ;
INV     gate2342  (.A(II6820), .Z(g3084) ) ;
INV     gate2343  (.A(g1945), .Z(g3085) ) ;
INV     gate2344  (.A(g1852), .Z(g3086) ) ;
INV     gate2345  (.A(g1603), .Z(g3091) ) ;
INV     gate2346  (.A(g2185), .Z(II6826) ) ;
INV     gate2347  (.A(II6826), .Z(g3092) ) ;
INV     gate2348  (.A(g1686), .Z(g3093) ) ;
INV     gate2349  (.A(g2185), .Z(II6831) ) ;
INV     gate2350  (.A(II6831), .Z(g3095) ) ;
INV     gate2351  (.A(g287), .Z(II6834) ) ;
INV     gate2352  (.A(g1857), .Z(g3124) ) ;
INV     gate2353  (.A(g2185), .Z(II6839) ) ;
INV     gate2354  (.A(II6839), .Z(g3128) ) ;
INV     gate2355  (.A(g368), .Z(II6849) ) ;
INV     gate2356  (.A(g2185), .Z(II6853) ) ;
INV     gate2357  (.A(II6853), .Z(g3158) ) ;
INV     gate2358  (.A(g449), .Z(II6856) ) ;
INV     gate2359  (.A(g2185), .Z(II6860) ) ;
INV     gate2360  (.A(II6860), .Z(g3187) ) ;
INV     gate2361  (.A(g2528), .Z(II6864) ) ;
INV     gate2362  (.A(II6864), .Z(g3189) ) ;
INV     gate2363  (.A(g530), .Z(II6868) ) ;
INV     gate2364  (.A(g2185), .Z(II6872) ) ;
INV     gate2365  (.A(II6872), .Z(g3219) ) ;
INV     gate2366  (.A(g1889), .Z(g3220) ) ;
INV     gate2367  (.A(g2528), .Z(II6887) ) ;
INV     gate2368  (.A(II6887), .Z(g3230) ) ;
INV     gate2369  (.A(g1863), .Z(II6894) ) ;
INV     gate2370  (.A(II6894), .Z(g3238) ) ;
INV     gate2371  (.A(g1866), .Z(II6900) ) ;
INV     gate2372  (.A(II6900), .Z(g3264) ) ;
INV     gate2373  (.A(g1689), .Z(g3285) ) ;
INV     gate2374  (.A(g1869), .Z(II6911) ) ;
INV     gate2375  (.A(II6911), .Z(g3287) ) ;
INV     gate2376  (.A(g1876), .Z(II6930) ) ;
INV     gate2377  (.A(II6930), .Z(g3316) ) ;
INV     gate2378  (.A(g1901), .Z(g3338) ) ;
NAND2   gate2379  (.A(g1405), .B(g1412), .Z(g2474) ) ;
INV     gate2380  (.A(g2474), .Z(g3340) ) ;
INV     gate2381  (.A(g1878), .Z(II6936) ) ;
INV     gate2382  (.A(II6936), .Z(g3341) ) ;
INV     gate2383  (.A(g1887), .Z(II6946) ) ;
INV     gate2384  (.A(II6946), .Z(g3359) ) ;
INV     gate2385  (.A(g2148), .Z(II6949) ) ;
INV     gate2386  (.A(II6949), .Z(g3390) ) ;
INV     gate2387  (.A(g1896), .Z(II6952) ) ;
INV     gate2388  (.A(II6952), .Z(g3398) ) ;
INV     gate2389  (.A(g1907), .Z(II6956) ) ;
INV     gate2390  (.A(II6956), .Z(g3430) ) ;
INV     gate2391  (.A(g1558), .Z(II6959) ) ;
INV     gate2392  (.A(II6959), .Z(g3461) ) ;
INV     gate2393  (.A(g1743), .Z(g3462) ) ;
INV     gate2394  (.A(g1558), .Z(II6963) ) ;
INV     gate2395  (.A(II6963), .Z(g3465) ) ;
INV     gate2396  (.A(g1737), .Z(g3485) ) ;
INV     gate2397  (.A(g1727), .Z(g3488) ) ;
INV     gate2398  (.A(g1800), .Z(g3491) ) ;
OR4     gate2399  (.A(g971), .B(g962), .C(g972), .D(II5757), .Z(g1872) ) ;
INV     gate2400  (.A(g1872), .Z(II6970) ) ;
INV     gate2401  (.A(II6970), .Z(g3492) ) ;
INV     gate2402  (.A(g1616), .Z(g3495) ) ;
INV     gate2403  (.A(g2528), .Z(II6974) ) ;
INV     gate2404  (.A(II6974), .Z(g3496) ) ;
INV     gate2405  (.A(g2185), .Z(g3497) ) ;
INV     gate2406  (.A(g1616), .Z(g3498) ) ;
INV     gate2407  (.A(g2185), .Z(g3499) ) ;
INV     gate2408  (.A(g1616), .Z(g3500) ) ;
INV     gate2409  (.A(g2185), .Z(g3501) ) ;
INV     gate2410  (.A(g1616), .Z(g3502) ) ;
INV     gate2411  (.A(g2407), .Z(g3503) ) ;
INV     gate2412  (.A(g1781), .Z(g3506) ) ;
INV     gate2413  (.A(g2185), .Z(g3510) ) ;
INV     gate2414  (.A(g1616), .Z(g3511) ) ;
INV     gate2415  (.A(g1616), .Z(g3512) ) ;
INV     gate2416  (.A(g2407), .Z(g3513) ) ;
INV     gate2417  (.A(g2424), .Z(g3514) ) ;
INV     gate2418  (.A(g2283), .Z(g3517) ) ;
INV     gate2419  (.A(g2185), .Z(g3519) ) ;
INV     gate2420  (.A(g1616), .Z(g3520) ) ;
INV     gate2421  (.A(g2185), .Z(g3521) ) ;
INV     gate2422  (.A(g2407), .Z(g3522) ) ;
INV     gate2423  (.A(g2407), .Z(g3523) ) ;
INV     gate2424  (.A(g2306), .Z(g3524) ) ;
INV     gate2425  (.A(g2185), .Z(g3526) ) ;
INV     gate2426  (.A(g1616), .Z(g3527) ) ;
INV     gate2427  (.A(g2323), .Z(g3529) ) ;
INV     gate2428  (.A(g2185), .Z(g3530) ) ;
INV     gate2429  (.A(g1616), .Z(g3531) ) ;
INV     gate2430  (.A(g2407), .Z(g3532) ) ;
INV     gate2431  (.A(g2397), .Z(g3533) ) ;
INV     gate2432  (.A(g2424), .Z(g3539) ) ;
INV     gate2433  (.A(g2424), .Z(g3540) ) ;
INV     gate2434  (.A(g1777), .Z(g3542) ) ;
INV     gate2435  (.A(g2344), .Z(g3545) ) ;
INV     gate2436  (.A(g2392), .Z(II7029) ) ;
INV     gate2437  (.A(II7029), .Z(g3546) ) ;
INV     gate2438  (.A(g2345), .Z(g3547) ) ;
INV     gate2439  (.A(g2185), .Z(g3548) ) ;
INV     gate2440  (.A(g2404), .Z(g3549) ) ;
INV     gate2441  (.A(g2454), .Z(II7036) ) ;
INV     gate2442  (.A(II7036), .Z(g3556) ) ;
INV     gate2443  (.A(g1773), .Z(g3557) ) ;
INV     gate2444  (.A(g2361), .Z(g3560) ) ;
INV     gate2445  (.A(g2401), .Z(II7041) ) ;
INV     gate2446  (.A(II7041), .Z(g3561) ) ;
INV     gate2447  (.A(g2402), .Z(II7044) ) ;
INV     gate2448  (.A(II7044), .Z(g3562) ) ;
INV     gate2449  (.A(g2007), .Z(g3563) ) ;
INV     gate2450  (.A(g2407), .Z(g3567) ) ;
INV     gate2451  (.A(g1935), .Z(g3568) ) ;
INV     gate2452  (.A(g2424), .Z(g3573) ) ;
INV     gate2453  (.A(g1771), .Z(g3574) ) ;
INV     gate2454  (.A(g2372), .Z(g3577) ) ;
INV     gate2455  (.A(g2452), .Z(II7053) ) ;
INV     gate2456  (.A(II7053), .Z(g3578) ) ;
INV     gate2457  (.A(g1929), .Z(g3579) ) ;
INV     gate2458  (.A(g2407), .Z(g3582) ) ;
INV     gate2459  (.A(g2128), .Z(g3583) ) ;
NOR2    gate2460  (.A(g1428), .B(g1429), .Z(g1964) ) ;
INV     gate2461  (.A(g1964), .Z(g3587) ) ;
INV     gate2462  (.A(g2379), .Z(g3588) ) ;
INV     gate2463  (.A(g2457), .Z(II7061) ) ;
INV     gate2464  (.A(II7061), .Z(g3589) ) ;
INV     gate2465  (.A(g2458), .Z(II7064) ) ;
INV     gate2466  (.A(II7064), .Z(g3590) ) ;
INV     gate2467  (.A(g1789), .Z(g3591) ) ;
INV     gate2468  (.A(g2092), .Z(g3603) ) ;
INV     gate2469  (.A(g2407), .Z(g3604) ) ;
INV     gate2470  (.A(g1938), .Z(g3605) ) ;
INV     gate2471  (.A(g2424), .Z(g3610) ) ;
INV     gate2472  (.A(g2532), .Z(II7079) ) ;
INV     gate2473  (.A(II7079), .Z(g3611) ) ;
INV     gate2474  (.A(g2470), .Z(II7082) ) ;
INV     gate2475  (.A(II7082), .Z(g3612) ) ;
INV     gate2476  (.A(g1655), .Z(g3617) ) ;
INV     gate2477  (.A(g2424), .Z(g3629) ) ;
INV     gate2478  (.A(g2539), .Z(II7095) ) ;
INV     gate2479  (.A(II7095), .Z(g3630) ) ;
INV     gate2480  (.A(g2477), .Z(II7098) ) ;
INV     gate2481  (.A(II7098), .Z(g3631) ) ;
INV     gate2482  (.A(g2478), .Z(II7101) ) ;
INV     gate2483  (.A(II7101), .Z(g3632) ) ;
INV     gate2484  (.A(g2479), .Z(II7104) ) ;
INV     gate2485  (.A(II7104), .Z(g3633) ) ;
INV     gate2486  (.A(g2480), .Z(II7107) ) ;
INV     gate2487  (.A(II7107), .Z(g3634) ) ;
INV     gate2488  (.A(g1949), .Z(g3635) ) ;
INV     gate2489  (.A(g2424), .Z(g3639) ) ;
INV     gate2490  (.A(g2546), .Z(II7112) ) ;
INV     gate2491  (.A(II7112), .Z(g3640) ) ;
INV     gate2492  (.A(g2547), .Z(II7115) ) ;
INV     gate2493  (.A(II7115), .Z(g3641) ) ;
INV     gate2494  (.A(g2484), .Z(II7118) ) ;
INV     gate2495  (.A(II7118), .Z(g3642) ) ;
INV     gate2496  (.A(g2453), .Z(g3643) ) ;
INV     gate2497  (.A(g2131), .Z(g3644) ) ;
INV     gate2498  (.A(g2424), .Z(g3647) ) ;
INV     gate2499  (.A(g2424), .Z(g3648) ) ;
INV     gate2500  (.A(g2424), .Z(g3649) ) ;
INV     gate2501  (.A(g2494), .Z(II7126) ) ;
INV     gate2502  (.A(II7126), .Z(g3650) ) ;
INV     gate2503  (.A(g2495), .Z(II7129) ) ;
INV     gate2504  (.A(II7129), .Z(g3651) ) ;
INV     gate2505  (.A(g2554), .Z(II7132) ) ;
INV     gate2506  (.A(II7132), .Z(g3652) ) ;
INV     gate2507  (.A(g2459), .Z(g3653) ) ;
NOR2    gate2508  (.A(g65), .B(g62), .Z(g2521) ) ;
INV     gate2509  (.A(g2521), .Z(g3654) ) ;
AND2    gate2510  (.A(g792), .B(g795), .Z(g1844) ) ;
INV     gate2511  (.A(g1844), .Z(g3655) ) ;
INV     gate2512  (.A(g2501), .Z(II7145) ) ;
INV     gate2513  (.A(II7145), .Z(g3657) ) ;
INV     gate2514  (.A(g2293), .Z(g3659) ) ;
INV     gate2515  (.A(g2134), .Z(g3666) ) ;
INV     gate2516  (.A(g2157), .Z(II7164) ) ;
INV     gate2517  (.A(II7164), .Z(g3674) ) ;
INV     gate2518  (.A(g2505), .Z(II7167) ) ;
INV     gate2519  (.A(II7167), .Z(g3675) ) ;
INV     gate2520  (.A(g2380), .Z(g3676) ) ;
INV     gate2521  (.A(g2485), .Z(g3677) ) ;
INV     gate2522  (.A(g2180), .Z(g3684) ) ;
INV     gate2523  (.A(g1795), .Z(II7195) ) ;
INV     gate2524  (.A(II7195), .Z(g3691) ) ;
INV     gate2525  (.A(g2509), .Z(II7198) ) ;
INV     gate2526  (.A(II7198), .Z(g3692) ) ;
INV     gate2527  (.A(g2424), .Z(g3693) ) ;
INV     gate2528  (.A(g2174), .Z(g3694) ) ;
INV     gate2529  (.A(g2514), .Z(g3700) ) ;
INV     gate2530  (.A(g2520), .Z(II7204) ) ;
INV     gate2531  (.A(II7204), .Z(g3705) ) ;
INV     gate2532  (.A(g2226), .Z(g3707) ) ;
INV     gate2533  (.A(g1952), .Z(g3712) ) ;
INV     gate2534  (.A(g2522), .Z(g3716) ) ;
INV     gate2535  (.A(g1742), .Z(II7211) ) ;
INV     gate2536  (.A(II7211), .Z(g3721) ) ;
INV     gate2537  (.A(g2096), .Z(g3723) ) ;
INV     gate2538  (.A(g2202), .Z(g3728) ) ;
INV     gate2539  (.A(g2533), .Z(g3732) ) ;
INV     gate2540  (.A(g1961), .Z(g3735) ) ;
INV     gate2541  (.A(g2536), .Z(g3739) ) ;
INV     gate2542  (.A(g1776), .Z(g3743) ) ;
INV     gate2543  (.A(g2100), .Z(g3746) ) ;
INV     gate2544  (.A(g2177), .Z(g3750) ) ;
INV     gate2545  (.A(g2540), .Z(g3753) ) ;
INV     gate2546  (.A(g2543), .Z(g3754) ) ;
INV     gate2547  (.A(g1977), .Z(g3757) ) ;
INV     gate2548  (.A(g1772), .Z(g3761) ) ;
INV     gate2549  (.A(g2039), .Z(g3764) ) ;
INV     gate2550  (.A(g2253), .Z(g3768) ) ;
INV     gate2551  (.A(g2548), .Z(g3769) ) ;
INV     gate2552  (.A(g2551), .Z(g3770) ) ;
INV     gate2553  (.A(g1853), .Z(g3771) ) ;
INV     gate2554  (.A(g1770), .Z(g3774) ) ;
INV     gate2555  (.A(g2170), .Z(g3777) ) ;
INV     gate2556  (.A(g2145), .Z(g3778) ) ;
INV     gate2557  (.A(g2511), .Z(g3779) ) ;
INV     gate2558  (.A(g1847), .Z(g3780) ) ;
INV     gate2559  (.A(g1955), .Z(II7255) ) ;
INV     gate2560  (.A(II7255), .Z(g3783) ) ;
INV     gate2561  (.A(g1768), .Z(g3784) ) ;
INV     gate2562  (.A(g1842), .Z(g3787) ) ;
INV     gate2563  (.A(g1757), .Z(g3798) ) ;
INV     gate2564  (.A(g2514), .Z(II7262) ) ;
INV     gate2565  (.A(II7262), .Z(g3801) ) ;
INV     gate2566  (.A(g1832), .Z(g3802) ) ;
INV     gate2567  (.A(g1752), .Z(g3805) ) ;
INV     gate2568  (.A(g1827), .Z(g3808) ) ;
INV     gate2569  (.A(g1750), .Z(g3812) ) ;
INV     gate2570  (.A(g1822), .Z(g3815) ) ;
INV     gate2571  (.A(g1748), .Z(g3819) ) ;
INV     gate2572  (.A(g1815), .Z(g3822) ) ;
INV     gate2573  (.A(g1826), .Z(g3825) ) ;
INV     gate2574  (.A(g2561), .Z(II7287) ) ;
INV     gate2575  (.A(II7287), .Z(g3828) ) ;
INV     gate2576  (.A(g2936), .Z(II7290) ) ;
INV     gate2577  (.A(g2955), .Z(II7293) ) ;
INV     gate2578  (.A(g2915), .Z(II7296) ) ;
INV     gate2579  (.A(g2961), .Z(II7299) ) ;
INV     gate2580  (.A(g2825), .Z(II7302) ) ;
INV     gate2581  (.A(g3048), .Z(II7305) ) ;
INV     gate2582  (.A(g3074), .Z(II7308) ) ;
INV     gate2583  (.A(g2879), .Z(II7311) ) ;
INV     gate2584  (.A(g2916), .Z(II7314) ) ;
INV     gate2585  (.A(g2893), .Z(II7317) ) ;
INV     gate2586  (.A(g2927), .Z(II7320) ) ;
INV     gate2587  (.A(g2905), .Z(II7323) ) ;
INV     gate2588  (.A(g2940), .Z(II7326) ) ;
INV     gate2589  (.A(g2920), .Z(II7329) ) ;
INV     gate2590  (.A(g2947), .Z(II7332) ) ;
INV     gate2591  (.A(g2910), .Z(II7335) ) ;
INV     gate2592  (.A(g2923), .Z(II7338) ) ;
INV     gate2593  (.A(g2931), .Z(II7341) ) ;
INV     gate2594  (.A(g2964), .Z(II7344) ) ;
INV     gate2595  (.A(g2985), .Z(II7347) ) ;
INV     gate2596  (.A(g2971), .Z(II7350) ) ;
INV     gate2597  (.A(g2833), .Z(II7353) ) ;
INV     gate2598  (.A(g2843), .Z(II7356) ) ;
INV     gate2599  (.A(g2871), .Z(II7359) ) ;
INV     gate2600  (.A(g2933), .Z(II7362) ) ;
INV     gate2601  (.A(g3061), .Z(II7365) ) ;
INV     gate2602  (.A(g3018), .Z(II7368) ) ;
INV     gate2603  (.A(g3050), .Z(II7371) ) ;
INV     gate2604  (.A(g3084), .Z(II7374) ) ;
INV     gate2605  (.A(g3189), .Z(II7377) ) ;
INV     gate2606  (.A(g3461), .Z(II7380) ) ;
INV     gate2607  (.A(g3465), .Z(II7383) ) ;
INV     gate2608  (.A(g3013), .Z(II7386) ) ;
INV     gate2609  (.A(g3496), .Z(II7389) ) ;
INV     gate2610  (.A(g3230), .Z(II7392) ) ;
INV     gate2611  (.A(g2943), .Z(g3864) ) ;
INV     gate2612  (.A(g2944), .Z(g3865) ) ;
INV     gate2613  (.A(g2945), .Z(g3866) ) ;
INV     gate2614  (.A(g2946), .Z(g3867) ) ;
INV     gate2615  (.A(g2948), .Z(g3868) ) ;
INV     gate2616  (.A(g3075), .Z(II7400) ) ;
INV     gate2617  (.A(II7400), .Z(g3869) ) ;
AND2    gate2618  (.A(g936), .B(g2557), .Z(g3466) ) ;
INV     gate2619  (.A(g3466), .Z(g3870) ) ;
INV     gate2620  (.A(g2953), .Z(g3871) ) ;
INV     gate2621  (.A(g2954), .Z(g3872) ) ;
INV     gate2622  (.A(g2956), .Z(g3873) ) ;
INV     gate2623  (.A(g2957), .Z(g3874) ) ;
INV     gate2624  (.A(g2958), .Z(g3875) ) ;
INV     gate2625  (.A(g3466), .Z(g3876) ) ;
INV     gate2626  (.A(g2960), .Z(g3877) ) ;
INV     gate2627  (.A(g2962), .Z(g3878) ) ;
INV     gate2628  (.A(g2963), .Z(g3879) ) ;
INV     gate2629  (.A(g2965), .Z(g3880) ) ;
INV     gate2630  (.A(g2969), .Z(g3881) ) ;
INV     gate2631  (.A(g2970), .Z(g3882) ) ;
INV     gate2632  (.A(g3659), .Z(II7417) ) ;
INV     gate2633  (.A(II7417), .Z(g3884) ) ;
OR2     gate2634  (.A(g1746), .B(g287), .Z(g3097) ) ;
INV     gate2635  (.A(g3097), .Z(g3888) ) ;
INV     gate2636  (.A(g3097), .Z(g3891) ) ;
OR2     gate2637  (.A(g1749), .B(g368), .Z(g3131) ) ;
INV     gate2638  (.A(g3131), .Z(g3892) ) ;
INV     gate2639  (.A(g3546), .Z(II7473) ) ;
INV     gate2640  (.A(II7473), .Z(g3896) ) ;
INV     gate2641  (.A(g3131), .Z(g3897) ) ;
OR2     gate2642  (.A(g1751), .B(g449), .Z(g3160) ) ;
INV     gate2643  (.A(g3160), .Z(g3898) ) ;
INV     gate2644  (.A(g3561), .Z(II7492) ) ;
INV     gate2645  (.A(II7492), .Z(g3901) ) ;
INV     gate2646  (.A(g3562), .Z(II7495) ) ;
INV     gate2647  (.A(II7495), .Z(g3902) ) ;
INV     gate2648  (.A(g2752), .Z(II7498) ) ;
INV     gate2649  (.A(II7498), .Z(g3903) ) ;
INV     gate2650  (.A(g3160), .Z(g3904) ) ;
OR2     gate2651  (.A(g1756), .B(g530), .Z(g3192) ) ;
INV     gate2652  (.A(g3192), .Z(g3905) ) ;
INV     gate2653  (.A(g3578), .Z(II7517) ) ;
INV     gate2654  (.A(II7517), .Z(g3908) ) ;
INV     gate2655  (.A(g2734), .Z(II7520) ) ;
INV     gate2656  (.A(II7520), .Z(g3909) ) ;
INV     gate2657  (.A(g2562), .Z(II7523) ) ;
INV     gate2658  (.A(II7523), .Z(g3910) ) ;
INV     gate2659  (.A(g2752), .Z(II7526) ) ;
INV     gate2660  (.A(II7526), .Z(g3911) ) ;
INV     gate2661  (.A(g3192), .Z(g3912) ) ;
INV     gate2662  (.A(g2834), .Z(g3913) ) ;
INV     gate2663  (.A(g3589), .Z(II7545) ) ;
INV     gate2664  (.A(II7545), .Z(g3916) ) ;
INV     gate2665  (.A(g3590), .Z(II7548) ) ;
INV     gate2666  (.A(II7548), .Z(g3917) ) ;
INV     gate2667  (.A(g2712), .Z(II7551) ) ;
INV     gate2668  (.A(II7551), .Z(g3918) ) ;
INV     gate2669  (.A(g2573), .Z(II7554) ) ;
INV     gate2670  (.A(II7554), .Z(g3919) ) ;
INV     gate2671  (.A(g3097), .Z(g3920) ) ;
INV     gate2672  (.A(g2734), .Z(II7558) ) ;
INV     gate2673  (.A(II7558), .Z(g3921) ) ;
INV     gate2674  (.A(g2562), .Z(II7561) ) ;
INV     gate2675  (.A(II7561), .Z(g3922) ) ;
INV     gate2676  (.A(g2752), .Z(II7564) ) ;
INV     gate2677  (.A(II7564), .Z(g3923) ) ;
INV     gate2678  (.A(g3612), .Z(II7581) ) ;
INV     gate2679  (.A(II7581), .Z(g3926) ) ;
INV     gate2680  (.A(g3062), .Z(II7584) ) ;
INV     gate2681  (.A(II7584), .Z(g3927) ) ;
INV     gate2682  (.A(g3097), .Z(g3928) ) ;
INV     gate2683  (.A(g2584), .Z(II7588) ) ;
INV     gate2684  (.A(II7588), .Z(g3929) ) ;
INV     gate2685  (.A(g3097), .Z(g3930) ) ;
INV     gate2686  (.A(g2712), .Z(II7592) ) ;
INV     gate2687  (.A(II7592), .Z(g3931) ) ;
INV     gate2688  (.A(g2573), .Z(II7595) ) ;
INV     gate2689  (.A(II7595), .Z(g3932) ) ;
INV     gate2690  (.A(g3131), .Z(g3933) ) ;
INV     gate2691  (.A(g2734), .Z(II7599) ) ;
INV     gate2692  (.A(II7599), .Z(g3934) ) ;
INV     gate2693  (.A(g2562), .Z(II7602) ) ;
INV     gate2694  (.A(II7602), .Z(g3935) ) ;
INV     gate2695  (.A(g2752), .Z(II7605) ) ;
INV     gate2696  (.A(II7605), .Z(g3936) ) ;
OR2     gate2697  (.A(g1877), .B(g576), .Z(g2845) ) ;
INV     gate2698  (.A(g2845), .Z(g3937) ) ;
INV     gate2699  (.A(g3631), .Z(II7623) ) ;
INV     gate2700  (.A(II7623), .Z(g3940) ) ;
INV     gate2701  (.A(g3632), .Z(II7626) ) ;
INV     gate2702  (.A(II7626), .Z(g3941) ) ;
INV     gate2703  (.A(g3633), .Z(II7629) ) ;
INV     gate2704  (.A(II7629), .Z(g3942) ) ;
INV     gate2705  (.A(g3634), .Z(II7632) ) ;
INV     gate2706  (.A(II7632), .Z(g3943) ) ;
INV     gate2707  (.A(g3052), .Z(II7635) ) ;
INV     gate2708  (.A(II7635), .Z(g3944) ) ;
INV     gate2709  (.A(g3097), .Z(g3945) ) ;
INV     gate2710  (.A(g3097), .Z(g3946) ) ;
INV     gate2711  (.A(g3062), .Z(II7640) ) ;
INV     gate2712  (.A(II7640), .Z(g3947) ) ;
INV     gate2713  (.A(g3131), .Z(g3948) ) ;
INV     gate2714  (.A(g2584), .Z(II7644) ) ;
INV     gate2715  (.A(II7644), .Z(g3949) ) ;
INV     gate2716  (.A(g3131), .Z(g3950) ) ;
INV     gate2717  (.A(g2712), .Z(II7648) ) ;
INV     gate2718  (.A(II7648), .Z(g3951) ) ;
INV     gate2719  (.A(g2573), .Z(II7651) ) ;
INV     gate2720  (.A(II7651), .Z(g3952) ) ;
INV     gate2721  (.A(g3160), .Z(g3953) ) ;
INV     gate2722  (.A(g2734), .Z(II7655) ) ;
INV     gate2723  (.A(II7655), .Z(g3954) ) ;
INV     gate2724  (.A(g2562), .Z(II7658) ) ;
INV     gate2725  (.A(II7658), .Z(g3955) ) ;
INV     gate2726  (.A(g2845), .Z(g3956) ) ;
INV     gate2727  (.A(g3642), .Z(II7662) ) ;
INV     gate2728  (.A(II7662), .Z(g3957) ) ;
INV     gate2729  (.A(g3097), .Z(g3958) ) ;
INV     gate2730  (.A(g3097), .Z(g3959) ) ;
INV     gate2731  (.A(g3052), .Z(II7667) ) ;
INV     gate2732  (.A(II7667), .Z(g3960) ) ;
INV     gate2733  (.A(g3131), .Z(g3961) ) ;
INV     gate2734  (.A(g3131), .Z(g3962) ) ;
INV     gate2735  (.A(g3062), .Z(II7672) ) ;
INV     gate2736  (.A(II7672), .Z(g3963) ) ;
INV     gate2737  (.A(g3160), .Z(g3964) ) ;
INV     gate2738  (.A(g2584), .Z(II7676) ) ;
INV     gate2739  (.A(II7676), .Z(g3965) ) ;
INV     gate2740  (.A(g3160), .Z(g3966) ) ;
INV     gate2741  (.A(g2712), .Z(II7680) ) ;
INV     gate2742  (.A(II7680), .Z(g3967) ) ;
INV     gate2743  (.A(g2573), .Z(II7683) ) ;
INV     gate2744  (.A(II7683), .Z(g3968) ) ;
INV     gate2745  (.A(g3192), .Z(g3969) ) ;
INV     gate2746  (.A(g2845), .Z(g3970) ) ;
INV     gate2747  (.A(g3650), .Z(II7688) ) ;
INV     gate2748  (.A(II7688), .Z(g3971) ) ;
INV     gate2749  (.A(g3651), .Z(II7691) ) ;
INV     gate2750  (.A(II7691), .Z(g3972) ) ;
INV     gate2751  (.A(g3097), .Z(g3973) ) ;
INV     gate2752  (.A(g3131), .Z(g3974) ) ;
INV     gate2753  (.A(g3131), .Z(g3975) ) ;
INV     gate2754  (.A(g3052), .Z(II7697) ) ;
INV     gate2755  (.A(II7697), .Z(g3976) ) ;
INV     gate2756  (.A(g3160), .Z(g3977) ) ;
INV     gate2757  (.A(g3160), .Z(g3978) ) ;
INV     gate2758  (.A(g3062), .Z(II7702) ) ;
INV     gate2759  (.A(II7702), .Z(g3979) ) ;
INV     gate2760  (.A(g3192), .Z(g3980) ) ;
INV     gate2761  (.A(g2584), .Z(II7706) ) ;
INV     gate2762  (.A(II7706), .Z(g3981) ) ;
INV     gate2763  (.A(g3192), .Z(g3982) ) ;
INV     gate2764  (.A(g2845), .Z(g3983) ) ;
INV     gate2765  (.A(g3657), .Z(II7712) ) ;
INV     gate2766  (.A(II7712), .Z(g3985) ) ;
INV     gate2767  (.A(g3038), .Z(II7716) ) ;
INV     gate2768  (.A(II7716), .Z(g3987) ) ;
INV     gate2769  (.A(g3097), .Z(g3988) ) ;
INV     gate2770  (.A(g3131), .Z(g3989) ) ;
INV     gate2771  (.A(g3160), .Z(g3990) ) ;
INV     gate2772  (.A(g3160), .Z(g3991) ) ;
INV     gate2773  (.A(g3052), .Z(II7723) ) ;
INV     gate2774  (.A(II7723), .Z(g3992) ) ;
INV     gate2775  (.A(g3192), .Z(g3993) ) ;
INV     gate2776  (.A(g3192), .Z(g3994) ) ;
INV     gate2777  (.A(g3675), .Z(II7728) ) ;
INV     gate2778  (.A(II7728), .Z(g3995) ) ;
INV     gate2779  (.A(g3029), .Z(II7731) ) ;
INV     gate2780  (.A(II7731), .Z(g3996) ) ;
INV     gate2781  (.A(g2595), .Z(II7734) ) ;
INV     gate2782  (.A(II7734), .Z(g3997) ) ;
INV     gate2783  (.A(g3097), .Z(g3998) ) ;
INV     gate2784  (.A(g3038), .Z(II7738) ) ;
INV     gate2785  (.A(II7738), .Z(g3999) ) ;
INV     gate2786  (.A(g3131), .Z(g4000) ) ;
INV     gate2787  (.A(g3160), .Z(g4001) ) ;
INV     gate2788  (.A(g3192), .Z(g4002) ) ;
INV     gate2789  (.A(g3192), .Z(g4003) ) ;
INV     gate2790  (.A(g2845), .Z(g4004) ) ;
INV     gate2791  (.A(g3591), .Z(II7746) ) ;
INV     gate2792  (.A(II7746), .Z(g4005) ) ;
INV     gate2793  (.A(g3692), .Z(II7749) ) ;
INV     gate2794  (.A(II7749), .Z(g4006) ) ;
INV     gate2795  (.A(g3591), .Z(II7752) ) ;
INV     gate2796  (.A(II7752), .Z(g4007) ) ;
INV     gate2797  (.A(g3019), .Z(II7755) ) ;
INV     gate2798  (.A(II7755), .Z(g4008) ) ;
INV     gate2799  (.A(g2605), .Z(II7758) ) ;
INV     gate2800  (.A(II7758), .Z(g4009) ) ;
INV     gate2801  (.A(g3097), .Z(g4010) ) ;
INV     gate2802  (.A(g3029), .Z(II7762) ) ;
INV     gate2803  (.A(II7762), .Z(g4011) ) ;
INV     gate2804  (.A(g2595), .Z(II7765) ) ;
INV     gate2805  (.A(II7765), .Z(g4012) ) ;
INV     gate2806  (.A(g3131), .Z(g4013) ) ;
INV     gate2807  (.A(g3038), .Z(II7769) ) ;
INV     gate2808  (.A(II7769), .Z(g4014) ) ;
INV     gate2809  (.A(g3160), .Z(g4015) ) ;
INV     gate2810  (.A(g3192), .Z(g4016) ) ;
INV     gate2811  (.A(g2845), .Z(g4017) ) ;
INV     gate2812  (.A(g3705), .Z(II7775) ) ;
INV     gate2813  (.A(II7775), .Z(g4018) ) ;
INV     gate2814  (.A(g3019), .Z(II7778) ) ;
INV     gate2815  (.A(II7778), .Z(g4019) ) ;
INV     gate2816  (.A(g2605), .Z(II7781) ) ;
INV     gate2817  (.A(II7781), .Z(g4020) ) ;
INV     gate2818  (.A(g3131), .Z(g4021) ) ;
INV     gate2819  (.A(g3029), .Z(II7785) ) ;
INV     gate2820  (.A(II7785), .Z(g4022) ) ;
INV     gate2821  (.A(g2595), .Z(II7788) ) ;
INV     gate2822  (.A(II7788), .Z(g4023) ) ;
INV     gate2823  (.A(g3160), .Z(g4024) ) ;
INV     gate2824  (.A(g3038), .Z(II7792) ) ;
INV     gate2825  (.A(II7792), .Z(g4025) ) ;
INV     gate2826  (.A(g3192), .Z(g4026) ) ;
INV     gate2827  (.A(g2845), .Z(g4027) ) ;
INV     gate2828  (.A(g3019), .Z(II7797) ) ;
INV     gate2829  (.A(II7797), .Z(g4028) ) ;
INV     gate2830  (.A(g2605), .Z(II7800) ) ;
INV     gate2831  (.A(II7800), .Z(g4029) ) ;
INV     gate2832  (.A(g3160), .Z(g4030) ) ;
INV     gate2833  (.A(g3029), .Z(II7804) ) ;
INV     gate2834  (.A(II7804), .Z(g4031) ) ;
INV     gate2835  (.A(g2595), .Z(II7807) ) ;
INV     gate2836  (.A(II7807), .Z(g4032) ) ;
INV     gate2837  (.A(g3192), .Z(g4033) ) ;
INV     gate2838  (.A(g3019), .Z(II7811) ) ;
INV     gate2839  (.A(II7811), .Z(g4034) ) ;
INV     gate2840  (.A(g2605), .Z(II7814) ) ;
INV     gate2841  (.A(II7814), .Z(g4035) ) ;
INV     gate2842  (.A(g3192), .Z(g4036) ) ;
INV     gate2843  (.A(g2845), .Z(g4037) ) ;
INV     gate2844  (.A(g2605), .Z(g4041) ) ;
INV     gate2845  (.A(g2595), .Z(g4044) ) ;
INV     gate2846  (.A(g3080), .Z(g4050) ) ;
INV     gate2847  (.A(g3093), .Z(g4051) ) ;
INV     gate2848  (.A(g3082), .Z(g4056) ) ;
AND2    gate2849  (.A(g1597), .B(g973), .Z(g2768) ) ;
INV     gate2850  (.A(g2768), .Z(II7832) ) ;
INV     gate2851  (.A(II7832), .Z(g4057) ) ;
AND2    gate2852  (.A(g1600), .B(g976), .Z(g2781) ) ;
INV     gate2853  (.A(g2781), .Z(II7838) ) ;
INV     gate2854  (.A(II7838), .Z(g4065) ) ;
INV     gate2855  (.A(g3784), .Z(II7844) ) ;
INV     gate2856  (.A(II7844), .Z(g4069) ) ;
INV     gate2857  (.A(g3798), .Z(II7847) ) ;
INV     gate2858  (.A(II7847), .Z(g4070) ) ;
INV     gate2859  (.A(g2795), .Z(II7850) ) ;
INV     gate2860  (.A(II7850), .Z(g4071) ) ;
INV     gate2861  (.A(g3805), .Z(II7856) ) ;
INV     gate2862  (.A(II7856), .Z(g4075) ) ;
INV     gate2863  (.A(g2804), .Z(II7859) ) ;
INV     gate2864  (.A(II7859), .Z(g4076) ) ;
INV     gate2865  (.A(g3812), .Z(II7864) ) ;
INV     gate2866  (.A(II7864), .Z(g4079) ) ;
INV     gate2867  (.A(g2818), .Z(II7867) ) ;
INV     gate2868  (.A(II7867), .Z(g4080) ) ;
AND2    gate2869  (.A(g1889), .B(g1690), .Z(g2827) ) ;
INV     gate2870  (.A(g2827), .Z(II7870) ) ;
INV     gate2871  (.A(II7870), .Z(g4081) ) ;
INV     gate2872  (.A(g3819), .Z(II7875) ) ;
INV     gate2873  (.A(II7875), .Z(g4084) ) ;
INV     gate2874  (.A(g2829), .Z(II7878) ) ;
INV     gate2875  (.A(II7878), .Z(g4085) ) ;
INV     gate2876  (.A(g2700), .Z(II7882) ) ;
INV     gate2877  (.A(II7882), .Z(g4087) ) ;
INV     gate2878  (.A(g2837), .Z(II7885) ) ;
INV     gate2879  (.A(II7885), .Z(g4088) ) ;
NOR2    gate2880  (.A(g2263), .B(g1395), .Z(g3505) ) ;
INV     gate2881  (.A(g3505), .Z(II7888) ) ;
INV     gate2882  (.A(II7888), .Z(g4089) ) ;
INV     gate2883  (.A(g3743), .Z(II7899) ) ;
INV     gate2884  (.A(II7899), .Z(g4092) ) ;
INV     gate2885  (.A(g2709), .Z(II7902) ) ;
INV     gate2886  (.A(II7902), .Z(g4093) ) ;
INV     gate2887  (.A(g2863), .Z(II7905) ) ;
INV     gate2888  (.A(II7905), .Z(g4094) ) ;
NOR2    gate2889  (.A(g2282), .B(g1401), .Z(g3516) ) ;
INV     gate2890  (.A(g3516), .Z(II7908) ) ;
INV     gate2891  (.A(II7908), .Z(g4095) ) ;
INV     gate2892  (.A(g2767), .Z(II7911) ) ;
INV     gate2893  (.A(II7911), .Z(g4096) ) ;
INV     gate2894  (.A(g3761), .Z(II7919) ) ;
INV     gate2895  (.A(II7919), .Z(g4102) ) ;
INV     gate2896  (.A(g3462), .Z(II7922) ) ;
INV     gate2897  (.A(II7922), .Z(g4103) ) ;
INV     gate2898  (.A(g2761), .Z(II7925) ) ;
INV     gate2899  (.A(II7925), .Z(g4104) ) ;
INV     gate2900  (.A(g2873), .Z(II7928) ) ;
INV     gate2901  (.A(II7928), .Z(g4105) ) ;
INV     gate2902  (.A(g2780), .Z(II7931) ) ;
INV     gate2903  (.A(II7931), .Z(g4106) ) ;
INV     gate2904  (.A(g3774), .Z(II7944) ) ;
INV     gate2905  (.A(II7944), .Z(g4111) ) ;
INV     gate2906  (.A(g3485), .Z(II7947) ) ;
INV     gate2907  (.A(II7947), .Z(g4112) ) ;
INV     gate2908  (.A(g2774), .Z(II7950) ) ;
INV     gate2909  (.A(II7950), .Z(g4113) ) ;
INV     gate2910  (.A(g3542), .Z(II7953) ) ;
INV     gate2911  (.A(II7953), .Z(g4114) ) ;
INV     gate2912  (.A(g2810), .Z(II7956) ) ;
INV     gate2913  (.A(II7956), .Z(g4115) ) ;
INV     gate2914  (.A(g2793), .Z(II7959) ) ;
INV     gate2915  (.A(II7959), .Z(g4116) ) ;
INV     gate2916  (.A(g3488), .Z(II7964) ) ;
INV     gate2917  (.A(II7964), .Z(g4119) ) ;
INV     gate2918  (.A(g2787), .Z(II7967) ) ;
INV     gate2919  (.A(II7967), .Z(g4120) ) ;
INV     gate2920  (.A(g3557), .Z(II7970) ) ;
INV     gate2921  (.A(II7970), .Z(g4121) ) ;
INV     gate2922  (.A(g3071), .Z(II7973) ) ;
INV     gate2923  (.A(II7973), .Z(g4122) ) ;
INV     gate2924  (.A(g3574), .Z(II7978) ) ;
INV     gate2925  (.A(II7978), .Z(g4125) ) ;
NOR2    gate2926  (.A(g2359), .B(g1398), .Z(g3555) ) ;
INV     gate2927  (.A(g3555), .Z(II7981) ) ;
INV     gate2928  (.A(II7981), .Z(g4126) ) ;
NOR2    gate2929  (.A(g2343), .B(g1391), .Z(g3528) ) ;
INV     gate2930  (.A(g3528), .Z(II7987) ) ;
INV     gate2931  (.A(II7987), .Z(g4130) ) ;
INV     gate2932  (.A(g3676), .Z(g4134) ) ;
NOR3    gate2933  (.A(g1021), .B(g1025), .C(g1889), .Z(g3225) ) ;
INV     gate2934  (.A(g3225), .Z(II8011) ) ;
INV     gate2935  (.A(II8011), .Z(g4146) ) ;
INV     gate2936  (.A(g3076), .Z(II8024) ) ;
INV     gate2937  (.A(II8024), .Z(g4153) ) ;
NAND2   gate2938  (.A(g1556), .B(g2510), .Z(g3706) ) ;
INV     gate2939  (.A(g3706), .Z(II8084) ) ;
INV     gate2940  (.A(II8084), .Z(g4191) ) ;
INV     gate2941  (.A(g2976), .Z(II8094) ) ;
INV     gate2942  (.A(II8094), .Z(g4195) ) ;
NOR3    gate2943  (.A(g1444), .B(g1838), .C(g1454), .Z(g3237) ) ;
INV     gate2944  (.A(g3237), .Z(II8097) ) ;
INV     gate2945  (.A(II8097), .Z(g4196) ) ;
INV     gate2946  (.A(g3591), .Z(g4197) ) ;
AND2    gate2947  (.A(g1976), .B(g1960), .Z(g3259) ) ;
INV     gate2948  (.A(g3259), .Z(II8101) ) ;
INV     gate2949  (.A(II8101), .Z(g4198) ) ;
OR2     gate2950  (.A(g1424), .B(g2014), .Z(g3339) ) ;
INV     gate2951  (.A(g3339), .Z(II8105) ) ;
INV     gate2952  (.A(II8105), .Z(g4200) ) ;
INV     gate2953  (.A(g2810), .Z(g4202) ) ;
INV     gate2954  (.A(g3591), .Z(g4226) ) ;
AND3    gate2955  (.A(g1454), .B(g1838), .C(g1444), .Z(g3429) ) ;
INV     gate2956  (.A(g3429), .Z(II8140) ) ;
INV     gate2957  (.A(II8140), .Z(g4229) ) ;
INV     gate2958  (.A(g3517), .Z(II8161) ) ;
INV     gate2959  (.A(II8161), .Z(g4242) ) ;
INV     gate2960  (.A(g3524), .Z(II8172) ) ;
INV     gate2961  (.A(II8172), .Z(g4245) ) ;
INV     gate2962  (.A(g2810), .Z(II8177) ) ;
INV     gate2963  (.A(II8177), .Z(g4250) ) ;
INV     gate2964  (.A(g3529), .Z(II8180) ) ;
INV     gate2965  (.A(II8180), .Z(g4251) ) ;
INV     gate2966  (.A(g2734), .Z(g4253) ) ;
INV     gate2967  (.A(g3545), .Z(II8190) ) ;
INV     gate2968  (.A(II8190), .Z(g4257) ) ;
INV     gate2969  (.A(g3547), .Z(II8193) ) ;
INV     gate2970  (.A(II8193), .Z(g4258) ) ;
INV     gate2971  (.A(g3654), .Z(II8196) ) ;
INV     gate2972  (.A(II8196), .Z(g4259) ) ;
INV     gate2973  (.A(g3591), .Z(g4265) ) ;
INV     gate2974  (.A(g3560), .Z(II8202) ) ;
INV     gate2975  (.A(II8202), .Z(g4266) ) ;
INV     gate2976  (.A(g2655), .Z(II8205) ) ;
INV     gate2977  (.A(g2573), .Z(g4270) ) ;
INV     gate2978  (.A(g3577), .Z(II8215) ) ;
INV     gate2979  (.A(II8215), .Z(g4273) ) ;
AND2    gate2980  (.A(g871), .B(g1834), .Z(g3002) ) ;
INV     gate2981  (.A(g3002), .Z(II8218) ) ;
INV     gate2982  (.A(II8218), .Z(g4274) ) ;
NOR3    gate2983  (.A(g985), .B(g990), .C(g2295), .Z(g3790) ) ;
INV     gate2984  (.A(g3790), .Z(g4275) ) ;
INV     gate2985  (.A(g3340), .Z(g4279) ) ;
INV     gate2986  (.A(g2562), .Z(g4281) ) ;
INV     gate2987  (.A(g3588), .Z(II8233) ) ;
INV     gate2988  (.A(II8233), .Z(g4285) ) ;
INV     gate2989  (.A(g3790), .Z(g4286) ) ;
INV     gate2990  (.A(g3790), .Z(g4296) ) ;
INV     gate2991  (.A(g3643), .Z(II8261) ) ;
INV     gate2992  (.A(II8261), .Z(g4300) ) ;
INV     gate2993  (.A(g3653), .Z(II8264) ) ;
INV     gate2994  (.A(II8264), .Z(g4301) ) ;
NAND2   gate2995  (.A(II6539), .B(II6540), .Z(g2801) ) ;
INV     gate2996  (.A(g2801), .Z(II8268) ) ;
INV     gate2997  (.A(II8268), .Z(g4303) ) ;
INV     gate2998  (.A(g2976), .Z(II8273) ) ;
INV     gate2999  (.A(II8273), .Z(g4306) ) ;
INV     gate3000  (.A(g3700), .Z(g4307) ) ;
NOR4    gate3001  (.A(g1375), .B(g2229), .C(g2213), .D(g2206), .Z(g3504) ) ;
INV     gate3002  (.A(g3504), .Z(II8277) ) ;
INV     gate3003  (.A(II8277), .Z(g4308) ) ;
NOR4    gate3004  (.A(g1388), .B(g2262), .C(g2230), .D(g2214), .Z(g3515) ) ;
INV     gate3005  (.A(g3515), .Z(II8282) ) ;
INV     gate3006  (.A(II8282), .Z(g4311) ) ;
INV     gate3007  (.A(g878), .Z(II8291) ) ;
INV     gate3008  (.A(g3086), .Z(g4328) ) ;
INV     gate3009  (.A(g3659), .Z(g4335) ) ;
INV     gate3010  (.A(g3674), .Z(II8308) ) ;
INV     gate3011  (.A(II8308), .Z(g4341) ) ;
INV     gate3012  (.A(g3124), .Z(g4344) ) ;
INV     gate3013  (.A(g3691), .Z(II8315) ) ;
INV     gate3014  (.A(II8315), .Z(g4350) ) ;
NAND2   gate3015  (.A(II7157), .B(II7158), .Z(g3665) ) ;
INV     gate3016  (.A(g3665), .Z(g4353) ) ;
NAND2   gate3017  (.A(II7180), .B(II7181), .Z(g3679) ) ;
INV     gate3018  (.A(g3679), .Z(g4357) ) ;
NAND2   gate3019  (.A(II7187), .B(II7188), .Z(g3680) ) ;
INV     gate3020  (.A(g3680), .Z(g4358) ) ;
INV     gate3021  (.A(g3721), .Z(II8333) ) ;
INV     gate3022  (.A(II8333), .Z(g4360) ) ;
INV     gate3023  (.A(g2810), .Z(g4362) ) ;
INV     gate3024  (.A(g1160), .Z(II8351) ) ;
INV     gate3025  (.A(g1163), .Z(II8354) ) ;
INV     gate3026  (.A(g1182), .Z(II8357) ) ;
INV     gate3027  (.A(g1186), .Z(II8360) ) ;
INV     gate3028  (.A(g3466), .Z(g4381) ) ;
INV     gate3029  (.A(g3783), .Z(II8373) ) ;
INV     gate3030  (.A(II8373), .Z(g4382) ) ;
INV     gate3031  (.A(g3611), .Z(II8428) ) ;
INV     gate3032  (.A(II8428), .Z(g4426) ) ;
INV     gate3033  (.A(g3014), .Z(II8446) ) ;
INV     gate3034  (.A(II8446), .Z(g4438) ) ;
INV     gate3035  (.A(g3630), .Z(II8449) ) ;
INV     gate3036  (.A(II8449), .Z(g4443) ) ;
INV     gate3037  (.A(g2816), .Z(II8452) ) ;
INV     gate3038  (.A(II8452), .Z(g4444) ) ;
NAND2   gate3039  (.A(II7269), .B(II7270), .Z(g3811) ) ;
INV     gate3040  (.A(g3811), .Z(g4455) ) ;
INV     gate3041  (.A(g3014), .Z(II8477) ) ;
INV     gate3042  (.A(II8477), .Z(g4457) ) ;
INV     gate3043  (.A(g3640), .Z(II8480) ) ;
INV     gate3044  (.A(II8480), .Z(g4462) ) ;
INV     gate3045  (.A(g3641), .Z(II8483) ) ;
INV     gate3046  (.A(II8483), .Z(g4463) ) ;
INV     gate3047  (.A(g2824), .Z(II8486) ) ;
INV     gate3048  (.A(II8486), .Z(g4464) ) ;
INV     gate3049  (.A(g3677), .Z(g4465) ) ;
NAND2   gate3050  (.A(II7278), .B(II7279), .Z(g3818) ) ;
INV     gate3051  (.A(g3818), .Z(g4475) ) ;
INV     gate3052  (.A(g3014), .Z(II8517) ) ;
INV     gate3053  (.A(II8517), .Z(g4477) ) ;
INV     gate3054  (.A(g3652), .Z(II8520) ) ;
INV     gate3055  (.A(II8520), .Z(g4482) ) ;
INV     gate3056  (.A(g2826), .Z(g4489) ) ;
INV     gate3057  (.A(g2810), .Z(II8543) ) ;
INV     gate3058  (.A(II8543), .Z(g4493) ) ;
INV     gate3059  (.A(g2832), .Z(g4500) ) ;
INV     gate3060  (.A(g2801), .Z(g4501) ) ;
INV     gate3061  (.A(g3071), .Z(II8565) ) ;
INV     gate3062  (.A(II8565), .Z(g4503) ) ;
INV     gate3063  (.A(g2840), .Z(g4510) ) ;
INV     gate3064  (.A(g2841), .Z(g4511) ) ;
INV     gate3065  (.A(g2842), .Z(g4512) ) ;
INV     gate3066  (.A(g2866), .Z(g4521) ) ;
INV     gate3067  (.A(g2867), .Z(g4522) ) ;
INV     gate3068  (.A(g2868), .Z(g4523) ) ;
INV     gate3069  (.A(g2869), .Z(g4524) ) ;
INV     gate3070  (.A(g2870), .Z(g4525) ) ;
INV     gate3071  (.A(g3466), .Z(g4527) ) ;
INV     gate3072  (.A(g2876), .Z(g4535) ) ;
INV     gate3073  (.A(g2877), .Z(g4536) ) ;
INV     gate3074  (.A(g2878), .Z(g4537) ) ;
INV     gate3075  (.A(g2880), .Z(g4538) ) ;
INV     gate3076  (.A(g2881), .Z(g4539) ) ;
INV     gate3077  (.A(g2882), .Z(g4540) ) ;
INV     gate3078  (.A(g2883), .Z(g4541) ) ;
INV     gate3079  (.A(g2884), .Z(g4542) ) ;
INV     gate3080  (.A(g2885), .Z(g4543) ) ;
INV     gate3081  (.A(g2886), .Z(g4544) ) ;
INV     gate3082  (.A(g2887), .Z(g4545) ) ;
INV     gate3083  (.A(g3466), .Z(g4547) ) ;
INV     gate3084  (.A(g2890), .Z(g4552) ) ;
INV     gate3085  (.A(g2891), .Z(g4553) ) ;
INV     gate3086  (.A(g2892), .Z(g4554) ) ;
INV     gate3087  (.A(g2894), .Z(g4555) ) ;
INV     gate3088  (.A(g2895), .Z(g4556) ) ;
INV     gate3089  (.A(g2896), .Z(g4557) ) ;
INV     gate3090  (.A(g2897), .Z(g4558) ) ;
INV     gate3091  (.A(g2898), .Z(g4559) ) ;
INV     gate3092  (.A(g2899), .Z(g4560) ) ;
INV     gate3093  (.A(g2900), .Z(g4561) ) ;
INV     gate3094  (.A(g3466), .Z(g4562) ) ;
INV     gate3095  (.A(g3051), .Z(II8665) ) ;
INV     gate3096  (.A(II8665), .Z(g4564) ) ;
INV     gate3097  (.A(g2901), .Z(g4565) ) ;
INV     gate3098  (.A(g2902), .Z(g4566) ) ;
INV     gate3099  (.A(g2903), .Z(g4567) ) ;
INV     gate3100  (.A(g2904), .Z(g4568) ) ;
INV     gate3101  (.A(g2906), .Z(g4569) ) ;
INV     gate3102  (.A(g2907), .Z(g4570) ) ;
INV     gate3103  (.A(g2908), .Z(g4571) ) ;
INV     gate3104  (.A(g2909), .Z(g4572) ) ;
INV     gate3105  (.A(g2911), .Z(g4573) ) ;
INV     gate3106  (.A(g3466), .Z(g4574) ) ;
INV     gate3107  (.A(g2913), .Z(g4576) ) ;
INV     gate3108  (.A(g2914), .Z(g4577) ) ;
INV     gate3109  (.A(g2917), .Z(g4578) ) ;
INV     gate3110  (.A(g2918), .Z(g4579) ) ;
INV     gate3111  (.A(g2919), .Z(g4580) ) ;
INV     gate3112  (.A(g2921), .Z(g4581) ) ;
INV     gate3113  (.A(g2922), .Z(g4582) ) ;
INV     gate3114  (.A(g2924), .Z(g4583) ) ;
INV     gate3115  (.A(g3466), .Z(g4584) ) ;
INV     gate3116  (.A(g2925), .Z(g4585) ) ;
INV     gate3117  (.A(g2926), .Z(g4586) ) ;
INV     gate3118  (.A(g2928), .Z(g4587) ) ;
INV     gate3119  (.A(g2929), .Z(g4588) ) ;
INV     gate3120  (.A(g2930), .Z(g4589) ) ;
INV     gate3121  (.A(g2932), .Z(g4590) ) ;
INV     gate3122  (.A(g2937), .Z(g4591) ) ;
INV     gate3123  (.A(g2938), .Z(g4592) ) ;
INV     gate3124  (.A(g2939), .Z(g4593) ) ;
INV     gate3125  (.A(g2941), .Z(g4594) ) ;
INV     gate3126  (.A(g2942), .Z(g4595) ) ;
INV     gate3127  (.A(g3466), .Z(g4596) ) ;
INV     gate3128  (.A(g3828), .Z(II8706) ) ;
INV     gate3129  (.A(II8706), .Z(g4597) ) ;
INV     gate3130  (.A(g4191), .Z(II8709) ) ;
INV     gate3131  (.A(g4007), .Z(II8712) ) ;
INV     gate3132  (.A(g3903), .Z(II8715) ) ;
INV     gate3133  (.A(g3909), .Z(II8718) ) ;
INV     gate3134  (.A(g3918), .Z(II8721) ) ;
INV     gate3135  (.A(g3927), .Z(II8724) ) ;
INV     gate3136  (.A(g3944), .Z(II8727) ) ;
INV     gate3137  (.A(g3987), .Z(II8730) ) ;
INV     gate3138  (.A(g3996), .Z(II8733) ) ;
INV     gate3139  (.A(g4008), .Z(II8736) ) ;
INV     gate3140  (.A(g3910), .Z(II8739) ) ;
INV     gate3141  (.A(g3919), .Z(II8742) ) ;
INV     gate3142  (.A(g3929), .Z(II8745) ) ;
INV     gate3143  (.A(g3997), .Z(II8748) ) ;
INV     gate3144  (.A(g4009), .Z(II8751) ) ;
INV     gate3145  (.A(g3911), .Z(II8754) ) ;
INV     gate3146  (.A(g3921), .Z(II8757) ) ;
INV     gate3147  (.A(g3931), .Z(II8760) ) ;
INV     gate3148  (.A(g3947), .Z(II8763) ) ;
INV     gate3149  (.A(g3960), .Z(II8766) ) ;
INV     gate3150  (.A(g3999), .Z(II8769) ) ;
INV     gate3151  (.A(g4011), .Z(II8772) ) ;
INV     gate3152  (.A(g4019), .Z(II8775) ) ;
INV     gate3153  (.A(g3922), .Z(II8778) ) ;
INV     gate3154  (.A(g3932), .Z(II8781) ) ;
INV     gate3155  (.A(g3949), .Z(II8784) ) ;
INV     gate3156  (.A(g4012), .Z(II8787) ) ;
INV     gate3157  (.A(g4020), .Z(II8790) ) ;
INV     gate3158  (.A(g3923), .Z(II8793) ) ;
INV     gate3159  (.A(g3934), .Z(II8796) ) ;
INV     gate3160  (.A(g3951), .Z(II8799) ) ;
INV     gate3161  (.A(g3963), .Z(II8802) ) ;
INV     gate3162  (.A(g3976), .Z(II8805) ) ;
INV     gate3163  (.A(g4014), .Z(II8808) ) ;
INV     gate3164  (.A(g4022), .Z(II8811) ) ;
INV     gate3165  (.A(g4028), .Z(II8814) ) ;
INV     gate3166  (.A(g3935), .Z(II8817) ) ;
INV     gate3167  (.A(g3952), .Z(II8820) ) ;
INV     gate3168  (.A(g3965), .Z(II8823) ) ;
INV     gate3169  (.A(g4023), .Z(II8826) ) ;
INV     gate3170  (.A(g4029), .Z(II8829) ) ;
INV     gate3171  (.A(g3936), .Z(II8832) ) ;
INV     gate3172  (.A(g3954), .Z(II8835) ) ;
INV     gate3173  (.A(g3967), .Z(II8838) ) ;
INV     gate3174  (.A(g3979), .Z(II8841) ) ;
INV     gate3175  (.A(g3992), .Z(II8844) ) ;
INV     gate3176  (.A(g4025), .Z(II8847) ) ;
INV     gate3177  (.A(g4031), .Z(II8850) ) ;
INV     gate3178  (.A(g4034), .Z(II8853) ) ;
INV     gate3179  (.A(g3955), .Z(II8856) ) ;
INV     gate3180  (.A(g3968), .Z(II8859) ) ;
INV     gate3181  (.A(g3981), .Z(II8862) ) ;
INV     gate3182  (.A(g4032), .Z(II8865) ) ;
INV     gate3183  (.A(g4035), .Z(II8868) ) ;
INV     gate3184  (.A(g3869), .Z(II8871) ) ;
INV     gate3185  (.A(g3884), .Z(II8874) ) ;
INV     gate3186  (.A(g4274), .Z(II8877) ) ;
INV     gate3187  (.A(g4303), .Z(II8880) ) ;
INV     gate3188  (.A(g4198), .Z(II8883) ) ;
INV     gate3189  (.A(g4308), .Z(II8886) ) ;
INV     gate3190  (.A(g4311), .Z(II8889) ) ;
INV     gate3191  (.A(g4115), .Z(II8892) ) ;
INV     gate3192  (.A(g4130), .Z(II8895) ) ;
INV     gate3193  (.A(g4089), .Z(II8898) ) ;
INV     gate3194  (.A(g4122), .Z(II8901) ) ;
INV     gate3195  (.A(g4126), .Z(II8904) ) ;
INV     gate3196  (.A(g4095), .Z(II8907) ) ;
INV     gate3197  (.A(g4200), .Z(II8910) ) ;
INV     gate3198  (.A(g4306), .Z(II8913) ) ;
INV     gate3199  (.A(g4195), .Z(II8916) ) ;
INV     gate3200  (.A(g4196), .Z(II8919) ) ;
INV     gate3201  (.A(g4229), .Z(II8922) ) ;
INV     gate3202  (.A(g4482), .Z(II8925) ) ;
INV     gate3203  (.A(II8925), .Z(g4670) ) ;
INV     gate3204  (.A(g4153), .Z(II8928) ) ;
INV     gate3205  (.A(II8928), .Z(g4673) ) ;
INV     gate3206  (.A(g4096), .Z(II8932) ) ;
INV     gate3207  (.A(II8932), .Z(g4677) ) ;
INV     gate3208  (.A(g4005), .Z(II8935) ) ;
INV     gate3209  (.A(II8935), .Z(g4678) ) ;
INV     gate3210  (.A(g4106), .Z(II8945) ) ;
INV     gate3211  (.A(II8945), .Z(g4680) ) ;
INV     gate3212  (.A(g4116), .Z(II8949) ) ;
INV     gate3213  (.A(II8949), .Z(g4684) ) ;
INV     gate3214  (.A(g4197), .Z(II8952) ) ;
INV     gate3215  (.A(II8952), .Z(g4685) ) ;
INV     gate3216  (.A(g4553), .Z(II8962) ) ;
INV     gate3217  (.A(II8962), .Z(g4687) ) ;
INV     gate3218  (.A(g4444), .Z(II8966) ) ;
INV     gate3219  (.A(II8966), .Z(g4689) ) ;
INV     gate3220  (.A(g4464), .Z(II8971) ) ;
INV     gate3221  (.A(II8971), .Z(g4692) ) ;
INV     gate3222  (.A(g3871), .Z(II8974) ) ;
INV     gate3223  (.A(II8974), .Z(g4693) ) ;
INV     gate3224  (.A(g3877), .Z(II8977) ) ;
INV     gate3225  (.A(II8977), .Z(g4694) ) ;
INV     gate3226  (.A(g4535), .Z(II8980) ) ;
INV     gate3227  (.A(II8980), .Z(g4695) ) ;
INV     gate3228  (.A(g4536), .Z(II8983) ) ;
INV     gate3229  (.A(II8983), .Z(g4696) ) ;
INV     gate3230  (.A(g4552), .Z(II8986) ) ;
INV     gate3231  (.A(II8986), .Z(g4697) ) ;
INV     gate3232  (.A(g4537), .Z(II8989) ) ;
INV     gate3233  (.A(II8989), .Z(g4698) ) ;
INV     gate3234  (.A(g4565), .Z(II8994) ) ;
INV     gate3235  (.A(II8994), .Z(g4701) ) ;
INV     gate3236  (.A(g4576), .Z(II8998) ) ;
INV     gate3237  (.A(II8998), .Z(g4703) ) ;
INV     gate3238  (.A(g4577), .Z(II9001) ) ;
INV     gate3239  (.A(II9001), .Z(g4704) ) ;
INV     gate3240  (.A(g4585), .Z(II9005) ) ;
INV     gate3241  (.A(II9005), .Z(g4706) ) ;
INV     gate3242  (.A(g4591), .Z(II9009) ) ;
INV     gate3243  (.A(II9009), .Z(g4710) ) ;
INV     gate3244  (.A(g3864), .Z(II9014) ) ;
INV     gate3245  (.A(II9014), .Z(g4713) ) ;
INV     gate3246  (.A(g3872), .Z(II9018) ) ;
INV     gate3247  (.A(II9018), .Z(g4718) ) ;
INV     gate3248  (.A(g4489), .Z(II9021) ) ;
INV     gate3249  (.A(II9021), .Z(g4719) ) ;
INV     gate3250  (.A(g4462), .Z(II9025) ) ;
INV     gate3251  (.A(II9025), .Z(g4721) ) ;
AND4    gate3252  (.A(g878), .B(g3086), .C(g1857), .D(g3659), .Z(g4317) ) ;
INV     gate3253  (.A(g4317), .Z(II9034) ) ;
INV     gate3254  (.A(II9034), .Z(g4732) ) ;
INV     gate3255  (.A(g4202), .Z(g4733) ) ;
INV     gate3256  (.A(g3881), .Z(II9050) ) ;
INV     gate3257  (.A(II9050), .Z(g4738) ) ;
AND2    gate3258  (.A(g2959), .B(g1867), .Z(g4327) ) ;
INV     gate3259  (.A(g4327), .Z(II9053) ) ;
INV     gate3260  (.A(II9053), .Z(g4739) ) ;
AND3    gate3261  (.A(g3086), .B(g3659), .C(g3124), .Z(g4302) ) ;
INV     gate3262  (.A(g4302), .Z(II9064) ) ;
INV     gate3263  (.A(II9064), .Z(g4742) ) ;
INV     gate3264  (.A(g4353), .Z(II9076) ) ;
INV     gate3265  (.A(II9076), .Z(g4746) ) ;
INV     gate3266  (.A(g4465), .Z(g4748) ) ;
INV     gate3267  (.A(g4357), .Z(II9081) ) ;
INV     gate3268  (.A(II9081), .Z(g4776) ) ;
INV     gate3269  (.A(g4358), .Z(II9084) ) ;
INV     gate3270  (.A(II9084), .Z(g4777) ) ;
INV     gate3271  (.A(g4566), .Z(II9089) ) ;
INV     gate3272  (.A(II9089), .Z(g4780) ) ;
OR2     gate3273  (.A(g3587), .B(g2665), .Z(g4283) ) ;
INV     gate3274  (.A(g4283), .Z(II9095) ) ;
INV     gate3275  (.A(II9095), .Z(g4784) ) ;
OR4     gate3276  (.A(g1182), .B(g1186), .C(g1179), .D(II8363), .Z(g4374) ) ;
INV     gate3277  (.A(g4374), .Z(II9103) ) ;
INV     gate3278  (.A(II9103), .Z(g4788) ) ;
NOR2    gate3279  (.A(g1934), .B(g3591), .Z(g4232) ) ;
INV     gate3280  (.A(g4232), .Z(II9111) ) ;
INV     gate3281  (.A(II9111), .Z(g4792) ) ;
OR2     gate3282  (.A(g3617), .B(g3602), .Z(g4297) ) ;
INV     gate3283  (.A(g4297), .Z(II9116) ) ;
INV     gate3284  (.A(II9116), .Z(g4795) ) ;
INV     gate3285  (.A(g4455), .Z(II9123) ) ;
INV     gate3286  (.A(II9123), .Z(g4800) ) ;
INV     gate3287  (.A(g3870), .Z(II9126) ) ;
INV     gate3288  (.A(II9126), .Z(g4801) ) ;
INV     gate3289  (.A(g4475), .Z(II9129) ) ;
INV     gate3290  (.A(II9129), .Z(g4802) ) ;
AND2    gate3291  (.A(g3260), .B(g3314), .Z(g4284) ) ;
INV     gate3292  (.A(g4284), .Z(II9132) ) ;
INV     gate3293  (.A(II9132), .Z(g4803) ) ;
OR2     gate3294  (.A(II8224), .B(II8225), .Z(g4280) ) ;
INV     gate3295  (.A(g4280), .Z(II9136) ) ;
INV     gate3296  (.A(II9136), .Z(g4805) ) ;
OR2     gate3297  (.A(g2952), .B(g1725), .Z(g4364) ) ;
INV     gate3298  (.A(g4364), .Z(II9139) ) ;
INV     gate3299  (.A(II9139), .Z(g4806) ) ;
AND2    gate3300  (.A(g3260), .B(g3221), .Z(g4236) ) ;
INV     gate3301  (.A(g4236), .Z(II9142) ) ;
INV     gate3302  (.A(II9142), .Z(g4807) ) ;
OR2     gate3303  (.A(g2490), .B(g3315), .Z(g4264) ) ;
INV     gate3304  (.A(g4264), .Z(II9145) ) ;
INV     gate3305  (.A(II9145), .Z(g4808) ) ;
NOR2    gate3306  (.A(g1424), .B(g3541), .Z(g4354) ) ;
INV     gate3307  (.A(g4354), .Z(II9148) ) ;
INV     gate3308  (.A(II9148), .Z(g4809) ) ;
NAND2   gate3309  (.A(g3233), .B(g1444), .Z(g4256) ) ;
INV     gate3310  (.A(g4256), .Z(II9158) ) ;
INV     gate3311  (.A(II9158), .Z(g4811) ) ;
AND2    gate3312  (.A(g3233), .B(g3286), .Z(g4272) ) ;
INV     gate3313  (.A(g4272), .Z(II9162) ) ;
INV     gate3314  (.A(II9162), .Z(g4813) ) ;
AND2    gate3315  (.A(g3233), .B(g3358), .Z(g4299) ) ;
INV     gate3316  (.A(g4299), .Z(II9177) ) ;
INV     gate3317  (.A(II9177), .Z(g4822) ) ;
INV     gate3318  (.A(g4250), .Z(g4841) ) ;
NOR2    gate3319  (.A(g2496), .B(g3310), .Z(g4349) ) ;
INV     gate3320  (.A(g4349), .Z(II9209) ) ;
INV     gate3321  (.A(II9209), .Z(g4867) ) ;
INV     gate3322  (.A(g4443), .Z(II9217) ) ;
INV     gate3323  (.A(II9217), .Z(g4873) ) ;
INV     gate3324  (.A(g4069), .Z(g4882) ) ;
INV     gate3325  (.A(g4070), .Z(g4885) ) ;
INV     gate3326  (.A(g4071), .Z(g4886) ) ;
INV     gate3327  (.A(g4075), .Z(g4890) ) ;
INV     gate3328  (.A(g4076), .Z(g4891) ) ;
INV     gate3329  (.A(g4134), .Z(II9250) ) ;
INV     gate3330  (.A(II9250), .Z(g4892) ) ;
AND4    gate3331  (.A(g3753), .B(g3732), .C(g3712), .D(g3700), .Z(g4078) ) ;
INV     gate3332  (.A(g4078), .Z(g4895) ) ;
INV     gate3333  (.A(g4079), .Z(g4898) ) ;
INV     gate3334  (.A(g4080), .Z(g4899) ) ;
OR2     gate3335  (.A(g3617), .B(g1639), .Z(g4249) ) ;
INV     gate3336  (.A(g4249), .Z(II9258) ) ;
INV     gate3337  (.A(II9258), .Z(g4900) ) ;
INV     gate3338  (.A(g4084), .Z(g4903) ) ;
INV     gate3339  (.A(g4085), .Z(g4904) ) ;
INV     gate3340  (.A(g4087), .Z(g4907) ) ;
INV     gate3341  (.A(g4088), .Z(g4908) ) ;
NAND2   gate3342  (.A(g3260), .B(g1435), .Z(g4263) ) ;
INV     gate3343  (.A(g4263), .Z(II9271) ) ;
INV     gate3344  (.A(II9271), .Z(g4909) ) ;
INV     gate3345  (.A(g4092), .Z(g4913) ) ;
INV     gate3346  (.A(g4093), .Z(g4914) ) ;
INV     gate3347  (.A(g4094), .Z(g4915) ) ;
INV     gate3348  (.A(g4202), .Z(g4916) ) ;
INV     gate3349  (.A(g4102), .Z(g4917) ) ;
INV     gate3350  (.A(g4103), .Z(g4918) ) ;
INV     gate3351  (.A(g4104), .Z(g4919) ) ;
INV     gate3352  (.A(g4105), .Z(g4920) ) ;
INV     gate3353  (.A(g4202), .Z(g4921) ) ;
INV     gate3354  (.A(g4111), .Z(g4922) ) ;
INV     gate3355  (.A(g4112), .Z(g4923) ) ;
INV     gate3356  (.A(g4113), .Z(g4924) ) ;
INV     gate3357  (.A(g4114), .Z(g4925) ) ;
INV     gate3358  (.A(g4202), .Z(g4926) ) ;
INV     gate3359  (.A(g4119), .Z(g4928) ) ;
INV     gate3360  (.A(g4120), .Z(g4929) ) ;
INV     gate3361  (.A(g4121), .Z(g4930) ) ;
OR2     gate3362  (.A(g2828), .B(g2668), .Z(g4295) ) ;
INV     gate3363  (.A(g4295), .Z(II9301) ) ;
INV     gate3364  (.A(II9301), .Z(g4931) ) ;
INV     gate3365  (.A(g4202), .Z(g4932) ) ;
INV     gate3366  (.A(g4125), .Z(g4934) ) ;
INV     gate3367  (.A(g4202), .Z(g4935) ) ;
AND2    gate3368  (.A(g2216), .B(g2655), .Z(g4268) ) ;
INV     gate3369  (.A(g4268), .Z(II9310) ) ;
INV     gate3370  (.A(II9310), .Z(g4938) ) ;
INV     gate3371  (.A(g4259), .Z(g4960) ) ;
INV     gate3372  (.A(g4328), .Z(g4963) ) ;
INV     gate3373  (.A(g4242), .Z(II9325) ) ;
INV     gate3374  (.A(II9325), .Z(g5000) ) ;
INV     gate3375  (.A(g4335), .Z(g5002) ) ;
INV     gate3376  (.A(g4245), .Z(II9333) ) ;
INV     gate3377  (.A(II9333), .Z(g5006) ) ;
INV     gate3378  (.A(g4493), .Z(II9336) ) ;
INV     gate3379  (.A(II9336), .Z(g5007) ) ;
INV     gate3380  (.A(g4344), .Z(g5009) ) ;
INV     gate3381  (.A(g4251), .Z(II9341) ) ;
INV     gate3382  (.A(II9341), .Z(g5013) ) ;
INV     gate3383  (.A(g4341), .Z(II9344) ) ;
INV     gate3384  (.A(II9344), .Z(g5014) ) ;
INV     gate3385  (.A(g3896), .Z(II9347) ) ;
INV     gate3386  (.A(II9347), .Z(g5015) ) ;
INV     gate3387  (.A(g4503), .Z(II9350) ) ;
INV     gate3388  (.A(II9350), .Z(g5016) ) ;
INV     gate3389  (.A(g4438), .Z(g5022) ) ;
INV     gate3390  (.A(g4257), .Z(II9360) ) ;
INV     gate3391  (.A(II9360), .Z(g5024) ) ;
INV     gate3392  (.A(g4258), .Z(II9363) ) ;
INV     gate3393  (.A(II9363), .Z(g5025) ) ;
INV     gate3394  (.A(g4350), .Z(II9366) ) ;
INV     gate3395  (.A(II9366), .Z(g5026) ) ;
INV     gate3396  (.A(g3901), .Z(II9369) ) ;
INV     gate3397  (.A(II9369), .Z(g5027) ) ;
INV     gate3398  (.A(g3902), .Z(II9372) ) ;
INV     gate3399  (.A(II9372), .Z(g5028) ) ;
INV     gate3400  (.A(g4438), .Z(g5037) ) ;
INV     gate3401  (.A(g4457), .Z(g5038) ) ;
INV     gate3402  (.A(g4266), .Z(II9393) ) ;
INV     gate3403  (.A(II9393), .Z(g5041) ) ;
INV     gate3404  (.A(g3908), .Z(II9396) ) ;
INV     gate3405  (.A(II9396), .Z(g5042) ) ;
INV     gate3406  (.A(g4232), .Z(II9407) ) ;
INV     gate3407  (.A(II9407), .Z(g5051) ) ;
INV     gate3408  (.A(g4438), .Z(g5053) ) ;
INV     gate3409  (.A(g4457), .Z(g5054) ) ;
INV     gate3410  (.A(g4477), .Z(g5055) ) ;
INV     gate3411  (.A(g4273), .Z(II9416) ) ;
INV     gate3412  (.A(II9416), .Z(g5058) ) ;
INV     gate3413  (.A(g3916), .Z(II9419) ) ;
INV     gate3414  (.A(II9419), .Z(g5059) ) ;
INV     gate3415  (.A(g4360), .Z(II9422) ) ;
INV     gate3416  (.A(II9422), .Z(g5060) ) ;
INV     gate3417  (.A(g3917), .Z(II9425) ) ;
INV     gate3418  (.A(II9425), .Z(g5061) ) ;
INV     gate3419  (.A(g4438), .Z(g5071) ) ;
INV     gate3420  (.A(g4457), .Z(g5072) ) ;
INV     gate3421  (.A(g4477), .Z(g5073) ) ;
INV     gate3422  (.A(g4285), .Z(II9440) ) ;
INV     gate3423  (.A(II9440), .Z(g5074) ) ;
INV     gate3424  (.A(g4564), .Z(II9443) ) ;
INV     gate3425  (.A(II9443), .Z(g5075) ) ;
INV     gate3426  (.A(g3926), .Z(II9446) ) ;
INV     gate3427  (.A(II9446), .Z(g5076) ) ;
INV     gate3428  (.A(g4457), .Z(g5083) ) ;
INV     gate3429  (.A(g4477), .Z(g5084) ) ;
INV     gate3430  (.A(g3940), .Z(II9457) ) ;
INV     gate3431  (.A(II9457), .Z(g5085) ) ;
INV     gate3432  (.A(g3941), .Z(II9460) ) ;
INV     gate3433  (.A(II9460), .Z(g5086) ) ;
INV     gate3434  (.A(g3942), .Z(II9463) ) ;
INV     gate3435  (.A(II9463), .Z(g5087) ) ;
INV     gate3436  (.A(g3943), .Z(II9466) ) ;
INV     gate3437  (.A(II9466), .Z(g5088) ) ;
INV     gate3438  (.A(g4477), .Z(g5099) ) ;
INV     gate3439  (.A(g3957), .Z(II9484) ) ;
INV     gate3440  (.A(II9484), .Z(g5100) ) ;
INV     gate3441  (.A(g4259), .Z(g5101) ) ;
INV     gate3442  (.A(g4426), .Z(II9493) ) ;
INV     gate3443  (.A(II9493), .Z(g5109) ) ;
INV     gate3444  (.A(g3971), .Z(II9496) ) ;
INV     gate3445  (.A(II9496), .Z(g5112) ) ;
INV     gate3446  (.A(g4382), .Z(II9499) ) ;
INV     gate3447  (.A(II9499), .Z(g5113) ) ;
INV     gate3448  (.A(g3972), .Z(II9502) ) ;
INV     gate3449  (.A(II9502), .Z(g5114) ) ;
INV     gate3450  (.A(g4300), .Z(II9505) ) ;
INV     gate3451  (.A(II9505), .Z(g5115) ) ;
INV     gate3452  (.A(g3985), .Z(II9512) ) ;
INV     gate3453  (.A(II9512), .Z(g5120) ) ;
INV     gate3454  (.A(g4301), .Z(II9515) ) ;
INV     gate3455  (.A(II9515), .Z(g5121) ) ;
INV     gate3456  (.A(g3995), .Z(II9520) ) ;
INV     gate3457  (.A(II9520), .Z(g5124) ) ;
OR2     gate3458  (.A(g2371), .B(g3285), .Z(g4413) ) ;
INV     gate3459  (.A(g4413), .Z(II9525) ) ;
INV     gate3460  (.A(II9525), .Z(g5127) ) ;
INV     gate3461  (.A(g4006), .Z(II9528) ) ;
INV     gate3462  (.A(II9528), .Z(g5128) ) ;
INV     gate3463  (.A(g4463), .Z(II9531) ) ;
INV     gate3464  (.A(II9531), .Z(g5129) ) ;
INV     gate3465  (.A(g4018), .Z(II9539) ) ;
INV     gate3466  (.A(II9539), .Z(g5137) ) ;
INV     gate3467  (.A(g4279), .Z(II9543) ) ;
INV     gate3468  (.A(II9543), .Z(g5139) ) ;
INV     gate3469  (.A(g4892), .Z(II9555) ) ;
INV     gate3470  (.A(g4597), .Z(II9558) ) ;
INV     gate3471  (.A(II9558), .Z(g5144) ) ;
INV     gate3472  (.A(g4695), .Z(II9561) ) ;
INV     gate3473  (.A(g4703), .Z(II9564) ) ;
INV     gate3474  (.A(g4693), .Z(II9567) ) ;
INV     gate3475  (.A(g4696), .Z(II9570) ) ;
INV     gate3476  (.A(g4701), .Z(II9573) ) ;
INV     gate3477  (.A(g4706), .Z(II9576) ) ;
INV     gate3478  (.A(g4713), .Z(II9579) ) ;
INV     gate3479  (.A(g4694), .Z(II9582) ) ;
INV     gate3480  (.A(g4697), .Z(II9585) ) ;
INV     gate3481  (.A(g4704), .Z(II9588) ) ;
INV     gate3482  (.A(g4710), .Z(II9591) ) ;
INV     gate3483  (.A(g4718), .Z(II9594) ) ;
INV     gate3484  (.A(g4738), .Z(II9597) ) ;
INV     gate3485  (.A(g4698), .Z(II9600) ) ;
INV     gate3486  (.A(g4719), .Z(II9603) ) ;
INV     gate3487  (.A(g4687), .Z(II9606) ) ;
INV     gate3488  (.A(g4780), .Z(II9609) ) ;
INV     gate3489  (.A(g4776), .Z(II9612) ) ;
INV     gate3490  (.A(g4739), .Z(II9615) ) ;
INV     gate3491  (.A(g4742), .Z(II9618) ) ;
INV     gate3492  (.A(g4732), .Z(II9621) ) ;
INV     gate3493  (.A(g4746), .Z(II9624) ) ;
INV     gate3494  (.A(g4777), .Z(II9627) ) ;
INV     gate3495  (.A(g4867), .Z(II9630) ) ;
INV     gate3496  (.A(g4800), .Z(II9633) ) ;
INV     gate3497  (.A(g4802), .Z(II9636) ) ;
INV     gate3498  (.A(g4685), .Z(II9639) ) ;
INV     gate3499  (.A(g4788), .Z(II9642) ) ;
INV     gate3500  (.A(g4900), .Z(II9645) ) ;
INV     gate3501  (.A(g4795), .Z(II9648) ) ;
INV     gate3502  (.A(g4805), .Z(II9651) ) ;
INV     gate3503  (.A(g4792), .Z(II9654) ) ;
INV     gate3504  (.A(g4784), .Z(II9657) ) ;
INV     gate3505  (.A(g4806), .Z(II9660) ) ;
INV     gate3506  (.A(g4809), .Z(II9663) ) ;
INV     gate3507  (.A(g4931), .Z(II9666) ) ;
INV     gate3508  (.A(g4909), .Z(II9669) ) ;
INV     gate3509  (.A(g4803), .Z(II9672) ) ;
INV     gate3510  (.A(g4807), .Z(II9675) ) ;
INV     gate3511  (.A(g4808), .Z(II9678) ) ;
INV     gate3512  (.A(g4811), .Z(II9681) ) ;
INV     gate3513  (.A(g4813), .Z(II9684) ) ;
INV     gate3514  (.A(g4822), .Z(II9687) ) ;
INV     gate3515  (.A(g4938), .Z(g5190) ) ;
AND2    gate3516  (.A(g4362), .B(g2216), .Z(g4969) ) ;
INV     gate3517  (.A(g4969), .Z(g5191) ) ;
INV     gate3518  (.A(g4841), .Z(g5192) ) ;
INV     gate3519  (.A(g4938), .Z(g5197) ) ;
INV     gate3520  (.A(g4969), .Z(g5198) ) ;
INV     gate3521  (.A(g4841), .Z(g5199) ) ;
INV     gate3522  (.A(g4938), .Z(g5206) ) ;
INV     gate3523  (.A(g4673), .Z(g5207) ) ;
INV     gate3524  (.A(g5114), .Z(g5224) ) ;
AND2    gate3525  (.A(g190), .B(g3986), .Z(g4705) ) ;
INV     gate3526  (.A(g4705), .Z(II9752) ) ;
INV     gate3527  (.A(II9752), .Z(g5240) ) ;
AND2    gate3528  (.A(g4517), .B(g1760), .Z(g4838) ) ;
INV     gate3529  (.A(g4838), .Z(II9760) ) ;
INV     gate3530  (.A(II9760), .Z(g5246) ) ;
INV     gate3531  (.A(g4678), .Z(II9774) ) ;
INV     gate3532  (.A(II9774), .Z(g5258) ) ;
INV     gate3533  (.A(g4748), .Z(g5261) ) ;
AND2    gate3534  (.A(g190), .B(g4055), .Z(g4720) ) ;
INV     gate3535  (.A(g4720), .Z(II9782) ) ;
INV     gate3536  (.A(II9782), .Z(g5266) ) ;
OR2     gate3537  (.A(g3984), .B(g2912), .Z(g4747) ) ;
INV     gate3538  (.A(g4747), .Z(II9785) ) ;
INV     gate3539  (.A(II9785), .Z(g5267) ) ;
AND2    gate3540  (.A(g190), .B(g4072), .Z(g4711) ) ;
INV     gate3541  (.A(g4711), .Z(II9788) ) ;
INV     gate3542  (.A(II9788), .Z(g5268) ) ;
AND2    gate3543  (.A(g4176), .B(g1760), .Z(g4779) ) ;
INV     gate3544  (.A(g4779), .Z(II9791) ) ;
INV     gate3545  (.A(II9791), .Z(g5269) ) ;
AND2    gate3546  (.A(g4169), .B(g1760), .Z(g4778) ) ;
INV     gate3547  (.A(g4778), .Z(II9794) ) ;
INV     gate3548  (.A(II9794), .Z(g5278) ) ;
INV     gate3549  (.A(g4841), .Z(g5285) ) ;
NAND3   gate3550  (.A(g4344), .B(g4335), .C(g4328), .Z(g4714) ) ;
INV     gate3551  (.A(g4714), .Z(g5286) ) ;
INV     gate3552  (.A(g5087), .Z(g5294) ) ;
INV     gate3553  (.A(g5113), .Z(II9804) ) ;
INV     gate3554  (.A(II9804), .Z(g5299) ) ;
INV     gate3555  (.A(g5028), .Z(g5302) ) ;
INV     gate3556  (.A(g4969), .Z(g5309) ) ;
INV     gate3557  (.A(g4938), .Z(g5311) ) ;
INV     gate3558  (.A(g4677), .Z(g5335) ) ;
AND2    gate3559  (.A(g4219), .B(g1690), .Z(g4691) ) ;
INV     gate3560  (.A(g4691), .Z(II9819) ) ;
INV     gate3561  (.A(II9819), .Z(g5344) ) ;
OR2     gate3562  (.A(g4108), .B(g3049), .Z(g5138) ) ;
INV     gate3563  (.A(g5138), .Z(II9823) ) ;
INV     gate3564  (.A(II9823), .Z(g5362) ) ;
INV     gate3565  (.A(g5124), .Z(g5364) ) ;
AND2    gate3566  (.A(g4187), .B(g1760), .Z(g4782) ) ;
INV     gate3567  (.A(g4782), .Z(II9834) ) ;
INV     gate3568  (.A(II9834), .Z(g5367) ) ;
AND2    gate3569  (.A(g4182), .B(g1760), .Z(g4781) ) ;
INV     gate3570  (.A(g4781), .Z(II9837) ) ;
INV     gate3571  (.A(II9837), .Z(g5384) ) ;
AND2    gate3572  (.A(g4243), .B(g1690), .Z(g4702) ) ;
INV     gate3573  (.A(g4702), .Z(II9840) ) ;
INV     gate3574  (.A(II9840), .Z(g5395) ) ;
INV     gate3575  (.A(g4692), .Z(g5396) ) ;
INV     gate3576  (.A(g5076), .Z(g5397) ) ;
AND2    gate3577  (.A(g190), .B(g4179), .Z(g4728) ) ;
INV     gate3578  (.A(g4728), .Z(II9845) ) ;
INV     gate3579  (.A(II9845), .Z(g5401) ) ;
INV     gate3580  (.A(g5000), .Z(g5402) ) ;
INV     gate3581  (.A(g5088), .Z(g5403) ) ;
AND2    gate3582  (.A(g4216), .B(g1760), .Z(g4798) ) ;
INV     gate3583  (.A(g4798), .Z(II9850) ) ;
INV     gate3584  (.A(II9850), .Z(g5412) ) ;
INV     gate3585  (.A(g5006), .Z(g5417) ) ;
INV     gate3586  (.A(g5100), .Z(g5418) ) ;
INV     gate3587  (.A(g5013), .Z(g5426) ) ;
INV     gate3588  (.A(g5115), .Z(g5427) ) ;
INV     gate3589  (.A(g5024), .Z(g5433) ) ;
INV     gate3590  (.A(g5112), .Z(g5434) ) ;
INV     gate3591  (.A(g5121), .Z(g5435) ) ;
INV     gate3592  (.A(g5041), .Z(g5437) ) ;
INV     gate3593  (.A(g5058), .Z(g5439) ) ;
INV     gate3594  (.A(g5074), .Z(g5444) ) ;
INV     gate3595  (.A(g5059), .Z(g5445) ) ;
INV     gate3596  (.A(g5137), .Z(g5448) ) ;
INV     gate3597  (.A(g4680), .Z(g5453) ) ;
INV     gate3598  (.A(g4882), .Z(g5459) ) ;
INV     gate3599  (.A(g4684), .Z(g5460) ) ;
INV     gate3600  (.A(g4885), .Z(g5461) ) ;
INV     gate3601  (.A(g4886), .Z(g5462) ) ;
INV     gate3602  (.A(g5085), .Z(g5463) ) ;
INV     gate3603  (.A(g4890), .Z(g5466) ) ;
INV     gate3604  (.A(g4891), .Z(g5467) ) ;
AND2    gate3605  (.A(g4227), .B(g4160), .Z(g4868) ) ;
INV     gate3606  (.A(g4868), .Z(II9884) ) ;
INV     gate3607  (.A(II9884), .Z(g5468) ) ;
INV     gate3608  (.A(g4898), .Z(g5469) ) ;
INV     gate3609  (.A(g4899), .Z(g5470) ) ;
AND3    gate3610  (.A(g2573), .B(g2562), .C(II9166), .Z(g4819) ) ;
INV     gate3611  (.A(g4819), .Z(II9889) ) ;
INV     gate3612  (.A(II9889), .Z(g5471) ) ;
NAND4   gate3613  (.A(g2595), .B(g2584), .C(g4270), .D(g4281), .Z(g4879) ) ;
INV     gate3614  (.A(g4879), .Z(II9892) ) ;
INV     gate3615  (.A(II9892), .Z(g5472) ) ;
INV     gate3616  (.A(g4903), .Z(g5473) ) ;
INV     gate3617  (.A(g4904), .Z(g5474) ) ;
INV     gate3618  (.A(g4907), .Z(g5476) ) ;
INV     gate3619  (.A(g4908), .Z(g5477) ) ;
INV     gate3620  (.A(g5025), .Z(g5478) ) ;
INV     gate3621  (.A(g4913), .Z(g5480) ) ;
INV     gate3622  (.A(g4914), .Z(g5481) ) ;
INV     gate3623  (.A(g4915), .Z(g5482) ) ;
AND3    gate3624  (.A(g2573), .B(g2562), .C(II9202), .Z(g4837) ) ;
INV     gate3625  (.A(g4837), .Z(II9907) ) ;
INV     gate3626  (.A(II9907), .Z(g5487) ) ;
AND2    gate3627  (.A(g4255), .B(g3533), .Z(g4681) ) ;
INV     gate3628  (.A(g4681), .Z(II9910) ) ;
INV     gate3629  (.A(II9910), .Z(g5488) ) ;
INV     gate3630  (.A(g4917), .Z(g5490) ) ;
INV     gate3631  (.A(g4918), .Z(g5491) ) ;
INV     gate3632  (.A(g4919), .Z(g5492) ) ;
INV     gate3633  (.A(g4920), .Z(g5493) ) ;
AND2    gate3634  (.A(g4403), .B(g1760), .Z(g4968) ) ;
INV     gate3635  (.A(g4968), .Z(II9918) ) ;
INV     gate3636  (.A(II9918), .Z(g5494) ) ;
INV     gate3637  (.A(g4922), .Z(g5514) ) ;
INV     gate3638  (.A(g4923), .Z(g5515) ) ;
INV     gate3639  (.A(g4924), .Z(g5516) ) ;
INV     gate3640  (.A(g4925), .Z(g5517) ) ;
OR2     gate3641  (.A(g4049), .B(g4054), .Z(g5052) ) ;
INV     gate3642  (.A(g5052), .Z(II9929) ) ;
INV     gate3643  (.A(II9929), .Z(g5519) ) ;
INV     gate3644  (.A(g4928), .Z(g5520) ) ;
INV     gate3645  (.A(g4929), .Z(g5521) ) ;
INV     gate3646  (.A(g4930), .Z(g5522) ) ;
OR2     gate3647  (.A(g2490), .B(g4237), .Z(g4812) ) ;
INV     gate3648  (.A(g4812), .Z(II9935) ) ;
INV     gate3649  (.A(II9935), .Z(g5523) ) ;
AND3    gate3650  (.A(g2573), .B(g2562), .C(II9222), .Z(g4878) ) ;
INV     gate3651  (.A(g4878), .Z(II9938) ) ;
INV     gate3652  (.A(II9938), .Z(g5524) ) ;
INV     gate3653  (.A(g4934), .Z(g5525) ) ;
INV     gate3654  (.A(g5086), .Z(g5526) ) ;
INV     gate3655  (.A(g4689), .Z(g5529) ) ;
AND2    gate3656  (.A(g150), .B(g4265), .Z(g4814) ) ;
INV     gate3657  (.A(g4814), .Z(g5541) ) ;
INV     gate3658  (.A(g5061), .Z(g5542) ) ;
NOR2    gate3659  (.A(g3885), .B(g3094), .Z(g4676) ) ;
INV     gate3660  (.A(g4676), .Z(II9974) ) ;
INV     gate3661  (.A(II9974), .Z(g5551) ) ;
AND2    gate3662  (.A(g4228), .B(g1964), .Z(g4825) ) ;
INV     gate3663  (.A(g4825), .Z(II10028) ) ;
INV     gate3664  (.A(II10028), .Z(g5569) ) ;
INV     gate3665  (.A(g1236), .Z(II10032) ) ;
INV     gate3666  (.A(g4969), .Z(g5574) ) ;
AND2    gate3667  (.A(g4235), .B(g1980), .Z(g4840) ) ;
INV     gate3668  (.A(g4840), .Z(II10046) ) ;
INV     gate3669  (.A(II10046), .Z(g5577) ) ;
INV     gate3670  (.A(g4841), .Z(g5578) ) ;
INV     gate3671  (.A(g4938), .Z(g5580) ) ;
INV     gate3672  (.A(g4969), .Z(g5581) ) ;
INV     gate3673  (.A(g4969), .Z(g5582) ) ;
INV     gate3674  (.A(g4841), .Z(g5584) ) ;
INV     gate3675  (.A(g4938), .Z(g5586) ) ;
INV     gate3676  (.A(g4938), .Z(g5587) ) ;
INV     gate3677  (.A(g4841), .Z(g5591) ) ;
INV     gate3678  (.A(g4969), .Z(g5592) ) ;
INV     gate3679  (.A(g4841), .Z(g5596) ) ;
INV     gate3680  (.A(g4969), .Z(g5597) ) ;
INV     gate3681  (.A(g4938), .Z(g5598) ) ;
INV     gate3682  (.A(g5128), .Z(g5600) ) ;
INV     gate3683  (.A(g4938), .Z(g5603) ) ;
INV     gate3684  (.A(g4969), .Z(g5604) ) ;
INV     gate3685  (.A(g4748), .Z(g5606) ) ;
INV     gate3686  (.A(g4938), .Z(g5607) ) ;
INV     gate3687  (.A(g4969), .Z(g5608) ) ;
INV     gate3688  (.A(g4748), .Z(g5609) ) ;
INV     gate3689  (.A(g4938), .Z(g5610) ) ;
INV     gate3690  (.A(g4969), .Z(g5611) ) ;
INV     gate3691  (.A(g4814), .Z(g5612) ) ;
INV     gate3692  (.A(g4748), .Z(g5613) ) ;
INV     gate3693  (.A(g4938), .Z(g5616) ) ;
INV     gate3694  (.A(g4969), .Z(g5617) ) ;
INV     gate3695  (.A(g5015), .Z(g5618) ) ;
INV     gate3696  (.A(g4748), .Z(g5621) ) ;
INV     gate3697  (.A(g4938), .Z(g5622) ) ;
INV     gate3698  (.A(g4969), .Z(g5623) ) ;
INV     gate3699  (.A(g4748), .Z(g5626) ) ;
INV     gate3700  (.A(g4673), .Z(g5627) ) ;
INV     gate3701  (.A(g4748), .Z(g5628) ) ;
INV     gate3702  (.A(g4938), .Z(g5631) ) ;
INV     gate3703  (.A(g4895), .Z(g5633) ) ;
INV     gate3704  (.A(g4748), .Z(g5638) ) ;
INV     gate3705  (.A(g4748), .Z(g5639) ) ;
INV     gate3706  (.A(g5127), .Z(II10125) ) ;
INV     gate3707  (.A(II10125), .Z(g5642) ) ;
OR2     gate3708  (.A(g4193), .B(g3190), .Z(g4688) ) ;
INV     gate3709  (.A(g4688), .Z(II10128) ) ;
INV     gate3710  (.A(II10128), .Z(g5643) ) ;
INV     gate3711  (.A(g4748), .Z(g5644) ) ;
INV     gate3712  (.A(g4748), .Z(g5645) ) ;
INV     gate3713  (.A(g4748), .Z(g5648) ) ;
INV     gate3714  (.A(g4748), .Z(g5649) ) ;
INV     gate3715  (.A(g4960), .Z(II10135) ) ;
INV     gate3716  (.A(II10135), .Z(g5652) ) ;
INV     gate3717  (.A(g4748), .Z(g5653) ) ;
INV     gate3718  (.A(g4748), .Z(g5654) ) ;
INV     gate3719  (.A(g4748), .Z(g5658) ) ;
INV     gate3720  (.A(g5027), .Z(g5662) ) ;
INV     gate3721  (.A(g4748), .Z(g5665) ) ;
INV     gate3722  (.A(g5007), .Z(II10151) ) ;
INV     gate3723  (.A(II10151), .Z(g5668) ) ;
INV     gate3724  (.A(g5109), .Z(II10154) ) ;
INV     gate3725  (.A(g5109), .Z(II10157) ) ;
INV     gate3726  (.A(II10157), .Z(g5670) ) ;
INV     gate3727  (.A(g5139), .Z(II10160) ) ;
INV     gate3728  (.A(II10160), .Z(g5671) ) ;
INV     gate3729  (.A(g5042), .Z(g5674) ) ;
INV     gate3730  (.A(g5016), .Z(II10166) ) ;
INV     gate3731  (.A(II10166), .Z(g5677) ) ;
INV     gate3732  (.A(g4873), .Z(II10169) ) ;
INV     gate3733  (.A(g4873), .Z(II10172) ) ;
INV     gate3734  (.A(II10172), .Z(g5679) ) ;
INV     gate3735  (.A(g5101), .Z(g5680) ) ;
INV     gate3736  (.A(g4721), .Z(II10177) ) ;
INV     gate3737  (.A(g4721), .Z(II10180) ) ;
INV     gate3738  (.A(II10180), .Z(g5683) ) ;
INV     gate3739  (.A(g5129), .Z(II10183) ) ;
INV     gate3740  (.A(g5129), .Z(II10186) ) ;
INV     gate3741  (.A(II10186), .Z(g5685) ) ;
INV     gate3742  (.A(g4670), .Z(II10190) ) ;
INV     gate3743  (.A(g4670), .Z(II10193) ) ;
INV     gate3744  (.A(II10193), .Z(g5688) ) ;
INV     gate3745  (.A(g4748), .Z(g5690) ) ;
INV     gate3746  (.A(g5060), .Z(II10204) ) ;
INV     gate3747  (.A(II10204), .Z(g5693) ) ;
INV     gate3748  (.A(g5075), .Z(II10207) ) ;
INV     gate3749  (.A(II10207), .Z(g5696) ) ;
INV     gate3750  (.A(g5120), .Z(g5701) ) ;
INV     gate3751  (.A(g4841), .Z(g5705) ) ;
INV     gate3752  (.A(g4841), .Z(g5709) ) ;
INV     gate3753  (.A(g4841), .Z(g5713) ) ;
INV     gate3754  (.A(g4969), .Z(g5717) ) ;
INV     gate3755  (.A(g4841), .Z(g5718) ) ;
INV     gate3756  (.A(g5014), .Z(II10236) ) ;
INV     gate3757  (.A(II10236), .Z(g5719) ) ;
INV     gate3758  (.A(g4938), .Z(g5723) ) ;
INV     gate3759  (.A(g4969), .Z(g5724) ) ;
INV     gate3760  (.A(g4841), .Z(g5725) ) ;
INV     gate3761  (.A(g5026), .Z(II10243) ) ;
INV     gate3762  (.A(II10243), .Z(g5726) ) ;
INV     gate3763  (.A(g5266), .Z(II10247) ) ;
INV     gate3764  (.A(g5268), .Z(II10250) ) ;
INV     gate3765  (.A(g5240), .Z(II10253) ) ;
INV     gate3766  (.A(g5401), .Z(II10256) ) ;
INV     gate3767  (.A(g5362), .Z(II10259) ) ;
INV     gate3768  (.A(g5551), .Z(II10262) ) ;
INV     gate3769  (.A(g5468), .Z(II10265) ) ;
INV     gate3770  (.A(g5471), .Z(II10268) ) ;
INV     gate3771  (.A(g5487), .Z(II10271) ) ;
INV     gate3772  (.A(g5524), .Z(II10274) ) ;
INV     gate3773  (.A(g5472), .Z(II10277) ) ;
INV     gate3774  (.A(g5488), .Z(II10280) ) ;
INV     gate3775  (.A(g5643), .Z(II10283) ) ;
INV     gate3776  (.A(g5519), .Z(II10286) ) ;
INV     gate3777  (.A(g5569), .Z(II10289) ) ;
INV     gate3778  (.A(g5577), .Z(II10292) ) ;
INV     gate3779  (.A(g5523), .Z(II10295) ) ;
INV     gate3780  (.A(g5207), .Z(g5749) ) ;
INV     gate3781  (.A(g5403), .Z(g5754) ) ;
INV     gate3782  (.A(g5494), .Z(g5755) ) ;
OR2     gate3783  (.A(g4936), .B(g4334), .Z(g5704) ) ;
INV     gate3784  (.A(g5704), .Z(II10343) ) ;
INV     gate3785  (.A(II10343), .Z(g5756) ) ;
INV     gate3786  (.A(g5261), .Z(g5757) ) ;
OR2     gate3787  (.A(g4955), .B(g4342), .Z(g5706) ) ;
INV     gate3788  (.A(g5706), .Z(II10347) ) ;
INV     gate3789  (.A(II10347), .Z(g5758) ) ;
OR2     gate3790  (.A(g4956), .B(g4343), .Z(g5707) ) ;
INV     gate3791  (.A(g5707), .Z(II10350) ) ;
INV     gate3792  (.A(II10350), .Z(g5759) ) ;
OR2     gate3793  (.A(g4958), .B(g4351), .Z(g5710) ) ;
INV     gate3794  (.A(g5710), .Z(II10353) ) ;
INV     gate3795  (.A(II10353), .Z(g5760) ) ;
OR2     gate3796  (.A(g4959), .B(g4352), .Z(g5711) ) ;
INV     gate3797  (.A(g5711), .Z(II10356) ) ;
INV     gate3798  (.A(II10356), .Z(g5761) ) ;
OR2     gate3799  (.A(g4961), .B(g4355), .Z(g5715) ) ;
INV     gate3800  (.A(g5715), .Z(II10366) ) ;
INV     gate3801  (.A(II10366), .Z(g5763) ) ;
OR2     gate3802  (.A(g4962), .B(g4356), .Z(g5716) ) ;
INV     gate3803  (.A(g5716), .Z(II10369) ) ;
INV     gate3804  (.A(II10369), .Z(g5764) ) ;
OR2     gate3805  (.A(g5001), .B(g4361), .Z(g5722) ) ;
INV     gate3806  (.A(g5722), .Z(II10373) ) ;
INV     gate3807  (.A(II10373), .Z(g5766) ) ;
OR2     gate3808  (.A(g5008), .B(g4365), .Z(g5188) ) ;
INV     gate3809  (.A(g5188), .Z(II10377) ) ;
INV     gate3810  (.A(II10377), .Z(g5768) ) ;
INV     gate3811  (.A(g5448), .Z(II10380) ) ;
INV     gate3812  (.A(II10380), .Z(g5769) ) ;
OR2     gate3813  (.A(g5017), .B(g4366), .Z(g5193) ) ;
INV     gate3814  (.A(g5193), .Z(II10384) ) ;
INV     gate3815  (.A(II10384), .Z(g5779) ) ;
OR2     gate3816  (.A(g5018), .B(g4367), .Z(g5194) ) ;
INV     gate3817  (.A(g5194), .Z(II10387) ) ;
INV     gate3818  (.A(II10387), .Z(g5780) ) ;
OR2     gate3819  (.A(g5019), .B(g4368), .Z(g5195) ) ;
INV     gate3820  (.A(g5195), .Z(II10390) ) ;
INV     gate3821  (.A(II10390), .Z(g5781) ) ;
OR2     gate3822  (.A(g5020), .B(g4369), .Z(g5196) ) ;
INV     gate3823  (.A(g5196), .Z(II10393) ) ;
INV     gate3824  (.A(II10393), .Z(g5782) ) ;
OR2     gate3825  (.A(g5029), .B(g4375), .Z(g5200) ) ;
INV     gate3826  (.A(g5200), .Z(II10397) ) ;
INV     gate3827  (.A(II10397), .Z(g5784) ) ;
OR2     gate3828  (.A(g5030), .B(g4376), .Z(g5201) ) ;
INV     gate3829  (.A(g5201), .Z(II10400) ) ;
INV     gate3830  (.A(II10400), .Z(g5785) ) ;
OR2     gate3831  (.A(g5031), .B(g4377), .Z(g5202) ) ;
INV     gate3832  (.A(g5202), .Z(II10403) ) ;
INV     gate3833  (.A(II10403), .Z(g5786) ) ;
OR2     gate3834  (.A(g5032), .B(g4378), .Z(g5203) ) ;
INV     gate3835  (.A(g5203), .Z(II10406) ) ;
INV     gate3836  (.A(II10406), .Z(g5787) ) ;
OR2     gate3837  (.A(g5033), .B(g4379), .Z(g5204) ) ;
INV     gate3838  (.A(g5204), .Z(II10409) ) ;
INV     gate3839  (.A(II10409), .Z(g5788) ) ;
OR2     gate3840  (.A(g5034), .B(g4380), .Z(g5205) ) ;
INV     gate3841  (.A(g5205), .Z(II10412) ) ;
INV     gate3842  (.A(II10412), .Z(g5789) ) ;
INV     gate3843  (.A(g5397), .Z(II10415) ) ;
INV     gate3844  (.A(II10415), .Z(g5790) ) ;
INV     gate3845  (.A(g5453), .Z(II10418) ) ;
INV     gate3846  (.A(II10418), .Z(g5793) ) ;
OR2     gate3847  (.A(g5043), .B(g4383), .Z(g5208) ) ;
INV     gate3848  (.A(g5208), .Z(II10421) ) ;
INV     gate3849  (.A(II10421), .Z(g5794) ) ;
OR2     gate3850  (.A(g5044), .B(g4384), .Z(g5209) ) ;
INV     gate3851  (.A(g5209), .Z(II10424) ) ;
INV     gate3852  (.A(II10424), .Z(g5795) ) ;
OR2     gate3853  (.A(g5045), .B(g4385), .Z(g5210) ) ;
INV     gate3854  (.A(g5210), .Z(II10427) ) ;
INV     gate3855  (.A(II10427), .Z(g5796) ) ;
OR2     gate3856  (.A(g5046), .B(g4386), .Z(g5211) ) ;
INV     gate3857  (.A(g5211), .Z(II10430) ) ;
INV     gate3858  (.A(II10430), .Z(g5797) ) ;
OR2     gate3859  (.A(g5047), .B(g4387), .Z(g5212) ) ;
INV     gate3860  (.A(g5212), .Z(II10433) ) ;
INV     gate3861  (.A(II10433), .Z(g5798) ) ;
OR2     gate3862  (.A(g5048), .B(g4388), .Z(g5213) ) ;
INV     gate3863  (.A(g5213), .Z(II10436) ) ;
INV     gate3864  (.A(II10436), .Z(g5799) ) ;
OR2     gate3865  (.A(g5049), .B(g4389), .Z(g5214) ) ;
INV     gate3866  (.A(g5214), .Z(II10439) ) ;
INV     gate3867  (.A(II10439), .Z(g5800) ) ;
OR2     gate3868  (.A(g5050), .B(g4390), .Z(g5215) ) ;
INV     gate3869  (.A(g5215), .Z(II10442) ) ;
INV     gate3870  (.A(II10442), .Z(g5801) ) ;
INV     gate3871  (.A(g5418), .Z(II10445) ) ;
INV     gate3872  (.A(II10445), .Z(g5802) ) ;
INV     gate3873  (.A(g5335), .Z(II10448) ) ;
INV     gate3874  (.A(II10448), .Z(g5805) ) ;
OR2     gate3875  (.A(g5062), .B(g4391), .Z(g5216) ) ;
INV     gate3876  (.A(g5216), .Z(II10451) ) ;
INV     gate3877  (.A(II10451), .Z(g5806) ) ;
OR2     gate3878  (.A(g5063), .B(g4392), .Z(g5217) ) ;
INV     gate3879  (.A(g5217), .Z(II10454) ) ;
INV     gate3880  (.A(II10454), .Z(g5807) ) ;
OR2     gate3881  (.A(g5064), .B(g4393), .Z(g5218) ) ;
INV     gate3882  (.A(g5218), .Z(II10457) ) ;
INV     gate3883  (.A(II10457), .Z(g5808) ) ;
OR2     gate3884  (.A(g5065), .B(g4394), .Z(g5219) ) ;
INV     gate3885  (.A(g5219), .Z(II10460) ) ;
INV     gate3886  (.A(II10460), .Z(g5809) ) ;
OR2     gate3887  (.A(g5066), .B(g4395), .Z(g5220) ) ;
INV     gate3888  (.A(g5220), .Z(II10463) ) ;
INV     gate3889  (.A(II10463), .Z(g5810) ) ;
OR2     gate3890  (.A(g5067), .B(g4396), .Z(g5221) ) ;
INV     gate3891  (.A(g5221), .Z(II10466) ) ;
INV     gate3892  (.A(II10466), .Z(g5811) ) ;
OR2     gate3893  (.A(g5068), .B(g4397), .Z(g5222) ) ;
INV     gate3894  (.A(g5222), .Z(II10469) ) ;
INV     gate3895  (.A(II10469), .Z(g5812) ) ;
OR2     gate3896  (.A(g5069), .B(g4398), .Z(g5223) ) ;
INV     gate3897  (.A(g5223), .Z(II10472) ) ;
INV     gate3898  (.A(II10472), .Z(g5813) ) ;
INV     gate3899  (.A(g5529), .Z(II10475) ) ;
INV     gate3900  (.A(II10475), .Z(g5814) ) ;
OR2     gate3901  (.A(g5077), .B(g4407), .Z(g5227) ) ;
INV     gate3902  (.A(g5227), .Z(II10479) ) ;
INV     gate3903  (.A(II10479), .Z(g5818) ) ;
OR2     gate3904  (.A(g5078), .B(g4408), .Z(g5228) ) ;
INV     gate3905  (.A(g5228), .Z(II10482) ) ;
INV     gate3906  (.A(II10482), .Z(g5819) ) ;
OR2     gate3907  (.A(g5079), .B(g4409), .Z(g5229) ) ;
INV     gate3908  (.A(g5229), .Z(II10485) ) ;
INV     gate3909  (.A(II10485), .Z(g5820) ) ;
OR2     gate3910  (.A(g5080), .B(g4410), .Z(g5230) ) ;
INV     gate3911  (.A(g5230), .Z(II10488) ) ;
INV     gate3912  (.A(II10488), .Z(g5821) ) ;
OR2     gate3913  (.A(g5081), .B(g4411), .Z(g5231) ) ;
INV     gate3914  (.A(g5231), .Z(II10491) ) ;
INV     gate3915  (.A(II10491), .Z(g5822) ) ;
OR2     gate3916  (.A(g5082), .B(g4412), .Z(g5232) ) ;
INV     gate3917  (.A(g5232), .Z(II10494) ) ;
INV     gate3918  (.A(II10494), .Z(g5823) ) ;
OR2     gate3919  (.A(g5089), .B(g4420), .Z(g5233) ) ;
INV     gate3920  (.A(g5233), .Z(II10497) ) ;
INV     gate3921  (.A(II10497), .Z(g5824) ) ;
OR2     gate3922  (.A(g5090), .B(g4421), .Z(g5234) ) ;
INV     gate3923  (.A(g5234), .Z(II10500) ) ;
INV     gate3924  (.A(II10500), .Z(g5825) ) ;
OR2     gate3925  (.A(g5091), .B(g4422), .Z(g5235) ) ;
INV     gate3926  (.A(g5235), .Z(II10503) ) ;
INV     gate3927  (.A(II10503), .Z(g5826) ) ;
OR2     gate3928  (.A(g5092), .B(g4423), .Z(g5236) ) ;
INV     gate3929  (.A(g5236), .Z(II10506) ) ;
INV     gate3930  (.A(II10506), .Z(g5827) ) ;
OR2     gate3931  (.A(g5093), .B(g4424), .Z(g5237) ) ;
INV     gate3932  (.A(g5237), .Z(II10509) ) ;
INV     gate3933  (.A(II10509), .Z(g5828) ) ;
OR2     gate3934  (.A(g5094), .B(g4425), .Z(g5238) ) ;
INV     gate3935  (.A(g5238), .Z(II10512) ) ;
INV     gate3936  (.A(II10512), .Z(g5829) ) ;
OR2     gate3937  (.A(g5104), .B(g4433), .Z(g5241) ) ;
INV     gate3938  (.A(g5241), .Z(II10516) ) ;
INV     gate3939  (.A(II10516), .Z(g5831) ) ;
OR2     gate3940  (.A(g5105), .B(g4434), .Z(g5242) ) ;
INV     gate3941  (.A(g5242), .Z(II10519) ) ;
INV     gate3942  (.A(II10519), .Z(g5832) ) ;
OR2     gate3943  (.A(g5106), .B(g4435), .Z(g5243) ) ;
INV     gate3944  (.A(g5243), .Z(II10522) ) ;
INV     gate3945  (.A(II10522), .Z(g5833) ) ;
OR2     gate3946  (.A(g5107), .B(g4436), .Z(g5244) ) ;
INV     gate3947  (.A(g5244), .Z(II10525) ) ;
INV     gate3948  (.A(II10525), .Z(g5834) ) ;
OR2     gate3949  (.A(g5108), .B(g4437), .Z(g5245) ) ;
INV     gate3950  (.A(g5245), .Z(II10528) ) ;
INV     gate3951  (.A(II10528), .Z(g5835) ) ;
INV     gate3952  (.A(g5529), .Z(g5836) ) ;
OR2     gate3953  (.A(g5116), .B(g4451), .Z(g5253) ) ;
INV     gate3954  (.A(g5253), .Z(II10532) ) ;
INV     gate3955  (.A(II10532), .Z(g5839) ) ;
OR2     gate3956  (.A(g5117), .B(g4452), .Z(g5254) ) ;
INV     gate3957  (.A(g5254), .Z(II10535) ) ;
INV     gate3958  (.A(II10535), .Z(g5840) ) ;
OR2     gate3959  (.A(g5118), .B(g4453), .Z(g5255) ) ;
INV     gate3960  (.A(g5255), .Z(II10538) ) ;
INV     gate3961  (.A(II10538), .Z(g5841) ) ;
OR2     gate3962  (.A(g5119), .B(g4454), .Z(g5256) ) ;
INV     gate3963  (.A(g5256), .Z(II10541) ) ;
INV     gate3964  (.A(II10541), .Z(g5842) ) ;
INV     gate3965  (.A(g5367), .Z(g5843) ) ;
OR2     gate3966  (.A(g5122), .B(g4472), .Z(g5259) ) ;
INV     gate3967  (.A(g5259), .Z(II10545) ) ;
INV     gate3968  (.A(II10545), .Z(g5844) ) ;
OR2     gate3969  (.A(g5123), .B(g4473), .Z(g5260) ) ;
INV     gate3970  (.A(g5260), .Z(II10548) ) ;
INV     gate3971  (.A(II10548), .Z(g5845) ) ;
INV     gate3972  (.A(g5367), .Z(g5846) ) ;
INV     gate3973  (.A(g5396), .Z(II10552) ) ;
INV     gate3974  (.A(II10552), .Z(g5847) ) ;
INV     gate3975  (.A(g5529), .Z(II10555) ) ;
INV     gate3976  (.A(II10555), .Z(g5868) ) ;
OR2     gate3977  (.A(g5125), .B(g4490), .Z(g5264) ) ;
INV     gate3978  (.A(g5264), .Z(II10558) ) ;
INV     gate3979  (.A(II10558), .Z(g5871) ) ;
OR2     gate3980  (.A(g5126), .B(g4491), .Z(g5265) ) ;
INV     gate3981  (.A(g5265), .Z(II10561) ) ;
INV     gate3982  (.A(II10561), .Z(g5872) ) ;
INV     gate3983  (.A(g5367), .Z(g5873) ) ;
INV     gate3984  (.A(g5402), .Z(II10565) ) ;
INV     gate3985  (.A(II10565), .Z(g5874) ) ;
INV     gate3986  (.A(g5417), .Z(II10569) ) ;
INV     gate3987  (.A(II10569), .Z(g5897) ) ;
INV     gate3988  (.A(g5384), .Z(g5916) ) ;
INV     gate3989  (.A(g5412), .Z(g5917) ) ;
INV     gate3990  (.A(g5426), .Z(II10574) ) ;
INV     gate3991  (.A(II10574), .Z(g5918) ) ;
INV     gate3992  (.A(g5412), .Z(g5938) ) ;
INV     gate3993  (.A(g5433), .Z(II10579) ) ;
INV     gate3994  (.A(II10579), .Z(g5939) ) ;
INV     gate3995  (.A(g5437), .Z(II10582) ) ;
INV     gate3996  (.A(II10582), .Z(g5956) ) ;
INV     gate3997  (.A(g5439), .Z(II10587) ) ;
INV     gate3998  (.A(II10587), .Z(g5971) ) ;
INV     gate3999  (.A(g5294), .Z(g5987) ) ;
INV     gate4000  (.A(g5444), .Z(II10592) ) ;
INV     gate4001  (.A(II10592), .Z(g5988) ) ;
INV     gate4002  (.A(g5494), .Z(g6004) ) ;
INV     gate4003  (.A(g5494), .Z(g6007) ) ;
INV     gate4004  (.A(g5367), .Z(g6008) ) ;
OR2     gate4005  (.A(g4790), .B(g4786), .Z(g5440) ) ;
INV     gate4006  (.A(g5440), .Z(II10605) ) ;
INV     gate4007  (.A(II10605), .Z(g6009) ) ;
INV     gate4008  (.A(g5701), .Z(II10608) ) ;
INV     gate4009  (.A(II10608), .Z(g6010) ) ;
INV     gate4010  (.A(g5494), .Z(g6011) ) ;
INV     gate4011  (.A(g5367), .Z(g6012) ) ;
INV     gate4012  (.A(g5302), .Z(II10614) ) ;
INV     gate4013  (.A(II10614), .Z(g6014) ) ;
INV     gate4014  (.A(g5677), .Z(II10617) ) ;
INV     gate4015  (.A(II10617), .Z(g6015) ) ;
INV     gate4016  (.A(g5494), .Z(g6018) ) ;
INV     gate4017  (.A(g5367), .Z(g6019) ) ;
INV     gate4018  (.A(g5367), .Z(g6020) ) ;
INV     gate4019  (.A(g5494), .Z(g6024) ) ;
INV     gate4020  (.A(g5367), .Z(g6025) ) ;
INV     gate4021  (.A(g5384), .Z(g6026) ) ;
INV     gate4022  (.A(g5384), .Z(g6027) ) ;
INV     gate4023  (.A(g5529), .Z(g6028) ) ;
INV     gate4024  (.A(g5494), .Z(g6032) ) ;
INV     gate4025  (.A(g5384), .Z(g6033) ) ;
INV     gate4026  (.A(g5224), .Z(II10639) ) ;
INV     gate4027  (.A(II10639), .Z(g6034) ) ;
INV     gate4028  (.A(g5494), .Z(g6035) ) ;
INV     gate4029  (.A(g5267), .Z(II10643) ) ;
INV     gate4030  (.A(II10643), .Z(g6036) ) ;
INV     gate4031  (.A(g5364), .Z(II10646) ) ;
INV     gate4032  (.A(II10646), .Z(g6037) ) ;
NAND2   gate4033  (.A(g5021), .B(g4381), .Z(g5657) ) ;
INV     gate4034  (.A(g5657), .Z(II10649) ) ;
INV     gate4035  (.A(II10649), .Z(g6038) ) ;
INV     gate4036  (.A(g5246), .Z(g6048) ) ;
INV     gate4037  (.A(g5246), .Z(g6050) ) ;
INV     gate4038  (.A(g5246), .Z(g6051) ) ;
OR3     gate4039  (.A(g4727), .B(g4737), .C(g4735), .Z(g5317) ) ;
INV     gate4040  (.A(g5317), .Z(g6059) ) ;
INV     gate4041  (.A(g5662), .Z(II10675) ) ;
INV     gate4042  (.A(II10675), .Z(g6062) ) ;
OR2     gate4043  (.A(g3617), .B(g4810), .Z(g5566) ) ;
INV     gate4044  (.A(g5566), .Z(II10678) ) ;
INV     gate4045  (.A(II10678), .Z(g6063) ) ;
NAND2   gate4046  (.A(g5132), .B(g1263), .Z(g5686) ) ;
INV     gate4047  (.A(g5686), .Z(II10681) ) ;
INV     gate4048  (.A(II10681), .Z(g6064) ) ;
INV     gate4049  (.A(g5258), .Z(II10684) ) ;
INV     gate4050  (.A(II10684), .Z(g6065) ) ;
INV     gate4051  (.A(g5674), .Z(II10687) ) ;
INV     gate4052  (.A(II10687), .Z(g6068) ) ;
NAND2   gate4053  (.A(g5132), .B(g1266), .Z(g5538) ) ;
INV     gate4054  (.A(g5538), .Z(II10690) ) ;
INV     gate4055  (.A(II10690), .Z(g6069) ) ;
INV     gate4056  (.A(g5317), .Z(g6070) ) ;
INV     gate4057  (.A(g5445), .Z(II10694) ) ;
INV     gate4058  (.A(II10694), .Z(g6071) ) ;
OR2     gate4059  (.A(g4736), .B(g4734), .Z(g5345) ) ;
INV     gate4060  (.A(g5345), .Z(g6072) ) ;
INV     gate4061  (.A(g5384), .Z(g6073) ) ;
INV     gate4062  (.A(g5317), .Z(g6074) ) ;
INV     gate4063  (.A(g5345), .Z(g6075) ) ;
AND2    gate4064  (.A(g786), .B(g4724), .Z(g5287) ) ;
INV     gate4065  (.A(g5287), .Z(g6076) ) ;
INV     gate4066  (.A(g5529), .Z(II10702) ) ;
INV     gate4067  (.A(II10702), .Z(g6083) ) ;
INV     gate4068  (.A(g5463), .Z(II10705) ) ;
INV     gate4069  (.A(II10705), .Z(g6087) ) ;
OR2     gate4070  (.A(g3617), .B(g4824), .Z(g5545) ) ;
INV     gate4071  (.A(g5545), .Z(II10708) ) ;
INV     gate4072  (.A(II10708), .Z(g6088) ) ;
INV     gate4073  (.A(g5317), .Z(g6089) ) ;
INV     gate4074  (.A(g5529), .Z(g6090) ) ;
INV     gate4075  (.A(g5317), .Z(g6092) ) ;
INV     gate4076  (.A(g5345), .Z(g6093) ) ;
OR2     gate4077  (.A(g3617), .B(g4835), .Z(g5537) ) ;
INV     gate4078  (.A(g5537), .Z(II10716) ) ;
INV     gate4079  (.A(II10716), .Z(g6094) ) ;
NAND2   gate4080  (.A(g5132), .B(g1257), .Z(g5559) ) ;
INV     gate4081  (.A(g5559), .Z(II10719) ) ;
INV     gate4082  (.A(II10719), .Z(g6095) ) ;
INV     gate4083  (.A(g5317), .Z(g6096) ) ;
INV     gate4084  (.A(g5345), .Z(g6097) ) ;
INV     gate4085  (.A(g5317), .Z(g6101) ) ;
INV     gate4086  (.A(g5345), .Z(g6102) ) ;
INV     gate4087  (.A(g5317), .Z(g6103) ) ;
INV     gate4088  (.A(g5345), .Z(g6104) ) ;
INV     gate4089  (.A(g5345), .Z(g6106) ) ;
INV     gate4090  (.A(g5345), .Z(g6108) ) ;
INV     gate4091  (.A(g5335), .Z(g6110) ) ;
INV     gate4092  (.A(g5453), .Z(g6111) ) ;
OR2     gate4093  (.A(g5051), .B(g1236), .Z(g5572) ) ;
INV     gate4094  (.A(g5572), .Z(II10739) ) ;
INV     gate4095  (.A(II10739), .Z(g6117) ) ;
OR2     gate4096  (.A(g2935), .B(g4712), .Z(g5549) ) ;
INV     gate4097  (.A(g5549), .Z(g6118) ) ;
INV     gate4098  (.A(g5618), .Z(II10752) ) ;
INV     gate4099  (.A(II10752), .Z(g6122) ) ;
INV     gate4100  (.A(g5662), .Z(II10758) ) ;
INV     gate4101  (.A(II10758), .Z(g6129) ) ;
INV     gate4102  (.A(g5302), .Z(II10761) ) ;
INV     gate4103  (.A(II10761), .Z(g6130) ) ;
INV     gate4104  (.A(g5529), .Z(g6131) ) ;
INV     gate4105  (.A(g5674), .Z(II10766) ) ;
INV     gate4106  (.A(II10766), .Z(g6133) ) ;
AND2    gate4107  (.A(g775), .B(g4707), .Z(g5428) ) ;
INV     gate4108  (.A(g5428), .Z(g6134) ) ;
AND2    gate4109  (.A(g4870), .B(g3497), .Z(g5441) ) ;
INV     gate4110  (.A(g5441), .Z(II10770) ) ;
INV     gate4111  (.A(II10770), .Z(g6135) ) ;
OR2     gate4112  (.A(g2889), .B(g4699), .Z(g5708) ) ;
INV     gate4113  (.A(g5708), .Z(II10773) ) ;
INV     gate4114  (.A(II10773), .Z(g6136) ) ;
NAND3   gate4115  (.A(g4894), .B(g4888), .C(g4884), .Z(g5576) ) ;
INV     gate4116  (.A(g5576), .Z(II10776) ) ;
INV     gate4117  (.A(II10776), .Z(g6137) ) ;
INV     gate4118  (.A(g5445), .Z(II10780) ) ;
INV     gate4119  (.A(II10780), .Z(g6139) ) ;
INV     gate4120  (.A(g5542), .Z(II10783) ) ;
INV     gate4121  (.A(II10783), .Z(g6140) ) ;
AND2    gate4122  (.A(g4876), .B(g3499), .Z(g5452) ) ;
INV     gate4123  (.A(g5452), .Z(II10786) ) ;
INV     gate4124  (.A(II10786), .Z(g6141) ) ;
INV     gate4125  (.A(g5397), .Z(II10796) ) ;
INV     gate4126  (.A(II10796), .Z(g6143) ) ;
INV     gate4127  (.A(g5463), .Z(II10801) ) ;
INV     gate4128  (.A(II10801), .Z(g6146) ) ;
INV     gate4129  (.A(g5526), .Z(II10804) ) ;
INV     gate4130  (.A(II10804), .Z(g6147) ) ;
INV     gate4131  (.A(g5294), .Z(II10807) ) ;
INV     gate4132  (.A(II10807), .Z(g6148) ) ;
INV     gate4133  (.A(g5403), .Z(II10810) ) ;
INV     gate4134  (.A(II10810), .Z(g6149) ) ;
INV     gate4135  (.A(g5287), .Z(g6150) ) ;
INV     gate4136  (.A(g5418), .Z(II10815) ) ;
INV     gate4137  (.A(II10815), .Z(g6152) ) ;
INV     gate4138  (.A(g5434), .Z(II10826) ) ;
INV     gate4139  (.A(II10826), .Z(g6155) ) ;
INV     gate4140  (.A(g5224), .Z(II10829) ) ;
INV     gate4141  (.A(II10829), .Z(g6156) ) ;
INV     gate4142  (.A(g5701), .Z(II10842) ) ;
INV     gate4143  (.A(II10842), .Z(g6161) ) ;
INV     gate4144  (.A(g5364), .Z(II10862) ) ;
INV     gate4145  (.A(II10862), .Z(g6167) ) ;
INV     gate4146  (.A(g5600), .Z(II10882) ) ;
INV     gate4147  (.A(II10882), .Z(g6173) ) ;
AND2    gate4148  (.A(g3801), .B(g5022), .Z(g5475) ) ;
INV     gate4149  (.A(g5475), .Z(II10896) ) ;
INV     gate4150  (.A(II10896), .Z(g6179) ) ;
INV     gate4151  (.A(g5448), .Z(II10914) ) ;
INV     gate4152  (.A(II10914), .Z(g6183) ) ;
AND2    gate4153  (.A(g5141), .B(g5037), .Z(g5479) ) ;
INV     gate4154  (.A(g5479), .Z(II10919) ) ;
INV     gate4155  (.A(II10919), .Z(g6186) ) ;
INV     gate4156  (.A(g5600), .Z(II10930) ) ;
INV     gate4157  (.A(II10930), .Z(g6189) ) ;
INV     gate4158  (.A(g5668), .Z(II10933) ) ;
INV     gate4159  (.A(II10933), .Z(g6190) ) ;
AND2    gate4160  (.A(g3390), .B(g5036), .Z(g5560) ) ;
INV     gate4161  (.A(g5560), .Z(II10937) ) ;
INV     gate4162  (.A(II10937), .Z(g6194) ) ;
AND2    gate4163  (.A(g4912), .B(g5053), .Z(g5489) ) ;
INV     gate4164  (.A(g5489), .Z(II10940) ) ;
INV     gate4165  (.A(II10940), .Z(g6195) ) ;
INV     gate4166  (.A(g5335), .Z(g6198) ) ;
AND2    gate4167  (.A(g3390), .B(g5070), .Z(g5563) ) ;
INV     gate4168  (.A(g5563), .Z(II10946) ) ;
INV     gate4169  (.A(II10946), .Z(g6201) ) ;
AND2    gate4170  (.A(g4889), .B(g5071), .Z(g5513) ) ;
INV     gate4171  (.A(g5513), .Z(II10949) ) ;
INV     gate4172  (.A(II10949), .Z(g6202) ) ;
INV     gate4173  (.A(g5628), .Z(g6205) ) ;
INV     gate4174  (.A(g5639), .Z(g6206) ) ;
INV     gate4175  (.A(g5719), .Z(II10962) ) ;
INV     gate4176  (.A(g5719), .Z(II10965) ) ;
INV     gate4177  (.A(II10965), .Z(g6208) ) ;
INV     gate4178  (.A(g5606), .Z(II10969) ) ;
INV     gate4179  (.A(II10969), .Z(g6210) ) ;
INV     gate4180  (.A(g5645), .Z(g6211) ) ;
INV     gate4181  (.A(g5726), .Z(II10973) ) ;
INV     gate4182  (.A(g5726), .Z(II10976) ) ;
INV     gate4183  (.A(II10976), .Z(g6213) ) ;
INV     gate4184  (.A(g5609), .Z(II10987) ) ;
INV     gate4185  (.A(II10987), .Z(g6216) ) ;
INV     gate4186  (.A(g5649), .Z(g6217) ) ;
NAND3   gate4187  (.A(g5056), .B(g5039), .C(g5023), .Z(g5672) ) ;
INV     gate4188  (.A(g5672), .Z(II10998) ) ;
INV     gate4189  (.A(II10998), .Z(g6219) ) ;
OR2     gate4190  (.A(g5057), .B(g5040), .Z(g5698) ) ;
INV     gate4191  (.A(g5698), .Z(II11001) ) ;
INV     gate4192  (.A(II11001), .Z(g6220) ) ;
INV     gate4193  (.A(g5613), .Z(II11004) ) ;
INV     gate4194  (.A(II11004), .Z(g6221) ) ;
INV     gate4195  (.A(g5654), .Z(g6222) ) ;
INV     gate4196  (.A(g5693), .Z(II11008) ) ;
INV     gate4197  (.A(g5693), .Z(II11011) ) ;
INV     gate4198  (.A(II11011), .Z(g6224) ) ;
INV     gate4199  (.A(g5621), .Z(II11014) ) ;
INV     gate4200  (.A(II11014), .Z(g6225) ) ;
INV     gate4201  (.A(g5658), .Z(g6226) ) ;
INV     gate4202  (.A(g5626), .Z(II11018) ) ;
INV     gate4203  (.A(II11018), .Z(g6227) ) ;
INV     gate4204  (.A(g5627), .Z(II11021) ) ;
INV     gate4205  (.A(II11021), .Z(g6228) ) ;
INV     gate4206  (.A(g5665), .Z(g6229) ) ;
INV     gate4207  (.A(g5638), .Z(II11025) ) ;
INV     gate4208  (.A(II11025), .Z(g6230) ) ;
INV     gate4209  (.A(g5642), .Z(II11028) ) ;
INV     gate4210  (.A(II11028), .Z(g6231) ) ;
INV     gate4211  (.A(g5335), .Z(II11031) ) ;
INV     gate4212  (.A(II11031), .Z(g6232) ) ;
INV     gate4213  (.A(g5644), .Z(II11034) ) ;
INV     gate4214  (.A(II11034), .Z(g6235) ) ;
INV     gate4215  (.A(g5299), .Z(II11037) ) ;
INV     gate4216  (.A(g5299), .Z(II11040) ) ;
INV     gate4217  (.A(II11040), .Z(g6237) ) ;
INV     gate4218  (.A(g5648), .Z(II11043) ) ;
INV     gate4219  (.A(II11043), .Z(g6238) ) ;
INV     gate4220  (.A(g5653), .Z(II11047) ) ;
INV     gate4221  (.A(II11047), .Z(g6242) ) ;
INV     gate4222  (.A(g5335), .Z(II11050) ) ;
INV     gate4223  (.A(II11050), .Z(g6243) ) ;
INV     gate4224  (.A(g5670), .Z(g6244) ) ;
INV     gate4225  (.A(g5690), .Z(g6245) ) ;
INV     gate4226  (.A(g5696), .Z(II11055) ) ;
INV     gate4227  (.A(II11055), .Z(g6246) ) ;
INV     gate4228  (.A(g5679), .Z(g6250) ) ;
INV     gate4229  (.A(g5453), .Z(II11060) ) ;
INV     gate4230  (.A(II11060), .Z(g6251) ) ;
INV     gate4231  (.A(g5418), .Z(g6252) ) ;
INV     gate4232  (.A(g5403), .Z(g6253) ) ;
INV     gate4233  (.A(g5683), .Z(g6254) ) ;
INV     gate4234  (.A(g5460), .Z(II11066) ) ;
INV     gate4235  (.A(II11066), .Z(g6255) ) ;
INV     gate4236  (.A(g5671), .Z(II11069) ) ;
INV     gate4237  (.A(II11069), .Z(g6256) ) ;
INV     gate4238  (.A(g5685), .Z(g6257) ) ;
INV     gate4239  (.A(g5427), .Z(g6258) ) ;
INV     gate4240  (.A(g5688), .Z(g6263) ) ;
INV     gate4241  (.A(g5403), .Z(g6264) ) ;
INV     gate4242  (.A(g5397), .Z(II11086) ) ;
INV     gate4243  (.A(II11086), .Z(g6267) ) ;
INV     gate4244  (.A(g1000), .Z(II11090) ) ;
INV     gate4245  (.A(g5418), .Z(II11129) ) ;
INV     gate4246  (.A(II11129), .Z(g6278) ) ;
AND2    gate4247  (.A(g5140), .B(g2794), .Z(g5624) ) ;
INV     gate4248  (.A(g5624), .Z(II11132) ) ;
INV     gate4249  (.A(II11132), .Z(g6279) ) ;
INV     gate4250  (.A(g6155), .Z(II11191) ) ;
INV     gate4251  (.A(g6243), .Z(II11194) ) ;
INV     gate4252  (.A(g6122), .Z(II11197) ) ;
INV     gate4253  (.A(g6251), .Z(II11200) ) ;
INV     gate4254  (.A(g6129), .Z(II11203) ) ;
INV     gate4255  (.A(g6133), .Z(II11206) ) ;
INV     gate4256  (.A(g6139), .Z(II11209) ) ;
INV     gate4257  (.A(g6146), .Z(II11212) ) ;
INV     gate4258  (.A(g6156), .Z(II11215) ) ;
INV     gate4259  (.A(g6161), .Z(II11218) ) ;
INV     gate4260  (.A(g6167), .Z(II11221) ) ;
INV     gate4261  (.A(g6255), .Z(II11224) ) ;
INV     gate4262  (.A(g6130), .Z(II11227) ) ;
INV     gate4263  (.A(g6140), .Z(II11230) ) ;
INV     gate4264  (.A(g6147), .Z(II11233) ) ;
INV     gate4265  (.A(g6148), .Z(II11236) ) ;
INV     gate4266  (.A(g6173), .Z(II11239) ) ;
INV     gate4267  (.A(g6183), .Z(II11242) ) ;
INV     gate4268  (.A(g6143), .Z(II11245) ) ;
INV     gate4269  (.A(g6149), .Z(II11248) ) ;
INV     gate4270  (.A(g6152), .Z(II11251) ) ;
INV     gate4271  (.A(g5793), .Z(II11254) ) ;
INV     gate4272  (.A(g5805), .Z(II11257) ) ;
INV     gate4273  (.A(g5779), .Z(II11260) ) ;
INV     gate4274  (.A(g5784), .Z(II11263) ) ;
INV     gate4275  (.A(g5794), .Z(II11266) ) ;
INV     gate4276  (.A(g5756), .Z(II11269) ) ;
INV     gate4277  (.A(g5758), .Z(II11272) ) ;
INV     gate4278  (.A(g5768), .Z(II11275) ) ;
INV     gate4279  (.A(g5780), .Z(II11278) ) ;
INV     gate4280  (.A(g5785), .Z(II11281) ) ;
INV     gate4281  (.A(g5795), .Z(II11284) ) ;
INV     gate4282  (.A(g5806), .Z(II11287) ) ;
INV     gate4283  (.A(g5818), .Z(II11290) ) ;
INV     gate4284  (.A(g5824), .Z(II11293) ) ;
INV     gate4285  (.A(g5831), .Z(II11296) ) ;
INV     gate4286  (.A(g5786), .Z(II11299) ) ;
INV     gate4287  (.A(g5796), .Z(II11302) ) ;
INV     gate4288  (.A(g5807), .Z(II11305) ) ;
INV     gate4289  (.A(g5759), .Z(II11308) ) ;
INV     gate4290  (.A(g5760), .Z(II11311) ) ;
INV     gate4291  (.A(g5781), .Z(II11314) ) ;
INV     gate4292  (.A(g5787), .Z(II11317) ) ;
INV     gate4293  (.A(g5797), .Z(II11320) ) ;
INV     gate4294  (.A(g5808), .Z(II11323) ) ;
INV     gate4295  (.A(g5819), .Z(II11326) ) ;
INV     gate4296  (.A(g5825), .Z(II11329) ) ;
INV     gate4297  (.A(g5832), .Z(II11332) ) ;
INV     gate4298  (.A(g5839), .Z(II11335) ) ;
INV     gate4299  (.A(g5798), .Z(II11338) ) ;
INV     gate4300  (.A(g5809), .Z(II11341) ) ;
INV     gate4301  (.A(g5820), .Z(II11344) ) ;
INV     gate4302  (.A(g5761), .Z(II11347) ) ;
INV     gate4303  (.A(g5763), .Z(II11350) ) ;
INV     gate4304  (.A(g5788), .Z(II11353) ) ;
INV     gate4305  (.A(g5799), .Z(II11356) ) ;
INV     gate4306  (.A(g5810), .Z(II11359) ) ;
INV     gate4307  (.A(g5821), .Z(II11362) ) ;
INV     gate4308  (.A(g5826), .Z(II11365) ) ;
INV     gate4309  (.A(g5833), .Z(II11368) ) ;
INV     gate4310  (.A(g5840), .Z(II11371) ) ;
INV     gate4311  (.A(g5844), .Z(II11374) ) ;
INV     gate4312  (.A(g5811), .Z(II11377) ) ;
INV     gate4313  (.A(g5822), .Z(II11380) ) ;
INV     gate4314  (.A(g5827), .Z(II11383) ) ;
INV     gate4315  (.A(g5764), .Z(II11386) ) ;
INV     gate4316  (.A(g5766), .Z(II11389) ) ;
INV     gate4317  (.A(g5800), .Z(II11392) ) ;
INV     gate4318  (.A(g5812), .Z(II11395) ) ;
INV     gate4319  (.A(g5823), .Z(II11398) ) ;
INV     gate4320  (.A(g5828), .Z(II11401) ) ;
INV     gate4321  (.A(g5834), .Z(II11404) ) ;
INV     gate4322  (.A(g5841), .Z(II11407) ) ;
INV     gate4323  (.A(g5845), .Z(II11410) ) ;
INV     gate4324  (.A(g5871), .Z(II11413) ) ;
INV     gate4325  (.A(g5829), .Z(II11416) ) ;
INV     gate4326  (.A(g5835), .Z(II11419) ) ;
INV     gate4327  (.A(g5842), .Z(II11422) ) ;
INV     gate4328  (.A(g5872), .Z(II11425) ) ;
INV     gate4329  (.A(g5813), .Z(II11428) ) ;
INV     gate4330  (.A(g5782), .Z(II11431) ) ;
INV     gate4331  (.A(g5789), .Z(II11434) ) ;
INV     gate4332  (.A(g5801), .Z(II11437) ) ;
INV     gate4333  (.A(g6009), .Z(II11440) ) ;
INV     gate4334  (.A(g6038), .Z(II11443) ) ;
INV     gate4335  (.A(g6062), .Z(II11446) ) ;
INV     gate4336  (.A(g6068), .Z(II11449) ) ;
INV     gate4337  (.A(g6071), .Z(II11452) ) ;
INV     gate4338  (.A(g6087), .Z(II11455) ) ;
INV     gate4339  (.A(g6063), .Z(II11458) ) ;
INV     gate4340  (.A(g6094), .Z(II11461) ) ;
INV     gate4341  (.A(g6088), .Z(II11464) ) ;
INV     gate4342  (.A(g6064), .Z(II11467) ) ;
INV     gate4343  (.A(g6095), .Z(II11470) ) ;
INV     gate4344  (.A(g6069), .Z(II11473) ) ;
INV     gate4345  (.A(g6194), .Z(II11476) ) ;
INV     gate4346  (.A(g6201), .Z(II11479) ) ;
INV     gate4347  (.A(g6117), .Z(II11482) ) ;
INV     gate4348  (.A(g6137), .Z(II11485) ) ;
INV     gate4349  (.A(g6034), .Z(II11488) ) ;
INV     gate4350  (.A(g6010), .Z(II11491) ) ;
INV     gate4351  (.A(g6037), .Z(II11494) ) ;
INV     gate4352  (.A(g6014), .Z(II11497) ) ;
INV     gate4353  (.A(g6219), .Z(II11500) ) ;
INV     gate4354  (.A(g6220), .Z(II11503) ) ;
INV     gate4355  (.A(g6189), .Z(II11506) ) ;
INV     gate4356  (.A(g5874), .Z(II11512) ) ;
INV     gate4357  (.A(II11512), .Z(g6397) ) ;
INV     gate4358  (.A(g5897), .Z(II11515) ) ;
INV     gate4359  (.A(II11515), .Z(g6398) ) ;
INV     gate4360  (.A(g5847), .Z(II11522) ) ;
INV     gate4361  (.A(II11522), .Z(g6403) ) ;
INV     gate4362  (.A(g5874), .Z(II11525) ) ;
INV     gate4363  (.A(II11525), .Z(g6404) ) ;
INV     gate4364  (.A(g5847), .Z(II11533) ) ;
INV     gate4365  (.A(II11533), .Z(g6410) ) ;
INV     gate4366  (.A(g6065), .Z(II11556) ) ;
INV     gate4367  (.A(g6065), .Z(II11559) ) ;
INV     gate4368  (.A(II11559), .Z(g6426) ) ;
INV     gate4369  (.A(g5939), .Z(II11562) ) ;
INV     gate4370  (.A(II11562), .Z(g6427) ) ;
INV     gate4371  (.A(g6279), .Z(II11569) ) ;
INV     gate4372  (.A(II11569), .Z(g6432) ) ;
INV     gate4373  (.A(g6256), .Z(II11586) ) ;
INV     gate4374  (.A(II11586), .Z(g6441) ) ;
INV     gate4375  (.A(g5814), .Z(II11591) ) ;
INV     gate4376  (.A(II11591), .Z(g6446) ) ;
INV     gate4377  (.A(g6228), .Z(II11596) ) ;
INV     gate4378  (.A(II11596), .Z(g6449) ) ;
AND2    gate4379  (.A(g5344), .B(g3079), .Z(g5767) ) ;
INV     gate4380  (.A(g5767), .Z(II11607) ) ;
INV     gate4381  (.A(II11607), .Z(g6461) ) ;
INV     gate4382  (.A(g5847), .Z(II11622) ) ;
INV     gate4383  (.A(II11622), .Z(g6468) ) ;
INV     gate4384  (.A(g5874), .Z(II11627) ) ;
INV     gate4385  (.A(II11627), .Z(g6471) ) ;
INV     gate4386  (.A(g5897), .Z(II11633) ) ;
INV     gate4387  (.A(II11633), .Z(g6475) ) ;
INV     gate4388  (.A(g5847), .Z(II11638) ) ;
INV     gate4389  (.A(II11638), .Z(g6478) ) ;
INV     gate4390  (.A(g5918), .Z(II11641) ) ;
INV     gate4391  (.A(II11641), .Z(g6481) ) ;
INV     gate4392  (.A(g5874), .Z(II11645) ) ;
INV     gate4393  (.A(II11645), .Z(g6483) ) ;
INV     gate4394  (.A(g6028), .Z(II11648) ) ;
INV     gate4395  (.A(II11648), .Z(g6486) ) ;
INV     gate4396  (.A(g5939), .Z(II11652) ) ;
INV     gate4397  (.A(II11652), .Z(g6488) ) ;
NOR2    gate4398  (.A(g5428), .B(g1888), .Z(g5772) ) ;
INV     gate4399  (.A(g5772), .Z(II11656) ) ;
INV     gate4400  (.A(II11656), .Z(g6490) ) ;
INV     gate4401  (.A(g5897), .Z(II11659) ) ;
INV     gate4402  (.A(II11659), .Z(g6493) ) ;
INV     gate4403  (.A(g5956), .Z(II11662) ) ;
INV     gate4404  (.A(II11662), .Z(g6496) ) ;
INV     gate4405  (.A(g5772), .Z(II11666) ) ;
INV     gate4406  (.A(II11666), .Z(g6498) ) ;
INV     gate4407  (.A(g5918), .Z(II11669) ) ;
INV     gate4408  (.A(II11669), .Z(g6501) ) ;
INV     gate4409  (.A(g5971), .Z(II11672) ) ;
INV     gate4410  (.A(II11672), .Z(g6502) ) ;
INV     gate4411  (.A(g6076), .Z(II11677) ) ;
INV     gate4412  (.A(II11677), .Z(g6505) ) ;
INV     gate4413  (.A(g5939), .Z(II11680) ) ;
INV     gate4414  (.A(II11680), .Z(g6506) ) ;
INV     gate4415  (.A(g5988), .Z(II11683) ) ;
INV     gate4416  (.A(II11683), .Z(g6507) ) ;
INV     gate4417  (.A(g6076), .Z(II11686) ) ;
INV     gate4418  (.A(II11686), .Z(g6508) ) ;
INV     gate4419  (.A(g5956), .Z(II11689) ) ;
INV     gate4420  (.A(II11689), .Z(g6509) ) ;
INV     gate4421  (.A(g6076), .Z(II11693) ) ;
INV     gate4422  (.A(II11693), .Z(g6511) ) ;
INV     gate4423  (.A(g5971), .Z(II11696) ) ;
INV     gate4424  (.A(II11696), .Z(g6514) ) ;
AND2    gate4425  (.A(g5548), .B(g4202), .Z(g6125) ) ;
INV     gate4426  (.A(g6125), .Z(g6515) ) ;
INV     gate4427  (.A(g5772), .Z(II11701) ) ;
INV     gate4428  (.A(II11701), .Z(g6517) ) ;
INV     gate4429  (.A(g6076), .Z(II11704) ) ;
INV     gate4430  (.A(II11704), .Z(g6520) ) ;
INV     gate4431  (.A(g5988), .Z(II11707) ) ;
INV     gate4432  (.A(II11707), .Z(g6523) ) ;
AND2    gate4433  (.A(g5681), .B(g1247), .Z(g6098) ) ;
INV     gate4434  (.A(g6098), .Z(II11710) ) ;
INV     gate4435  (.A(II11710), .Z(g6524) ) ;
INV     gate4436  (.A(g5772), .Z(II11714) ) ;
INV     gate4437  (.A(II11714), .Z(g6538) ) ;
OR2     gate4438  (.A(g3617), .B(g5558), .Z(g6115) ) ;
INV     gate4439  (.A(g6115), .Z(II11718) ) ;
INV     gate4440  (.A(II11718), .Z(g6542) ) ;
INV     gate4441  (.A(g5772), .Z(II11722) ) ;
INV     gate4442  (.A(II11722), .Z(g6552) ) ;
INV     gate4443  (.A(g6036), .Z(II11725) ) ;
INV     gate4444  (.A(II11725), .Z(g6553) ) ;
INV     gate4445  (.A(g5772), .Z(II11729) ) ;
INV     gate4446  (.A(II11729), .Z(g6555) ) ;
INV     gate4447  (.A(g6076), .Z(II11732) ) ;
INV     gate4448  (.A(II11732), .Z(g6556) ) ;
INV     gate4449  (.A(g6076), .Z(II11736) ) ;
INV     gate4450  (.A(II11736), .Z(g6562) ) ;
INV     gate4451  (.A(g6136), .Z(II11740) ) ;
INV     gate4452  (.A(II11740), .Z(g6566) ) ;
OR2     gate4453  (.A(g3617), .B(g5555), .Z(g6120) ) ;
INV     gate4454  (.A(g6120), .Z(II11744) ) ;
INV     gate4455  (.A(II11744), .Z(g6568) ) ;
OR2     gate4456  (.A(g3617), .B(g5556), .Z(g6123) ) ;
INV     gate4457  (.A(g6123), .Z(II11747) ) ;
INV     gate4458  (.A(II11747), .Z(g6569) ) ;
AND3    gate4459  (.A(g3760), .B(g5286), .C(g1695), .Z(g6056) ) ;
INV     gate4460  (.A(g6056), .Z(II11764) ) ;
INV     gate4461  (.A(II11764), .Z(g6572) ) ;
INV     gate4462  (.A(g5868), .Z(g6573) ) ;
OR2     gate4463  (.A(g4074), .B(g5334), .Z(g6262) ) ;
INV     gate4464  (.A(g6262), .Z(II11773) ) ;
INV     gate4465  (.A(II11773), .Z(g6581) ) ;
NAND2   gate4466  (.A(II10900), .B(II10901), .Z(g6180) ) ;
INV     gate4467  (.A(g6180), .Z(II11778) ) ;
INV     gate4468  (.A(II11778), .Z(g6586) ) ;
NAND2   gate4469  (.A(II11164), .B(II11165), .Z(g6284) ) ;
INV     gate4470  (.A(g6284), .Z(II11781) ) ;
INV     gate4471  (.A(II11781), .Z(g6587) ) ;
INV     gate4472  (.A(g5836), .Z(g6588) ) ;
INV     gate4473  (.A(g6083), .Z(g6589) ) ;
NAND2   gate4474  (.A(II11095), .B(II11096), .Z(g6273) ) ;
INV     gate4475  (.A(g6273), .Z(II11787) ) ;
INV     gate4476  (.A(II11787), .Z(g6591) ) ;
NAND2   gate4477  (.A(II11150), .B(II11151), .Z(g6282) ) ;
INV     gate4478  (.A(g6282), .Z(II11790) ) ;
INV     gate4479  (.A(II11790), .Z(g6592) ) ;
NAND2   gate4480  (.A(II10924), .B(II10925), .Z(g6188) ) ;
INV     gate4481  (.A(g6188), .Z(II11793) ) ;
INV     gate4482  (.A(II11793), .Z(g6593) ) ;
NAND2   gate4483  (.A(II11185), .B(II11186), .Z(g6287) ) ;
INV     gate4484  (.A(g6287), .Z(II11796) ) ;
INV     gate4485  (.A(II11796), .Z(g6594) ) ;
INV     gate4486  (.A(g6083), .Z(g6595) ) ;
NAND2   gate4487  (.A(II10848), .B(II10849), .Z(g6164) ) ;
INV     gate4488  (.A(g6164), .Z(II11800) ) ;
INV     gate4489  (.A(II11800), .Z(g6596) ) ;
NAND2   gate4490  (.A(II11136), .B(II11137), .Z(g6280) ) ;
INV     gate4491  (.A(g6280), .Z(II11803) ) ;
INV     gate4492  (.A(II11803), .Z(g6597) ) ;
NAND2   gate4493  (.A(II11109), .B(II11110), .Z(g6275) ) ;
INV     gate4494  (.A(g6275), .Z(II11806) ) ;
INV     gate4495  (.A(II11806), .Z(g6598) ) ;
NAND2   gate4496  (.A(II11171), .B(II11172), .Z(g6285) ) ;
INV     gate4497  (.A(g6285), .Z(II11809) ) ;
INV     gate4498  (.A(II11809), .Z(g6599) ) ;
INV     gate4499  (.A(g6083), .Z(g6601) ) ;
NAND2   gate4500  (.A(II10867), .B(II10868), .Z(g6169) ) ;
INV     gate4501  (.A(g6169), .Z(II11815) ) ;
INV     gate4502  (.A(II11815), .Z(g6603) ) ;
NAND2   gate4503  (.A(II11116), .B(II11117), .Z(g6276) ) ;
INV     gate4504  (.A(g6276), .Z(II11818) ) ;
INV     gate4505  (.A(II11818), .Z(g6604) ) ;
NAND2   gate4506  (.A(II10874), .B(II10875), .Z(g6170) ) ;
INV     gate4507  (.A(g6170), .Z(II11821) ) ;
INV     gate4508  (.A(II11821), .Z(g6605) ) ;
NAND2   gate4509  (.A(II11157), .B(II11158), .Z(g6283) ) ;
INV     gate4510  (.A(g6283), .Z(II11824) ) ;
INV     gate4511  (.A(II11824), .Z(g6606) ) ;
INV     gate4512  (.A(g6231), .Z(II11827) ) ;
INV     gate4513  (.A(II11827), .Z(g6607) ) ;
NAND2   gate4514  (.A(II11102), .B(II11103), .Z(g6274) ) ;
INV     gate4515  (.A(g6274), .Z(II11832) ) ;
INV     gate4516  (.A(II11832), .Z(g6612) ) ;
NAND2   gate4517  (.A(II10907), .B(II10908), .Z(g6181) ) ;
INV     gate4518  (.A(g6181), .Z(II11835) ) ;
INV     gate4519  (.A(II11835), .Z(g6613) ) ;
NAND2   gate4520  (.A(II11143), .B(II11144), .Z(g6281) ) ;
INV     gate4521  (.A(g6281), .Z(II11838) ) ;
INV     gate4522  (.A(II11838), .Z(g6614) ) ;
NAND2   gate4523  (.A(II10835), .B(II10836), .Z(g6159) ) ;
INV     gate4524  (.A(g6159), .Z(II11848) ) ;
INV     gate4525  (.A(II11848), .Z(g6616) ) ;
NAND2   gate4526  (.A(II11123), .B(II11124), .Z(g6277) ) ;
INV     gate4527  (.A(g6277), .Z(II11851) ) ;
INV     gate4528  (.A(II11851), .Z(g6617) ) ;
AND3    gate4529  (.A(g3716), .B(g5633), .C(II10597), .Z(g6003) ) ;
INV     gate4530  (.A(g6003), .Z(g6618) ) ;
NAND2   gate4531  (.A(II10321), .B(II10322), .Z(g5751) ) ;
INV     gate4532  (.A(g5751), .Z(II11855) ) ;
INV     gate4533  (.A(II11855), .Z(g6621) ) ;
NAND2   gate4534  (.A(II10855), .B(II10856), .Z(g6165) ) ;
INV     gate4535  (.A(g6165), .Z(II11858) ) ;
INV     gate4536  (.A(II11858), .Z(g6622) ) ;
NAND2   gate4537  (.A(II10299), .B(II10300), .Z(g5747) ) ;
INV     gate4538  (.A(g5747), .Z(II11861) ) ;
INV     gate4539  (.A(II11861), .Z(g6623) ) ;
NAND2   gate4540  (.A(II10335), .B(II10336), .Z(g5753) ) ;
INV     gate4541  (.A(g5753), .Z(II11864) ) ;
INV     gate4542  (.A(II11864), .Z(g6624) ) ;
NAND2   gate4543  (.A(II11178), .B(II11179), .Z(g6286) ) ;
INV     gate4544  (.A(g6286), .Z(II11867) ) ;
INV     gate4545  (.A(II11867), .Z(g6625) ) ;
NAND2   gate4546  (.A(II10328), .B(II10329), .Z(g5752) ) ;
INV     gate4547  (.A(g5752), .Z(II11870) ) ;
INV     gate4548  (.A(II11870), .Z(g6626) ) ;
NAND2   gate4549  (.A(II10306), .B(II10307), .Z(g5748) ) ;
INV     gate4550  (.A(g5748), .Z(II11880) ) ;
INV     gate4551  (.A(II11880), .Z(g6628) ) ;
AND2    gate4552  (.A(g5712), .B(g5038), .Z(g6091) ) ;
INV     gate4553  (.A(g6091), .Z(II11884) ) ;
INV     gate4554  (.A(II11884), .Z(g6630) ) ;
INV     gate4555  (.A(g5918), .Z(II11887) ) ;
INV     gate4556  (.A(II11887), .Z(g6631) ) ;
INV     gate4557  (.A(g6135), .Z(II11890) ) ;
INV     gate4558  (.A(II11890), .Z(g6632) ) ;
INV     gate4559  (.A(g5956), .Z(II11894) ) ;
INV     gate4560  (.A(II11894), .Z(g6634) ) ;
INV     gate4561  (.A(g6141), .Z(II11897) ) ;
INV     gate4562  (.A(II11897), .Z(g6635) ) ;
INV     gate4563  (.A(g5847), .Z(II11900) ) ;
INV     gate4564  (.A(II11900), .Z(g6636) ) ;
INV     gate4565  (.A(g5939), .Z(II11903) ) ;
INV     gate4566  (.A(II11903), .Z(g6637) ) ;
INV     gate4567  (.A(g6198), .Z(g6639) ) ;
INV     gate4568  (.A(g5918), .Z(II11908) ) ;
INV     gate4569  (.A(II11908), .Z(g6640) ) ;
INV     gate4570  (.A(g5897), .Z(II11912) ) ;
INV     gate4571  (.A(II11912), .Z(g6642) ) ;
INV     gate4572  (.A(g6208), .Z(g6644) ) ;
INV     gate4573  (.A(g5897), .Z(II11917) ) ;
INV     gate4574  (.A(II11917), .Z(g6645) ) ;
INV     gate4575  (.A(g5874), .Z(II11920) ) ;
INV     gate4576  (.A(II11920), .Z(g6646) ) ;
INV     gate4577  (.A(g5939), .Z(II11923) ) ;
INV     gate4578  (.A(II11923), .Z(g6647) ) ;
INV     gate4579  (.A(g6190), .Z(II11926) ) ;
INV     gate4580  (.A(g6190), .Z(II11929) ) ;
INV     gate4581  (.A(II11929), .Z(g6649) ) ;
INV     gate4582  (.A(g6213), .Z(g6650) ) ;
INV     gate4583  (.A(g5847), .Z(II11933) ) ;
INV     gate4584  (.A(II11933), .Z(g6651) ) ;
INV     gate4585  (.A(g5918), .Z(II11936) ) ;
INV     gate4586  (.A(II11936), .Z(g6652) ) ;
INV     gate4587  (.A(g6015), .Z(II11939) ) ;
INV     gate4588  (.A(g6015), .Z(II11942) ) ;
INV     gate4589  (.A(II11942), .Z(g6654) ) ;
INV     gate4590  (.A(g5874), .Z(II11945) ) ;
INV     gate4591  (.A(II11945), .Z(g6655) ) ;
INV     gate4592  (.A(g5897), .Z(II11948) ) ;
INV     gate4593  (.A(II11948), .Z(g6656) ) ;
INV     gate4594  (.A(g5847), .Z(II11951) ) ;
INV     gate4595  (.A(II11951), .Z(g6657) ) ;
INV     gate4596  (.A(g6224), .Z(g6658) ) ;
INV     gate4597  (.A(g5988), .Z(II11955) ) ;
INV     gate4598  (.A(II11955), .Z(g6659) ) ;
INV     gate4599  (.A(g5874), .Z(II11958) ) ;
INV     gate4600  (.A(II11958), .Z(g6660) ) ;
INV     gate4601  (.A(g5988), .Z(II11961) ) ;
INV     gate4602  (.A(II11961), .Z(g6661) ) ;
INV     gate4603  (.A(g5971), .Z(II11964) ) ;
INV     gate4604  (.A(II11964), .Z(g6662) ) ;
INV     gate4605  (.A(g5971), .Z(II11967) ) ;
INV     gate4606  (.A(II11967), .Z(g6663) ) ;
INV     gate4607  (.A(g6179), .Z(II11971) ) ;
INV     gate4608  (.A(II11971), .Z(g6671) ) ;
INV     gate4609  (.A(g5956), .Z(II11974) ) ;
INV     gate4610  (.A(II11974), .Z(g6672) ) ;
INV     gate4611  (.A(g6186), .Z(II11978) ) ;
INV     gate4612  (.A(II11978), .Z(g6674) ) ;
INV     gate4613  (.A(g6246), .Z(II11981) ) ;
INV     gate4614  (.A(g6246), .Z(II11984) ) ;
INV     gate4615  (.A(II11984), .Z(g6676) ) ;
INV     gate4616  (.A(g6278), .Z(II11987) ) ;
INV     gate4617  (.A(II11987), .Z(g6677) ) ;
INV     gate4618  (.A(g5939), .Z(II11991) ) ;
INV     gate4619  (.A(II11991), .Z(g6681) ) ;
INV     gate4620  (.A(g6195), .Z(II11994) ) ;
INV     gate4621  (.A(II11994), .Z(g6682) ) ;
INV     gate4622  (.A(g6237), .Z(g6683) ) ;
INV     gate4623  (.A(g5918), .Z(II11998) ) ;
INV     gate4624  (.A(II11998), .Z(g6684) ) ;
INV     gate4625  (.A(g6202), .Z(II12003) ) ;
INV     gate4626  (.A(II12003), .Z(g6687) ) ;
INV     gate4627  (.A(g5897), .Z(II12008) ) ;
INV     gate4628  (.A(II12008), .Z(g6692) ) ;
INV     gate4629  (.A(g5939), .Z(II12011) ) ;
INV     gate4630  (.A(II12011), .Z(g6693) ) ;
INV     gate4631  (.A(g5874), .Z(II12022) ) ;
INV     gate4632  (.A(II12022), .Z(g6696) ) ;
INV     gate4633  (.A(g5918), .Z(II12025) ) ;
INV     gate4634  (.A(II12025), .Z(g6697) ) ;
INV     gate4635  (.A(g6244), .Z(g6700) ) ;
INV     gate4636  (.A(g5847), .Z(II12038) ) ;
INV     gate4637  (.A(II12038), .Z(g6702) ) ;
INV     gate4638  (.A(g5897), .Z(II12041) ) ;
INV     gate4639  (.A(II12041), .Z(g6703) ) ;
INV     gate4640  (.A(g5847), .Z(II12044) ) ;
INV     gate4641  (.A(II12044), .Z(g6704) ) ;
INV     gate4642  (.A(g6250), .Z(g6708) ) ;
INV     gate4643  (.A(g5874), .Z(II12059) ) ;
INV     gate4644  (.A(II12059), .Z(g6711) ) ;
INV     gate4645  (.A(g5988), .Z(II12062) ) ;
INV     gate4646  (.A(II12062), .Z(g6712) ) ;
INV     gate4647  (.A(g5897), .Z(II12065) ) ;
INV     gate4648  (.A(II12065), .Z(g6713) ) ;
INV     gate4649  (.A(g5847), .Z(II12068) ) ;
INV     gate4650  (.A(II12068), .Z(g6714) ) ;
INV     gate4651  (.A(g6254), .Z(g6720) ) ;
INV     gate4652  (.A(g6257), .Z(g6721) ) ;
INV     gate4653  (.A(g5971), .Z(II12085) ) ;
INV     gate4654  (.A(II12085), .Z(g6723) ) ;
INV     gate4655  (.A(g5874), .Z(II12088) ) ;
INV     gate4656  (.A(II12088), .Z(g6724) ) ;
INV     gate4657  (.A(g5988), .Z(II12091) ) ;
INV     gate4658  (.A(II12091), .Z(g6725) ) ;
INV     gate4659  (.A(g6263), .Z(g6729) ) ;
INV     gate4660  (.A(g5956), .Z(II12098) ) ;
INV     gate4661  (.A(II12098), .Z(g6730) ) ;
INV     gate4662  (.A(g5971), .Z(II12101) ) ;
INV     gate4663  (.A(II12101), .Z(g6731) ) ;
INV     gate4664  (.A(g5939), .Z(II12108) ) ;
INV     gate4665  (.A(II12108), .Z(g6736) ) ;
INV     gate4666  (.A(g5956), .Z(II12111) ) ;
INV     gate4667  (.A(II12111), .Z(g6737) ) ;
INV     gate4668  (.A(g5918), .Z(II12117) ) ;
INV     gate4669  (.A(II12117), .Z(g6741) ) ;
INV     gate4670  (.A(g5939), .Z(II12120) ) ;
INV     gate4671  (.A(II12120), .Z(g6742) ) ;
INV     gate4672  (.A(g5847), .Z(II12124) ) ;
INV     gate4673  (.A(II12124), .Z(g6744) ) ;
INV     gate4674  (.A(g5897), .Z(II12128) ) ;
INV     gate4675  (.A(II12128), .Z(g6751) ) ;
INV     gate4676  (.A(g5918), .Z(II12131) ) ;
INV     gate4677  (.A(II12131), .Z(g6752) ) ;
INV     gate4678  (.A(g5988), .Z(II12135) ) ;
INV     gate4679  (.A(II12135), .Z(g6754) ) ;
INV     gate4680  (.A(g5874), .Z(II12138) ) ;
INV     gate4681  (.A(II12138), .Z(g6755) ) ;
INV     gate4682  (.A(g5897), .Z(II12141) ) ;
INV     gate4683  (.A(II12141), .Z(g6756) ) ;
INV     gate4684  (.A(g5971), .Z(II12145) ) ;
INV     gate4685  (.A(II12145), .Z(g6758) ) ;
INV     gate4686  (.A(g5988), .Z(II12148) ) ;
INV     gate4687  (.A(II12148), .Z(g6759) ) ;
INV     gate4688  (.A(g5847), .Z(II12151) ) ;
INV     gate4689  (.A(II12151), .Z(g6760) ) ;
INV     gate4690  (.A(g5874), .Z(II12154) ) ;
INV     gate4691  (.A(II12154), .Z(g6761) ) ;
INV     gate4692  (.A(g5956), .Z(II12158) ) ;
INV     gate4693  (.A(II12158), .Z(g6763) ) ;
INV     gate4694  (.A(g5971), .Z(II12161) ) ;
INV     gate4695  (.A(II12161), .Z(g6764) ) ;
INV     gate4696  (.A(g5847), .Z(II12164) ) ;
INV     gate4697  (.A(II12164), .Z(g6765) ) ;
INV     gate4698  (.A(g5939), .Z(II12167) ) ;
INV     gate4699  (.A(II12167), .Z(g6766) ) ;
INV     gate4700  (.A(g5956), .Z(II12170) ) ;
INV     gate4701  (.A(II12170), .Z(g6767) ) ;
INV     gate4702  (.A(g5918), .Z(II12173) ) ;
INV     gate4703  (.A(II12173), .Z(g6768) ) ;
INV     gate4704  (.A(g5939), .Z(II12176) ) ;
INV     gate4705  (.A(II12176), .Z(g6769) ) ;
INV     gate4706  (.A(g5897), .Z(II12187) ) ;
INV     gate4707  (.A(II12187), .Z(g6772) ) ;
INV     gate4708  (.A(g5918), .Z(II12190) ) ;
INV     gate4709  (.A(II12190), .Z(g6773) ) ;
INV     gate4710  (.A(g6468), .Z(II12193) ) ;
INV     gate4711  (.A(g6471), .Z(II12196) ) ;
INV     gate4712  (.A(g6475), .Z(II12199) ) ;
INV     gate4713  (.A(g6481), .Z(II12202) ) ;
INV     gate4714  (.A(g6488), .Z(II12205) ) ;
INV     gate4715  (.A(g6496), .Z(II12208) ) ;
INV     gate4716  (.A(g6502), .Z(II12211) ) ;
INV     gate4717  (.A(g6507), .Z(II12214) ) ;
INV     gate4718  (.A(g6631), .Z(II12217) ) ;
INV     gate4719  (.A(g6645), .Z(II12220) ) ;
INV     gate4720  (.A(g6655), .Z(II12223) ) ;
INV     gate4721  (.A(g6636), .Z(II12226) ) ;
INV     gate4722  (.A(g6659), .Z(II12229) ) ;
INV     gate4723  (.A(g6662), .Z(II12232) ) ;
INV     gate4724  (.A(g6634), .Z(II12235) ) ;
INV     gate4725  (.A(g6637), .Z(II12238) ) ;
INV     gate4726  (.A(g6640), .Z(II12241) ) ;
INV     gate4727  (.A(g6642), .Z(II12244) ) ;
INV     gate4728  (.A(g6646), .Z(II12247) ) ;
INV     gate4729  (.A(g6651), .Z(II12250) ) ;
INV     gate4730  (.A(g6427), .Z(II12253) ) ;
INV     gate4731  (.A(g6647), .Z(II12256) ) ;
INV     gate4732  (.A(g6652), .Z(II12259) ) ;
INV     gate4733  (.A(g6656), .Z(II12262) ) ;
INV     gate4734  (.A(g6660), .Z(II12265) ) ;
INV     gate4735  (.A(g6661), .Z(II12268) ) ;
INV     gate4736  (.A(g6663), .Z(II12271) ) ;
INV     gate4737  (.A(g6672), .Z(II12274) ) ;
INV     gate4738  (.A(g6681), .Z(II12277) ) ;
INV     gate4739  (.A(g6684), .Z(II12280) ) ;
INV     gate4740  (.A(g6692), .Z(II12283) ) ;
INV     gate4741  (.A(g6696), .Z(II12286) ) ;
INV     gate4742  (.A(g6702), .Z(II12289) ) ;
INV     gate4743  (.A(g6657), .Z(II12292) ) ;
INV     gate4744  (.A(g6693), .Z(II12295) ) ;
INV     gate4745  (.A(g6697), .Z(II12298) ) ;
INV     gate4746  (.A(g6703), .Z(II12301) ) ;
INV     gate4747  (.A(g6711), .Z(II12304) ) ;
INV     gate4748  (.A(g6712), .Z(II12307) ) ;
INV     gate4749  (.A(g6723), .Z(II12310) ) ;
INV     gate4750  (.A(g6730), .Z(II12313) ) ;
INV     gate4751  (.A(g6736), .Z(II12316) ) ;
INV     gate4752  (.A(g6741), .Z(II12319) ) ;
INV     gate4753  (.A(g6751), .Z(II12322) ) ;
INV     gate4754  (.A(g6755), .Z(II12325) ) ;
INV     gate4755  (.A(g6760), .Z(II12328) ) ;
INV     gate4756  (.A(g6704), .Z(II12331) ) ;
INV     gate4757  (.A(g6713), .Z(II12334) ) ;
INV     gate4758  (.A(g6724), .Z(II12337) ) ;
INV     gate4759  (.A(g6725), .Z(II12340) ) ;
INV     gate4760  (.A(g6731), .Z(II12343) ) ;
INV     gate4761  (.A(g6737), .Z(II12346) ) ;
INV     gate4762  (.A(g6742), .Z(II12349) ) ;
INV     gate4763  (.A(g6752), .Z(II12352) ) ;
INV     gate4764  (.A(g6756), .Z(II12355) ) ;
INV     gate4765  (.A(g6761), .Z(II12358) ) ;
INV     gate4766  (.A(g6765), .Z(II12361) ) ;
INV     gate4767  (.A(g6714), .Z(II12364) ) ;
INV     gate4768  (.A(g6754), .Z(II12367) ) ;
INV     gate4769  (.A(g6758), .Z(II12370) ) ;
INV     gate4770  (.A(g6763), .Z(II12373) ) ;
INV     gate4771  (.A(g6766), .Z(II12376) ) ;
INV     gate4772  (.A(g6768), .Z(II12379) ) ;
INV     gate4773  (.A(g6772), .Z(II12382) ) ;
INV     gate4774  (.A(g6397), .Z(II12385) ) ;
INV     gate4775  (.A(g6403), .Z(II12388) ) ;
INV     gate4776  (.A(g6744), .Z(II12391) ) ;
INV     gate4777  (.A(g6759), .Z(II12394) ) ;
INV     gate4778  (.A(g6764), .Z(II12397) ) ;
INV     gate4779  (.A(g6767), .Z(II12400) ) ;
INV     gate4780  (.A(g6769), .Z(II12403) ) ;
INV     gate4781  (.A(g6773), .Z(II12406) ) ;
INV     gate4782  (.A(g6398), .Z(II12409) ) ;
INV     gate4783  (.A(g6404), .Z(II12412) ) ;
INV     gate4784  (.A(g6410), .Z(II12415) ) ;
INV     gate4785  (.A(g6572), .Z(II12418) ) ;
INV     gate4786  (.A(g6486), .Z(II12421) ) ;
INV     gate4787  (.A(g6446), .Z(II12424) ) ;
INV     gate4788  (.A(g6553), .Z(II12427) ) ;
INV     gate4789  (.A(g6432), .Z(II12430) ) ;
INV     gate4790  (.A(g6632), .Z(II12433) ) ;
INV     gate4791  (.A(g6635), .Z(II12436) ) ;
INV     gate4792  (.A(g6566), .Z(II12439) ) ;
INV     gate4793  (.A(g6542), .Z(II12442) ) ;
INV     gate4794  (.A(g6568), .Z(II12445) ) ;
INV     gate4795  (.A(g6569), .Z(II12448) ) ;
INV     gate4796  (.A(g6524), .Z(II12451) ) ;
INV     gate4797  (.A(g6581), .Z(II12454) ) ;
INV     gate4798  (.A(g6671), .Z(II12457) ) ;
INV     gate4799  (.A(g6674), .Z(II12460) ) ;
INV     gate4800  (.A(g6682), .Z(II12463) ) ;
INV     gate4801  (.A(g6687), .Z(II12466) ) ;
INV     gate4802  (.A(g6586), .Z(II12469) ) ;
INV     gate4803  (.A(g6591), .Z(II12472) ) ;
INV     gate4804  (.A(g6596), .Z(II12475) ) ;
INV     gate4805  (.A(g6603), .Z(II12478) ) ;
INV     gate4806  (.A(g6616), .Z(II12481) ) ;
INV     gate4807  (.A(g6621), .Z(II12484) ) ;
INV     gate4808  (.A(g6623), .Z(II12487) ) ;
INV     gate4809  (.A(g6625), .Z(II12490) ) ;
INV     gate4810  (.A(g6587), .Z(II12493) ) ;
INV     gate4811  (.A(g6592), .Z(II12496) ) ;
INV     gate4812  (.A(g6597), .Z(II12499) ) ;
INV     gate4813  (.A(g6604), .Z(II12502) ) ;
INV     gate4814  (.A(g6612), .Z(II12505) ) ;
INV     gate4815  (.A(g6593), .Z(II12508) ) ;
INV     gate4816  (.A(g6598), .Z(II12511) ) ;
INV     gate4817  (.A(g6605), .Z(II12514) ) ;
INV     gate4818  (.A(g6613), .Z(II12517) ) ;
INV     gate4819  (.A(g6622), .Z(II12520) ) ;
INV     gate4820  (.A(g6624), .Z(II12523) ) ;
INV     gate4821  (.A(g6626), .Z(II12526) ) ;
INV     gate4822  (.A(g6628), .Z(II12529) ) ;
INV     gate4823  (.A(g6594), .Z(II12532) ) ;
INV     gate4824  (.A(g6599), .Z(II12535) ) ;
INV     gate4825  (.A(g6606), .Z(II12538) ) ;
INV     gate4826  (.A(g6614), .Z(II12541) ) ;
INV     gate4827  (.A(g6617), .Z(II12544) ) ;
INV     gate4828  (.A(g6708), .Z(II12547) ) ;
INV     gate4829  (.A(II12547), .Z(g6892) ) ;
OR2     gate4830  (.A(g6112), .B(g5547), .Z(g6525) ) ;
INV     gate4831  (.A(g6525), .Z(g6894) ) ;
INV     gate4832  (.A(g6449), .Z(II12558) ) ;
INV     gate4833  (.A(g6449), .Z(II12561) ) ;
INV     gate4834  (.A(II12561), .Z(g6896) ) ;
INV     gate4835  (.A(g6720), .Z(II12564) ) ;
INV     gate4836  (.A(II12564), .Z(g6897) ) ;
INV     gate4837  (.A(g6721), .Z(II12567) ) ;
INV     gate4838  (.A(II12567), .Z(g6898) ) ;
INV     gate4839  (.A(g6525), .Z(g6899) ) ;
INV     gate4840  (.A(g6729), .Z(II12571) ) ;
INV     gate4841  (.A(II12571), .Z(g6900) ) ;
INV     gate4842  (.A(g6525), .Z(g6901) ) ;
AND2    gate4843  (.A(g1872), .B(g6198), .Z(g6745) ) ;
INV     gate4844  (.A(g6745), .Z(II12582) ) ;
INV     gate4845  (.A(II12582), .Z(g6903) ) ;
INV     gate4846  (.A(g6426), .Z(g6904) ) ;
AND2    gate4847  (.A(g1860), .B(g5868), .Z(g6643) ) ;
INV     gate4848  (.A(g6643), .Z(II12586) ) ;
INV     gate4849  (.A(II12586), .Z(g6905) ) ;
INV     gate4850  (.A(g1008), .Z(II12592) ) ;
NAND2   gate4851  (.A(II11758), .B(II11759), .Z(g6571) ) ;
INV     gate4852  (.A(g6571), .Z(II12609) ) ;
INV     gate4853  (.A(II12609), .Z(g6918) ) ;
INV     gate4854  (.A(g6525), .Z(g6922) ) ;
INV     gate4855  (.A(g6523), .Z(II12629) ) ;
INV     gate4856  (.A(II12629), .Z(g6936) ) ;
INV     gate4857  (.A(g6514), .Z(II12632) ) ;
INV     gate4858  (.A(II12632), .Z(g6937) ) ;
INV     gate4859  (.A(g6509), .Z(II12635) ) ;
INV     gate4860  (.A(II12635), .Z(g6938) ) ;
OR2     gate4861  (.A(g6125), .B(g1553), .Z(g6543) ) ;
INV     gate4862  (.A(g6543), .Z(g6939) ) ;
INV     gate4863  (.A(g6506), .Z(II12639) ) ;
INV     gate4864  (.A(II12639), .Z(g6940) ) ;
INV     gate4865  (.A(g6501), .Z(II12643) ) ;
INV     gate4866  (.A(II12643), .Z(g6944) ) ;
INV     gate4867  (.A(g6493), .Z(II12646) ) ;
INV     gate4868  (.A(II12646), .Z(g6945) ) ;
OR3     gate4869  (.A(g6196), .B(g6209), .C(g4937), .Z(g6457) ) ;
INV     gate4870  (.A(g6457), .Z(II12649) ) ;
INV     gate4871  (.A(II12649), .Z(g6946) ) ;
NOR3    gate4872  (.A(g5836), .B(g1901), .C(g1788), .Z(g6664) ) ;
INV     gate4873  (.A(g6664), .Z(II12652) ) ;
INV     gate4874  (.A(II12652), .Z(g6947) ) ;
OR4     gate4875  (.A(g6184), .B(g6259), .C(g6174), .D(g6214), .Z(g6458) ) ;
INV     gate4876  (.A(g6458), .Z(II12655) ) ;
INV     gate4877  (.A(II12655), .Z(g6948) ) ;
OR3     gate4878  (.A(g6259), .B(g6185), .C(II11603), .Z(g6459) ) ;
INV     gate4879  (.A(g6459), .Z(II12659) ) ;
INV     gate4880  (.A(II12659), .Z(g6950) ) ;
INV     gate4881  (.A(g6745), .Z(g6953) ) ;
NAND2   gate4882  (.A(g5939), .B(g5269), .Z(g6476) ) ;
INV     gate4883  (.A(g6476), .Z(II12666) ) ;
INV     gate4884  (.A(II12666), .Z(g6955) ) ;
NAND2   gate4885  (.A(g5269), .B(g5918), .Z(g6477) ) ;
INV     gate4886  (.A(g6477), .Z(II12669) ) ;
INV     gate4887  (.A(II12669), .Z(g6956) ) ;
NAND2   gate4888  (.A(g5269), .B(g5988), .Z(g6473) ) ;
INV     gate4889  (.A(g6473), .Z(II12672) ) ;
INV     gate4890  (.A(II12672), .Z(g6957) ) ;
NAND2   gate4891  (.A(g5278), .B(g5874), .Z(g6510) ) ;
INV     gate4892  (.A(g6510), .Z(II12675) ) ;
INV     gate4893  (.A(II12675), .Z(g6958) ) ;
NAND2   gate4894  (.A(g5897), .B(g5278), .Z(g6516) ) ;
INV     gate4895  (.A(g6516), .Z(II12678) ) ;
INV     gate4896  (.A(II12678), .Z(g6959) ) ;
NAND2   gate4897  (.A(g5918), .B(g5278), .Z(g6469) ) ;
INV     gate4898  (.A(g6469), .Z(II12681) ) ;
INV     gate4899  (.A(II12681), .Z(g6960) ) ;
NAND2   gate4900  (.A(g5971), .B(g5269), .Z(g6472) ) ;
INV     gate4901  (.A(g6472), .Z(II12684) ) ;
INV     gate4902  (.A(II12684), .Z(g6961) ) ;
INV     gate4903  (.A(g6745), .Z(II12687) ) ;
INV     gate4904  (.A(II12687), .Z(g6962) ) ;
NAND2   gate4905  (.A(g5956), .B(g5269), .Z(g6467) ) ;
INV     gate4906  (.A(g6467), .Z(II12690) ) ;
INV     gate4907  (.A(II12690), .Z(g6963) ) ;
NAND2   gate4908  (.A(g5269), .B(g5897), .Z(g6503) ) ;
INV     gate4909  (.A(g6503), .Z(II12696) ) ;
INV     gate4910  (.A(II12696), .Z(g6967) ) ;
NAND2   gate4911  (.A(g5269), .B(g5874), .Z(g6504) ) ;
INV     gate4912  (.A(g6504), .Z(II12699) ) ;
INV     gate4913  (.A(II12699), .Z(g6968) ) ;
NAND2   gate4914  (.A(g5278), .B(g5847), .Z(g6497) ) ;
INV     gate4915  (.A(g6497), .Z(II12702) ) ;
INV     gate4916  (.A(II12702), .Z(g6969) ) ;
NAND2   gate4917  (.A(g5269), .B(g5847), .Z(g6482) ) ;
INV     gate4918  (.A(g6482), .Z(II12708) ) ;
INV     gate4919  (.A(II12708), .Z(g6973) ) ;
INV     gate4920  (.A(g6543), .Z(II12712) ) ;
INV     gate4921  (.A(II12712), .Z(g6975) ) ;
INV     gate4922  (.A(g6664), .Z(g6977) ) ;
INV     gate4923  (.A(g6543), .Z(II12717) ) ;
INV     gate4924  (.A(II12717), .Z(g6978) ) ;
AND2    gate4925  (.A(g3390), .B(g6249), .Z(g6611) ) ;
INV     gate4926  (.A(g6611), .Z(II12722) ) ;
INV     gate4927  (.A(II12722), .Z(g6983) ) ;
OR3     gate4928  (.A(g2396), .B(g6131), .C(g1603), .Z(g6565) ) ;
INV     gate4929  (.A(g6565), .Z(II12725) ) ;
INV     gate4930  (.A(II12725), .Z(g6984) ) ;
OR2     gate4931  (.A(g6098), .B(g1975), .Z(g6579) ) ;
INV     gate4932  (.A(g6579), .Z(II12731) ) ;
INV     gate4933  (.A(II12731), .Z(g6993) ) ;
AND2    gate4934  (.A(g6178), .B(g2424), .Z(g6460) ) ;
INV     gate4935  (.A(g6460), .Z(II12737) ) ;
INV     gate4936  (.A(II12737), .Z(g6997) ) ;
OR2     gate4937  (.A(g3617), .B(g6153), .Z(g6590) ) ;
INV     gate4938  (.A(g6590), .Z(II12742) ) ;
INV     gate4939  (.A(II12742), .Z(g7000) ) ;
OR2     gate4940  (.A(g3617), .B(g6119), .Z(g6585) ) ;
INV     gate4941  (.A(g6585), .Z(II12748) ) ;
INV     gate4942  (.A(II12748), .Z(g7006) ) ;
OR2     gate4943  (.A(g6105), .B(g6107), .Z(g6445) ) ;
INV     gate4944  (.A(g6445), .Z(II12753) ) ;
INV     gate4945  (.A(II12753), .Z(g7009) ) ;
AND2    gate4946  (.A(g6142), .B(g4160), .Z(g6577) ) ;
INV     gate4947  (.A(g6577), .Z(II12757) ) ;
INV     gate4948  (.A(II12757), .Z(g7013) ) ;
OR2     gate4949  (.A(g4067), .B(g5969), .Z(g6685) ) ;
INV     gate4950  (.A(g6685), .Z(II12760) ) ;
INV     gate4951  (.A(II12760), .Z(g7014) ) ;
OR2     gate4952  (.A(g4068), .B(g5970), .Z(g6686) ) ;
INV     gate4953  (.A(g6686), .Z(II12763) ) ;
INV     gate4954  (.A(II12763), .Z(g7015) ) ;
OR2     gate4955  (.A(g4083), .B(g6006), .Z(g6718) ) ;
INV     gate4956  (.A(g6718), .Z(II12768) ) ;
INV     gate4957  (.A(II12768), .Z(g7018) ) ;
OR2     gate4958  (.A(g4091), .B(g6013), .Z(g6735) ) ;
INV     gate4959  (.A(g6735), .Z(II12771) ) ;
INV     gate4960  (.A(II12771), .Z(g7019) ) ;
OR2     gate4961  (.A(g4099), .B(g6021), .Z(g6739) ) ;
INV     gate4962  (.A(g6739), .Z(II12776) ) ;
INV     gate4963  (.A(II12776), .Z(g7022) ) ;
OR2     gate4964  (.A(g4100), .B(g6022), .Z(g6740) ) ;
INV     gate4965  (.A(g6740), .Z(II12779) ) ;
INV     gate4966  (.A(II12779), .Z(g7023) ) ;
NAND2   gate4967  (.A(g5918), .B(g5278), .Z(g6463) ) ;
INV     gate4968  (.A(g6463), .Z(II12782) ) ;
INV     gate4969  (.A(II12782), .Z(g7024) ) ;
INV     gate4970  (.A(g6525), .Z(g7028) ) ;
INV     gate4971  (.A(g6525), .Z(g7032) ) ;
INV     gate4972  (.A(g6525), .Z(g7034) ) ;
INV     gate4973  (.A(g6543), .Z(g7035) ) ;
INV     gate4974  (.A(g6525), .Z(g7037) ) ;
INV     gate4975  (.A(g6543), .Z(g7039) ) ;
INV     gate4976  (.A(g6543), .Z(g7042) ) ;
INV     gate4977  (.A(g6543), .Z(g7043) ) ;
INV     gate4978  (.A(g6543), .Z(g7044) ) ;
INV     gate4979  (.A(g6490), .Z(g7045) ) ;
OR2     gate4980  (.A(g6058), .B(g3092), .Z(g6602) ) ;
INV     gate4981  (.A(g6602), .Z(II12806) ) ;
INV     gate4982  (.A(II12806), .Z(g7046) ) ;
INV     gate4983  (.A(g6498), .Z(g7047) ) ;
INV     gate4984  (.A(g6607), .Z(II12810) ) ;
INV     gate4985  (.A(g6607), .Z(II12813) ) ;
INV     gate4986  (.A(II12813), .Z(g7049) ) ;
INV     gate4987  (.A(g6618), .Z(g7050) ) ;
INV     gate4988  (.A(g6511), .Z(g7054) ) ;
INV     gate4989  (.A(g6517), .Z(g7055) ) ;
INV     gate4990  (.A(g6520), .Z(g7056) ) ;
INV     gate4991  (.A(g6644), .Z(g7057) ) ;
INV     gate4992  (.A(g6649), .Z(g7058) ) ;
INV     gate4993  (.A(g6538), .Z(g7059) ) ;
INV     gate4994  (.A(g6654), .Z(g7060) ) ;
INV     gate4995  (.A(g6650), .Z(g7061) ) ;
INV     gate4996  (.A(g6441), .Z(II12826) ) ;
INV     gate4997  (.A(g6441), .Z(II12829) ) ;
INV     gate4998  (.A(II12829), .Z(g7064) ) ;
INV     gate4999  (.A(g6630), .Z(II12839) ) ;
INV     gate5000  (.A(II12839), .Z(g7066) ) ;
INV     gate5001  (.A(g6658), .Z(g7067) ) ;
INV     gate5002  (.A(g6556), .Z(g7068) ) ;
INV     gate5003  (.A(g6562), .Z(g7070) ) ;
INV     gate5004  (.A(g6676), .Z(g7077) ) ;
INV     gate5005  (.A(g6683), .Z(g7078) ) ;
INV     gate5006  (.A(g6525), .Z(g7090) ) ;
INV     gate5007  (.A(g6525), .Z(g7091) ) ;
INV     gate5008  (.A(g6483), .Z(II12866) ) ;
INV     gate5009  (.A(II12866), .Z(g7092) ) ;
INV     gate5010  (.A(g6525), .Z(g7094) ) ;
INV     gate5011  (.A(g6700), .Z(II12877) ) ;
INV     gate5012  (.A(II12877), .Z(g7095) ) ;
INV     gate5013  (.A(g6478), .Z(II12881) ) ;
INV     gate5014  (.A(II12881), .Z(g7097) ) ;
INV     gate5015  (.A(g6525), .Z(g7098) ) ;
INV     gate5016  (.A(g6946), .Z(II12885) ) ;
INV     gate5017  (.A(g6948), .Z(II12888) ) ;
INV     gate5018  (.A(g6950), .Z(II12891) ) ;
INV     gate5019  (.A(g7009), .Z(II12894) ) ;
INV     gate5020  (.A(g6962), .Z(II12897) ) ;
INV     gate5021  (.A(g6947), .Z(II12900) ) ;
INV     gate5022  (.A(g6905), .Z(II12903) ) ;
INV     gate5023  (.A(g6918), .Z(II12906) ) ;
INV     gate5024  (.A(g7046), .Z(II12909) ) ;
INV     gate5025  (.A(g7006), .Z(II12912) ) ;
INV     gate5026  (.A(g7000), .Z(II12915) ) ;
INV     gate5027  (.A(g7013), .Z(II12918) ) ;
INV     gate5028  (.A(g6993), .Z(II12921) ) ;
INV     gate5029  (.A(g6983), .Z(II12924) ) ;
INV     gate5030  (.A(g7014), .Z(II12927) ) ;
INV     gate5031  (.A(g7019), .Z(II12930) ) ;
INV     gate5032  (.A(g7018), .Z(II12933) ) ;
INV     gate5033  (.A(g7015), .Z(II12936) ) ;
INV     gate5034  (.A(g7022), .Z(II12939) ) ;
INV     gate5035  (.A(g7023), .Z(II12942) ) ;
INV     gate5036  (.A(g7066), .Z(II12945) ) ;
OR2     gate5037  (.A(g6771), .B(g6394), .Z(g6919) ) ;
INV     gate5038  (.A(g6919), .Z(II12948) ) ;
INV     gate5039  (.A(II12948), .Z(g7120) ) ;
OR2     gate5040  (.A(g6395), .B(g6399), .Z(g6920) ) ;
INV     gate5041  (.A(g6920), .Z(II12958) ) ;
INV     gate5042  (.A(II12958), .Z(g7122) ) ;
OR2     gate5043  (.A(g6396), .B(g6401), .Z(g6921) ) ;
INV     gate5044  (.A(g6921), .Z(II12961) ) ;
INV     gate5045  (.A(II12961), .Z(g7123) ) ;
INV     gate5046  (.A(g6896), .Z(g7124) ) ;
OR2     gate5047  (.A(g6400), .B(g6405), .Z(g6924) ) ;
INV     gate5048  (.A(g6924), .Z(II12965) ) ;
INV     gate5049  (.A(II12965), .Z(g7125) ) ;
OR2     gate5050  (.A(g6402), .B(g6407), .Z(g6925) ) ;
INV     gate5051  (.A(g6925), .Z(II12968) ) ;
INV     gate5052  (.A(II12968), .Z(g7126) ) ;
AND2    gate5053  (.A(g3613), .B(g6505), .Z(g6974) ) ;
INV     gate5054  (.A(g6974), .Z(g7127) ) ;
OR2     gate5055  (.A(g6408), .B(g6413), .Z(g6927) ) ;
INV     gate5056  (.A(g6927), .Z(II12973) ) ;
INV     gate5057  (.A(II12973), .Z(g7129) ) ;
OR2     gate5058  (.A(g6409), .B(g6415), .Z(g6928) ) ;
INV     gate5059  (.A(g6928), .Z(II12976) ) ;
INV     gate5060  (.A(II12976), .Z(g7130) ) ;
AND2    gate5061  (.A(g4399), .B(g6508), .Z(g6976) ) ;
INV     gate5062  (.A(g6976), .Z(g7131) ) ;
OR2     gate5063  (.A(g6412), .B(g6418), .Z(g6929) ) ;
INV     gate5064  (.A(g6929), .Z(II12980) ) ;
INV     gate5065  (.A(II12980), .Z(g7132) ) ;
OR2     gate5066  (.A(g6414), .B(g6420), .Z(g6930) ) ;
INV     gate5067  (.A(g6930), .Z(II12983) ) ;
INV     gate5068  (.A(II12983), .Z(g7133) ) ;
OR2     gate5069  (.A(g6416), .B(g6421), .Z(g6931) ) ;
INV     gate5070  (.A(g6931), .Z(II12986) ) ;
INV     gate5071  (.A(II12986), .Z(g7134) ) ;
OR2     gate5072  (.A(g6417), .B(g6423), .Z(g6932) ) ;
INV     gate5073  (.A(g6932), .Z(II12989) ) ;
INV     gate5074  (.A(II12989), .Z(g7135) ) ;
OR2     gate5075  (.A(g6419), .B(g6428), .Z(g6933) ) ;
INV     gate5076  (.A(g6933), .Z(II12993) ) ;
INV     gate5077  (.A(II12993), .Z(g7137) ) ;
OR2     gate5078  (.A(g6422), .B(g6430), .Z(g6934) ) ;
INV     gate5079  (.A(g6934), .Z(II12996) ) ;
INV     gate5080  (.A(II12996), .Z(g7138) ) ;
OR2     gate5081  (.A(g6433), .B(g5765), .Z(g7029) ) ;
INV     gate5082  (.A(g7029), .Z(II12999) ) ;
INV     gate5083  (.A(II12999), .Z(g7139) ) ;
OR2     gate5084  (.A(g6429), .B(g6431), .Z(g6935) ) ;
INV     gate5085  (.A(g6935), .Z(II13009) ) ;
INV     gate5086  (.A(II13009), .Z(g7141) ) ;
AND2    gate5087  (.A(g6639), .B(g1872), .Z(g7071) ) ;
INV     gate5088  (.A(g7071), .Z(II13012) ) ;
INV     gate5089  (.A(II13012), .Z(g7142) ) ;
AND2    gate5090  (.A(g3678), .B(g6552), .Z(g6996) ) ;
INV     gate5091  (.A(g6996), .Z(g7143) ) ;
OR2     gate5092  (.A(g6439), .B(g5783), .Z(g7040) ) ;
INV     gate5093  (.A(g7040), .Z(II13023) ) ;
INV     gate5094  (.A(II13023), .Z(g7145) ) ;
AND2    gate5095  (.A(g4474), .B(g6555), .Z(g6998) ) ;
INV     gate5096  (.A(g6998), .Z(g7146) ) ;
INV     gate5097  (.A(g6904), .Z(g7147) ) ;
AND2    gate5098  (.A(g6440), .B(g5311), .Z(g7087) ) ;
INV     gate5099  (.A(g7087), .Z(II13028) ) ;
INV     gate5100  (.A(II13028), .Z(g7148) ) ;
INV     gate5101  (.A(g6984), .Z(II13031) ) ;
INV     gate5102  (.A(II13031), .Z(g7149) ) ;
OR2     gate5103  (.A(g6633), .B(g6204), .Z(g6952) ) ;
INV     gate5104  (.A(g6952), .Z(g7150) ) ;
OR2     gate5105  (.A(g6447), .B(g6448), .Z(g6964) ) ;
INV     gate5106  (.A(g6964), .Z(II13035) ) ;
INV     gate5107  (.A(II13035), .Z(g7151) ) ;
INV     gate5108  (.A(g6961), .Z(II13039) ) ;
INV     gate5109  (.A(II13039), .Z(g7155) ) ;
INV     gate5110  (.A(g6963), .Z(II13042) ) ;
INV     gate5111  (.A(II13042), .Z(g7156) ) ;
INV     gate5112  (.A(g6955), .Z(II13045) ) ;
INV     gate5113  (.A(II13045), .Z(g7157) ) ;
INV     gate5114  (.A(g6956), .Z(II13048) ) ;
INV     gate5115  (.A(II13048), .Z(g7158) ) ;
INV     gate5116  (.A(g6967), .Z(II13051) ) ;
INV     gate5117  (.A(II13051), .Z(g7159) ) ;
INV     gate5118  (.A(g6960), .Z(II13054) ) ;
INV     gate5119  (.A(II13054), .Z(g7160) ) ;
INV     gate5120  (.A(g6968), .Z(II13057) ) ;
INV     gate5121  (.A(II13057), .Z(g7161) ) ;
INV     gate5122  (.A(g6959), .Z(II13060) ) ;
INV     gate5123  (.A(II13060), .Z(g7162) ) ;
INV     gate5124  (.A(g6973), .Z(II13063) ) ;
INV     gate5125  (.A(II13063), .Z(g7163) ) ;
INV     gate5126  (.A(g6957), .Z(II13066) ) ;
INV     gate5127  (.A(II13066), .Z(g7164) ) ;
INV     gate5128  (.A(g6969), .Z(II13072) ) ;
INV     gate5129  (.A(II13072), .Z(g7168) ) ;
INV     gate5130  (.A(g6958), .Z(II13075) ) ;
INV     gate5131  (.A(II13075), .Z(g7169) ) ;
INV     gate5132  (.A(g7071), .Z(g7171) ) ;
INV     gate5133  (.A(g7092), .Z(g7172) ) ;
OR2     gate5134  (.A(g6745), .B(g6028), .Z(g6980) ) ;
INV     gate5135  (.A(g6980), .Z(g7173) ) ;
INV     gate5136  (.A(g7097), .Z(g7174) ) ;
INV     gate5137  (.A(g7071), .Z(II13084) ) ;
INV     gate5138  (.A(II13084), .Z(g7176) ) ;
INV     gate5139  (.A(g7045), .Z(II13088) ) ;
INV     gate5140  (.A(II13088), .Z(g7178) ) ;
INV     gate5141  (.A(g7047), .Z(II13092) ) ;
INV     gate5142  (.A(II13092), .Z(g7180) ) ;
INV     gate5143  (.A(g7054), .Z(II13099) ) ;
INV     gate5144  (.A(II13099), .Z(g7185) ) ;
INV     gate5145  (.A(g7055), .Z(II13103) ) ;
INV     gate5146  (.A(II13103), .Z(g7187) ) ;
INV     gate5147  (.A(g7056), .Z(II13106) ) ;
INV     gate5148  (.A(II13106), .Z(g7188) ) ;
INV     gate5149  (.A(g7059), .Z(II13109) ) ;
INV     gate5150  (.A(II13109), .Z(g7189) ) ;
AND2    gate5151  (.A(g3390), .B(g6673), .Z(g7021) ) ;
INV     gate5152  (.A(g7021), .Z(II13112) ) ;
INV     gate5153  (.A(II13112), .Z(g7190) ) ;
INV     gate5154  (.A(g7068), .Z(II13118) ) ;
INV     gate5155  (.A(II13118), .Z(g7194) ) ;
INV     gate5156  (.A(g7070), .Z(II13122) ) ;
INV     gate5157  (.A(II13122), .Z(g7196) ) ;
AND2    gate5158  (.A(g5483), .B(g6589), .Z(g6949) ) ;
INV     gate5159  (.A(g6949), .Z(II13126) ) ;
INV     gate5160  (.A(II13126), .Z(g7198) ) ;
AND2    gate5161  (.A(g5511), .B(g6595), .Z(g6951) ) ;
INV     gate5162  (.A(g6951), .Z(II13131) ) ;
INV     gate5163  (.A(II13131), .Z(g7205) ) ;
AND2    gate5164  (.A(g3390), .B(g6706), .Z(g7017) ) ;
INV     gate5165  (.A(g7017), .Z(II13134) ) ;
INV     gate5166  (.A(II13134), .Z(g7206) ) ;
AND2    gate5167  (.A(g3390), .B(g6698), .Z(g7027) ) ;
INV     gate5168  (.A(g7027), .Z(II13137) ) ;
INV     gate5169  (.A(II13137), .Z(g7207) ) ;
AND2    gate5170  (.A(g5518), .B(g6601), .Z(g6954) ) ;
INV     gate5171  (.A(g6954), .Z(II13140) ) ;
INV     gate5172  (.A(II13140), .Z(g7208) ) ;
AND2    gate5173  (.A(g3390), .B(g6717), .Z(g7031) ) ;
INV     gate5174  (.A(g7031), .Z(II13144) ) ;
INV     gate5175  (.A(II13144), .Z(g7210) ) ;
INV     gate5176  (.A(g7024), .Z(II13147) ) ;
INV     gate5177  (.A(II13147), .Z(g7211) ) ;
AND2    gate5178  (.A(g6580), .B(g5580), .Z(g6966) ) ;
INV     gate5179  (.A(g6966), .Z(II13152) ) ;
INV     gate5180  (.A(II13152), .Z(g7216) ) ;
INV     gate5181  (.A(g6997), .Z(II13157) ) ;
INV     gate5182  (.A(II13157), .Z(g7221) ) ;
OR2     gate5183  (.A(g4086), .B(g6462), .Z(g7080) ) ;
INV     gate5184  (.A(g7080), .Z(II13161) ) ;
INV     gate5185  (.A(II13161), .Z(g7223) ) ;
OR2     gate5186  (.A(g4101), .B(g6464), .Z(g7086) ) ;
INV     gate5187  (.A(g7086), .Z(II13164) ) ;
INV     gate5188  (.A(II13164), .Z(g7224) ) ;
INV     gate5189  (.A(g6936), .Z(g7225) ) ;
INV     gate5190  (.A(g6937), .Z(g7226) ) ;
INV     gate5191  (.A(g6938), .Z(g7229) ) ;
OR2     gate5192  (.A(g4128), .B(g6474), .Z(g7089) ) ;
INV     gate5193  (.A(g7089), .Z(II13173) ) ;
INV     gate5194  (.A(II13173), .Z(g7231) ) ;
INV     gate5195  (.A(g6940), .Z(g7233) ) ;
INV     gate5196  (.A(g6944), .Z(g7236) ) ;
INV     gate5197  (.A(g6945), .Z(g7239) ) ;
OR2     gate5198  (.A(g3617), .B(g6578), .Z(g7020) ) ;
INV     gate5199  (.A(g7020), .Z(II13185) ) ;
INV     gate5200  (.A(II13185), .Z(g7241) ) ;
AND2    gate5201  (.A(g6770), .B(g5054), .Z(g7002) ) ;
INV     gate5202  (.A(g7002), .Z(II13189) ) ;
INV     gate5203  (.A(II13189), .Z(g7243) ) ;
AND2    gate5204  (.A(g6627), .B(g5072), .Z(g7007) ) ;
INV     gate5205  (.A(g7007), .Z(II13193) ) ;
INV     gate5206  (.A(II13193), .Z(g7245) ) ;
AND2    gate5207  (.A(g6615), .B(g5083), .Z(g7008) ) ;
INV     gate5208  (.A(g7008), .Z(II13196) ) ;
INV     gate5209  (.A(II13196), .Z(g7246) ) ;
OR2     gate5210  (.A(g6541), .B(g3095), .Z(g7025) ) ;
INV     gate5211  (.A(g7025), .Z(II13199) ) ;
INV     gate5212  (.A(II13199), .Z(g7247) ) ;
OR2     gate5213  (.A(g6638), .B(g6641), .Z(g7088) ) ;
INV     gate5214  (.A(g7088), .Z(II13203) ) ;
INV     gate5215  (.A(II13203), .Z(g7251) ) ;
INV     gate5216  (.A(g7049), .Z(g7253) ) ;
OR2     gate5217  (.A(g4199), .B(g6567), .Z(g6912) ) ;
INV     gate5218  (.A(g6912), .Z(II13209) ) ;
INV     gate5219  (.A(II13209), .Z(g7255) ) ;
INV     gate5220  (.A(g7058), .Z(g7256) ) ;
INV     gate5221  (.A(g7060), .Z(g7259) ) ;
INV     gate5222  (.A(g7064), .Z(g7260) ) ;
INV     gate5223  (.A(g7095), .Z(II13225) ) ;
INV     gate5224  (.A(II13225), .Z(g7261) ) ;
INV     gate5225  (.A(g6892), .Z(II13228) ) ;
INV     gate5226  (.A(II13228), .Z(g7262) ) ;
INV     gate5227  (.A(g6897), .Z(II13231) ) ;
INV     gate5228  (.A(II13231), .Z(g7263) ) ;
INV     gate5229  (.A(g6898), .Z(II13234) ) ;
INV     gate5230  (.A(II13234), .Z(g7264) ) ;
INV     gate5231  (.A(g7077), .Z(g7265) ) ;
INV     gate5232  (.A(g6900), .Z(II13238) ) ;
INV     gate5233  (.A(II13238), .Z(g7266) ) ;
AND2    gate5234  (.A(g6705), .B(g5723), .Z(g7030) ) ;
INV     gate5235  (.A(g7030), .Z(II13241) ) ;
INV     gate5236  (.A(II13241), .Z(g7267) ) ;
AND2    gate5237  (.A(g6716), .B(g5190), .Z(g7033) ) ;
INV     gate5238  (.A(g7033), .Z(II13244) ) ;
INV     gate5239  (.A(II13244), .Z(g7268) ) ;
OR2     gate5240  (.A(g6715), .B(g6726), .Z(g6906) ) ;
INV     gate5241  (.A(g6906), .Z(II13247) ) ;
INV     gate5242  (.A(II13247), .Z(g7269) ) ;
AND2    gate5243  (.A(g6728), .B(g5197), .Z(g7036) ) ;
INV     gate5244  (.A(g7036), .Z(II13250) ) ;
INV     gate5245  (.A(II13250), .Z(g7270) ) ;
INV     gate5246  (.A(g7057), .Z(II13255) ) ;
INV     gate5247  (.A(II13255), .Z(g7273) ) ;
OR2     gate5248  (.A(g6727), .B(g6732), .Z(g6907) ) ;
INV     gate5249  (.A(g6907), .Z(II13258) ) ;
INV     gate5250  (.A(II13258), .Z(g7274) ) ;
AND2    gate5251  (.A(g6734), .B(g5206), .Z(g7041) ) ;
INV     gate5252  (.A(g7041), .Z(II13261) ) ;
INV     gate5253  (.A(II13261), .Z(g7275) ) ;
INV     gate5254  (.A(g7061), .Z(II13264) ) ;
INV     gate5255  (.A(II13264), .Z(g7276) ) ;
OR2     gate5256  (.A(g6733), .B(g6738), .Z(g6913) ) ;
INV     gate5257  (.A(g6913), .Z(II13267) ) ;
INV     gate5258  (.A(II13267), .Z(g7277) ) ;
INV     gate5259  (.A(g7067), .Z(II13271) ) ;
INV     gate5260  (.A(II13271), .Z(g7279) ) ;
OR2     gate5261  (.A(g6743), .B(g6753), .Z(g6917) ) ;
INV     gate5262  (.A(g6917), .Z(II13274) ) ;
INV     gate5263  (.A(II13274), .Z(g7280) ) ;
INV     gate5264  (.A(g7078), .Z(II13277) ) ;
INV     gate5265  (.A(II13277), .Z(g7281) ) ;
INV     gate5266  (.A(g7155), .Z(II13281) ) ;
INV     gate5267  (.A(g7156), .Z(II13284) ) ;
INV     gate5268  (.A(g7157), .Z(II13287) ) ;
INV     gate5269  (.A(g7158), .Z(II13290) ) ;
INV     gate5270  (.A(g7159), .Z(II13293) ) ;
INV     gate5271  (.A(g7161), .Z(II13296) ) ;
INV     gate5272  (.A(g7163), .Z(II13299) ) ;
INV     gate5273  (.A(g7164), .Z(II13302) ) ;
INV     gate5274  (.A(g7168), .Z(II13305) ) ;
INV     gate5275  (.A(g7169), .Z(II13308) ) ;
INV     gate5276  (.A(g7162), .Z(II13311) ) ;
INV     gate5277  (.A(g7160), .Z(II13314) ) ;
INV     gate5278  (.A(g7211), .Z(II13317) ) ;
INV     gate5279  (.A(g7139), .Z(II13320) ) ;
INV     gate5280  (.A(g7145), .Z(II13323) ) ;
INV     gate5281  (.A(g7176), .Z(II13326) ) ;
INV     gate5282  (.A(g7247), .Z(II13329) ) ;
INV     gate5283  (.A(g7241), .Z(II13332) ) ;
INV     gate5284  (.A(g7206), .Z(II13335) ) ;
INV     gate5285  (.A(g7190), .Z(II13338) ) ;
INV     gate5286  (.A(g7207), .Z(II13341) ) ;
INV     gate5287  (.A(g7210), .Z(II13344) ) ;
INV     gate5288  (.A(g7224), .Z(II13347) ) ;
INV     gate5289  (.A(g7223), .Z(II13350) ) ;
INV     gate5290  (.A(g7231), .Z(II13353) ) ;
INV     gate5291  (.A(g7221), .Z(II13356) ) ;
INV     gate5292  (.A(g7255), .Z(II13359) ) ;
INV     gate5293  (.A(g7265), .Z(II13362) ) ;
INV     gate5294  (.A(II13362), .Z(g7310) ) ;
INV     gate5295  (.A(g7267), .Z(II13365) ) ;
INV     gate5296  (.A(II13365), .Z(g7311) ) ;
INV     gate5297  (.A(g7268), .Z(II13369) ) ;
INV     gate5298  (.A(II13369), .Z(g7313) ) ;
INV     gate5299  (.A(g7270), .Z(II13373) ) ;
INV     gate5300  (.A(II13373), .Z(g7315) ) ;
INV     gate5301  (.A(g7275), .Z(II13383) ) ;
INV     gate5302  (.A(II13383), .Z(g7317) ) ;
INV     gate5303  (.A(g7124), .Z(g7319) ) ;
INV     gate5304  (.A(g7149), .Z(II13388) ) ;
INV     gate5305  (.A(II13388), .Z(g7320) ) ;
INV     gate5306  (.A(g7269), .Z(II13403) ) ;
INV     gate5307  (.A(II13403), .Z(g7327) ) ;
AND2    gate5308  (.A(g6436), .B(g6922), .Z(g7271) ) ;
INV     gate5309  (.A(g7271), .Z(II13407) ) ;
INV     gate5310  (.A(II13407), .Z(g7329) ) ;
INV     gate5311  (.A(g7274), .Z(II13410) ) ;
INV     gate5312  (.A(II13410), .Z(g7330) ) ;
INV     gate5313  (.A(g7127), .Z(II13413) ) ;
INV     gate5314  (.A(II13413), .Z(g7331) ) ;
OR2     gate5315  (.A(g6434), .B(g6908), .Z(g7165) ) ;
INV     gate5316  (.A(g7165), .Z(II13416) ) ;
INV     gate5317  (.A(II13416), .Z(g7332) ) ;
INV     gate5318  (.A(g7277), .Z(II13419) ) ;
INV     gate5319  (.A(II13419), .Z(g7333) ) ;
INV     gate5320  (.A(g7131), .Z(II13422) ) ;
INV     gate5321  (.A(II13422), .Z(g7334) ) ;
OR2     gate5322  (.A(g6437), .B(g6914), .Z(g7166) ) ;
INV     gate5323  (.A(g7166), .Z(II13425) ) ;
INV     gate5324  (.A(II13425), .Z(g7335) ) ;
OR2     gate5325  (.A(g6438), .B(g6915), .Z(g7167) ) ;
INV     gate5326  (.A(g7167), .Z(II13428) ) ;
INV     gate5327  (.A(II13428), .Z(g7336) ) ;
INV     gate5328  (.A(g7280), .Z(II13432) ) ;
INV     gate5329  (.A(II13432), .Z(g7338) ) ;
OR2     gate5330  (.A(g6916), .B(g6444), .Z(g7170) ) ;
INV     gate5331  (.A(g7170), .Z(II13435) ) ;
INV     gate5332  (.A(II13435), .Z(g7339) ) ;
INV     gate5333  (.A(g7143), .Z(II13438) ) ;
INV     gate5334  (.A(II13438), .Z(g7340) ) ;
INV     gate5335  (.A(g7146), .Z(II13441) ) ;
INV     gate5336  (.A(II13441), .Z(g7341) ) ;
AND2    gate5337  (.A(g5830), .B(g6939), .Z(g7282) ) ;
INV     gate5338  (.A(g7282), .Z(II13444) ) ;
INV     gate5339  (.A(II13444), .Z(g7342) ) ;
INV     gate5340  (.A(g7261), .Z(II13447) ) ;
INV     gate5341  (.A(II13447), .Z(g7343) ) ;
INV     gate5342  (.A(g7150), .Z(g7344) ) ;
INV     gate5343  (.A(g7262), .Z(II13451) ) ;
INV     gate5344  (.A(II13451), .Z(g7345) ) ;
INV     gate5345  (.A(g7147), .Z(II13454) ) ;
INV     gate5346  (.A(II13454), .Z(g7346) ) ;
INV     gate5347  (.A(g7120), .Z(II13457) ) ;
INV     gate5348  (.A(II13457), .Z(g7347) ) ;
INV     gate5349  (.A(g7263), .Z(II13460) ) ;
INV     gate5350  (.A(II13460), .Z(g7348) ) ;
INV     gate5351  (.A(g7264), .Z(II13463) ) ;
INV     gate5352  (.A(II13463), .Z(g7349) ) ;
INV     gate5353  (.A(g7122), .Z(II13466) ) ;
INV     gate5354  (.A(II13466), .Z(g7350) ) ;
INV     gate5355  (.A(g7123), .Z(II13469) ) ;
INV     gate5356  (.A(II13469), .Z(g7351) ) ;
INV     gate5357  (.A(g7266), .Z(II13472) ) ;
INV     gate5358  (.A(II13472), .Z(g7352) ) ;
INV     gate5359  (.A(g7125), .Z(II13475) ) ;
INV     gate5360  (.A(II13475), .Z(g7353) ) ;
INV     gate5361  (.A(g7126), .Z(II13478) ) ;
INV     gate5362  (.A(II13478), .Z(g7354) ) ;
OR2     gate5363  (.A(g6923), .B(g5298), .Z(g7254) ) ;
INV     gate5364  (.A(g7254), .Z(II13481) ) ;
INV     gate5365  (.A(II13481), .Z(g7355) ) ;
AND2    gate5366  (.A(g6926), .B(g3047), .Z(g7128) ) ;
INV     gate5367  (.A(g7128), .Z(II13484) ) ;
INV     gate5368  (.A(II13484), .Z(g7356) ) ;
INV     gate5369  (.A(g7129), .Z(II13487) ) ;
INV     gate5370  (.A(II13487), .Z(g7357) ) ;
INV     gate5371  (.A(g7130), .Z(II13490) ) ;
INV     gate5372  (.A(II13490), .Z(g7358) ) ;
INV     gate5373  (.A(g7132), .Z(II13493) ) ;
INV     gate5374  (.A(II13493), .Z(g7359) ) ;
INV     gate5375  (.A(g7133), .Z(II13496) ) ;
INV     gate5376  (.A(II13496), .Z(g7360) ) ;
INV     gate5377  (.A(g7134), .Z(II13499) ) ;
INV     gate5378  (.A(II13499), .Z(g7361) ) ;
INV     gate5379  (.A(g7135), .Z(II13502) ) ;
INV     gate5380  (.A(II13502), .Z(g7362) ) ;
INV     gate5381  (.A(g7148), .Z(II13506) ) ;
INV     gate5382  (.A(II13506), .Z(g7364) ) ;
INV     gate5383  (.A(g7137), .Z(II13509) ) ;
INV     gate5384  (.A(II13509), .Z(g7365) ) ;
INV     gate5385  (.A(g7138), .Z(II13512) ) ;
INV     gate5386  (.A(II13512), .Z(g7366) ) ;
NOR3    gate5387  (.A(g6253), .B(g7083), .C(g5418), .Z(g7152) ) ;
INV     gate5388  (.A(g7152), .Z(II13515) ) ;
INV     gate5389  (.A(II13515), .Z(g7367) ) ;
INV     gate5390  (.A(g7141), .Z(II13518) ) ;
INV     gate5391  (.A(II13518), .Z(g7405) ) ;
OR2     gate5392  (.A(g6028), .B(g7071), .Z(g7202) ) ;
INV     gate5393  (.A(g7202), .Z(g7411) ) ;
INV     gate5394  (.A(g7151), .Z(II13524) ) ;
INV     gate5395  (.A(II13524), .Z(g7413) ) ;
AND2    gate5396  (.A(g1142), .B(g6941), .Z(g7217) ) ;
INV     gate5397  (.A(g7217), .Z(II13527) ) ;
INV     gate5398  (.A(II13527), .Z(g7414) ) ;
OR2     gate5399  (.A(g1304), .B(g7062), .Z(g7220) ) ;
INV     gate5400  (.A(g7220), .Z(II13533) ) ;
INV     gate5401  (.A(II13533), .Z(g7418) ) ;
INV     gate5402  (.A(g7152), .Z(II13537) ) ;
INV     gate5403  (.A(II13537), .Z(g7420) ) ;
NOR3    gate5404  (.A(g1789), .B(g146), .C(g6984), .Z(g7209) ) ;
INV     gate5405  (.A(g7209), .Z(II13541) ) ;
INV     gate5406  (.A(II13541), .Z(g7422) ) ;
INV     gate5407  (.A(g1167), .Z(II13544) ) ;
INV     gate5408  (.A(g1170), .Z(II13547) ) ;
INV     gate5409  (.A(g1173), .Z(II13550) ) ;
AND2    gate5410  (.A(g7016), .B(g5586), .Z(g7177) ) ;
INV     gate5411  (.A(g7177), .Z(II13559) ) ;
INV     gate5412  (.A(II13559), .Z(g7432) ) ;
AND2    gate5413  (.A(g6121), .B(g7035), .Z(g7179) ) ;
INV     gate5414  (.A(g7179), .Z(II13562) ) ;
INV     gate5415  (.A(II13562), .Z(g7433) ) ;
AND2    gate5416  (.A(g6124), .B(g7039), .Z(g7181) ) ;
INV     gate5417  (.A(g7181), .Z(II13565) ) ;
INV     gate5418  (.A(II13565), .Z(g7434) ) ;
INV     gate5419  (.A(g7198), .Z(II13570) ) ;
INV     gate5420  (.A(II13570), .Z(g7437) ) ;
INV     gate5421  (.A(g7205), .Z(II13574) ) ;
INV     gate5422  (.A(II13574), .Z(g7439) ) ;
AND2    gate5423  (.A(g6600), .B(g7044), .Z(g7186) ) ;
INV     gate5424  (.A(g7186), .Z(II13577) ) ;
INV     gate5425  (.A(II13577), .Z(g7440) ) ;
INV     gate5426  (.A(g7208), .Z(II13580) ) ;
INV     gate5427  (.A(II13580), .Z(g7441) ) ;
AND2    gate5428  (.A(g3591), .B(g6977), .Z(g7252) ) ;
INV     gate5429  (.A(g7252), .Z(II13583) ) ;
INV     gate5430  (.A(II13583), .Z(g7442) ) ;
INV     gate5431  (.A(g7216), .Z(II13595) ) ;
INV     gate5432  (.A(II13595), .Z(g7446) ) ;
AND2    gate5433  (.A(g7093), .B(g5055), .Z(g7197) ) ;
INV     gate5434  (.A(g7197), .Z(II13605) ) ;
INV     gate5435  (.A(II13605), .Z(g7448) ) ;
OR2     gate5436  (.A(g6992), .B(g3128), .Z(g7227) ) ;
INV     gate5437  (.A(g7227), .Z(II13610) ) ;
INV     gate5438  (.A(II13610), .Z(g7454) ) ;
INV     gate5439  (.A(g7273), .Z(II13613) ) ;
INV     gate5440  (.A(II13613), .Z(g7455) ) ;
INV     gate5441  (.A(g7174), .Z(g7456) ) ;
INV     gate5442  (.A(g7276), .Z(II13617) ) ;
INV     gate5443  (.A(II13617), .Z(g7459) ) ;
INV     gate5444  (.A(g7172), .Z(g7460) ) ;
INV     gate5445  (.A(g7239), .Z(g7463) ) ;
INV     gate5446  (.A(g7279), .Z(II13622) ) ;
INV     gate5447  (.A(II13622), .Z(g7466) ) ;
INV     gate5448  (.A(g7236), .Z(g7467) ) ;
INV     gate5449  (.A(g7253), .Z(g7470) ) ;
INV     gate5450  (.A(g7233), .Z(g7471) ) ;
OR2     gate5451  (.A(g7079), .B(g5652), .Z(g7248) ) ;
INV     gate5452  (.A(g7248), .Z(II13628) ) ;
INV     gate5453  (.A(g7248), .Z(II13631) ) ;
INV     gate5454  (.A(II13631), .Z(g7475) ) ;
INV     gate5455  (.A(g7229), .Z(g7476) ) ;
INV     gate5456  (.A(g7243), .Z(II13635) ) ;
INV     gate5457  (.A(II13635), .Z(g7479) ) ;
INV     gate5458  (.A(g7226), .Z(g7483) ) ;
INV     gate5459  (.A(g7245), .Z(II13646) ) ;
INV     gate5460  (.A(II13646), .Z(g7486) ) ;
INV     gate5461  (.A(g7281), .Z(II13649) ) ;
INV     gate5462  (.A(II13649), .Z(g7487) ) ;
INV     gate5463  (.A(g7225), .Z(g7488) ) ;
INV     gate5464  (.A(g7246), .Z(II13653) ) ;
INV     gate5465  (.A(II13653), .Z(g7491) ) ;
AND2    gate5466  (.A(g6688), .B(g7090), .Z(g7228) ) ;
INV     gate5467  (.A(g7228), .Z(II13656) ) ;
INV     gate5468  (.A(II13656), .Z(g7492) ) ;
AND2    gate5469  (.A(g6694), .B(g7091), .Z(g7232) ) ;
INV     gate5470  (.A(g7232), .Z(II13659) ) ;
INV     gate5471  (.A(II13659), .Z(g7493) ) ;
INV     gate5472  (.A(g7260), .Z(g7494) ) ;
AND2    gate5473  (.A(g6699), .B(g7094), .Z(g7235) ) ;
INV     gate5474  (.A(g7235), .Z(II13663) ) ;
INV     gate5475  (.A(II13663), .Z(g7495) ) ;
AND2    gate5476  (.A(g6707), .B(g7098), .Z(g7238) ) ;
INV     gate5477  (.A(g7238), .Z(II13666) ) ;
INV     gate5478  (.A(II13666), .Z(g7496) ) ;
AND2    gate5479  (.A(g6719), .B(g6894), .Z(g7240) ) ;
INV     gate5480  (.A(g7240), .Z(II13669) ) ;
INV     gate5481  (.A(II13669), .Z(g7497) ) ;
AND2    gate5482  (.A(g7081), .B(g6899), .Z(g7242) ) ;
INV     gate5483  (.A(g7242), .Z(II13672) ) ;
INV     gate5484  (.A(II13672), .Z(g7498) ) ;
OR3     gate5485  (.A(g7083), .B(g5403), .C(II13220), .Z(g7258) ) ;
INV     gate5486  (.A(g7258), .Z(g7499) ) ;
INV     gate5487  (.A(g7256), .Z(II13676) ) ;
INV     gate5488  (.A(II13676), .Z(g7500) ) ;
INV     gate5489  (.A(g7259), .Z(II13679) ) ;
INV     gate5490  (.A(II13679), .Z(g7501) ) ;
INV     gate5491  (.A(g7251), .Z(II13682) ) ;
INV     gate5492  (.A(II13682), .Z(g7502) ) ;
INV     gate5493  (.A(g7343), .Z(II13692) ) ;
INV     gate5494  (.A(g7345), .Z(II13695) ) ;
INV     gate5495  (.A(g7348), .Z(II13698) ) ;
INV     gate5496  (.A(g7349), .Z(II13701) ) ;
INV     gate5497  (.A(g7352), .Z(II13704) ) ;
INV     gate5498  (.A(g7420), .Z(II13707) ) ;
INV     gate5499  (.A(g7340), .Z(II13710) ) ;
INV     gate5500  (.A(g7341), .Z(II13713) ) ;
INV     gate5501  (.A(g7331), .Z(II13716) ) ;
INV     gate5502  (.A(g7334), .Z(II13719) ) ;
INV     gate5503  (.A(g7442), .Z(II13722) ) ;
INV     gate5504  (.A(g7437), .Z(II13725) ) ;
INV     gate5505  (.A(g7439), .Z(II13728) ) ;
INV     gate5506  (.A(g7441), .Z(II13731) ) ;
INV     gate5507  (.A(g7422), .Z(II13734) ) ;
INV     gate5508  (.A(g7446), .Z(II13737) ) ;
INV     gate5509  (.A(g7364), .Z(II13740) ) ;
INV     gate5510  (.A(g7454), .Z(II13743) ) ;
INV     gate5511  (.A(g7311), .Z(II13746) ) ;
INV     gate5512  (.A(g7313), .Z(II13749) ) ;
INV     gate5513  (.A(g7315), .Z(II13752) ) ;
INV     gate5514  (.A(g7317), .Z(II13755) ) ;
INV     gate5515  (.A(g7414), .Z(II13758) ) ;
INV     gate5516  (.A(g7418), .Z(II13761) ) ;
INV     gate5517  (.A(g7479), .Z(II13764) ) ;
INV     gate5518  (.A(g7486), .Z(II13767) ) ;
INV     gate5519  (.A(g7491), .Z(II13770) ) ;
INV     gate5520  (.A(g7496), .Z(II13773) ) ;
INV     gate5521  (.A(II13773), .Z(g7531) ) ;
INV     gate5522  (.A(g7497), .Z(II13776) ) ;
INV     gate5523  (.A(II13776), .Z(g7532) ) ;
NOR2    gate5524  (.A(g7191), .B(g1600), .Z(g7406) ) ;
INV     gate5525  (.A(g7406), .Z(II13779) ) ;
INV     gate5526  (.A(II13779), .Z(g7533) ) ;
INV     gate5527  (.A(g7498), .Z(II13782) ) ;
INV     gate5528  (.A(II13782), .Z(g7534) ) ;
INV     gate5529  (.A(g7346), .Z(II13794) ) ;
INV     gate5530  (.A(II13794), .Z(g7538) ) ;
INV     gate5531  (.A(g7502), .Z(II13797) ) ;
INV     gate5532  (.A(II13797), .Z(g7539) ) ;
INV     gate5533  (.A(g7320), .Z(II13807) ) ;
INV     gate5534  (.A(II13807), .Z(g7541) ) ;
NOR2    gate5535  (.A(g7178), .B(g6970), .Z(g7312) ) ;
INV     gate5536  (.A(g7312), .Z(II13810) ) ;
INV     gate5537  (.A(II13810), .Z(g7542) ) ;
NOR2    gate5538  (.A(g7180), .B(g6972), .Z(g7314) ) ;
INV     gate5539  (.A(g7314), .Z(II13813) ) ;
INV     gate5540  (.A(II13813), .Z(g7543) ) ;
INV     gate5541  (.A(g7455), .Z(II13816) ) ;
INV     gate5542  (.A(II13816), .Z(g7544) ) ;
OR3     gate5543  (.A(g1173), .B(g7217), .C(II13553), .Z(g7426) ) ;
INV     gate5544  (.A(g7426), .Z(II13819) ) ;
INV     gate5545  (.A(II13819), .Z(g7545) ) ;
INV     gate5546  (.A(g7459), .Z(II13822) ) ;
INV     gate5547  (.A(II13822), .Z(g7546) ) ;
NOR2    gate5548  (.A(g7185), .B(g6979), .Z(g7318) ) ;
INV     gate5549  (.A(g7318), .Z(II13825) ) ;
INV     gate5550  (.A(II13825), .Z(g7547) ) ;
NOR2    gate5551  (.A(g7187), .B(g6990), .Z(g7321) ) ;
INV     gate5552  (.A(g7321), .Z(II13828) ) ;
INV     gate5553  (.A(II13828), .Z(g7548) ) ;
NOR2    gate5554  (.A(g7188), .B(g6991), .Z(g7322) ) ;
INV     gate5555  (.A(g7322), .Z(II13831) ) ;
INV     gate5556  (.A(II13831), .Z(g7549) ) ;
INV     gate5557  (.A(g7466), .Z(II13834) ) ;
INV     gate5558  (.A(II13834), .Z(g7550) ) ;
NOR2    gate5559  (.A(g7189), .B(g6994), .Z(g7324) ) ;
INV     gate5560  (.A(g7324), .Z(II13837) ) ;
INV     gate5561  (.A(II13837), .Z(g7551) ) ;
NOR2    gate5562  (.A(g7194), .B(g6999), .Z(g7326) ) ;
INV     gate5563  (.A(g7326), .Z(II13843) ) ;
INV     gate5564  (.A(II13843), .Z(g7555) ) ;
INV     gate5565  (.A(g7487), .Z(II13846) ) ;
INV     gate5566  (.A(II13846), .Z(g7556) ) ;
NOR2    gate5567  (.A(g7196), .B(g7001), .Z(g7328) ) ;
INV     gate5568  (.A(g7328), .Z(II13850) ) ;
INV     gate5569  (.A(II13850), .Z(g7558) ) ;
INV     gate5570  (.A(g7327), .Z(II13854) ) ;
INV     gate5571  (.A(II13854), .Z(g7560) ) ;
INV     gate5572  (.A(g7329), .Z(II13858) ) ;
INV     gate5573  (.A(II13858), .Z(g7562) ) ;
INV     gate5574  (.A(g7330), .Z(II13861) ) ;
INV     gate5575  (.A(II13861), .Z(g7563) ) ;
INV     gate5576  (.A(g7333), .Z(II13865) ) ;
INV     gate5577  (.A(II13865), .Z(g7565) ) ;
INV     gate5578  (.A(g7338), .Z(II13869) ) ;
INV     gate5579  (.A(II13869), .Z(g7574) ) ;
INV     gate5580  (.A(g7342), .Z(II13873) ) ;
INV     gate5581  (.A(II13873), .Z(g7576) ) ;
INV     gate5582  (.A(g7347), .Z(II13876) ) ;
INV     gate5583  (.A(II13876), .Z(g7577) ) ;
INV     gate5584  (.A(g7332), .Z(II13879) ) ;
INV     gate5585  (.A(II13879), .Z(g7578) ) ;
INV     gate5586  (.A(g7350), .Z(II13882) ) ;
INV     gate5587  (.A(II13882), .Z(g7579) ) ;
INV     gate5588  (.A(g7351), .Z(II13885) ) ;
INV     gate5589  (.A(II13885), .Z(g7580) ) ;
INV     gate5590  (.A(g7335), .Z(II13888) ) ;
INV     gate5591  (.A(II13888), .Z(g7581) ) ;
INV     gate5592  (.A(g7336), .Z(II13891) ) ;
INV     gate5593  (.A(II13891), .Z(g7582) ) ;
INV     gate5594  (.A(g7353), .Z(II13894) ) ;
INV     gate5595  (.A(II13894), .Z(g7583) ) ;
INV     gate5596  (.A(g7354), .Z(II13897) ) ;
INV     gate5597  (.A(II13897), .Z(g7584) ) ;
INV     gate5598  (.A(g7356), .Z(II13900) ) ;
INV     gate5599  (.A(II13900), .Z(g7585) ) ;
INV     gate5600  (.A(g7357), .Z(II13903) ) ;
INV     gate5601  (.A(II13903), .Z(g7586) ) ;
INV     gate5602  (.A(g7358), .Z(II13906) ) ;
INV     gate5603  (.A(II13906), .Z(g7587) ) ;
INV     gate5604  (.A(g7339), .Z(II13909) ) ;
INV     gate5605  (.A(II13909), .Z(g7588) ) ;
INV     gate5606  (.A(g7359), .Z(II13912) ) ;
INV     gate5607  (.A(II13912), .Z(g7589) ) ;
INV     gate5608  (.A(g7360), .Z(II13915) ) ;
INV     gate5609  (.A(II13915), .Z(g7590) ) ;
INV     gate5610  (.A(g7361), .Z(II13918) ) ;
INV     gate5611  (.A(II13918), .Z(g7591) ) ;
INV     gate5612  (.A(g7362), .Z(II13921) ) ;
INV     gate5613  (.A(II13921), .Z(g7592) ) ;
INV     gate5614  (.A(g7365), .Z(II13924) ) ;
INV     gate5615  (.A(II13924), .Z(g7593) ) ;
INV     gate5616  (.A(g7366), .Z(II13927) ) ;
INV     gate5617  (.A(II13927), .Z(g7594) ) ;
INV     gate5618  (.A(g7405), .Z(II13930) ) ;
INV     gate5619  (.A(II13930), .Z(g7595) ) ;
OR2     gate5620  (.A(g6090), .B(g7195), .Z(g7450) ) ;
INV     gate5621  (.A(g7450), .Z(g7599) ) ;
INV     gate5622  (.A(g7450), .Z(g7601) ) ;
INV     gate5623  (.A(g7355), .Z(II13940) ) ;
INV     gate5624  (.A(II13940), .Z(g7603) ) ;
INV     gate5625  (.A(g7450), .Z(g7610) ) ;
INV     gate5626  (.A(g7499), .Z(II13956) ) ;
INV     gate5627  (.A(II13956), .Z(g7627) ) ;
INV     gate5628  (.A(g7413), .Z(II13962) ) ;
INV     gate5629  (.A(II13962), .Z(g7633) ) ;
AND2    gate5630  (.A(g7222), .B(g5603), .Z(g7415) ) ;
INV     gate5631  (.A(g7415), .Z(II13979) ) ;
INV     gate5632  (.A(II13979), .Z(g7686) ) ;
INV     gate5633  (.A(g7406), .Z(g7688) ) ;
INV     gate5634  (.A(g7432), .Z(II13997) ) ;
INV     gate5635  (.A(II13997), .Z(g7702) ) ;
INV     gate5636  (.A(g7433), .Z(II14001) ) ;
INV     gate5637  (.A(II14001), .Z(g7704) ) ;
INV     gate5638  (.A(g7434), .Z(II14005) ) ;
INV     gate5639  (.A(II14005), .Z(g7708) ) ;
OR2     gate5640  (.A(g7183), .B(g6975), .Z(g7436) ) ;
INV     gate5641  (.A(g7436), .Z(II14009) ) ;
INV     gate5642  (.A(II14009), .Z(g7710) ) ;
OR2     gate5643  (.A(g7184), .B(g6978), .Z(g7438) ) ;
INV     gate5644  (.A(g7438), .Z(II14012) ) ;
INV     gate5645  (.A(II14012), .Z(g7711) ) ;
INV     gate5646  (.A(g7440), .Z(II14015) ) ;
INV     gate5647  (.A(II14015), .Z(g7712) ) ;
NAND2   gate5648  (.A(II13639), .B(II13640), .Z(g7480) ) ;
INV     gate5649  (.A(g7480), .Z(II14019) ) ;
INV     gate5650  (.A(II14019), .Z(g7714) ) ;
OR2     gate5651  (.A(g7192), .B(g3158), .Z(g7443) ) ;
INV     gate5652  (.A(g7443), .Z(II14022) ) ;
INV     gate5653  (.A(II14022), .Z(g7715) ) ;
INV     gate5654  (.A(g7500), .Z(II14025) ) ;
INV     gate5655  (.A(II14025), .Z(g7716) ) ;
INV     gate5656  (.A(g7501), .Z(II14028) ) ;
INV     gate5657  (.A(II14028), .Z(g7717) ) ;
INV     gate5658  (.A(g7448), .Z(II14031) ) ;
INV     gate5659  (.A(II14031), .Z(g7718) ) ;
INV     gate5660  (.A(g7475), .Z(g7719) ) ;
INV     gate5661  (.A(g7310), .Z(II14035) ) ;
INV     gate5662  (.A(II14035), .Z(g7720) ) ;
INV     gate5663  (.A(g7344), .Z(g7721) ) ;
AND2    gate5664  (.A(g7272), .B(g6901), .Z(g7449) ) ;
INV     gate5665  (.A(g7449), .Z(II14039) ) ;
INV     gate5666  (.A(II14039), .Z(g7722) ) ;
INV     gate5667  (.A(g7470), .Z(II14042) ) ;
INV     gate5668  (.A(II14042), .Z(g7723) ) ;
INV     gate5669  (.A(g7492), .Z(II14046) ) ;
INV     gate5670  (.A(II14046), .Z(g7725) ) ;
INV     gate5671  (.A(g7493), .Z(II14049) ) ;
INV     gate5672  (.A(II14049), .Z(g7726) ) ;
INV     gate5673  (.A(g7494), .Z(II14052) ) ;
INV     gate5674  (.A(II14052), .Z(g7727) ) ;
INV     gate5675  (.A(g7495), .Z(II14055) ) ;
INV     gate5676  (.A(II14055), .Z(g7728) ) ;
INV     gate5677  (.A(g7544), .Z(II14058) ) ;
INV     gate5678  (.A(g7546), .Z(II14061) ) ;
INV     gate5679  (.A(g7556), .Z(II14064) ) ;
INV     gate5680  (.A(g7550), .Z(II14067) ) ;
INV     gate5681  (.A(g7714), .Z(II14070) ) ;
INV     gate5682  (.A(g7627), .Z(II14073) ) ;
INV     gate5683  (.A(g7577), .Z(II14076) ) ;
INV     gate5684  (.A(g7579), .Z(II14079) ) ;
INV     gate5685  (.A(g7539), .Z(II14082) ) ;
INV     gate5686  (.A(g7583), .Z(II14085) ) ;
INV     gate5687  (.A(g7585), .Z(II14088) ) ;
INV     gate5688  (.A(g7589), .Z(II14091) ) ;
INV     gate5689  (.A(g7593), .Z(II14094) ) ;
INV     gate5690  (.A(g7595), .Z(II14097) ) ;
INV     gate5691  (.A(g7580), .Z(II14100) ) ;
INV     gate5692  (.A(g7584), .Z(II14103) ) ;
INV     gate5693  (.A(g7586), .Z(II14106) ) ;
INV     gate5694  (.A(g7590), .Z(II14109) ) ;
INV     gate5695  (.A(g7560), .Z(II14112) ) ;
INV     gate5696  (.A(g7563), .Z(II14115) ) ;
INV     gate5697  (.A(g7565), .Z(II14118) ) ;
INV     gate5698  (.A(g7587), .Z(II14121) ) ;
INV     gate5699  (.A(g7591), .Z(II14124) ) ;
INV     gate5700  (.A(g7594), .Z(II14127) ) ;
INV     gate5701  (.A(g7592), .Z(II14130) ) ;
INV     gate5702  (.A(g7574), .Z(II14133) ) ;
INV     gate5703  (.A(g7633), .Z(II14136) ) ;
INV     gate5704  (.A(g7548), .Z(II14139) ) ;
INV     gate5705  (.A(g7551), .Z(II14142) ) ;
INV     gate5706  (.A(g7542), .Z(II14145) ) ;
INV     gate5707  (.A(g7543), .Z(II14148) ) ;
INV     gate5708  (.A(g7555), .Z(II14151) ) ;
INV     gate5709  (.A(g7558), .Z(II14154) ) ;
INV     gate5710  (.A(g7547), .Z(II14157) ) ;
INV     gate5711  (.A(g7549), .Z(II14160) ) ;
INV     gate5712  (.A(g7533), .Z(II14163) ) ;
INV     gate5713  (.A(g7702), .Z(II14166) ) ;
INV     gate5714  (.A(g7715), .Z(II14169) ) ;
INV     gate5715  (.A(g7545), .Z(II14172) ) ;
INV     gate5716  (.A(g7718), .Z(II14175) ) ;
INV     gate5717  (.A(g7562), .Z(II14178) ) ;
INV     gate5718  (.A(g7725), .Z(II14181) ) ;
INV     gate5719  (.A(g7726), .Z(II14184) ) ;
INV     gate5720  (.A(g7728), .Z(II14187) ) ;
INV     gate5721  (.A(g7531), .Z(II14190) ) ;
INV     gate5722  (.A(g7532), .Z(II14193) ) ;
INV     gate5723  (.A(g7534), .Z(II14196) ) ;
INV     gate5724  (.A(g7704), .Z(II14199) ) ;
INV     gate5725  (.A(g7708), .Z(II14202) ) ;
INV     gate5726  (.A(g7710), .Z(II14205) ) ;
INV     gate5727  (.A(g7711), .Z(II14208) ) ;
INV     gate5728  (.A(g7712), .Z(II14211) ) ;
INV     gate5729  (.A(g7576), .Z(II14214) ) ;
INV     gate5730  (.A(g7722), .Z(II14224) ) ;
INV     gate5731  (.A(II14224), .Z(g7789) ) ;
AND2    gate5732  (.A(g7319), .B(g5749), .Z(g7552) ) ;
INV     gate5733  (.A(g7552), .Z(II14227) ) ;
INV     gate5734  (.A(II14227), .Z(g7790) ) ;
NOR2    gate5735  (.A(g7421), .B(g1597), .Z(g7566) ) ;
INV     gate5736  (.A(g7566), .Z(II14231) ) ;
INV     gate5737  (.A(II14231), .Z(g7792) ) ;
AND2    gate5738  (.A(g7367), .B(g4176), .Z(g7614) ) ;
INV     gate5739  (.A(g7614), .Z(II14234) ) ;
INV     gate5740  (.A(II14234), .Z(g7793) ) ;
AND2    gate5741  (.A(g7367), .B(g4169), .Z(g7608) ) ;
INV     gate5742  (.A(g7608), .Z(II14238) ) ;
INV     gate5743  (.A(II14238), .Z(g7811) ) ;
INV     gate5744  (.A(g7541), .Z(II14251) ) ;
INV     gate5745  (.A(II14251), .Z(g7829) ) ;
INV     gate5746  (.A(g7716), .Z(II14257) ) ;
INV     gate5747  (.A(II14257), .Z(g7835) ) ;
INV     gate5748  (.A(g7717), .Z(II14260) ) ;
INV     gate5749  (.A(II14260), .Z(g7836) ) ;
AND2    gate5750  (.A(g7367), .B(g4483), .Z(g7698) ) ;
INV     gate5751  (.A(g7698), .Z(II14264) ) ;
INV     gate5752  (.A(II14264), .Z(g7838) ) ;
AND2    gate5753  (.A(g7367), .B(g4466), .Z(g7695) ) ;
INV     gate5754  (.A(g7695), .Z(II14267) ) ;
INV     gate5755  (.A(II14267), .Z(g7855) ) ;
AND2    gate5756  (.A(g7367), .B(g4504), .Z(g7703) ) ;
INV     gate5757  (.A(g7703), .Z(II14270) ) ;
INV     gate5758  (.A(II14270), .Z(g7870) ) ;
AND2    gate5759  (.A(g7367), .B(g4187), .Z(g7631) ) ;
INV     gate5760  (.A(g7631), .Z(II14273) ) ;
INV     gate5761  (.A(II14273), .Z(g7887) ) ;
INV     gate5762  (.A(g7720), .Z(II14276) ) ;
INV     gate5763  (.A(II14276), .Z(g7904) ) ;
AND2    gate5764  (.A(g7367), .B(g4494), .Z(g7700) ) ;
INV     gate5765  (.A(g7700), .Z(II14279) ) ;
INV     gate5766  (.A(II14279), .Z(g7905) ) ;
AND2    gate5767  (.A(g7367), .B(g4529), .Z(g7709) ) ;
INV     gate5768  (.A(g7709), .Z(II14282) ) ;
INV     gate5769  (.A(II14282), .Z(g7920) ) ;
AND2    gate5770  (.A(g7367), .B(g4182), .Z(g7625) ) ;
INV     gate5771  (.A(g7625), .Z(II14285) ) ;
INV     gate5772  (.A(II14285), .Z(g7937) ) ;
AND2    gate5773  (.A(g7367), .B(g4514), .Z(g7705) ) ;
INV     gate5774  (.A(g7705), .Z(II14288) ) ;
INV     gate5775  (.A(II14288), .Z(g7951) ) ;
AND2    gate5776  (.A(g7367), .B(g4166), .Z(g7680) ) ;
INV     gate5777  (.A(g7680), .Z(II14291) ) ;
INV     gate5778  (.A(II14291), .Z(g7966) ) ;
AND2    gate5779  (.A(g7367), .B(g4135), .Z(g7553) ) ;
INV     gate5780  (.A(g7553), .Z(II14294) ) ;
INV     gate5781  (.A(II14294), .Z(g7983) ) ;
AND2    gate5782  (.A(g7367), .B(g4147), .Z(g7557) ) ;
INV     gate5783  (.A(g7557), .Z(g7992) ) ;
AND2    gate5784  (.A(g7367), .B(g4158), .Z(g7678) ) ;
INV     gate5785  (.A(g7678), .Z(II14298) ) ;
INV     gate5786  (.A(II14298), .Z(g7993) ) ;
AND2    gate5787  (.A(g7367), .B(g4155), .Z(g7559) ) ;
INV     gate5788  (.A(g7559), .Z(g8008) ) ;
AND2    gate5789  (.A(g7363), .B(g7411), .Z(g7537) ) ;
INV     gate5790  (.A(g7537), .Z(II14305) ) ;
INV     gate5791  (.A(II14305), .Z(g8012) ) ;
AND2    gate5792  (.A(g7367), .B(g4163), .Z(g7561) ) ;
INV     gate5793  (.A(g7561), .Z(g8013) ) ;
AND2    gate5794  (.A(g7367), .B(g4172), .Z(g7564) ) ;
INV     gate5795  (.A(g7564), .Z(g8014) ) ;
AND2    gate5796  (.A(g7367), .B(g4417), .Z(g7689) ) ;
INV     gate5797  (.A(g7689), .Z(g8015) ) ;
INV     gate5798  (.A(g7566), .Z(II14311) ) ;
INV     gate5799  (.A(II14311), .Z(g8016) ) ;
AND2    gate5800  (.A(g7367), .B(g4430), .Z(g7692) ) ;
INV     gate5801  (.A(g7692), .Z(g8017) ) ;
AND2    gate5802  (.A(g7367), .B(g4216), .Z(g7676) ) ;
INV     gate5803  (.A(g7676), .Z(II14315) ) ;
INV     gate5804  (.A(II14315), .Z(g8018) ) ;
AND2    gate5805  (.A(g7367), .B(g4201), .Z(g7657) ) ;
INV     gate5806  (.A(g7657), .Z(II14318) ) ;
INV     gate5807  (.A(II14318), .Z(g8029) ) ;
AND2    gate5808  (.A(g7367), .B(g4448), .Z(g7694) ) ;
INV     gate5809  (.A(g7694), .Z(g8038) ) ;
AND2    gate5810  (.A(g7367), .B(g4469), .Z(g7696) ) ;
INV     gate5811  (.A(g7696), .Z(g8039) ) ;
AND2    gate5812  (.A(g7367), .B(g4486), .Z(g7699) ) ;
INV     gate5813  (.A(g7699), .Z(g8040) ) ;
AND2    gate5814  (.A(g7367), .B(g4497), .Z(g7701) ) ;
INV     gate5815  (.A(g7701), .Z(g8041) ) ;
AND2    gate5816  (.A(g4403), .B(g7367), .Z(g7713) ) ;
INV     gate5817  (.A(g7713), .Z(II14325) ) ;
INV     gate5818  (.A(II14325), .Z(g8042) ) ;
INV     gate5819  (.A(g7538), .Z(II14330) ) ;
INV     gate5820  (.A(II14330), .Z(g8061) ) ;
INV     gate5821  (.A(g7578), .Z(II14334) ) ;
INV     gate5822  (.A(II14334), .Z(g8063) ) ;
INV     gate5823  (.A(g7581), .Z(II14338) ) ;
INV     gate5824  (.A(II14338), .Z(g8065) ) ;
INV     gate5825  (.A(g7582), .Z(II14342) ) ;
INV     gate5826  (.A(II14342), .Z(g8067) ) ;
INV     gate5827  (.A(g7588), .Z(II14349) ) ;
INV     gate5828  (.A(II14349), .Z(g8072) ) ;
INV     gate5829  (.A(g7603), .Z(II14370) ) ;
INV     gate5830  (.A(II14370), .Z(g8093) ) ;
INV     gate5831  (.A(g7705), .Z(g8094) ) ;
AND2    gate5832  (.A(g7367), .B(g4445), .Z(g7693) ) ;
INV     gate5833  (.A(g7693), .Z(II14374) ) ;
INV     gate5834  (.A(II14374), .Z(g8111) ) ;
AND2    gate5835  (.A(g7367), .B(g4427), .Z(g7691) ) ;
INV     gate5836  (.A(g7691), .Z(II14378) ) ;
INV     gate5837  (.A(II14378), .Z(g8131) ) ;
AND2    gate5838  (.A(g7428), .B(g7028), .Z(g7596) ) ;
INV     gate5839  (.A(g7596), .Z(II14381) ) ;
INV     gate5840  (.A(II14381), .Z(g8145) ) ;
AND2    gate5841  (.A(g7435), .B(g5607), .Z(g7605) ) ;
INV     gate5842  (.A(g7605), .Z(II14388) ) ;
INV     gate5843  (.A(II14388), .Z(g8152) ) ;
AND2    gate5844  (.A(g4414), .B(g7367), .Z(g7536) ) ;
INV     gate5845  (.A(g7536), .Z(II14394) ) ;
INV     gate5846  (.A(II14394), .Z(g8156) ) ;
INV     gate5847  (.A(g7686), .Z(II14397) ) ;
INV     gate5848  (.A(II14397), .Z(g8172) ) ;
AND2    gate5849  (.A(g7503), .B(g5073), .Z(g7677) ) ;
INV     gate5850  (.A(g7677), .Z(II14400) ) ;
INV     gate5851  (.A(II14400), .Z(g8173) ) ;
AND2    gate5852  (.A(g7447), .B(g5084), .Z(g7679) ) ;
INV     gate5853  (.A(g7679), .Z(II14403) ) ;
INV     gate5854  (.A(II14403), .Z(g8174) ) ;
AND2    gate5855  (.A(g7444), .B(g5099), .Z(g7681) ) ;
INV     gate5856  (.A(g7681), .Z(II14406) ) ;
INV     gate5857  (.A(II14406), .Z(g8175) ) ;
OR2     gate5858  (.A(g7419), .B(g3187), .Z(g7697) ) ;
INV     gate5859  (.A(g7697), .Z(II14410) ) ;
INV     gate5860  (.A(II14410), .Z(g8177) ) ;
INV     gate5861  (.A(g7723), .Z(II14413) ) ;
INV     gate5862  (.A(II14413), .Z(g8178) ) ;
INV     gate5863  (.A(g7727), .Z(II14416) ) ;
INV     gate5864  (.A(II14416), .Z(g8179) ) ;
INV     gate5865  (.A(g7719), .Z(g8180) ) ;
AND2    gate5866  (.A(g7367), .B(g4139), .Z(g7554) ) ;
INV     gate5867  (.A(g7554), .Z(II14420) ) ;
INV     gate5868  (.A(II14420), .Z(g8181) ) ;
INV     gate5869  (.A(g7721), .Z(g8198) ) ;
AND2    gate5870  (.A(g7367), .B(g4194), .Z(g7652) ) ;
INV     gate5871  (.A(g7652), .Z(II14424) ) ;
INV     gate5872  (.A(II14424), .Z(g8199) ) ;
INV     gate5873  (.A(g7835), .Z(II14427) ) ;
INV     gate5874  (.A(g7836), .Z(II14430) ) ;
INV     gate5875  (.A(g8061), .Z(II14433) ) ;
INV     gate5876  (.A(g7904), .Z(II14436) ) ;
INV     gate5877  (.A(g8063), .Z(II14439) ) ;
INV     gate5878  (.A(g8065), .Z(II14442) ) ;
INV     gate5879  (.A(g8067), .Z(II14445) ) ;
INV     gate5880  (.A(g7792), .Z(II14448) ) ;
INV     gate5881  (.A(g8172), .Z(II14451) ) ;
INV     gate5882  (.A(g8177), .Z(II14454) ) ;
INV     gate5883  (.A(g8093), .Z(II14457) ) ;
INV     gate5884  (.A(g7789), .Z(II14460) ) ;
INV     gate5885  (.A(g8072), .Z(II14463) ) ;
INV     gate5886  (.A(g7829), .Z(II14489) ) ;
INV     gate5887  (.A(g7829), .Z(II14492) ) ;
INV     gate5888  (.A(II14492), .Z(g8235) ) ;
INV     gate5889  (.A(g8178), .Z(II14531) ) ;
INV     gate5890  (.A(II14531), .Z(g8284) ) ;
INV     gate5891  (.A(g8179), .Z(II14573) ) ;
INV     gate5892  (.A(II14573), .Z(g8324) ) ;
INV     gate5893  (.A(g8008), .Z(g8342) ) ;
INV     gate5894  (.A(g7992), .Z(g8363) ) ;
AND2    gate5895  (.A(g7575), .B(g7173), .Z(g7827) ) ;
INV     gate5896  (.A(g7827), .Z(II14603) ) ;
INV     gate5897  (.A(II14603), .Z(g8381) ) ;
INV     gate5898  (.A(g8014), .Z(g8386) ) ;
AND2    gate5899  (.A(g5343), .B(g7599), .Z(g7832) ) ;
INV     gate5900  (.A(g7832), .Z(II14614) ) ;
INV     gate5901  (.A(II14614), .Z(g8406) ) ;
INV     gate5902  (.A(g8013), .Z(g8407) ) ;
INV     gate5903  (.A(g8017), .Z(g8421) ) ;
AND2    gate5904  (.A(g6461), .B(g7601), .Z(g7833) ) ;
INV     gate5905  (.A(g7833), .Z(II14623) ) ;
INV     gate5906  (.A(II14623), .Z(g8442) ) ;
INV     gate5907  (.A(g8015), .Z(g8443) ) ;
INV     gate5908  (.A(g8094), .Z(g8463) ) ;
INV     gate5909  (.A(g8039), .Z(g8464) ) ;
INV     gate5910  (.A(g8012), .Z(II14637) ) ;
INV     gate5911  (.A(II14637), .Z(g8481) ) ;
INV     gate5912  (.A(g8094), .Z(g8482) ) ;
INV     gate5913  (.A(g8038), .Z(g8483) ) ;
INV     gate5914  (.A(g8041), .Z(g8493) ) ;
AND2    gate5915  (.A(g6470), .B(g7610), .Z(g7837) ) ;
INV     gate5916  (.A(g7837), .Z(II14643) ) ;
INV     gate5917  (.A(II14643), .Z(g8510) ) ;
INV     gate5918  (.A(g7790), .Z(II14646) ) ;
INV     gate5919  (.A(II14646), .Z(g8511) ) ;
INV     gate5920  (.A(g8094), .Z(g8512) ) ;
INV     gate5921  (.A(g8040), .Z(g8514) ) ;
INV     gate5922  (.A(g7855), .Z(g8524) ) ;
INV     gate5923  (.A(g8094), .Z(g8541) ) ;
OR2     gate5924  (.A(g4783), .B(g7598), .Z(g7782) ) ;
INV     gate5925  (.A(g7782), .Z(II14657) ) ;
INV     gate5926  (.A(II14657), .Z(g8544) ) ;
INV     gate5927  (.A(g7905), .Z(g8545) ) ;
INV     gate5928  (.A(g8094), .Z(g8562) ) ;
OR2     gate5929  (.A(g4787), .B(g7600), .Z(g7783) ) ;
INV     gate5930  (.A(g7783), .Z(II14662) ) ;
INV     gate5931  (.A(II14662), .Z(g8563) ) ;
INV     gate5932  (.A(g7951), .Z(g8564) ) ;
INV     gate5933  (.A(g8094), .Z(g8581) ) ;
INV     gate5934  (.A(g8094), .Z(g8582) ) ;
OR2     gate5935  (.A(g4791), .B(g7602), .Z(g7787) ) ;
INV     gate5936  (.A(g7787), .Z(II14668) ) ;
INV     gate5937  (.A(II14668), .Z(g8583) ) ;
INV     gate5938  (.A(g7993), .Z(g8585) ) ;
INV     gate5939  (.A(g8094), .Z(g8602) ) ;
OR2     gate5940  (.A(g4794), .B(g7604), .Z(g7788) ) ;
INV     gate5941  (.A(g7788), .Z(II14674) ) ;
INV     gate5942  (.A(II14674), .Z(g8603) ) ;
OR2     gate5943  (.A(g4796), .B(g7606), .Z(g7791) ) ;
INV     gate5944  (.A(g7791), .Z(II14677) ) ;
INV     gate5945  (.A(II14677), .Z(g8604) ) ;
OR2     gate5946  (.A(g4799), .B(g7609), .Z(g7810) ) ;
INV     gate5947  (.A(g7810), .Z(II14680) ) ;
INV     gate5948  (.A(II14680), .Z(g8605) ) ;
OR2     gate5949  (.A(g4801), .B(g7615), .Z(g7825) ) ;
INV     gate5950  (.A(g7825), .Z(II14683) ) ;
INV     gate5951  (.A(II14683), .Z(g8606) ) ;
OR2     gate5952  (.A(g4804), .B(g7626), .Z(g7826) ) ;
INV     gate5953  (.A(g7826), .Z(II14687) ) ;
INV     gate5954  (.A(II14687), .Z(g8608) ) ;
INV     gate5955  (.A(g8016), .Z(II14695) ) ;
INV     gate5956  (.A(II14695), .Z(g8619) ) ;
INV     gate5957  (.A(g8198), .Z(II14709) ) ;
INV     gate5958  (.A(II14709), .Z(g8631) ) ;
AND2    gate5959  (.A(g7682), .B(g7032), .Z(g8059) ) ;
INV     gate5960  (.A(g8059), .Z(II14712) ) ;
INV     gate5961  (.A(II14712), .Z(g8632) ) ;
AND2    gate5962  (.A(g7687), .B(g5610), .Z(g8068) ) ;
INV     gate5963  (.A(g8068), .Z(II14718) ) ;
INV     gate5964  (.A(II14718), .Z(g8636) ) ;
AND2    gate5965  (.A(g7690), .B(g3521), .Z(g8076) ) ;
INV     gate5966  (.A(g8076), .Z(II14722) ) ;
INV     gate5967  (.A(II14722), .Z(g8638) ) ;
INV     gate5968  (.A(g8145), .Z(II14725) ) ;
INV     gate5969  (.A(II14725), .Z(g8639) ) ;
INV     gate5970  (.A(g8152), .Z(II14728) ) ;
INV     gate5971  (.A(II14728), .Z(g8640) ) ;
OR2     gate5972  (.A(g7632), .B(g3219), .Z(g8155) ) ;
INV     gate5973  (.A(g8155), .Z(II14732) ) ;
INV     gate5974  (.A(II14732), .Z(g8642) ) ;
INV     gate5975  (.A(g8173), .Z(II14739) ) ;
INV     gate5976  (.A(II14739), .Z(g8647) ) ;
INV     gate5977  (.A(g8174), .Z(II14743) ) ;
INV     gate5978  (.A(II14743), .Z(g8649) ) ;
INV     gate5979  (.A(g8175), .Z(II14747) ) ;
INV     gate5980  (.A(II14747), .Z(g8651) ) ;
OR2     gate5981  (.A(g7724), .B(g6762), .Z(g7834) ) ;
INV     gate5982  (.A(g7834), .Z(II14763) ) ;
INV     gate5983  (.A(II14763), .Z(g8657) ) ;
INV     gate5984  (.A(g8511), .Z(II14777) ) ;
INV     gate5985  (.A(g8284), .Z(II14780) ) ;
INV     gate5986  (.A(g8324), .Z(II14783) ) ;
INV     gate5987  (.A(g8606), .Z(II14786) ) ;
INV     gate5988  (.A(g8544), .Z(II14789) ) ;
INV     gate5989  (.A(g8583), .Z(II14792) ) ;
INV     gate5990  (.A(g8604), .Z(II14795) ) ;
INV     gate5991  (.A(g8605), .Z(II14798) ) ;
INV     gate5992  (.A(g8608), .Z(II14801) ) ;
INV     gate5993  (.A(g8563), .Z(II14804) ) ;
INV     gate5994  (.A(g8603), .Z(II14807) ) ;
INV     gate5995  (.A(g8481), .Z(II14810) ) ;
INV     gate5996  (.A(g8640), .Z(II14813) ) ;
INV     gate5997  (.A(g8642), .Z(II14816) ) ;
INV     gate5998  (.A(g8647), .Z(II14819) ) ;
INV     gate5999  (.A(g8649), .Z(II14822) ) ;
INV     gate6000  (.A(g8651), .Z(II14825) ) ;
INV     gate6001  (.A(g8639), .Z(II14828) ) ;
NOR4    gate6002  (.A(g6559), .B(g162), .C(g7784), .D(g3591), .Z(g8641) ) ;
INV     gate6003  (.A(g8641), .Z(II14844) ) ;
INV     gate6004  (.A(II14844), .Z(g8682) ) ;
INV     gate6005  (.A(g8235), .Z(g8683) ) ;
NOR4    gate6006  (.A(g1000), .B(g6573), .C(g1860), .D(g8009), .Z(g8625) ) ;
INV     gate6007  (.A(g8625), .Z(II14848) ) ;
INV     gate6008  (.A(II14848), .Z(g8684) ) ;
NOR4    gate6009  (.A(g6110), .B(g7784), .C(g3591), .D(g1864), .Z(g8630) ) ;
INV     gate6010  (.A(g8630), .Z(II14851) ) ;
INV     gate6011  (.A(II14851), .Z(g8685) ) ;
INV     gate6012  (.A(g8657), .Z(II14857) ) ;
INV     gate6013  (.A(II14857), .Z(g8689) ) ;
NOR2    gate6014  (.A(g6270), .B(g8009), .Z(g8629) ) ;
INV     gate6015  (.A(g8629), .Z(II14904) ) ;
INV     gate6016  (.A(II14904), .Z(g8734) ) ;
INV     gate6017  (.A(g8524), .Z(g8743) ) ;
INV     gate6018  (.A(g8524), .Z(g8746) ) ;
INV     gate6019  (.A(g8545), .Z(g8747) ) ;
INV     gate6020  (.A(g8524), .Z(g8750) ) ;
INV     gate6021  (.A(g8545), .Z(g8751) ) ;
INV     gate6022  (.A(g8564), .Z(g8752) ) ;
INV     gate6023  (.A(g8381), .Z(II14925) ) ;
INV     gate6024  (.A(II14925), .Z(g8753) ) ;
INV     gate6025  (.A(g8524), .Z(g8754) ) ;
INV     gate6026  (.A(g8545), .Z(g8755) ) ;
INV     gate6027  (.A(g8564), .Z(g8756) ) ;
INV     gate6028  (.A(g8585), .Z(g8757) ) ;
INV     gate6029  (.A(g8524), .Z(g8759) ) ;
INV     gate6030  (.A(g8545), .Z(g8760) ) ;
INV     gate6031  (.A(g8564), .Z(g8761) ) ;
INV     gate6032  (.A(g8585), .Z(g8762) ) ;
INV     gate6033  (.A(g8524), .Z(g8765) ) ;
INV     gate6034  (.A(g8545), .Z(g8766) ) ;
INV     gate6035  (.A(g8564), .Z(g8767) ) ;
INV     gate6036  (.A(g8585), .Z(g8768) ) ;
INV     gate6037  (.A(g8545), .Z(g8770) ) ;
INV     gate6038  (.A(g8564), .Z(g8771) ) ;
INV     gate6039  (.A(g8585), .Z(g8772) ) ;
INV     gate6040  (.A(g8406), .Z(II14964) ) ;
INV     gate6041  (.A(II14964), .Z(g8774) ) ;
INV     gate6042  (.A(g8564), .Z(g8775) ) ;
INV     gate6043  (.A(g8585), .Z(g8776) ) ;
INV     gate6044  (.A(g8442), .Z(II14974) ) ;
INV     gate6045  (.A(II14974), .Z(g8778) ) ;
INV     gate6046  (.A(g8524), .Z(g8780) ) ;
INV     gate6047  (.A(g8585), .Z(g8781) ) ;
INV     gate6048  (.A(g8524), .Z(g8783) ) ;
INV     gate6049  (.A(g8545), .Z(g8784) ) ;
INV     gate6050  (.A(g8545), .Z(g8786) ) ;
INV     gate6051  (.A(g8564), .Z(g8787) ) ;
INV     gate6052  (.A(g8564), .Z(g8789) ) ;
INV     gate6053  (.A(g8585), .Z(g8790) ) ;
INV     gate6054  (.A(g8585), .Z(g8791) ) ;
INV     gate6055  (.A(g8510), .Z(II14996) ) ;
INV     gate6056  (.A(II14996), .Z(g8792) ) ;
NAND2   gate6057  (.A(g8176), .B(g6232), .Z(g8633) ) ;
INV     gate6058  (.A(g8633), .Z(II15003) ) ;
INV     gate6059  (.A(II15003), .Z(g8797) ) ;
NAND2   gate6060  (.A(g6232), .B(g8091), .Z(g8627) ) ;
INV     gate6061  (.A(g8627), .Z(II15007) ) ;
INV     gate6062  (.A(II15007), .Z(g8799) ) ;
AND2    gate6063  (.A(g8146), .B(g7034), .Z(g8584) ) ;
INV     gate6064  (.A(g8584), .Z(II15010) ) ;
INV     gate6065  (.A(II15010), .Z(g8800) ) ;
AND2    gate6066  (.A(g8154), .B(g5616), .Z(g8607) ) ;
INV     gate6067  (.A(g8607), .Z(II15014) ) ;
INV     gate6068  (.A(II15014), .Z(g8802) ) ;
INV     gate6069  (.A(g8632), .Z(II15062) ) ;
INV     gate6070  (.A(II15062), .Z(g8808) ) ;
INV     gate6071  (.A(g8636), .Z(II15065) ) ;
INV     gate6072  (.A(II15065), .Z(g8809) ) ;
INV     gate6073  (.A(g8638), .Z(II15068) ) ;
INV     gate6074  (.A(II15068), .Z(g8810) ) ;
INV     gate6075  (.A(g8631), .Z(II15160) ) ;
INV     gate6076  (.A(II15160), .Z(g8856) ) ;
INV     gate6077  (.A(g8753), .Z(II15178) ) ;
INV     gate6078  (.A(g8734), .Z(II15181) ) ;
INV     gate6079  (.A(g8684), .Z(II15184) ) ;
INV     gate6080  (.A(g8682), .Z(II15187) ) ;
INV     gate6081  (.A(g8685), .Z(II15190) ) ;
INV     gate6082  (.A(g8774), .Z(II15193) ) ;
INV     gate6083  (.A(g8778), .Z(II15196) ) ;
INV     gate6084  (.A(g8792), .Z(II15199) ) ;
INV     gate6085  (.A(g8797), .Z(II15202) ) ;
INV     gate6086  (.A(g8809), .Z(II15205) ) ;
INV     gate6087  (.A(g8810), .Z(II15208) ) ;
INV     gate6088  (.A(g8808), .Z(II15211) ) ;
NOR2    gate6089  (.A(g8635), .B(g3790), .Z(g8801) ) ;
INV     gate6090  (.A(g8801), .Z(II15218) ) ;
INV     gate6091  (.A(II15218), .Z(g8880) ) ;
INV     gate6092  (.A(g8683), .Z(g8881) ) ;
OR2     gate6093  (.A(g7096), .B(g8229), .Z(g8834) ) ;
INV     gate6094  (.A(g8834), .Z(II15222) ) ;
INV     gate6095  (.A(II15222), .Z(g8882) ) ;
INV     gate6096  (.A(g8689), .Z(II15225) ) ;
INV     gate6097  (.A(II15225), .Z(g8883) ) ;
INV     gate6098  (.A(g8799), .Z(II15308) ) ;
INV     gate6099  (.A(II15308), .Z(g8898) ) ;
AND2    gate6100  (.A(g8619), .B(g3338), .Z(g8738) ) ;
INV     gate6101  (.A(g8738), .Z(II15315) ) ;
INV     gate6102  (.A(II15315), .Z(g8903) ) ;
AND2    gate6103  (.A(g8634), .B(g7037), .Z(g8779) ) ;
INV     gate6104  (.A(g8779), .Z(II15324) ) ;
INV     gate6105  (.A(II15324), .Z(g8910) ) ;
AND2    gate6106  (.A(g8637), .B(g5622), .Z(g8793) ) ;
INV     gate6107  (.A(g8793), .Z(II15329) ) ;
INV     gate6108  (.A(II15329), .Z(g8913) ) ;
INV     gate6109  (.A(g8800), .Z(II15334) ) ;
INV     gate6110  (.A(II15334), .Z(g8916) ) ;
INV     gate6111  (.A(g8802), .Z(II15337) ) ;
INV     gate6112  (.A(II15337), .Z(g8917) ) ;
INV     gate6113  (.A(g8856), .Z(II15340) ) ;
INV     gate6114  (.A(II15340), .Z(g8918) ) ;
INV     gate6115  (.A(g8882), .Z(II15379) ) ;
INV     gate6116  (.A(g8883), .Z(II15382) ) ;
INV     gate6117  (.A(g8880), .Z(II15385) ) ;
INV     gate6118  (.A(g8898), .Z(II15388) ) ;
INV     gate6119  (.A(g8917), .Z(II15391) ) ;
INV     gate6120  (.A(g8916), .Z(II15394) ) ;
OR2     gate6121  (.A(g8844), .B(g8654), .Z(g8902) ) ;
INV     gate6122  (.A(g8902), .Z(II15405) ) ;
INV     gate6123  (.A(II15405), .Z(g8967) ) ;
OR2     gate6124  (.A(g8828), .B(g8648), .Z(g8896) ) ;
INV     gate6125  (.A(g8896), .Z(II15408) ) ;
INV     gate6126  (.A(II15408), .Z(g8968) ) ;
OR2     gate6127  (.A(g8833), .B(g8650), .Z(g8897) ) ;
INV     gate6128  (.A(g8897), .Z(II15411) ) ;
INV     gate6129  (.A(II15411), .Z(g8969) ) ;
OR2     gate6130  (.A(g8840), .B(g8653), .Z(g8900) ) ;
INV     gate6131  (.A(g8900), .Z(II15414) ) ;
INV     gate6132  (.A(II15414), .Z(g8970) ) ;
OR2     gate6133  (.A(g8814), .B(g8643), .Z(g8893) ) ;
INV     gate6134  (.A(g8893), .Z(II15417) ) ;
INV     gate6135  (.A(II15417), .Z(g8971) ) ;
INV     gate6136  (.A(g8881), .Z(II15420) ) ;
INV     gate6137  (.A(II15420), .Z(g8972) ) ;
OR2     gate6138  (.A(g8817), .B(g8645), .Z(g8894) ) ;
INV     gate6139  (.A(g8894), .Z(II15423) ) ;
INV     gate6140  (.A(II15423), .Z(g8973) ) ;
OR2     gate6141  (.A(g8823), .B(g8646), .Z(g8895) ) ;
INV     gate6142  (.A(g8895), .Z(II15426) ) ;
INV     gate6143  (.A(II15426), .Z(g8974) ) ;
OR2     gate6144  (.A(g8839), .B(g8652), .Z(g8899) ) ;
INV     gate6145  (.A(g8899), .Z(II15429) ) ;
INV     gate6146  (.A(II15429), .Z(g8975) ) ;
AND2    gate6147  (.A(g8798), .B(g7688), .Z(g8911) ) ;
INV     gate6148  (.A(g8911), .Z(II15433) ) ;
INV     gate6149  (.A(II15433), .Z(g8977) ) ;
AND2    gate6150  (.A(g8804), .B(g5631), .Z(g8901) ) ;
INV     gate6151  (.A(g8901), .Z(II15475) ) ;
INV     gate6152  (.A(II15475), .Z(g9017) ) ;
INV     gate6153  (.A(g8910), .Z(II15478) ) ;
INV     gate6154  (.A(II15478), .Z(g9018) ) ;
INV     gate6155  (.A(g8913), .Z(II15481) ) ;
INV     gate6156  (.A(II15481), .Z(g9019) ) ;
INV     gate6157  (.A(g8918), .Z(II15484) ) ;
INV     gate6158  (.A(II15484), .Z(g9020) ) ;
INV     gate6159  (.A(g8971), .Z(II15492) ) ;
INV     gate6160  (.A(g8973), .Z(II15495) ) ;
INV     gate6161  (.A(g8974), .Z(II15498) ) ;
INV     gate6162  (.A(g8975), .Z(II15501) ) ;
INV     gate6163  (.A(g8967), .Z(II15504) ) ;
INV     gate6164  (.A(g8968), .Z(II15507) ) ;
INV     gate6165  (.A(g8969), .Z(II15510) ) ;
INV     gate6166  (.A(g8970), .Z(II15513) ) ;
INV     gate6167  (.A(g8977), .Z(II15516) ) ;
INV     gate6168  (.A(g9019), .Z(II15519) ) ;
INV     gate6169  (.A(g9018), .Z(II15522) ) ;
INV     gate6170  (.A(g9020), .Z(II15527) ) ;
INV     gate6171  (.A(II15527), .Z(g9039) ) ;
INV     gate6172  (.A(g8972), .Z(II15530) ) ;
INV     gate6173  (.A(II15530), .Z(g9042) ) ;
OR2     gate6174  (.A(g8942), .B(g8848), .Z(g9002) ) ;
INV     gate6175  (.A(g9002), .Z(II15533) ) ;
INV     gate6176  (.A(II15533), .Z(g9043) ) ;
OR2     gate6177  (.A(g8944), .B(g8851), .Z(g9004) ) ;
INV     gate6178  (.A(g9004), .Z(II15536) ) ;
INV     gate6179  (.A(II15536), .Z(g9044) ) ;
OR2     gate6180  (.A(g8945), .B(g8852), .Z(g9005) ) ;
INV     gate6181  (.A(g9005), .Z(II15539) ) ;
INV     gate6182  (.A(II15539), .Z(g9045) ) ;
OR2     gate6183  (.A(g8946), .B(g8853), .Z(g9006) ) ;
INV     gate6184  (.A(g9006), .Z(II15543) ) ;
INV     gate6185  (.A(II15543), .Z(g9047) ) ;
OR2     gate6186  (.A(g8947), .B(g8854), .Z(g9007) ) ;
INV     gate6187  (.A(g9007), .Z(II15546) ) ;
INV     gate6188  (.A(II15546), .Z(g9048) ) ;
OR2     gate6189  (.A(g8948), .B(g8857), .Z(g9008) ) ;
INV     gate6190  (.A(g9008), .Z(II15550) ) ;
INV     gate6191  (.A(II15550), .Z(g9050) ) ;
OR2     gate6192  (.A(g8949), .B(g8858), .Z(g9009) ) ;
INV     gate6193  (.A(g9009), .Z(II15553) ) ;
INV     gate6194  (.A(II15553), .Z(g9051) ) ;
OR2     gate6195  (.A(g8950), .B(g8860), .Z(g9010) ) ;
INV     gate6196  (.A(g9010), .Z(II15557) ) ;
INV     gate6197  (.A(II15557), .Z(g9053) ) ;
OR2     gate6198  (.A(g8919), .B(g8813), .Z(g8979) ) ;
INV     gate6199  (.A(g8979), .Z(II15562) ) ;
INV     gate6200  (.A(II15562), .Z(g9056) ) ;
OR2     gate6201  (.A(g8920), .B(g8815), .Z(g8980) ) ;
INV     gate6202  (.A(g8980), .Z(II15565) ) ;
INV     gate6203  (.A(II15565), .Z(g9057) ) ;
OR2     gate6204  (.A(g8921), .B(g8816), .Z(g8981) ) ;
INV     gate6205  (.A(g8981), .Z(II15568) ) ;
INV     gate6206  (.A(II15568), .Z(g9058) ) ;
OR2     gate6207  (.A(g8922), .B(g8820), .Z(g8982) ) ;
INV     gate6208  (.A(g8982), .Z(II15571) ) ;
INV     gate6209  (.A(II15571), .Z(g9059) ) ;
OR2     gate6210  (.A(g8923), .B(g8821), .Z(g8983) ) ;
INV     gate6211  (.A(g8983), .Z(II15574) ) ;
INV     gate6212  (.A(II15574), .Z(g9060) ) ;
OR2     gate6213  (.A(g8924), .B(g8822), .Z(g8984) ) ;
INV     gate6214  (.A(g8984), .Z(II15577) ) ;
INV     gate6215  (.A(II15577), .Z(g9061) ) ;
OR2     gate6216  (.A(g8925), .B(g8824), .Z(g8985) ) ;
INV     gate6217  (.A(g8985), .Z(II15580) ) ;
INV     gate6218  (.A(II15580), .Z(g9062) ) ;
OR2     gate6219  (.A(g8926), .B(g8825), .Z(g8986) ) ;
INV     gate6220  (.A(g8986), .Z(II15583) ) ;
INV     gate6221  (.A(II15583), .Z(g9063) ) ;
OR2     gate6222  (.A(g8927), .B(g8826), .Z(g8987) ) ;
INV     gate6223  (.A(g8987), .Z(II15586) ) ;
INV     gate6224  (.A(II15586), .Z(g9064) ) ;
OR2     gate6225  (.A(g8928), .B(g8827), .Z(g8988) ) ;
INV     gate6226  (.A(g8988), .Z(II15589) ) ;
INV     gate6227  (.A(II15589), .Z(g9065) ) ;
OR2     gate6228  (.A(g8929), .B(g8829), .Z(g8989) ) ;
INV     gate6229  (.A(g8989), .Z(II15592) ) ;
INV     gate6230  (.A(II15592), .Z(g9066) ) ;
OR2     gate6231  (.A(g8930), .B(g8830), .Z(g8990) ) ;
INV     gate6232  (.A(g8990), .Z(II15595) ) ;
INV     gate6233  (.A(II15595), .Z(g9067) ) ;
OR2     gate6234  (.A(g8931), .B(g8831), .Z(g8991) ) ;
INV     gate6235  (.A(g8991), .Z(II15598) ) ;
INV     gate6236  (.A(II15598), .Z(g9068) ) ;
OR2     gate6237  (.A(g8932), .B(g8832), .Z(g8992) ) ;
INV     gate6238  (.A(g8992), .Z(II15601) ) ;
INV     gate6239  (.A(II15601), .Z(g9069) ) ;
OR2     gate6240  (.A(g8933), .B(g8835), .Z(g8993) ) ;
INV     gate6241  (.A(g8993), .Z(II15604) ) ;
INV     gate6242  (.A(II15604), .Z(g9070) ) ;
OR2     gate6243  (.A(g8934), .B(g8836), .Z(g8994) ) ;
INV     gate6244  (.A(g8994), .Z(II15607) ) ;
INV     gate6245  (.A(II15607), .Z(g9071) ) ;
OR2     gate6246  (.A(g8935), .B(g8837), .Z(g8995) ) ;
INV     gate6247  (.A(g8995), .Z(II15610) ) ;
INV     gate6248  (.A(II15610), .Z(g9072) ) ;
OR2     gate6249  (.A(g8936), .B(g8838), .Z(g8996) ) ;
INV     gate6250  (.A(g8996), .Z(II15613) ) ;
INV     gate6251  (.A(II15613), .Z(g9073) ) ;
OR2     gate6252  (.A(g8937), .B(g8841), .Z(g8997) ) ;
INV     gate6253  (.A(g8997), .Z(II15616) ) ;
INV     gate6254  (.A(II15616), .Z(g9074) ) ;
OR2     gate6255  (.A(g8938), .B(g8842), .Z(g8998) ) ;
INV     gate6256  (.A(g8998), .Z(II15619) ) ;
INV     gate6257  (.A(II15619), .Z(g9075) ) ;
OR2     gate6258  (.A(g8939), .B(g8843), .Z(g8999) ) ;
INV     gate6259  (.A(g8999), .Z(II15622) ) ;
INV     gate6260  (.A(II15622), .Z(g9076) ) ;
OR2     gate6261  (.A(g8940), .B(g8845), .Z(g9000) ) ;
INV     gate6262  (.A(g9000), .Z(II15625) ) ;
INV     gate6263  (.A(II15625), .Z(g9077) ) ;
OR2     gate6264  (.A(g8941), .B(g8846), .Z(g9001) ) ;
INV     gate6265  (.A(g9001), .Z(II15628) ) ;
INV     gate6266  (.A(II15628), .Z(g9078) ) ;
OR2     gate6267  (.A(g8943), .B(g8849), .Z(g9003) ) ;
INV     gate6268  (.A(g9003), .Z(II15631) ) ;
INV     gate6269  (.A(II15631), .Z(g9079) ) ;
AND2    gate6270  (.A(g8903), .B(g6588), .Z(g8976) ) ;
INV     gate6271  (.A(g8976), .Z(II15635) ) ;
INV     gate6272  (.A(II15635), .Z(g9081) ) ;
AND2    gate6273  (.A(g8909), .B(g5587), .Z(g8978) ) ;
INV     gate6274  (.A(g8978), .Z(II15638) ) ;
INV     gate6275  (.A(II15638), .Z(g9082) ) ;
INV     gate6276  (.A(g9017), .Z(II15641) ) ;
INV     gate6277  (.A(II15641), .Z(g9083) ) ;
INV     gate6278  (.A(g9043), .Z(II15645) ) ;
INV     gate6279  (.A(g9044), .Z(II15648) ) ;
INV     gate6280  (.A(g9056), .Z(II15651) ) ;
INV     gate6281  (.A(g9057), .Z(II15654) ) ;
INV     gate6282  (.A(g9059), .Z(II15657) ) ;
INV     gate6283  (.A(g9062), .Z(II15660) ) ;
INV     gate6284  (.A(g9066), .Z(II15663) ) ;
INV     gate6285  (.A(g9070), .Z(II15666) ) ;
INV     gate6286  (.A(g9045), .Z(II15669) ) ;
INV     gate6287  (.A(g9047), .Z(II15672) ) ;
INV     gate6288  (.A(g9058), .Z(II15675) ) ;
INV     gate6289  (.A(g9060), .Z(II15678) ) ;
INV     gate6290  (.A(g9063), .Z(II15681) ) ;
INV     gate6291  (.A(g9067), .Z(II15684) ) ;
INV     gate6292  (.A(g9071), .Z(II15687) ) ;
INV     gate6293  (.A(g9074), .Z(II15690) ) ;
INV     gate6294  (.A(g9048), .Z(II15693) ) ;
INV     gate6295  (.A(g9050), .Z(II15696) ) ;
INV     gate6296  (.A(g9061), .Z(II15699) ) ;
INV     gate6297  (.A(g9064), .Z(II15702) ) ;
INV     gate6298  (.A(g9068), .Z(II15705) ) ;
INV     gate6299  (.A(g9072), .Z(II15708) ) ;
INV     gate6300  (.A(g9075), .Z(II15711) ) ;
INV     gate6301  (.A(g9077), .Z(II15714) ) ;
INV     gate6302  (.A(g9051), .Z(II15717) ) ;
INV     gate6303  (.A(g9053), .Z(II15720) ) ;
INV     gate6304  (.A(g9065), .Z(II15723) ) ;
INV     gate6305  (.A(g9069), .Z(II15726) ) ;
INV     gate6306  (.A(g9073), .Z(II15729) ) ;
INV     gate6307  (.A(g9076), .Z(II15732) ) ;
INV     gate6308  (.A(g9078), .Z(II15735) ) ;
INV     gate6309  (.A(g9079), .Z(II15738) ) ;
INV     gate6310  (.A(g9083), .Z(II15741) ) ;
INV     gate6311  (.A(g9042), .Z(II15747) ) ;
INV     gate6312  (.A(II15747), .Z(g9121) ) ;
AND2    gate6313  (.A(g9011), .B(g5598), .Z(g9080) ) ;
INV     gate6314  (.A(g9080), .Z(II15753) ) ;
INV     gate6315  (.A(II15753), .Z(g9125) ) ;
INV     gate6316  (.A(g9081), .Z(II15756) ) ;
INV     gate6317  (.A(II15756), .Z(g9126) ) ;
INV     gate6318  (.A(g9082), .Z(II15759) ) ;
INV     gate6319  (.A(II15759), .Z(g9127) ) ;
INV     gate6320  (.A(g9039), .Z(II15762) ) ;
INV     gate6321  (.A(g9039), .Z(II15765) ) ;
INV     gate6322  (.A(II15765), .Z(g9129) ) ;
INV     gate6323  (.A(g9121), .Z(II15770) ) ;
INV     gate6324  (.A(g9126), .Z(II15773) ) ;
INV     gate6325  (.A(g9127), .Z(II15776) ) ;
INV     gate6326  (.A(g9125), .Z(II15784) ) ;
INV     gate6327  (.A(II15784), .Z(g9140) ) ;
INV     gate6328  (.A(g9129), .Z(g9141) ) ;
INV     gate6329  (.A(g9140), .Z(II15791) ) ;
INV     gate6330  (.A(g9141), .Z(g9157) ) ;
OR2     gate6331  (.A(g9143), .B(g9024), .Z(g9148) ) ;
INV     gate6332  (.A(g9148), .Z(II15803) ) ;
INV     gate6333  (.A(II15803), .Z(g9161) ) ;
OR2     gate6334  (.A(g9144), .B(g8961), .Z(g9151) ) ;
INV     gate6335  (.A(g9151), .Z(II15811) ) ;
INV     gate6336  (.A(II15811), .Z(g9177) ) ;
OR2     gate6337  (.A(g9142), .B(g9021), .Z(g9154) ) ;
INV     gate6338  (.A(g9154), .Z(II15814) ) ;
INV     gate6339  (.A(II15814), .Z(g9178) ) ;
INV     gate6340  (.A(g9157), .Z(II15824) ) ;
INV     gate6341  (.A(II15824), .Z(g9180) ) ;
INV     gate6342  (.A(g9177), .Z(g9181) ) ;
INV     gate6343  (.A(g9178), .Z(g9182) ) ;
INV     gate6344  (.A(g9161), .Z(g9183) ) ;
INV     gate6345  (.A(g9180), .Z(II15830) ) ;
INV     gate6346  (.A(II15830), .Z(g9184) ) ;
OR2     gate6347  (.A(g9158), .B(g9022), .Z(g9162) ) ;
INV     gate6348  (.A(g9162), .Z(II15833) ) ;
INV     gate6349  (.A(II15833), .Z(g9185) ) ;
OR2     gate6350  (.A(g9159), .B(g9023), .Z(g9165) ) ;
INV     gate6351  (.A(g9165), .Z(II15836) ) ;
INV     gate6352  (.A(II15836), .Z(g9186) ) ;
OR2     gate6353  (.A(g9160), .B(g9025), .Z(g9168) ) ;
INV     gate6354  (.A(g9168), .Z(II15839) ) ;
INV     gate6355  (.A(II15839), .Z(g9187) ) ;
OR2     gate6356  (.A(g9146), .B(g8962), .Z(g9171) ) ;
INV     gate6357  (.A(g9171), .Z(II15842) ) ;
INV     gate6358  (.A(II15842), .Z(g9188) ) ;
OR2     gate6359  (.A(g9147), .B(g8963), .Z(g9174) ) ;
INV     gate6360  (.A(g9174), .Z(II15845) ) ;
INV     gate6361  (.A(II15845), .Z(g9189) ) ;
INV     gate6362  (.A(g9181), .Z(g9193) ) ;
INV     gate6363  (.A(g9182), .Z(g9194) ) ;
INV     gate6364  (.A(g9184), .Z(II15871) ) ;
INV     gate6365  (.A(II15871), .Z(g9195) ) ;
INV     gate6366  (.A(g9185), .Z(g9196) ) ;
INV     gate6367  (.A(g9186), .Z(g9197) ) ;
INV     gate6368  (.A(g9187), .Z(g9198) ) ;
INV     gate6369  (.A(g9188), .Z(g9199) ) ;
INV     gate6370  (.A(g9189), .Z(g9200) ) ;
INV     gate6371  (.A(g9183), .Z(g9201) ) ;
INV     gate6372  (.A(g9195), .Z(II15894) ) ;
INV     gate6373  (.A(g9196), .Z(g9206) ) ;
INV     gate6374  (.A(g9197), .Z(g9207) ) ;
INV     gate6375  (.A(g9198), .Z(g9208) ) ;
INV     gate6376  (.A(g9199), .Z(g9209) ) ;
INV     gate6377  (.A(g9200), .Z(g9210) ) ;
INV     gate6378  (.A(g9201), .Z(II15909) ) ;
INV     gate6379  (.A(II15909), .Z(g9211) ) ;
INV     gate6380  (.A(g9193), .Z(II15912) ) ;
INV     gate6381  (.A(II15912), .Z(g9212) ) ;
INV     gate6382  (.A(g9194), .Z(II15915) ) ;
INV     gate6383  (.A(II15915), .Z(g9213) ) ;
INV     gate6384  (.A(g9211), .Z(II15918) ) ;
INV     gate6385  (.A(II15918), .Z(g9214) ) ;
INV     gate6386  (.A(g9206), .Z(II15921) ) ;
INV     gate6387  (.A(II15921), .Z(g9215) ) ;
INV     gate6388  (.A(g9207), .Z(II15924) ) ;
INV     gate6389  (.A(II15924), .Z(g9216) ) ;
INV     gate6390  (.A(g9208), .Z(II15927) ) ;
INV     gate6391  (.A(II15927), .Z(g9217) ) ;
INV     gate6392  (.A(g9209), .Z(II15930) ) ;
INV     gate6393  (.A(II15930), .Z(g9218) ) ;
INV     gate6394  (.A(g9210), .Z(II15933) ) ;
INV     gate6395  (.A(II15933), .Z(g9219) ) ;
NAND2   gate6396  (.A(II15898), .B(II15899), .Z(g9205) ) ;
INV     gate6397  (.A(g9205), .Z(g9220) ) ;
INV     gate6398  (.A(g9212), .Z(II15937) ) ;
INV     gate6399  (.A(II15937), .Z(g9221) ) ;
INV     gate6400  (.A(g9213), .Z(II15940) ) ;
INV     gate6401  (.A(II15940), .Z(g9222) ) ;
INV     gate6402  (.A(g9214), .Z(II15943) ) ;
INV     gate6403  (.A(II15943), .Z(g9223) ) ;
INV     gate6404  (.A(g9221), .Z(II15947) ) ;
INV     gate6405  (.A(II15947), .Z(g9227) ) ;
INV     gate6406  (.A(g9222), .Z(II15950) ) ;
INV     gate6407  (.A(II15950), .Z(g9230) ) ;
INV     gate6408  (.A(g9215), .Z(II15953) ) ;
INV     gate6409  (.A(II15953), .Z(g9233) ) ;
INV     gate6410  (.A(g9216), .Z(II15956) ) ;
INV     gate6411  (.A(II15956), .Z(g9234) ) ;
INV     gate6412  (.A(g9217), .Z(II15959) ) ;
INV     gate6413  (.A(II15959), .Z(g9235) ) ;
INV     gate6414  (.A(g9218), .Z(II15962) ) ;
INV     gate6415  (.A(II15962), .Z(g9236) ) ;
INV     gate6416  (.A(g9219), .Z(II15965) ) ;
INV     gate6417  (.A(II15965), .Z(g9237) ) ;
INV     gate6418  (.A(g9233), .Z(II15971) ) ;
INV     gate6419  (.A(II15971), .Z(g9241) ) ;
INV     gate6420  (.A(g9234), .Z(II15974) ) ;
INV     gate6421  (.A(II15974), .Z(g9244) ) ;
INV     gate6422  (.A(g9235), .Z(II15978) ) ;
INV     gate6423  (.A(II15978), .Z(g9248) ) ;
INV     gate6424  (.A(g9236), .Z(II15982) ) ;
INV     gate6425  (.A(II15982), .Z(g9252) ) ;
INV     gate6426  (.A(g9237), .Z(II15985) ) ;
INV     gate6427  (.A(II15985), .Z(g9255) ) ;
OR2     gate6428  (.A(g7653), .B(g9226), .Z(g9239) ) ;
INV     gate6429  (.A(g9239), .Z(II15990) ) ;
INV     gate6430  (.A(II15990), .Z(g9260) ) ;
OR2     gate6431  (.A(g9238), .B(g6227), .Z(g9261) ) ;
INV     gate6432  (.A(g9261), .Z(II16006) ) ;
INV     gate6433  (.A(g9261), .Z(II16009) ) ;
INV     gate6434  (.A(II16009), .Z(g9281) ) ;
OR2     gate6435  (.A(g9247), .B(g6242), .Z(g9264) ) ;
INV     gate6436  (.A(g9264), .Z(II16017) ) ;
INV     gate6437  (.A(g9264), .Z(II16020) ) ;
INV     gate6438  (.A(II16020), .Z(g9298) ) ;
OR2     gate6439  (.A(g9251), .B(g6225), .Z(g9267) ) ;
INV     gate6440  (.A(g9267), .Z(II16023) ) ;
INV     gate6441  (.A(g9267), .Z(II16026) ) ;
INV     gate6442  (.A(II16026), .Z(g9300) ) ;
INV     gate6443  (.A(g9260), .Z(g9301) ) ;
INV     gate6444  (.A(g9281), .Z(g9302) ) ;
INV     gate6445  (.A(g9301), .Z(g9303) ) ;
INV     gate6446  (.A(g9298), .Z(g9304) ) ;
OR2     gate6447  (.A(g9270), .B(g6238), .Z(g9282) ) ;
INV     gate6448  (.A(g9282), .Z(II16033) ) ;
INV     gate6449  (.A(g9282), .Z(II16036) ) ;
INV     gate6450  (.A(II16036), .Z(g9306) ) ;
INV     gate6451  (.A(g9300), .Z(g9307) ) ;
OR2     gate6452  (.A(g9271), .B(g6221), .Z(g9285) ) ;
INV     gate6453  (.A(g9285), .Z(II16040) ) ;
INV     gate6454  (.A(g9285), .Z(II16043) ) ;
INV     gate6455  (.A(II16043), .Z(g9309) ) ;
OR2     gate6456  (.A(g9272), .B(g6235), .Z(g9288) ) ;
INV     gate6457  (.A(g9288), .Z(II16046) ) ;
INV     gate6458  (.A(g9288), .Z(II16049) ) ;
INV     gate6459  (.A(II16049), .Z(g9311) ) ;
OR2     gate6460  (.A(g9273), .B(g6216), .Z(g9291) ) ;
INV     gate6461  (.A(g9291), .Z(II16052) ) ;
INV     gate6462  (.A(g9291), .Z(II16055) ) ;
INV     gate6463  (.A(II16055), .Z(g9313) ) ;
OR2     gate6464  (.A(g9274), .B(g6230), .Z(g9294) ) ;
INV     gate6465  (.A(g9294), .Z(II16058) ) ;
INV     gate6466  (.A(g9294), .Z(II16061) ) ;
INV     gate6467  (.A(II16061), .Z(g9315) ) ;
INV     gate6468  (.A(g9302), .Z(g9316) ) ;
INV     gate6469  (.A(g9306), .Z(g9317) ) ;
INV     gate6470  (.A(g9304), .Z(g9318) ) ;
INV     gate6471  (.A(g9309), .Z(g9319) ) ;
INV     gate6472  (.A(g9307), .Z(g9320) ) ;
INV     gate6473  (.A(g9311), .Z(g9321) ) ;
INV     gate6474  (.A(g9313), .Z(g9322) ) ;
INV     gate6475  (.A(g9315), .Z(g9323) ) ;
INV     gate6476  (.A(g9303), .Z(II16072) ) ;
INV     gate6477  (.A(II16072), .Z(g9324) ) ;
INV     gate6478  (.A(g9317), .Z(g9329) ) ;
INV     gate6479  (.A(g9319), .Z(g9330) ) ;
INV     gate6480  (.A(g9321), .Z(g9331) ) ;
INV     gate6481  (.A(g9322), .Z(g9332) ) ;
INV     gate6482  (.A(g9323), .Z(g9333) ) ;
INV     gate6483  (.A(g9324), .Z(II16084) ) ;
INV     gate6484  (.A(II16084), .Z(g9336) ) ;
INV     gate6485  (.A(g9336), .Z(II16090) ) ;
INV     gate6486  (.A(II16090), .Z(g9340) ) ;
OR2     gate6487  (.A(g9258), .B(g9334), .Z(g9338) ) ;
INV     gate6488  (.A(g9338), .Z(II16100) ) ;
INV     gate6489  (.A(II16100), .Z(g9350) ) ;
OR2     gate6490  (.A(g9259), .B(g9335), .Z(g9339) ) ;
INV     gate6491  (.A(g9339), .Z(II16103) ) ;
INV     gate6492  (.A(II16103), .Z(g9351) ) ;
OR2     gate6493  (.A(g9240), .B(g9327), .Z(g9337) ) ;
INV     gate6494  (.A(g9337), .Z(II16107) ) ;
INV     gate6495  (.A(II16107), .Z(g9353) ) ;
INV     gate6496  (.A(g9350), .Z(II16116) ) ;
INV     gate6497  (.A(g9351), .Z(II16119) ) ;
INV     gate6498  (.A(g9353), .Z(II16122) ) ;
OR2     gate6499  (.A(g9275), .B(g9344), .Z(g9354) ) ;
INV     gate6500  (.A(g9354), .Z(II16126) ) ;
INV     gate6501  (.A(II16126), .Z(g9366) ) ;
OR2     gate6502  (.A(g9276), .B(g9345), .Z(g9355) ) ;
INV     gate6503  (.A(g9355), .Z(II16129) ) ;
INV     gate6504  (.A(II16129), .Z(g9367) ) ;
OR2     gate6505  (.A(g9277), .B(g9346), .Z(g9356) ) ;
INV     gate6506  (.A(g9356), .Z(II16132) ) ;
INV     gate6507  (.A(II16132), .Z(g9368) ) ;
OR2     gate6508  (.A(g9278), .B(g9347), .Z(g9357) ) ;
INV     gate6509  (.A(g9357), .Z(II16135) ) ;
INV     gate6510  (.A(II16135), .Z(g9369) ) ;
OR2     gate6511  (.A(g9279), .B(g9348), .Z(g9358) ) ;
INV     gate6512  (.A(g9358), .Z(II16138) ) ;
INV     gate6513  (.A(II16138), .Z(g9370) ) ;
INV     gate6514  (.A(g9366), .Z(II16142) ) ;
INV     gate6515  (.A(g9367), .Z(II16145) ) ;
INV     gate6516  (.A(g9368), .Z(II16148) ) ;
INV     gate6517  (.A(g9369), .Z(II16151) ) ;
INV     gate6518  (.A(g9370), .Z(II16154) ) ;
OR2     gate6519  (.A(g9359), .B(g6210), .Z(g9363) ) ;
INV     gate6520  (.A(g9363), .Z(II16158) ) ;
INV     gate6521  (.A(g9363), .Z(II16161) ) ;
INV     gate6522  (.A(II16161), .Z(g9379) ) ;
INV     gate6523  (.A(g9379), .Z(g9380) ) ;
OR2     gate6524  (.A(g9371), .B(g6757), .Z(g9377) ) ;
INV     gate6525  (.A(g9377), .Z(II16165) ) ;
INV     gate6526  (.A(II16165), .Z(g9381) ) ;
INV     gate6527  (.A(g9381), .Z(II16168) ) ;
INV     gate6528  (.A(II16168), .Z(g9382) ) ;
INV     gate6529  (.A(g9380), .Z(g9383) ) ;
INV     gate6530  (.A(g9382), .Z(II16173) ) ;
INV     gate6531  (.A(II16173), .Z(g9385) ) ;
INV     gate6532  (.A(g9385), .Z(II16176) ) ;
OR2     gate6533  (.A(g9349), .B(g9384), .Z(g9387) ) ;
INV     gate6534  (.A(g9387), .Z(II16180) ) ;
INV     gate6535  (.A(II16180), .Z(g9388) ) ;
INV     gate6536  (.A(g9388), .Z(II16183) ) ;
AND2    gate6537  (.A(g1454), .B(g1450), .Z(g1714) ) ;
AND2    gate6538  (.A(g1409), .B(g1416), .Z(g1725) ) ;
AND2    gate6539  (.A(g1432), .B(g1439), .Z(g1728) ) ;
AND2    gate6540  (.A(g1489), .B(g1481), .Z(g1733) ) ;
AND2    gate6541  (.A(g803), .B(g799), .Z(g1739) ) ;
AND2    gate6542  (.A(g819), .B(g815), .Z(g1753) ) ;
AND2    gate6543  (.A(g933), .B(g929), .Z(g1834) ) ;
AND2    gate6544  (.A(g959), .B(g955), .Z(g1898) ) ;
AND2    gate6545  (.A(g1528), .B(g1532), .Z(g1913) ) ;
AND2    gate6546  (.A(g1098), .B(g1087), .Z(g1919) ) ;
AND2    gate6547  (.A(g1130), .B(g1092), .Z(g2386) ) ;
OR3     gate6548  (.A(g1021), .B(g1025), .C(g1018), .Z(g1690) ) ;
AND2    gate6549  (.A(g1612), .B(g1077), .Z(g2889) ) ;
AND2    gate6550  (.A(g1080), .B(g1945), .Z(g2912) ) ;
AND2    gate6551  (.A(g1612), .B(g1077), .Z(g2935) ) ;
AND2    gate6552  (.A(g822), .B(g1753), .Z(g2949) ) ;
AND2    gate6553  (.A(g2474), .B(g2215), .Z(g2952) ) ;
AND2    gate6554  (.A(g2397), .B(g2407), .Z(g2972) ) ;
AND2    gate6555  (.A(g1494), .B(g1733), .Z(g2979) ) ;
AND2    gate6556  (.A(g806), .B(g1739), .Z(g2986) ) ;
AND2    gate6557  (.A(g2274), .B(g1844), .Z(g3049) ) ;
NAND2   gate6558  (.A(II5520), .B(II5521), .Z(g1682) ) ;
AND2    gate6559  (.A(g1682), .B(g1616), .Z(g3081) ) ;
AND2    gate6560  (.A(g945), .B(g1898), .Z(g3094) ) ;
AND2    gate6561  (.A(g2298), .B(g2316), .Z(g3188) ) ;
AND2    gate6562  (.A(g1658), .B(g2424), .Z(g3190) ) ;
AND2    gate6563  (.A(g1537), .B(g1913), .Z(g3222) ) ;
AND2    gate6564  (.A(g1102), .B(g1919), .Z(g3226) ) ;
AND2    gate6565  (.A(g1728), .B(g2015), .Z(g3229) ) ;
AND4    gate6566  (.A(g2298), .B(g2316), .C(g2334), .D(g2354), .Z(g3258) ) ;
AND3    gate6567  (.A(g2334), .B(g2316), .C(g2298), .Z(g3313) ) ;
AND2    gate6568  (.A(g1637), .B(g1616), .Z(g3509) ) ;
AND2    gate6569  (.A(g1134), .B(g2386), .Z(g3614) ) ;
AND2    gate6570  (.A(g2403), .B(g3085), .Z(g3984) ) ;
AND2    gate6571  (.A(g825), .B(g2949), .Z(g4038) ) ;
AND2    gate6572  (.A(g1272), .B(g3503), .Z(g4047) ) ;
AND2    gate6573  (.A(g1288), .B(g3513), .Z(g4048) ) ;
AND2    gate6574  (.A(g141), .B(g3514), .Z(g4049) ) ;
AND2    gate6575  (.A(g1276), .B(g3522), .Z(g4052) ) ;
AND2    gate6576  (.A(g1292), .B(g3523), .Z(g4053) ) ;
NAND2   gate6577  (.A(II7240), .B(II7241), .Z(g3767) ) ;
AND2    gate6578  (.A(g3767), .B(g2424), .Z(g4054) ) ;
NAND2   gate6579  (.A(II7139), .B(II7140), .Z(g3656) ) ;
AND2    gate6580  (.A(g3656), .B(g2407), .Z(g4058) ) ;
AND2    gate6581  (.A(g1499), .B(g2979), .Z(g4059) ) ;
AND2    gate6582  (.A(g809), .B(g2986), .Z(g4062) ) ;
AND2    gate6583  (.A(g1280), .B(g3532), .Z(g4066) ) ;
AND2    gate6584  (.A(g133), .B(g3539), .Z(g4067) ) ;
AND2    gate6585  (.A(g121), .B(g3540), .Z(g4068) ) ;
AND2    gate6586  (.A(g1300), .B(g3567), .Z(g4073) ) ;
AND2    gate6587  (.A(g137), .B(g3573), .Z(g4074) ) ;
AND2    gate6588  (.A(g1284), .B(g3582), .Z(g4077) ) ;
AND2    gate6589  (.A(g1296), .B(g3604), .Z(g4082) ) ;
AND2    gate6590  (.A(g125), .B(g3610), .Z(g4083) ) ;
AND2    gate6591  (.A(g103), .B(g3629), .Z(g4086) ) ;
AND2    gate6592  (.A(g129), .B(g3639), .Z(g4091) ) ;
AND2    gate6593  (.A(g2624), .B(g2614), .Z(g4097) ) ;
AND2    gate6594  (.A(g985), .B(g3790), .Z(g4098) ) ;
AND2    gate6595  (.A(g117), .B(g3647), .Z(g4099) ) ;
AND2    gate6596  (.A(g113), .B(g3648), .Z(g4100) ) ;
AND2    gate6597  (.A(g108), .B(g3649), .Z(g4101) ) ;
AND2    gate6598  (.A(g2625), .B(g2615), .Z(g4107) ) ;
AND2    gate6599  (.A(g782), .B(g3655), .Z(g4108) ) ;
AND2    gate6600  (.A(g990), .B(g3790), .Z(g4109) ) ;
AND2    gate6601  (.A(g2626), .B(g2616), .Z(g4117) ) ;
AND2    gate6602  (.A(g995), .B(g3790), .Z(g4118) ) ;
AND2    gate6603  (.A(g2627), .B(g2617), .Z(g4123) ) ;
AND2    gate6604  (.A(g2641), .B(g2640), .Z(g4124) ) ;
AND2    gate6605  (.A(g2628), .B(g2618), .Z(g4127) ) ;
AND2    gate6606  (.A(g98), .B(g3693), .Z(g4128) ) ;
AND2    gate6607  (.A(g2629), .B(g2621), .Z(g4129) ) ;
AND2    gate6608  (.A(g2630), .B(g2622), .Z(g4131) ) ;
AND2    gate6609  (.A(g2637), .B(g2633), .Z(g4132) ) ;
AND2    gate6610  (.A(g2631), .B(g2623), .Z(g4133) ) ;
AND4    gate6611  (.A(g3430), .B(g3398), .C(g3359), .D(g3341), .Z(II7994) ) ;
AND4    gate6612  (.A(g2074), .B(g3287), .C(g2020), .D(g3238), .Z(II7995) ) ;
AND2    gate6613  (.A(II7994), .B(II7995), .Z(g4135) ) ;
AND2    gate6614  (.A(g2638), .B(g2634), .Z(g4138) ) ;
AND4    gate6615  (.A(g3430), .B(g3398), .C(g3359), .D(g3341), .Z(II8000) ) ;
AND4    gate6616  (.A(g2074), .B(g3287), .C(g2020), .D(g1987), .Z(II8001) ) ;
AND2    gate6617  (.A(II8000), .B(II8001), .Z(g4139) ) ;
AND4    gate6618  (.A(g3430), .B(g3398), .C(g3359), .D(g2106), .Z(II8005) ) ;
AND4    gate6619  (.A(g2074), .B(g3287), .C(g2020), .D(g3238), .Z(II8006) ) ;
AND2    gate6620  (.A(II8005), .B(II8006), .Z(g4142) ) ;
AND2    gate6621  (.A(g2639), .B(g2635), .Z(g4145) ) ;
AND4    gate6622  (.A(g3430), .B(g3398), .C(g3359), .D(g3341), .Z(II8014) ) ;
AND4    gate6623  (.A(g2074), .B(g2057), .C(g3264), .D(g3238), .Z(II8015) ) ;
AND2    gate6624  (.A(II8014), .B(II8015), .Z(g4147) ) ;
AND4    gate6625  (.A(g3430), .B(g3398), .C(g3359), .D(g2106), .Z(II8019) ) ;
AND4    gate6626  (.A(g2074), .B(g3287), .C(g2020), .D(g1987), .Z(II8020) ) ;
AND2    gate6627  (.A(II8019), .B(II8020), .Z(g4150) ) ;
AND2    gate6628  (.A(g1098), .B(g3495), .Z(g4154) ) ;
AND4    gate6629  (.A(g3430), .B(g3398), .C(g3359), .D(g3341), .Z(II8028) ) ;
AND4    gate6630  (.A(g2074), .B(g2057), .C(g3264), .D(g1987), .Z(II8029) ) ;
AND2    gate6631  (.A(II8028), .B(II8029), .Z(g4155) ) ;
AND4    gate6632  (.A(g3430), .B(g3398), .C(g3359), .D(g2106), .Z(II8033) ) ;
AND4    gate6633  (.A(g2074), .B(g2057), .C(g3264), .D(g3238), .Z(II8034) ) ;
AND2    gate6634  (.A(II8033), .B(II8034), .Z(g4158) ) ;
AND2    gate6635  (.A(g1102), .B(g3498), .Z(g4159) ) ;
AND4    gate6636  (.A(g3430), .B(g3398), .C(g3359), .D(g3341), .Z(II8040) ) ;
AND4    gate6637  (.A(g2074), .B(g2057), .C(g2020), .D(g3238), .Z(II8041) ) ;
AND2    gate6638  (.A(II8040), .B(II8041), .Z(g4163) ) ;
AND4    gate6639  (.A(g3430), .B(g3398), .C(g3359), .D(g2106), .Z(II8045) ) ;
AND4    gate6640  (.A(g2074), .B(g2057), .C(g3264), .D(g1987), .Z(II8046) ) ;
AND2    gate6641  (.A(II8045), .B(II8046), .Z(g4166) ) ;
NAND2   gate6642  (.A(II6523), .B(II6524), .Z(g2783) ) ;
AND2    gate6643  (.A(g2783), .B(g1616), .Z(g4167) ) ;
AND2    gate6644  (.A(g1106), .B(g3500), .Z(g4168) ) ;
AND4    gate6645  (.A(g2162), .B(g2149), .C(g2137), .D(g2106), .Z(II8052) ) ;
AND4    gate6646  (.A(g3316), .B(g3287), .C(g3264), .D(g3238), .Z(II8053) ) ;
AND2    gate6647  (.A(II8052), .B(II8053), .Z(g4169) ) ;
AND4    gate6648  (.A(g3430), .B(g3398), .C(g3359), .D(g3341), .Z(II8057) ) ;
AND4    gate6649  (.A(g2074), .B(g2057), .C(g2020), .D(g1987), .Z(II8058) ) ;
AND2    gate6650  (.A(II8057), .B(II8058), .Z(g4172) ) ;
AND2    gate6651  (.A(g1110), .B(g3502), .Z(g4175) ) ;
AND4    gate6652  (.A(g2162), .B(g2149), .C(g2137), .D(g2106), .Z(II8063) ) ;
AND4    gate6653  (.A(g3316), .B(g3287), .C(g3264), .D(g1987), .Z(II8064) ) ;
AND2    gate6654  (.A(II8063), .B(II8064), .Z(g4176) ) ;
AND2    gate6655  (.A(g1114), .B(g3511), .Z(g4180) ) ;
AND2    gate6656  (.A(g1142), .B(g3512), .Z(g4181) ) ;
AND4    gate6657  (.A(g2162), .B(g2149), .C(g2137), .D(g2106), .Z(II8071) ) ;
AND4    gate6658  (.A(g3316), .B(g3287), .C(g2020), .D(g3238), .Z(II8072) ) ;
AND2    gate6659  (.A(II8071), .B(II8072), .Z(g4182) ) ;
AND2    gate6660  (.A(g2636), .B(g2632), .Z(g4185) ) ;
AND2    gate6661  (.A(g1118), .B(g3520), .Z(g4186) ) ;
AND4    gate6662  (.A(g2162), .B(g2149), .C(g2137), .D(g2106), .Z(II8078) ) ;
AND4    gate6663  (.A(g3316), .B(g3287), .C(g2020), .D(g1987), .Z(II8079) ) ;
AND2    gate6664  (.A(II8078), .B(II8079), .Z(g4187) ) ;
AND2    gate6665  (.A(g1122), .B(g3527), .Z(g4190) ) ;
AND2    gate6666  (.A(g1126), .B(g3531), .Z(g4192) ) ;
AND2    gate6667  (.A(g145), .B(g2727), .Z(g4193) ) ;
AND4    gate6668  (.A(g2162), .B(g2149), .C(g2137), .D(g2106), .Z(II8089) ) ;
AND4    gate6669  (.A(g3316), .B(g2057), .C(g2020), .D(g3238), .Z(II8090) ) ;
AND2    gate6670  (.A(II8089), .B(II8090), .Z(g4194) ) ;
AND2    gate6671  (.A(g93), .B(g2769), .Z(g4199) ) ;
AND4    gate6672  (.A(g2162), .B(g2149), .C(g2137), .D(g2106), .Z(II8108) ) ;
AND4    gate6673  (.A(g2074), .B(g3287), .C(g3264), .D(g3238), .Z(II8109) ) ;
AND2    gate6674  (.A(II8108), .B(II8109), .Z(g4201) ) ;
AND4    gate6675  (.A(g2162), .B(g2149), .C(g2137), .D(g2106), .Z(II8114) ) ;
AND4    gate6676  (.A(g2074), .B(g3287), .C(g3264), .D(g1987), .Z(II8115) ) ;
AND2    gate6677  (.A(II8114), .B(II8115), .Z(g4216) ) ;
AND4    gate6678  (.A(g3533), .B(g3549), .C(g3568), .D(g3583), .Z(g4220) ) ;
AND3    gate6679  (.A(g2699), .B(g2674), .C(g2677), .Z(II8127) ) ;
AND3    gate6680  (.A(g2680), .B(g2683), .C(II8127), .Z(g4224) ) ;
AND4    gate6681  (.A(g2686), .B(g2689), .C(g2692), .D(g2695), .Z(g4225) ) ;
AND3    gate6682  (.A(g2674), .B(g2677), .C(g2680), .Z(II8143) ) ;
AND3    gate6683  (.A(g2683), .B(g3491), .C(II8143), .Z(g4230) ) ;
NOR2    gate6684  (.A(g1728), .B(g2490), .Z(g3260) ) ;
NAND2   gate6685  (.A(II6877), .B(II6878), .Z(g3221) ) ;
AND3    gate6686  (.A(g2686), .B(g2689), .C(g2692), .Z(II8157) ) ;
AND3    gate6687  (.A(g2695), .B(g2698), .C(II8157), .Z(g4238) ) ;
AND2    gate6688  (.A(g1541), .B(g3222), .Z(g4239) ) ;
AND2    gate6689  (.A(g1106), .B(g3226), .Z(g4246) ) ;
AND3    gate6690  (.A(g3583), .B(g3568), .C(g3549), .Z(g4254) ) ;
AND4    gate6691  (.A(g3778), .B(g3549), .C(g3568), .D(g3583), .Z(II8186) ) ;
AND4    gate6692  (.A(g3605), .B(g3644), .C(g3635), .D(II8186), .Z(g4255) ) ;
AND3    gate6693  (.A(g2298), .B(g2316), .C(g2334), .Z(II8209) ) ;
AND3    gate6694  (.A(g2354), .B(g3563), .C(II8209), .Z(g4269) ) ;
AND2    gate6695  (.A(g3666), .B(g3684), .Z(g4271) ) ;
NOR2    gate6696  (.A(g1714), .B(g1459), .Z(g3233) ) ;
NAND2   gate6697  (.A(II6905), .B(II6906), .Z(g3286) ) ;
AND2    gate6698  (.A(g2216), .B(g2618), .Z(g4276) ) ;
AND2    gate6699  (.A(g3549), .B(g3568), .Z(g4282) ) ;
NAND2   gate6700  (.A(II6917), .B(II6918), .Z(g3314) ) ;
AND3    gate6701  (.A(g2298), .B(g2316), .C(g2354), .Z(II8237) ) ;
AND4    gate6702  (.A(g3563), .B(g2334), .C(g3579), .D(II8237), .Z(g4287) ) ;
AND4    gate6703  (.A(g2298), .B(g2316), .C(g2334), .D(g2354), .Z(II8240) ) ;
AND4    gate6704  (.A(g3563), .B(g3579), .C(g3603), .D(II8240), .Z(g4288) ) ;
NAND2   gate6705  (.A(II6940), .B(II6941), .Z(g3358) ) ;
AND2    gate6706  (.A(g2784), .B(g3779), .Z(g4304) ) ;
AND4    gate6707  (.A(g3666), .B(g3684), .C(g3694), .D(g3707), .Z(g4312) ) ;
AND3    gate6708  (.A(g3694), .B(g3684), .C(g3666), .Z(g4314) ) ;
AND3    gate6709  (.A(g3666), .B(g3684), .C(g3694), .Z(II8288) ) ;
AND3    gate6710  (.A(g3707), .B(g3728), .C(II8288), .Z(g4315) ) ;
AND3    gate6711  (.A(g3666), .B(g3684), .C(g3707), .Z(II8296) ) ;
AND4    gate6712  (.A(g3728), .B(g3694), .C(g3750), .D(II8296), .Z(g4319) ) ;
AND4    gate6713  (.A(g3666), .B(g3684), .C(g3694), .D(g3707), .Z(II8299) ) ;
AND4    gate6714  (.A(g3728), .B(g3750), .C(g3768), .D(II8299), .Z(g4320) ) ;
AND2    gate6715  (.A(g1087), .B(g2782), .Z(g4333) ) ;
AND2    gate6716  (.A(g225), .B(g3097), .Z(g4334) ) ;
AND2    gate6717  (.A(g228), .B(g3097), .Z(g4342) ) ;
AND2    gate6718  (.A(g306), .B(g3131), .Z(g4343) ) ;
AND2    gate6719  (.A(g309), .B(g3131), .Z(g4351) ) ;
AND2    gate6720  (.A(g387), .B(g3160), .Z(g4352) ) ;
AND2    gate6721  (.A(g390), .B(g3160), .Z(g4355) ) ;
AND2    gate6722  (.A(g468), .B(g3192), .Z(g4356) ) ;
AND2    gate6723  (.A(g471), .B(g3192), .Z(g4361) ) ;
AND2    gate6724  (.A(g237), .B(g3097), .Z(g4365) ) ;
AND2    gate6725  (.A(g216), .B(g3097), .Z(g4366) ) ;
AND2    gate6726  (.A(g240), .B(g3097), .Z(g4367) ) ;
AND2    gate6727  (.A(g318), .B(g3131), .Z(g4368) ) ;
AND2    gate6728  (.A(g580), .B(g2845), .Z(g4369) ) ;
AND2    gate6729  (.A(g219), .B(g3097), .Z(g4375) ) ;
AND2    gate6730  (.A(g243), .B(g3097), .Z(g4376) ) ;
AND2    gate6731  (.A(g297), .B(g3131), .Z(g4377) ) ;
AND2    gate6732  (.A(g321), .B(g3131), .Z(g4378) ) ;
AND2    gate6733  (.A(g399), .B(g3160), .Z(g4379) ) ;
AND2    gate6734  (.A(g584), .B(g2845), .Z(g4380) ) ;
AND2    gate6735  (.A(g222), .B(g3097), .Z(g4383) ) ;
AND2    gate6736  (.A(g246), .B(g3097), .Z(g4384) ) ;
AND2    gate6737  (.A(g300), .B(g3131), .Z(g4385) ) ;
AND2    gate6738  (.A(g324), .B(g3131), .Z(g4386) ) ;
AND2    gate6739  (.A(g378), .B(g3160), .Z(g4387) ) ;
AND2    gate6740  (.A(g402), .B(g3160), .Z(g4388) ) ;
AND2    gate6741  (.A(g480), .B(g3192), .Z(g4389) ) ;
AND2    gate6742  (.A(g560), .B(g2845), .Z(g4390) ) ;
AND2    gate6743  (.A(g249), .B(g3097), .Z(g4391) ) ;
AND2    gate6744  (.A(g303), .B(g3131), .Z(g4392) ) ;
AND2    gate6745  (.A(g327), .B(g3131), .Z(g4393) ) ;
AND2    gate6746  (.A(g381), .B(g3160), .Z(g4394) ) ;
AND2    gate6747  (.A(g405), .B(g3160), .Z(g4395) ) ;
AND2    gate6748  (.A(g459), .B(g3192), .Z(g4396) ) ;
AND2    gate6749  (.A(g483), .B(g3192), .Z(g4397) ) ;
AND2    gate6750  (.A(g567), .B(g2845), .Z(g4398) ) ;
AND2    gate6751  (.A(g1138), .B(g3614), .Z(g4400) ) ;
AND4    gate6752  (.A(g3430), .B(g3398), .C(g3359), .D(g3341), .Z(II8400) ) ;
AND4    gate6753  (.A(g3316), .B(g3287), .C(g3264), .D(g3238), .Z(II8401) ) ;
AND2    gate6754  (.A(II8400), .B(II8401), .Z(g4403) ) ;
AND2    gate6755  (.A(g252), .B(g3097), .Z(g4407) ) ;
AND2    gate6756  (.A(g330), .B(g3131), .Z(g4408) ) ;
AND2    gate6757  (.A(g384), .B(g3160), .Z(g4409) ) ;
AND2    gate6758  (.A(g408), .B(g3160), .Z(g4410) ) ;
AND2    gate6759  (.A(g462), .B(g3192), .Z(g4411) ) ;
AND2    gate6760  (.A(g486), .B(g3192), .Z(g4412) ) ;
AND4    gate6761  (.A(g3430), .B(g3398), .C(g3359), .D(g3341), .Z(II8412) ) ;
AND4    gate6762  (.A(g3316), .B(g3287), .C(g3264), .D(g1987), .Z(II8413) ) ;
AND2    gate6763  (.A(II8412), .B(II8413), .Z(g4414) ) ;
AND4    gate6764  (.A(g3430), .B(g3398), .C(g3359), .D(g2106), .Z(II8417) ) ;
AND4    gate6765  (.A(g3316), .B(g3287), .C(g3264), .D(g3238), .Z(II8418) ) ;
AND2    gate6766  (.A(II8417), .B(II8418), .Z(g4417) ) ;
AND2    gate6767  (.A(g275), .B(g3097), .Z(g4420) ) ;
AND2    gate6768  (.A(g333), .B(g3131), .Z(g4421) ) ;
AND2    gate6769  (.A(g411), .B(g3160), .Z(g4422) ) ;
AND2    gate6770  (.A(g465), .B(g3192), .Z(g4423) ) ;
AND2    gate6771  (.A(g489), .B(g3192), .Z(g4424) ) ;
AND2    gate6772  (.A(g536), .B(g2845), .Z(g4425) ) ;
AND4    gate6773  (.A(g3430), .B(g3398), .C(g3359), .D(g3341), .Z(II8431) ) ;
AND4    gate6774  (.A(g3316), .B(g3287), .C(g2020), .D(g3238), .Z(II8432) ) ;
AND2    gate6775  (.A(II8431), .B(II8432), .Z(g4427) ) ;
AND4    gate6776  (.A(g3430), .B(g3398), .C(g3359), .D(g2106), .Z(II8436) ) ;
AND4    gate6777  (.A(g3316), .B(g3287), .C(g3264), .D(g1987), .Z(II8437) ) ;
AND2    gate6778  (.A(II8436), .B(II8437), .Z(g4430) ) ;
AND2    gate6779  (.A(g278), .B(g3097), .Z(g4433) ) ;
AND2    gate6780  (.A(g356), .B(g3131), .Z(g4434) ) ;
AND2    gate6781  (.A(g414), .B(g3160), .Z(g4435) ) ;
AND2    gate6782  (.A(g492), .B(g3192), .Z(g4436) ) ;
AND2    gate6783  (.A(g540), .B(g2845), .Z(g4437) ) ;
AND4    gate6784  (.A(g3430), .B(g3398), .C(g3359), .D(g3341), .Z(II8455) ) ;
AND4    gate6785  (.A(g3316), .B(g3287), .C(g2020), .D(g1987), .Z(II8456) ) ;
AND2    gate6786  (.A(II8455), .B(II8456), .Z(g4445) ) ;
AND4    gate6787  (.A(g3430), .B(g3398), .C(g3359), .D(g2106), .Z(II8460) ) ;
AND4    gate6788  (.A(g3316), .B(g3287), .C(g2020), .D(g3238), .Z(II8461) ) ;
AND2    gate6789  (.A(II8460), .B(II8461), .Z(g4448) ) ;
AND2    gate6790  (.A(g359), .B(g3131), .Z(g4451) ) ;
AND2    gate6791  (.A(g437), .B(g3160), .Z(g4452) ) ;
AND2    gate6792  (.A(g495), .B(g3192), .Z(g4453) ) ;
AND2    gate6793  (.A(g544), .B(g2845), .Z(g4454) ) ;
AND4    gate6794  (.A(g3430), .B(g3398), .C(g3359), .D(g3341), .Z(II8490) ) ;
AND4    gate6795  (.A(g3316), .B(g2057), .C(g3264), .D(g3238), .Z(II8491) ) ;
AND2    gate6796  (.A(II8490), .B(II8491), .Z(g4466) ) ;
AND4    gate6797  (.A(g3430), .B(g3398), .C(g3359), .D(g2106), .Z(II8495) ) ;
AND4    gate6798  (.A(g3316), .B(g3287), .C(g2020), .D(g1987), .Z(II8496) ) ;
AND2    gate6799  (.A(II8495), .B(II8496), .Z(g4469) ) ;
AND2    gate6800  (.A(g440), .B(g3160), .Z(g4472) ) ;
AND2    gate6801  (.A(g518), .B(g3192), .Z(g4473) ) ;
AND4    gate6802  (.A(g3430), .B(g3398), .C(g3359), .D(g3341), .Z(II8523) ) ;
AND4    gate6803  (.A(g3316), .B(g2057), .C(g3264), .D(g1987), .Z(II8524) ) ;
AND2    gate6804  (.A(II8523), .B(II8524), .Z(g4483) ) ;
AND4    gate6805  (.A(g3430), .B(g3398), .C(g3359), .D(g2106), .Z(II8528) ) ;
AND4    gate6806  (.A(g3316), .B(g2057), .C(g3264), .D(g3238), .Z(II8529) ) ;
AND2    gate6807  (.A(II8528), .B(II8529), .Z(g4486) ) ;
AND2    gate6808  (.A(g521), .B(g3192), .Z(g4490) ) ;
AND2    gate6809  (.A(g557), .B(g2845), .Z(g4491) ) ;
AND4    gate6810  (.A(g3430), .B(g3398), .C(g3359), .D(g3341), .Z(II8546) ) ;
AND4    gate6811  (.A(g3316), .B(g2057), .C(g2020), .D(g3238), .Z(II8547) ) ;
AND2    gate6812  (.A(II8546), .B(II8547), .Z(g4494) ) ;
AND4    gate6813  (.A(g3430), .B(g3398), .C(g3359), .D(g2106), .Z(II8551) ) ;
AND4    gate6814  (.A(g3316), .B(g2057), .C(g3264), .D(g1987), .Z(II8552) ) ;
AND2    gate6815  (.A(II8551), .B(II8552), .Z(g4497) ) ;
AND4    gate6816  (.A(g3430), .B(g3398), .C(g3359), .D(g3341), .Z(II8568) ) ;
AND4    gate6817  (.A(g3316), .B(g2057), .C(g2020), .D(g1987), .Z(II8569) ) ;
AND2    gate6818  (.A(II8568), .B(II8569), .Z(g4504) ) ;
AND4    gate6819  (.A(g3430), .B(g3398), .C(g3359), .D(g2106), .Z(II8573) ) ;
AND4    gate6820  (.A(g3316), .B(g2057), .C(g2020), .D(g3238), .Z(II8574) ) ;
AND2    gate6821  (.A(II8573), .B(II8574), .Z(g4507) ) ;
AND4    gate6822  (.A(g3430), .B(g3398), .C(g3359), .D(g3341), .Z(II8588) ) ;
AND4    gate6823  (.A(g2074), .B(g3287), .C(g3264), .D(g3238), .Z(II8589) ) ;
AND2    gate6824  (.A(II8588), .B(II8589), .Z(g4514) ) ;
AND4    gate6825  (.A(g3430), .B(g3398), .C(g3359), .D(g2106), .Z(II8593) ) ;
AND4    gate6826  (.A(g3316), .B(g2057), .C(g2020), .D(g1987), .Z(II8594) ) ;
AND2    gate6827  (.A(II8593), .B(II8594), .Z(g4517) ) ;
AND2    gate6828  (.A(g2642), .B(g741), .Z(g4526) ) ;
AND4    gate6829  (.A(g3430), .B(g3398), .C(g3359), .D(g3341), .Z(II8612) ) ;
AND4    gate6830  (.A(g2074), .B(g3287), .C(g3264), .D(g1987), .Z(II8613) ) ;
AND2    gate6831  (.A(II8612), .B(II8613), .Z(g4529) ) ;
AND4    gate6832  (.A(g3430), .B(g3398), .C(g3359), .D(g2106), .Z(II8617) ) ;
AND4    gate6833  (.A(g2074), .B(g3287), .C(g3264), .D(g3238), .Z(II8618) ) ;
AND2    gate6834  (.A(II8617), .B(II8618), .Z(g4532) ) ;
AND2    gate6835  (.A(g2643), .B(g746), .Z(g4546) ) ;
AND4    gate6836  (.A(g3430), .B(g3398), .C(g3359), .D(g2106), .Z(II8642) ) ;
AND4    gate6837  (.A(g2074), .B(g3287), .C(g3264), .D(g1987), .Z(II8643) ) ;
AND2    gate6838  (.A(II8642), .B(II8643), .Z(g4549) ) ;
AND2    gate6839  (.A(g4081), .B(g3078), .Z(g4690) ) ;
NAND2   gate6840  (.A(II8120), .B(II8121), .Z(g4219) ) ;
AND2    gate6841  (.A(g1557), .B(g4276), .Z(g4699) ) ;
NAND2   gate6842  (.A(II8165), .B(II8166), .Z(g4243) ) ;
OR2     gate6843  (.A(g202), .B(g3129), .Z(g3986) ) ;
AND2    gate6844  (.A(g812), .B(g4062), .Z(g4707) ) ;
OR2     gate6845  (.A(g196), .B(g2995), .Z(g4072) ) ;
AND2    gate6846  (.A(g1179), .B(g4276), .Z(g4712) ) ;
OR2     gate6847  (.A(g187), .B(g3012), .Z(g4055) ) ;
AND2    gate6848  (.A(g828), .B(g4038), .Z(g4724) ) ;
OR2     gate6849  (.A(g207), .B(g3083), .Z(g4179) ) ;
AND2    gate6850  (.A(g1504), .B(g4059), .Z(g4729) ) ;
AND2    gate6851  (.A(g2242), .B(g4275), .Z(g4740) ) ;
NAND2   gate6852  (.A(II6997), .B(II6998), .Z(g3518) ) ;
AND2    gate6853  (.A(g3518), .B(g4286), .Z(g4743) ) ;
NAND2   gate6854  (.A(II7010), .B(II7011), .Z(g3525) ) ;
AND2    gate6855  (.A(g3525), .B(g4296), .Z(g4744) ) ;
AND2    gate6856  (.A(g948), .B(g4527), .Z(g4783) ) ;
NAND2   gate6857  (.A(II5506), .B(II5507), .Z(g1678) ) ;
AND2    gate6858  (.A(g1678), .B(g4202), .Z(g4785) ) ;
AND2    gate6859  (.A(g953), .B(g4547), .Z(g4787) ) ;
NAND2   gate6860  (.A(II6500), .B(II6501), .Z(g2751) ) ;
AND2    gate6861  (.A(g2751), .B(g4202), .Z(g4789) ) ;
AND2    gate6862  (.A(g949), .B(g4562), .Z(g4791) ) ;
NAND2   gate6863  (.A(II7429), .B(II7430), .Z(g3887) ) ;
AND2    gate6864  (.A(g3887), .B(g4202), .Z(g4793) ) ;
AND2    gate6865  (.A(g954), .B(g4574), .Z(g4794) ) ;
AND2    gate6866  (.A(g950), .B(g4584), .Z(g4796) ) ;
NAND2   gate6867  (.A(II7453), .B(II7454), .Z(g3893) ) ;
AND2    gate6868  (.A(g3893), .B(g1616), .Z(g4797) ) ;
AND2    gate6869  (.A(g951), .B(g4596), .Z(g4799) ) ;
AND2    gate6870  (.A(g952), .B(g3876), .Z(g4804) ) ;
AND3    gate6871  (.A(g4041), .B(g2595), .C(g2584), .Z(II9166) ) ;
AND3    gate6872  (.A(g4238), .B(g4230), .C(g174), .Z(g4823) ) ;
NAND2   gate6873  (.A(g1408), .B(g2665), .Z(g4228) ) ;
AND2    gate6874  (.A(g1545), .B(g4239), .Z(g4826) ) ;
AND2    gate6875  (.A(g4288), .B(g3723), .Z(g4830) ) ;
AND2    gate6876  (.A(g1110), .B(g4246), .Z(g4832) ) ;
AND3    gate6877  (.A(g2605), .B(g4044), .C(g2584), .Z(II9202) ) ;
NAND2   gate6878  (.A(g1415), .B(g2668), .Z(g4235) ) ;
NAND2   gate6879  (.A(II8133), .B(II8134), .Z(g4227) ) ;
NOR2    gate6880  (.A(g1231), .B(g2834), .Z(g4160) ) ;
AND3    gate6881  (.A(g1924), .B(g4225), .C(g4224), .Z(g4872) ) ;
AND4    gate6882  (.A(g3746), .B(g3723), .C(g4288), .D(g3764), .Z(g4877) ) ;
AND3    gate6883  (.A(g4041), .B(g4044), .C(g2584), .Z(II9222) ) ;
AND3    gate6884  (.A(g3746), .B(g3723), .C(g4288), .Z(g4883) ) ;
AND3    gate6885  (.A(g3777), .B(g3764), .C(g3746), .Z(II9261) ) ;
AND3    gate6886  (.A(g3723), .B(g4288), .C(II9261), .Z(g4901) ) ;
AND4    gate6887  (.A(g4304), .B(g2770), .C(g2746), .D(g2728), .Z(g4902) ) ;
AND2    gate6888  (.A(g4320), .B(g2728), .Z(g4906) ) ;
AND4    gate6889  (.A(g2746), .B(g2728), .C(g4320), .D(g2770), .Z(g4933) ) ;
AND2    gate6890  (.A(g214), .B(g3888), .Z(g4936) ) ;
NAND3   gate6891  (.A(g3002), .B(g3124), .C(g3659), .Z(g4309) ) ;
AND2    gate6892  (.A(g3086), .B(g4309), .Z(g4937) ) ;
AND2    gate6893  (.A(g215), .B(g3891), .Z(g4955) ) ;
AND2    gate6894  (.A(g295), .B(g3892), .Z(g4956) ) ;
AND3    gate6895  (.A(g2746), .B(g2728), .C(g4320), .Z(g4957) ) ;
AND2    gate6896  (.A(g296), .B(g3897), .Z(g4958) ) ;
AND2    gate6897  (.A(g376), .B(g3898), .Z(g4959) ) ;
AND2    gate6898  (.A(g377), .B(g3904), .Z(g4961) ) ;
AND2    gate6899  (.A(g457), .B(g3905), .Z(g4962) ) ;
AND2    gate6900  (.A(g458), .B(g3912), .Z(g5001) ) ;
AND3    gate6901  (.A(g2784), .B(g2770), .C(g2746), .Z(II9330) ) ;
AND3    gate6902  (.A(g2728), .B(g4320), .C(II9330), .Z(g5005) ) ;
AND2    gate6903  (.A(g231), .B(g3920), .Z(g5008) ) ;
AND2    gate6904  (.A(g211), .B(g3928), .Z(g5017) ) ;
AND2    gate6905  (.A(g232), .B(g3930), .Z(g5018) ) ;
AND2    gate6906  (.A(g312), .B(g3933), .Z(g5019) ) ;
AND2    gate6907  (.A(g579), .B(g3937), .Z(g5020) ) ;
AND2    gate6908  (.A(g212), .B(g3945), .Z(g5029) ) ;
AND2    gate6909  (.A(g233), .B(g3946), .Z(g5030) ) ;
AND2    gate6910  (.A(g292), .B(g3948), .Z(g5031) ) ;
AND2    gate6911  (.A(g313), .B(g3950), .Z(g5032) ) ;
AND2    gate6912  (.A(g393), .B(g3953), .Z(g5033) ) ;
AND2    gate6913  (.A(g583), .B(g3956), .Z(g5034) ) ;
AND2    gate6914  (.A(g213), .B(g3958), .Z(g5043) ) ;
AND2    gate6915  (.A(g234), .B(g3959), .Z(g5044) ) ;
AND2    gate6916  (.A(g293), .B(g3961), .Z(g5045) ) ;
AND2    gate6917  (.A(g314), .B(g3962), .Z(g5046) ) ;
AND2    gate6918  (.A(g373), .B(g3964), .Z(g5047) ) ;
AND2    gate6919  (.A(g394), .B(g3966), .Z(g5048) ) ;
AND2    gate6920  (.A(g474), .B(g3969), .Z(g5049) ) ;
AND2    gate6921  (.A(g587), .B(g3970), .Z(g5050) ) ;
AND2    gate6922  (.A(g235), .B(g3973), .Z(g5062) ) ;
AND2    gate6923  (.A(g294), .B(g3974), .Z(g5063) ) ;
AND2    gate6924  (.A(g315), .B(g3975), .Z(g5064) ) ;
AND2    gate6925  (.A(g374), .B(g3977), .Z(g5065) ) ;
AND2    gate6926  (.A(g395), .B(g3978), .Z(g5066) ) ;
AND2    gate6927  (.A(g454), .B(g3980), .Z(g5067) ) ;
AND2    gate6928  (.A(g475), .B(g3982), .Z(g5068) ) ;
AND2    gate6929  (.A(g566), .B(g3983), .Z(g5069) ) ;
AND2    gate6930  (.A(g236), .B(g3988), .Z(g5077) ) ;
AND2    gate6931  (.A(g316), .B(g3989), .Z(g5078) ) ;
AND2    gate6932  (.A(g375), .B(g3990), .Z(g5079) ) ;
AND2    gate6933  (.A(g396), .B(g3991), .Z(g5080) ) ;
AND2    gate6934  (.A(g455), .B(g3993), .Z(g5081) ) ;
AND2    gate6935  (.A(g476), .B(g3994), .Z(g5082) ) ;
AND2    gate6936  (.A(g273), .B(g3998), .Z(g5089) ) ;
AND2    gate6937  (.A(g317), .B(g4000), .Z(g5090) ) ;
AND2    gate6938  (.A(g397), .B(g4001), .Z(g5091) ) ;
AND2    gate6939  (.A(g456), .B(g4002), .Z(g5092) ) ;
AND2    gate6940  (.A(g477), .B(g4003), .Z(g5093) ) ;
AND2    gate6941  (.A(g535), .B(g4004), .Z(g5094) ) ;
AND2    gate6942  (.A(g1149), .B(g4400), .Z(g5096) ) ;
AND2    gate6943  (.A(g274), .B(g4010), .Z(g5104) ) ;
AND2    gate6944  (.A(g354), .B(g4013), .Z(g5105) ) ;
AND2    gate6945  (.A(g398), .B(g4015), .Z(g5106) ) ;
AND2    gate6946  (.A(g478), .B(g4016), .Z(g5107) ) ;
AND2    gate6947  (.A(g539), .B(g4017), .Z(g5108) ) ;
AND2    gate6948  (.A(g355), .B(g4021), .Z(g5116) ) ;
AND2    gate6949  (.A(g435), .B(g4024), .Z(g5117) ) ;
AND2    gate6950  (.A(g479), .B(g4026), .Z(g5118) ) ;
AND2    gate6951  (.A(g543), .B(g4027), .Z(g5119) ) ;
AND2    gate6952  (.A(g436), .B(g4030), .Z(g5122) ) ;
AND2    gate6953  (.A(g516), .B(g4033), .Z(g5123) ) ;
AND2    gate6954  (.A(g517), .B(g4036), .Z(g5125) ) ;
AND2    gate6955  (.A(g556), .B(g4037), .Z(g5126) ) ;
AND4    gate6956  (.A(g3019), .B(g3029), .C(g3038), .D(g3052), .Z(II9534) ) ;
AND4    gate6957  (.A(g3062), .B(g2712), .C(g4253), .D(g2752), .Z(II9535) ) ;
AND2    gate6958  (.A(II9534), .B(II9535), .Z(g5132) ) ;
AND2    gate6959  (.A(g1677), .B(g4202), .Z(g5142) ) ;
AND2    gate6960  (.A(g1912), .B(g4814), .Z(g5298) ) ;
NAND2   gate6961  (.A(II9170), .B(II9171), .Z(g4820) ) ;
AND2    gate6962  (.A(g4820), .B(g2407), .Z(g5313) ) ;
AND2    gate6963  (.A(g1509), .B(g4729), .Z(g5314) ) ;
NAND2   gate6964  (.A(II9234), .B(II9235), .Z(g4887) ) ;
AND2    gate6965  (.A(g4887), .B(g2424), .Z(g5334) ) ;
AND2    gate6966  (.A(g1528), .B(g4916), .Z(g5425) ) ;
AND2    gate6967  (.A(g1537), .B(g4921), .Z(g5432) ) ;
AND2    gate6968  (.A(g1541), .B(g4926), .Z(g5436) ) ;
AND2    gate6969  (.A(g1545), .B(g4932), .Z(g5438) ) ;
OR2     gate6970  (.A(g4154), .B(g3081), .Z(g4870) ) ;
NAND2   gate6971  (.A(II8939), .B(II8940), .Z(g4679) ) ;
AND2    gate6972  (.A(g4679), .B(g4202), .Z(g5442) ) ;
AND2    gate6973  (.A(g1549), .B(g4935), .Z(g5443) ) ;
OR2     gate6974  (.A(g4159), .B(g4167), .Z(g4876) ) ;
NAND2   gate6975  (.A(II8956), .B(II8957), .Z(g4686) ) ;
AND2    gate6976  (.A(g4686), .B(g1616), .Z(g5458) ) ;
NAND2   gate6977  (.A(II9548), .B(II9549), .Z(g5141) ) ;
AND2    gate6978  (.A(g1037), .B(g5096), .Z(g5484) ) ;
NAND2   gate6979  (.A(II9277), .B(II9278), .Z(g4912) ) ;
NAND2   gate6980  (.A(II9242), .B(II9243), .Z(g4889) ) ;
NAND2   gate6981  (.A(II5696), .B(II5697), .Z(g1819) ) ;
AND2    gate6982  (.A(g4814), .B(g1819), .Z(g5547) ) ;
AND2    gate6983  (.A(g1549), .B(g4826), .Z(g5548) ) ;
AND2    gate6984  (.A(g1114), .B(g4832), .Z(g5552) ) ;
OR2     gate6985  (.A(g4047), .B(g2972), .Z(g5036) ) ;
OR2     gate6986  (.A(g4052), .B(g4058), .Z(g5070) ) ;
NAND2   gate6987  (.A(II5599), .B(II5600), .Z(g1759) ) ;
AND2    gate6988  (.A(g1759), .B(g4841), .Z(g5570) ) ;
NAND2   gate6989  (.A(II6751), .B(II6752), .Z(g3011) ) ;
AND2    gate6990  (.A(g3011), .B(g4841), .Z(g5573) ) ;
NAND2   gate6991  (.A(II7892), .B(II7893), .Z(g4090) ) ;
AND2    gate6992  (.A(g4090), .B(g4841), .Z(g5579) ) ;
NAND2   gate6993  (.A(II5620), .B(II5621), .Z(g1775) ) ;
AND2    gate6994  (.A(g1775), .B(g4969), .Z(g5583) ) ;
NAND2   gate6995  (.A(II9058), .B(II9059), .Z(g4741) ) ;
AND2    gate6996  (.A(g4741), .B(g4841), .Z(g5585) ) ;
NAND2   gate6997  (.A(II6775), .B(II6776), .Z(g3028) ) ;
AND2    gate6998  (.A(g3028), .B(g4969), .Z(g5588) ) ;
NAND2   gate6999  (.A(II7938), .B(II7939), .Z(g4110) ) ;
AND2    gate7000  (.A(g4110), .B(g4969), .Z(g5593) ) ;
NAND2   gate7001  (.A(II9070), .B(II9071), .Z(g4745) ) ;
AND2    gate7002  (.A(g4745), .B(g4969), .Z(g5599) ) ;
OR2     gate7003  (.A(g4333), .B(g3509), .Z(g5140) ) ;
AND2    gate7004  (.A(g1667), .B(g4841), .Z(g5699) ) ;
AND2    gate7005  (.A(g1638), .B(g4969), .Z(g5700) ) ;
AND2    gate7006  (.A(g1532), .B(g4733), .Z(g5714) ) ;
AND2    gate7007  (.A(g1695), .B(g5428), .Z(g5765) ) ;
AND2    gate7008  (.A(g1897), .B(g5287), .Z(g5783) ) ;
AND2    gate7009  (.A(g5395), .B(g3091), .Z(g5817) ) ;
AND2    gate7010  (.A(g1118), .B(g5552), .Z(g5894) ) ;
NAND2   gate7011  (.A(II10010), .B(II10011), .Z(g5562) ) ;
AND2    gate7012  (.A(g5562), .B(g2407), .Z(g5937) ) ;
NAND2   gate7013  (.A(II10018), .B(II10019), .Z(g5564) ) ;
AND2    gate7014  (.A(g5564), .B(g2424), .Z(g5969) ) ;
NAND2   gate7015  (.A(II10093), .B(II10094), .Z(g5605) ) ;
AND2    gate7016  (.A(g5605), .B(g2424), .Z(g5970) ) ;
AND2    gate7017  (.A(g1041), .B(g5484), .Z(g5984) ) ;
NAND2   gate7018  (.A(II9954), .B(II9955), .Z(g5540) ) ;
AND2    gate7019  (.A(g5540), .B(g2407), .Z(g6001) ) ;
NAND2   gate7020  (.A(II9947), .B(II9948), .Z(g5539) ) ;
AND2    gate7021  (.A(g5539), .B(g2407), .Z(g6002) ) ;
AND3    gate7022  (.A(g3769), .B(g3754), .C(g3735), .Z(II10597) ) ;
NAND2   gate7023  (.A(II9993), .B(II9994), .Z(g5557) ) ;
AND2    gate7024  (.A(g5557), .B(g2407), .Z(g6005) ) ;
NAND2   gate7025  (.A(II10039), .B(II10040), .Z(g5575) ) ;
AND2    gate7026  (.A(g5575), .B(g2424), .Z(g6006) ) ;
NAND2   gate7027  (.A(II10061), .B(II10062), .Z(g5589) ) ;
AND2    gate7028  (.A(g5589), .B(g2424), .Z(g6013) ) ;
NAND2   gate7029  (.A(II10072), .B(II10073), .Z(g5594) ) ;
AND2    gate7030  (.A(g5594), .B(g2424), .Z(g6021) ) ;
NAND2   gate7031  (.A(II10079), .B(II10080), .Z(g5595) ) ;
AND2    gate7032  (.A(g5595), .B(g2424), .Z(g6022) ) ;
AND2    gate7033  (.A(g1037), .B(g5574), .Z(g6039) ) ;
AND2    gate7034  (.A(g1462), .B(g5578), .Z(g6040) ) ;
NAND2   gate7035  (.A(II9692), .B(II9693), .Z(g5189) ) ;
AND2    gate7036  (.A(g5189), .B(g4969), .Z(g6041) ) ;
AND2    gate7037  (.A(g1041), .B(g5581), .Z(g6042) ) ;
AND2    gate7038  (.A(g1069), .B(g5582), .Z(g6043) ) ;
AND2    gate7039  (.A(g1467), .B(g5584), .Z(g6044) ) ;
AND2    gate7040  (.A(g1472), .B(g5591), .Z(g6045) ) ;
AND2    gate7041  (.A(g1073), .B(g5592), .Z(g6046) ) ;
AND2    gate7042  (.A(g1477), .B(g5596), .Z(g6047) ) ;
AND2    gate7043  (.A(g1045), .B(g5597), .Z(g6049) ) ;
AND2    gate7044  (.A(g1049), .B(g5604), .Z(g6052) ) ;
AND2    gate7045  (.A(g1053), .B(g5608), .Z(g6053) ) ;
AND2    gate7046  (.A(g1057), .B(g5611), .Z(g6054) ) ;
NAND2   gate7047  (.A(II9746), .B(II9747), .Z(g5239) ) ;
AND2    gate7048  (.A(g5239), .B(g4202), .Z(g6055) ) ;
OR2     gate7049  (.A(II7232), .B(II7233), .Z(g3760) ) ;
AND2    gate7050  (.A(g1061), .B(g5617), .Z(g6057) ) ;
OR2     gate7051  (.A(g4168), .B(g4797), .Z(g5561) ) ;
AND2    gate7052  (.A(g5561), .B(g3501), .Z(g6058) ) ;
AND2    gate7053  (.A(g1065), .B(g5623), .Z(g6060) ) ;
NAND2   gate7054  (.A(II9768), .B(II9769), .Z(g5257) ) ;
AND2    gate7055  (.A(g5257), .B(g1616), .Z(g6061) ) ;
NAND2   gate7056  (.A(II10224), .B(II10225), .Z(g5712) ) ;
NAND2   gate7057  (.A(g5132), .B(g2043), .Z(g5681) ) ;
AND2    gate7058  (.A(g5618), .B(g2817), .Z(g6105) ) ;
AND2    gate7059  (.A(g5478), .B(g1849), .Z(g6107) ) ;
AND2    gate7060  (.A(g5453), .B(g5335), .Z(g6109) ) ;
OR2     gate7061  (.A(g4823), .B(g4872), .Z(g5673) ) ;
AND3    gate7062  (.A(g5673), .B(g4841), .C(g5541), .Z(g6112) ) ;
AND2    gate7063  (.A(g1489), .B(g5705), .Z(g6145) ) ;
AND2    gate7064  (.A(g1494), .B(g5709), .Z(g6151) ) ;
AND2    gate7065  (.A(g1499), .B(g5713), .Z(g6154) ) ;
AND2    gate7066  (.A(g1130), .B(g5717), .Z(g6157) ) ;
AND2    gate7067  (.A(g1504), .B(g5718), .Z(g6160) ) ;
AND2    gate7068  (.A(g1134), .B(g5724), .Z(g6162) ) ;
AND2    gate7069  (.A(g1509), .B(g5725), .Z(g6166) ) ;
AND2    gate7070  (.A(g1138), .B(g5191), .Z(g6168) ) ;
NAND2   gate7071  (.A(II9827), .B(II9828), .Z(g5363) ) ;
AND2    gate7072  (.A(g5363), .B(g4841), .Z(g6171) ) ;
AND2    gate7073  (.A(g1514), .B(g5192), .Z(g6172) ) ;
NAND2   gate7074  (.A(g3681), .B(g2368), .Z(g4332) ) ;
NOR3    gate7075  (.A(g3002), .B(g1590), .C(g4714), .Z(g5614) ) ;
AND2    gate7076  (.A(g4332), .B(g5614), .Z(g6175) ) ;
AND2    gate7077  (.A(g1149), .B(g5198), .Z(g6176) ) ;
AND2    gate7078  (.A(g1519), .B(g5199), .Z(g6182) ) ;
OR2     gate7079  (.A(g4318), .B(g1590), .Z(g4927) ) ;
NOR2    gate7080  (.A(g4714), .B(g3002), .Z(g5615) ) ;
AND2    gate7081  (.A(g4927), .B(g5615), .Z(g6196) ) ;
AND2    gate7082  (.A(g5542), .B(g5294), .Z(g6204) ) ;
AND2    gate7083  (.A(g1514), .B(g5314), .Z(g6239) ) ;
AND2    gate7084  (.A(g1481), .B(g5285), .Z(g6266) ) ;
AND2    gate7085  (.A(g1092), .B(g5309), .Z(g6268) ) ;
AND2    gate7086  (.A(g5988), .B(g5494), .Z(g6394) ) ;
AND2    gate7087  (.A(g2157), .B(g6007), .Z(g6395) ) ;
AND2    gate7088  (.A(g661), .B(g6008), .Z(g6396) ) ;
AND2    gate7089  (.A(g5971), .B(g5494), .Z(g6399) ) ;
AND2    gate7090  (.A(g150), .B(g6011), .Z(g6400) ) ;
AND2    gate7091  (.A(g5971), .B(g5367), .Z(g6401) ) ;
AND2    gate7092  (.A(g665), .B(g6012), .Z(g6402) ) ;
AND2    gate7093  (.A(g5956), .B(g5494), .Z(g6405) ) ;
AND2    gate7094  (.A(g154), .B(g6018), .Z(g6406) ) ;
AND2    gate7095  (.A(g5956), .B(g5367), .Z(g6407) ) ;
AND2    gate7096  (.A(g669), .B(g6019), .Z(g6408) ) ;
AND2    gate7097  (.A(g706), .B(g6020), .Z(g6409) ) ;
AND2    gate7098  (.A(g5918), .B(g5494), .Z(g6411) ) ;
AND2    gate7099  (.A(g158), .B(g6024), .Z(g6412) ) ;
AND2    gate7100  (.A(g5939), .B(g5367), .Z(g6413) ) ;
AND2    gate7101  (.A(g673), .B(g6025), .Z(g6414) ) ;
AND2    gate7102  (.A(g5988), .B(g5367), .Z(g6415) ) ;
AND2    gate7103  (.A(g710), .B(g6026), .Z(g6416) ) ;
AND2    gate7104  (.A(g718), .B(g6027), .Z(g6417) ) ;
AND2    gate7105  (.A(g5897), .B(g5494), .Z(g6418) ) ;
AND2    gate7106  (.A(g162), .B(g6032), .Z(g6419) ) ;
AND2    gate7107  (.A(g5918), .B(g5367), .Z(g6420) ) ;
AND2    gate7108  (.A(g5847), .B(g5384), .Z(g6421) ) ;
AND2    gate7109  (.A(g714), .B(g6033), .Z(g6422) ) ;
AND2    gate7110  (.A(g5897), .B(g5384), .Z(g6423) ) ;
AND2    gate7111  (.A(g5874), .B(g5494), .Z(g6428) ) ;
AND2    gate7112  (.A(g168), .B(g6035), .Z(g6429) ) ;
AND2    gate7113  (.A(g5874), .B(g5384), .Z(g6430) ) ;
AND2    gate7114  (.A(g5847), .B(g5494), .Z(g6431) ) ;
AND2    gate7115  (.A(g778), .B(g6134), .Z(g6433) ) ;
AND2    gate7116  (.A(g855), .B(g6048), .Z(g6434) ) ;
AND2    gate7117  (.A(g859), .B(g6050), .Z(g6437) ) ;
OR2     gate7118  (.A(g863), .B(g4051), .Z(g4829) ) ;
AND2    gate7119  (.A(g4829), .B(g6051), .Z(g6438) ) ;
AND2    gate7120  (.A(g789), .B(g6150), .Z(g6439) ) ;
AND2    gate7121  (.A(g1676), .B(g6125), .Z(g6444) ) ;
AND2    gate7122  (.A(g734), .B(g6073), .Z(g6447) ) ;
AND2    gate7123  (.A(g5918), .B(g5384), .Z(g6448) ) ;
OR2     gate7124  (.A(g5546), .B(g4681), .Z(g6116) ) ;
AND2    gate7125  (.A(g6116), .B(g2407), .Z(g6456) ) ;
NAND2   gate7126  (.A(g2205), .B(g5568), .Z(g6178) ) ;
NAND2   gate7127  (.A(II10981), .B(II10982), .Z(g6215) ) ;
AND2    gate7128  (.A(g6215), .B(g2424), .Z(g6462) ) ;
NAND2   gate7129  (.A(II10889), .B(II10890), .Z(g6177) ) ;
AND2    gate7130  (.A(g6177), .B(g2424), .Z(g6464) ) ;
NAND2   gate7131  (.A(II10953), .B(II10954), .Z(g6203) ) ;
AND2    gate7132  (.A(g6203), .B(g2424), .Z(g6474) ) ;
NAND2   gate7133  (.A(II10314), .B(II10315), .Z(g5750) ) ;
AND2    gate7134  (.A(g5750), .B(g4969), .Z(g6487) ) ;
OR2     gate7135  (.A(g4175), .B(g5458), .Z(g6144) ) ;
AND2    gate7136  (.A(g6144), .B(g3510), .Z(g6541) ) ;
NAND2   gate7137  (.A(II10360), .B(II10361), .Z(g5762) ) ;
AND2    gate7138  (.A(g5762), .B(g1616), .Z(g6554) ) ;
NAND2   gate7139  (.A(II11079), .B(II11080), .Z(g6265) ) ;
AND2    gate7140  (.A(g6265), .B(g2424), .Z(g6567) ) ;
AND2    gate7141  (.A(g1045), .B(g5984), .Z(g6574) ) ;
NAND2   gate7142  (.A(II10790), .B(II10791), .Z(g6142) ) ;
NAND2   gate7143  (.A(II10992), .B(II10993), .Z(g6218) ) ;
AND2    gate7144  (.A(g6218), .B(g3913), .Z(g6578) ) ;
AND2    gate7145  (.A(g1122), .B(g5894), .Z(g6582) ) ;
OR2     gate7146  (.A(g4066), .B(g5313), .Z(g6249) ) ;
NAND2   gate7147  (.A(II10626), .B(II10627), .Z(g6023) ) ;
AND2    gate7148  (.A(g6023), .B(g4841), .Z(g6629) ) ;
AND2    gate7149  (.A(g5526), .B(g5987), .Z(g6633) ) ;
AND2    gate7150  (.A(g174), .B(g5755), .Z(g6638) ) ;
AND2    gate7151  (.A(g5939), .B(g5494), .Z(g6641) ) ;
AND2    gate7152  (.A(g1519), .B(g6239), .Z(g6689) ) ;
AND2    gate7153  (.A(g677), .B(g5843), .Z(g6715) ) ;
AND2    gate7154  (.A(g5897), .B(g5367), .Z(g6726) ) ;
AND2    gate7155  (.A(g681), .B(g5846), .Z(g6727) ) ;
AND2    gate7156  (.A(g5874), .B(g5367), .Z(g6732) ) ;
AND2    gate7157  (.A(g685), .B(g5873), .Z(g6733) ) ;
AND2    gate7158  (.A(g5847), .B(g5367), .Z(g6738) ) ;
AND2    gate7159  (.A(g730), .B(g5916), .Z(g6743) ) ;
AND2    gate7160  (.A(g5939), .B(g5384), .Z(g6753) ) ;
AND2    gate7161  (.A(g5874), .B(g5412), .Z(g6757) ) ;
AND2    gate7162  (.A(g5847), .B(g5412), .Z(g6762) ) ;
AND2    gate7163  (.A(g146), .B(g6004), .Z(g6771) ) ;
AND2    gate7164  (.A(g6478), .B(g5246), .Z(g6908) ) ;
AND2    gate7165  (.A(g6483), .B(g5246), .Z(g6914) ) ;
AND2    gate7166  (.A(g6493), .B(g5246), .Z(g6915) ) ;
AND2    gate7167  (.A(g727), .B(g6515), .Z(g6916) ) ;
NAND2   gate7168  (.A(II11751), .B(II11752), .Z(g6570) ) ;
AND2    gate7169  (.A(g6570), .B(g5612), .Z(g6923) ) ;
AND2    gate7170  (.A(g1126), .B(g6582), .Z(g6941) ) ;
OR2     gate7171  (.A(g4740), .B(g4098), .Z(g5483) ) ;
OR2     gate7172  (.A(g4743), .B(g4109), .Z(g5511) ) ;
OR2     gate7173  (.A(g4744), .B(g4118), .Z(g5518) ) ;
NOR3    gate7174  (.A(g5802), .B(g5769), .C(g5790), .Z(g6489) ) ;
AND2    gate7175  (.A(g55), .B(g6489), .Z(g6965) ) ;
OR2     gate7176  (.A(g6039), .B(g6041), .Z(g6580) ) ;
NAND2   gate7177  (.A(II9382), .B(II9383), .Z(g5035) ) ;
AND2    gate7178  (.A(g5035), .B(g6490), .Z(g6970) ) ;
NAND2   gate7179  (.A(II11550), .B(II11551), .Z(g6424) ) ;
AND2    gate7180  (.A(g6424), .B(g4969), .Z(g6971) ) ;
NAND2   gate7181  (.A(II10143), .B(II10144), .Z(g5661) ) ;
AND2    gate7182  (.A(g5661), .B(g6498), .Z(g6972) ) ;
NAND2   gate7183  (.A(II7086), .B(II7087), .Z(g3613) ) ;
NAND2   gate7184  (.A(II8393), .B(II8394), .Z(g4399) ) ;
NAND2   gate7185  (.A(II9476), .B(II9477), .Z(g5095) ) ;
AND2    gate7186  (.A(g5095), .B(g6511), .Z(g6979) ) ;
AND2    gate7187  (.A(g799), .B(g6517), .Z(g6990) ) ;
NAND2   gate7188  (.A(II10197), .B(II10198), .Z(g5689) ) ;
AND2    gate7189  (.A(g5689), .B(g6520), .Z(g6991) ) ;
OR2     gate7190  (.A(g4180), .B(g6061), .Z(g6610) ) ;
AND2    gate7191  (.A(g6610), .B(g3519), .Z(g6992) ) ;
NAND2   gate7192  (.A(II7149), .B(II7150), .Z(g3658) ) ;
AND2    gate7193  (.A(g3658), .B(g6538), .Z(g6994) ) ;
NAND2   gate7194  (.A(II11575), .B(II11576), .Z(g6435) ) ;
AND2    gate7195  (.A(g6435), .B(g1616), .Z(g6995) ) ;
NAND2   gate7196  (.A(II7173), .B(II7174), .Z(g3678) ) ;
NAND2   gate7197  (.A(II8503), .B(II8504), .Z(g4474) ) ;
AND2    gate7198  (.A(g815), .B(g6556), .Z(g6999) ) ;
NAND2   gate7199  (.A(II7215), .B(II7216), .Z(g3722) ) ;
AND2    gate7200  (.A(g3722), .B(g6562), .Z(g7001) ) ;
NAND2   gate7201  (.A(II12180), .B(II12181), .Z(g6770) ) ;
AND2    gate7202  (.A(g1462), .B(g6689), .Z(g7003) ) ;
NAND2   gate7203  (.A(II11874), .B(II11875), .Z(g6627) ) ;
NAND2   gate7204  (.A(II11842), .B(II11843), .Z(g6615) ) ;
AND2    gate7205  (.A(g1049), .B(g6574), .Z(g7010) ) ;
OR2     gate7206  (.A(g4077), .B(g6002), .Z(g6706) ) ;
OR2     gate7207  (.A(g4053), .B(g5937), .Z(g6673) ) ;
OR2     gate7208  (.A(g4073), .B(g6001), .Z(g6698) ) ;
OR2     gate7209  (.A(g6157), .B(g5583), .Z(g6705) ) ;
OR2     gate7210  (.A(g4082), .B(g6005), .Z(g6717) ) ;
OR2     gate7211  (.A(g6162), .B(g5588), .Z(g6716) ) ;
OR2     gate7212  (.A(g6168), .B(g5593), .Z(g6728) ) ;
NAND2   gate7213  (.A(II11615), .B(II11616), .Z(g6466) ) ;
AND2    gate7214  (.A(g6466), .B(g4841), .Z(g7038) ) ;
OR2     gate7215  (.A(g6176), .B(g5599), .Z(g6734) ) ;
AND2    gate7216  (.A(g4259), .B(g6677), .Z(g7079) ) ;
OR2     gate7217  (.A(g6268), .B(g5700), .Z(g6440) ) ;
AND2    gate7218  (.A(g6677), .B(g5101), .Z(g7096) ) ;
OR2     gate7219  (.A(g6406), .B(g6411), .Z(g6926) ) ;
AND2    gate7220  (.A(g4057), .B(g6953), .Z(g7136) ) ;
NAND2   gate7221  (.A(II12551), .B(II12552), .Z(g6893) ) ;
AND2    gate7222  (.A(g6893), .B(g4841), .Z(g7175) ) ;
OR2     gate7223  (.A(g6042), .B(g6487), .Z(g7016) ) ;
OR2     gate7224  (.A(g5425), .B(g4785), .Z(g6121) ) ;
OR2     gate7225  (.A(g5432), .B(g4789), .Z(g6124) ) ;
NAND2   gate7226  (.A(II12576), .B(II12577), .Z(g6902) ) ;
AND2    gate7227  (.A(g6902), .B(g4969), .Z(g7182) ) ;
OR2     gate7228  (.A(g5436), .B(g4793), .Z(g6132) ) ;
AND2    gate7229  (.A(g6132), .B(g7042), .Z(g7183) ) ;
OR2     gate7230  (.A(g5438), .B(g5442), .Z(g6138) ) ;
AND2    gate7231  (.A(g6138), .B(g7043), .Z(g7184) ) ;
OR2     gate7232  (.A(g5443), .B(g6055), .Z(g6600) ) ;
OR2     gate7233  (.A(g4186), .B(g6554), .Z(g7026) ) ;
AND2    gate7234  (.A(g7026), .B(g3526), .Z(g7192) ) ;
NAND2   gate7235  (.A(II12597), .B(II12598), .Z(g6911) ) ;
AND2    gate7236  (.A(g6911), .B(g1616), .Z(g7193) ) ;
AND2    gate7237  (.A(g6984), .B(g4226), .Z(g7195) ) ;
NAND2   gate7238  (.A(II12870), .B(II12871), .Z(g7093) ) ;
AND2    gate7239  (.A(g1467), .B(g7003), .Z(g7199) ) ;
AND2    gate7240  (.A(g1053), .B(g7010), .Z(g7212) ) ;
AND2    gate7241  (.A(g6111), .B(g6984), .Z(g7215) ) ;
OR2     gate7242  (.A(g6145), .B(g5570), .Z(g6688) ) ;
OR2     gate7243  (.A(g6151), .B(g5573), .Z(g6694) ) ;
OR2     gate7244  (.A(g6154), .B(g5579), .Z(g6699) ) ;
OR2     gate7245  (.A(g6160), .B(g5585), .Z(g6707) ) ;
OR2     gate7246  (.A(g6166), .B(g6171), .Z(g6719) ) ;
OR2     gate7247  (.A(g6172), .B(g6629), .Z(g7081) ) ;
OR2     gate7248  (.A(g6266), .B(g5699), .Z(g6436) ) ;
AND2    gate7249  (.A(g6965), .B(g1745), .Z(g7278) ) ;
OR2     gate7250  (.A(g5714), .B(g5142), .Z(g5830) ) ;
AND2    gate7251  (.A(g4065), .B(g7171), .Z(g7323) ) ;
NAND2   gate7252  (.A(II12952), .B(II12953), .Z(g7121) ) ;
AND2    gate7253  (.A(g7121), .B(g4841), .Z(g7412) ) ;
OR2     gate7254  (.A(g6049), .B(g6971), .Z(g7222) ) ;
NAND2   gate7255  (.A(II13003), .B(II13004), .Z(g7140) ) ;
AND2    gate7256  (.A(g7140), .B(g4969), .Z(g7416) ) ;
NAND2   gate7257  (.A(II13017), .B(II13018), .Z(g7144) ) ;
AND2    gate7258  (.A(g7144), .B(g1616), .Z(g7417) ) ;
OR2     gate7259  (.A(g4190), .B(g6995), .Z(g7230) ) ;
AND2    gate7260  (.A(g7230), .B(g3530), .Z(g7419) ) ;
AND2    gate7261  (.A(g1472), .B(g7199), .Z(g7427) ) ;
AND2    gate7262  (.A(g1057), .B(g7212), .Z(g7429) ) ;
OR2     gate7263  (.A(g6182), .B(g7038), .Z(g7272) ) ;
OR2     gate7264  (.A(g7136), .B(g6903), .Z(g7363) ) ;
OR2     gate7265  (.A(g6040), .B(g7175), .Z(g7428) ) ;
NAND2   gate7266  (.A(II13377), .B(II13378), .Z(g7316) ) ;
AND2    gate7267  (.A(g7316), .B(g4841), .Z(g7597) ) ;
AND2    gate7268  (.A(g7483), .B(g3466), .Z(g7598) ) ;
AND2    gate7269  (.A(g7460), .B(g3466), .Z(g7600) ) ;
AND2    gate7270  (.A(g7476), .B(g3466), .Z(g7602) ) ;
AND2    gate7271  (.A(g7456), .B(g3466), .Z(g7604) ) ;
OR2     gate7272  (.A(g6052), .B(g7182), .Z(g7435) ) ;
AND2    gate7273  (.A(g7471), .B(g3466), .Z(g7606) ) ;
NAND2   gate7274  (.A(II13396), .B(II13397), .Z(g7325) ) ;
AND2    gate7275  (.A(g7325), .B(g4969), .Z(g7607) ) ;
AND2    gate7276  (.A(g7467), .B(g3466), .Z(g7609) ) ;
AND2    gate7277  (.A(g7367), .B(g4507), .Z(g7611) ) ;
AND2    gate7278  (.A(g7488), .B(g3466), .Z(g7615) ) ;
AND2    gate7279  (.A(g7367), .B(g4517), .Z(g7616) ) ;
AND2    gate7280  (.A(g7463), .B(g3466), .Z(g7626) ) ;
AND2    gate7281  (.A(g7367), .B(g4532), .Z(g7628) ) ;
OR2     gate7282  (.A(g4192), .B(g7193), .Z(g7445) ) ;
AND2    gate7283  (.A(g7445), .B(g3548), .Z(g7632) ) ;
AND2    gate7284  (.A(g7367), .B(g4549), .Z(g7634) ) ;
AND2    gate7285  (.A(g7480), .B(g5754), .Z(g7653) ) ;
AND2    gate7286  (.A(g7367), .B(g4142), .Z(g7654) ) ;
AND2    gate7287  (.A(g7367), .B(g4150), .Z(g7658) ) ;
NAND2   gate7288  (.A(II13686), .B(II13687), .Z(g7503) ) ;
NAND2   gate7289  (.A(II13599), .B(II13600), .Z(g7447) ) ;
NAND2   gate7290  (.A(II13588), .B(II13589), .Z(g7444) ) ;
AND2    gate7291  (.A(g1061), .B(g7429), .Z(g7683) ) ;
OR2     gate7292  (.A(g7278), .B(g4546), .Z(g7337) ) ;
AND2    gate7293  (.A(g7337), .B(g5938), .Z(g7724) ) ;
OR2     gate7294  (.A(g7323), .B(g7142), .Z(g7575) ) ;
OR2     gate7295  (.A(g4690), .B(g2862), .Z(g5343) ) ;
OR2     gate7296  (.A(g5817), .B(g2934), .Z(g6470) ) ;
OR2     gate7297  (.A(g6044), .B(g7412), .Z(g7682) ) ;
NAND2   gate7298  (.A(II13786), .B(II13787), .Z(g7535) ) ;
AND2    gate7299  (.A(g7535), .B(g4841), .Z(g8060) ) ;
AND2    gate7300  (.A(g7476), .B(g7634), .Z(g8062) ) ;
AND2    gate7301  (.A(g7483), .B(g7634), .Z(g8064) ) ;
AND2    gate7302  (.A(g7488), .B(g7634), .Z(g8066) ) ;
OR2     gate7303  (.A(g6053), .B(g7416), .Z(g7687) ) ;
AND2    gate7304  (.A(g7456), .B(g7634), .Z(g8069) ) ;
AND2    gate7305  (.A(g863), .B(g7616), .Z(g8070) ) ;
NAND2   gate7306  (.A(II13801), .B(II13802), .Z(g7540) ) ;
AND2    gate7307  (.A(g7540), .B(g4969), .Z(g8071) ) ;
AND2    gate7308  (.A(g855), .B(g7616), .Z(g8074) ) ;
AND2    gate7309  (.A(g7460), .B(g7634), .Z(g8075) ) ;
OR2     gate7310  (.A(g4181), .B(g7417), .Z(g7690) ) ;
AND2    gate7311  (.A(g859), .B(g7616), .Z(g8077) ) ;
AND2    gate7312  (.A(g7463), .B(g7634), .Z(g8078) ) ;
AND2    gate7313  (.A(g831), .B(g7658), .Z(g8079) ) ;
AND2    gate7314  (.A(g7467), .B(g7634), .Z(g8080) ) ;
AND2    gate7315  (.A(g834), .B(g7658), .Z(g8081) ) ;
AND2    gate7316  (.A(g7471), .B(g7634), .Z(g8087) ) ;
AND2    gate7317  (.A(g837), .B(g7658), .Z(g8088) ) ;
AND2    gate7318  (.A(g840), .B(g7658), .Z(g8089) ) ;
AND2    gate7319  (.A(g843), .B(g7658), .Z(g8090) ) ;
AND2    gate7320  (.A(g1065), .B(g7683), .Z(g8147) ) ;
AND2    gate7321  (.A(g846), .B(g7658), .Z(g8150) ) ;
AND2    gate7322  (.A(g849), .B(g7658), .Z(g8151) ) ;
AND2    gate7323  (.A(g852), .B(g7658), .Z(g8153) ) ;
AND2    gate7324  (.A(g8180), .B(g5680), .Z(g8229) ) ;
AND2    gate7325  (.A(g89), .B(g8131), .Z(g8237) ) ;
AND2    gate7326  (.A(g100), .B(g8131), .Z(g8238) ) ;
AND2    gate7327  (.A(g95), .B(g8131), .Z(g8256) ) ;
AND2    gate7328  (.A(g146), .B(g8042), .Z(g8257) ) ;
AND2    gate7329  (.A(g142), .B(g8111), .Z(g8258) ) ;
AND2    gate7330  (.A(g4538), .B(g7855), .Z(g8259) ) ;
AND2    gate7331  (.A(g138), .B(g8111), .Z(g8260) ) ;
AND2    gate7332  (.A(g174), .B(g8042), .Z(g8261) ) ;
AND2    gate7333  (.A(g4554), .B(g7855), .Z(g8262) ) ;
AND2    gate7334  (.A(g4555), .B(g7905), .Z(g8263) ) ;
AND2    gate7335  (.A(g105), .B(g8131), .Z(g8264) ) ;
AND2    gate7336  (.A(g134), .B(g8111), .Z(g8265) ) ;
AND2    gate7337  (.A(g2157), .B(g8042), .Z(g8266) ) ;
AND2    gate7338  (.A(g154), .B(g8042), .Z(g8267) ) ;
AND2    gate7339  (.A(g4568), .B(g7905), .Z(g8268) ) ;
AND2    gate7340  (.A(g4569), .B(g7951), .Z(g8269) ) ;
AND2    gate7341  (.A(g110), .B(g8131), .Z(g8270) ) ;
AND2    gate7342  (.A(g130), .B(g8111), .Z(g8271) ) ;
AND2    gate7343  (.A(g158), .B(g8042), .Z(g8272) ) ;
AND2    gate7344  (.A(g185), .B(g8156), .Z(g8273) ) ;
AND2    gate7345  (.A(g4580), .B(g7951), .Z(g8274) ) ;
AND2    gate7346  (.A(g4581), .B(g7993), .Z(g8275) ) ;
AND2    gate7347  (.A(g150), .B(g8042), .Z(g8276) ) ;
AND2    gate7348  (.A(g162), .B(g8042), .Z(g8277) ) ;
AND2    gate7349  (.A(g4589), .B(g7993), .Z(g8278) ) ;
AND2    gate7350  (.A(g114), .B(g8111), .Z(g8280) ) ;
AND2    gate7351  (.A(g168), .B(g8042), .Z(g8281) ) ;
AND2    gate7352  (.A(g179), .B(g8156), .Z(g8282) ) ;
AND2    gate7353  (.A(g267), .B(g7838), .Z(g8283) ) ;
AND2    gate7354  (.A(g118), .B(g8111), .Z(g8285) ) ;
AND2    gate7355  (.A(g180), .B(g8156), .Z(g8286) ) ;
AND2    gate7356  (.A(g4500), .B(g7855), .Z(g8287) ) ;
AND2    gate7357  (.A(g270), .B(g7838), .Z(g8288) ) ;
AND2    gate7358  (.A(g348), .B(g7870), .Z(g8289) ) ;
AND2    gate7359  (.A(g588), .B(g8181), .Z(g8290) ) ;
AND2    gate7360  (.A(g122), .B(g8111), .Z(g8291) ) ;
AND2    gate7361  (.A(g181), .B(g8156), .Z(g8292) ) ;
AND2    gate7362  (.A(g4510), .B(g7855), .Z(g8293) ) ;
AND2    gate7363  (.A(g281), .B(g7838), .Z(g8294) ) ;
AND2    gate7364  (.A(g4512), .B(g7905), .Z(g8295) ) ;
AND2    gate7365  (.A(g351), .B(g7870), .Z(g8296) ) ;
AND2    gate7366  (.A(g429), .B(g7920), .Z(g8297) ) ;
AND2    gate7367  (.A(g553), .B(g8181), .Z(g8298) ) ;
AND2    gate7368  (.A(g591), .B(g8181), .Z(g8299) ) ;
AND2    gate7369  (.A(g126), .B(g8111), .Z(g8300) ) ;
AND2    gate7370  (.A(g182), .B(g8156), .Z(g8301) ) ;
AND2    gate7371  (.A(g4521), .B(g7855), .Z(g8302) ) ;
AND2    gate7372  (.A(g284), .B(g7838), .Z(g8303) ) ;
AND2    gate7373  (.A(g4523), .B(g7905), .Z(g8304) ) ;
AND2    gate7374  (.A(g362), .B(g7870), .Z(g8305) ) ;
AND2    gate7375  (.A(g4525), .B(g7951), .Z(g8306) ) ;
AND2    gate7376  (.A(g432), .B(g7920), .Z(g8307) ) ;
AND2    gate7377  (.A(g510), .B(g7966), .Z(g8308) ) ;
AND2    gate7378  (.A(g550), .B(g8181), .Z(g8309) ) ;
AND2    gate7379  (.A(g573), .B(g8181), .Z(g8310) ) ;
AND2    gate7380  (.A(g4540), .B(g7905), .Z(g8311) ) ;
AND2    gate7381  (.A(g365), .B(g7870), .Z(g8312) ) ;
AND2    gate7382  (.A(g4542), .B(g7951), .Z(g8313) ) ;
AND2    gate7383  (.A(g443), .B(g7920), .Z(g8314) ) ;
AND2    gate7384  (.A(g4544), .B(g7993), .Z(g8315) ) ;
AND2    gate7385  (.A(g513), .B(g7966), .Z(g8316) ) ;
AND2    gate7386  (.A(g547), .B(g8181), .Z(g8317) ) ;
AND2    gate7387  (.A(g183), .B(g8156), .Z(g8318) ) ;
AND2    gate7388  (.A(g255), .B(g7838), .Z(g8319) ) ;
AND2    gate7389  (.A(g4557), .B(g7951), .Z(g8320) ) ;
AND2    gate7390  (.A(g446), .B(g7920), .Z(g8321) ) ;
AND2    gate7391  (.A(g4559), .B(g7993), .Z(g8322) ) ;
AND2    gate7392  (.A(g524), .B(g7966), .Z(g8323) ) ;
AND2    gate7393  (.A(g184), .B(g8156), .Z(g8325) ) ;
AND2    gate7394  (.A(g258), .B(g7838), .Z(g8326) ) ;
AND2    gate7395  (.A(g336), .B(g7870), .Z(g8327) ) ;
AND2    gate7396  (.A(g4571), .B(g7993), .Z(g8328) ) ;
AND2    gate7397  (.A(g527), .B(g7966), .Z(g8329) ) ;
AND2    gate7398  (.A(g261), .B(g7838), .Z(g8330) ) ;
AND2    gate7399  (.A(g339), .B(g7870), .Z(g8331) ) ;
AND2    gate7400  (.A(g417), .B(g7920), .Z(g8332) ) ;
AND2    gate7401  (.A(g563), .B(g8181), .Z(g8333) ) ;
AND2    gate7402  (.A(g264), .B(g7838), .Z(g8334) ) ;
AND2    gate7403  (.A(g342), .B(g7870), .Z(g8335) ) ;
AND2    gate7404  (.A(g420), .B(g7920), .Z(g8336) ) ;
AND2    gate7405  (.A(g498), .B(g7966), .Z(g8337) ) ;
AND2    gate7406  (.A(g570), .B(g8181), .Z(g8338) ) ;
AND2    gate7407  (.A(g345), .B(g7870), .Z(g8339) ) ;
AND2    gate7408  (.A(g423), .B(g7920), .Z(g8340) ) ;
AND2    gate7409  (.A(g501), .B(g7966), .Z(g8341) ) ;
AND2    gate7410  (.A(g642), .B(g7793), .Z(g8359) ) ;
AND2    gate7411  (.A(g426), .B(g7920), .Z(g8361) ) ;
AND2    gate7412  (.A(g504), .B(g7966), .Z(g8362) ) ;
AND2    gate7413  (.A(g507), .B(g7966), .Z(g8377) ) ;
AND2    gate7414  (.A(g677), .B(g7887), .Z(g8378) ) ;
AND2    gate7415  (.A(g691), .B(g7793), .Z(g8379) ) ;
AND2    gate7416  (.A(g681), .B(g7887), .Z(g8380) ) ;
AND2    gate7417  (.A(g685), .B(g7887), .Z(g8382) ) ;
AND2    gate7418  (.A(g730), .B(g7937), .Z(g8383) ) ;
AND2    gate7419  (.A(g636), .B(g7793), .Z(g8384) ) ;
AND2    gate7420  (.A(g695), .B(g7811), .Z(g8385) ) ;
AND2    gate7421  (.A(g639), .B(g7793), .Z(g8403) ) ;
AND2    gate7422  (.A(g710), .B(g7937), .Z(g8404) ) ;
AND2    gate7423  (.A(g741), .B(g8018), .Z(g8405) ) ;
AND2    gate7424  (.A(g649), .B(g7793), .Z(g8438) ) ;
AND2    gate7425  (.A(g699), .B(g7811), .Z(g8439) ) ;
AND2    gate7426  (.A(g714), .B(g7937), .Z(g8440) ) ;
AND2    gate7427  (.A(g746), .B(g8018), .Z(g8441) ) ;
AND2    gate7428  (.A(g652), .B(g7793), .Z(g8455) ) ;
AND2    gate7429  (.A(g703), .B(g7811), .Z(g8456) ) ;
AND2    gate7430  (.A(g724), .B(g7811), .Z(g8457) ) ;
AND2    gate7431  (.A(g756), .B(g8199), .Z(g8458) ) ;
AND2    gate7432  (.A(g655), .B(g7793), .Z(g8459) ) ;
AND2    gate7433  (.A(g757), .B(g8199), .Z(g8460) ) ;
AND2    gate7434  (.A(g658), .B(g7793), .Z(g8461) ) ;
AND2    gate7435  (.A(g49), .B(g8199), .Z(g8462) ) ;
AND2    gate7436  (.A(g718), .B(g7937), .Z(g8513) ) ;
AND2    gate7437  (.A(g661), .B(g7887), .Z(g8542) ) ;
AND2    gate7438  (.A(g706), .B(g7887), .Z(g8543) ) ;
OR2     gate7439  (.A(g6045), .B(g7597), .Z(g8146) ) ;
OR2     gate7440  (.A(g6054), .B(g7607), .Z(g8154) ) ;
NAND2   gate7441  (.A(II14245), .B(II14246), .Z(g7828) ) ;
AND2    gate7442  (.A(g7828), .B(g4969), .Z(g8609) ) ;
AND2    gate7443  (.A(g665), .B(g7887), .Z(g8610) ) ;
AND2    gate7444  (.A(g669), .B(g7887), .Z(g8611) ) ;
AND2    gate7445  (.A(g673), .B(g7887), .Z(g8612) ) ;
AND2    gate7446  (.A(g751), .B(g8199), .Z(g8620) ) ;
AND2    gate7447  (.A(g734), .B(g7937), .Z(g8621) ) ;
AND2    gate7448  (.A(g738), .B(g7811), .Z(g8622) ) ;
AND2    gate7449  (.A(g755), .B(g8199), .Z(g8623) ) ;
AND2    gate7450  (.A(g754), .B(g8199), .Z(g8624) ) ;
AND2    gate7451  (.A(g752), .B(g8199), .Z(g8626) ) ;
AND2    gate7452  (.A(g753), .B(g8199), .Z(g8628) ) ;
AND2    gate7453  (.A(g547), .B(g8094), .Z(g8643) ) ;
AND2    gate7454  (.A(g550), .B(g8094), .Z(g8645) ) ;
AND2    gate7455  (.A(g553), .B(g8094), .Z(g8646) ) ;
AND2    gate7456  (.A(g588), .B(g8094), .Z(g8648) ) ;
AND2    gate7457  (.A(g591), .B(g8094), .Z(g8650) ) ;
AND2    gate7458  (.A(g563), .B(g8094), .Z(g8652) ) ;
AND2    gate7459  (.A(g573), .B(g8094), .Z(g8653) ) ;
AND2    gate7460  (.A(g570), .B(g8094), .Z(g8654) ) ;
AND2    gate7461  (.A(g1069), .B(g8147), .Z(g8660) ) ;
AND2    gate7462  (.A(g3819), .B(g8342), .Z(g8686) ) ;
AND2    gate7463  (.A(g3488), .B(g8363), .Z(g8687) ) ;
AND2    gate7464  (.A(g3812), .B(g8342), .Z(g8688) ) ;
AND2    gate7465  (.A(g3485), .B(g8363), .Z(g8690) ) ;
AND2    gate7466  (.A(g3805), .B(g8342), .Z(g8691) ) ;
AND2    gate7467  (.A(g3462), .B(g8363), .Z(g8692) ) ;
AND2    gate7468  (.A(g3798), .B(g8342), .Z(g8693) ) ;
AND2    gate7469  (.A(g2709), .B(g8363), .Z(g8695) ) ;
AND2    gate7470  (.A(g3743), .B(g8342), .Z(g8696) ) ;
AND2    gate7471  (.A(g3761), .B(g8342), .Z(g8697) ) ;
AND2    gate7472  (.A(g3774), .B(g8342), .Z(g8698) ) ;
AND2    gate7473  (.A(g3784), .B(g8342), .Z(g8700) ) ;
AND2    gate7474  (.A(g2700), .B(g8363), .Z(g8701) ) ;
AND2    gate7475  (.A(g2837), .B(g8386), .Z(g8702) ) ;
AND2    gate7476  (.A(g3574), .B(g8407), .Z(g8703) ) ;
AND2    gate7477  (.A(g2829), .B(g8386), .Z(g8704) ) ;
AND2    gate7478  (.A(g2798), .B(g8421), .Z(g8705) ) ;
AND2    gate7479  (.A(g3557), .B(g8407), .Z(g8708) ) ;
AND2    gate7480  (.A(g2818), .B(g8386), .Z(g8709) ) ;
AND2    gate7481  (.A(g2790), .B(g8421), .Z(g8710) ) ;
AND2    gate7482  (.A(g3542), .B(g8407), .Z(g8711) ) ;
AND2    gate7483  (.A(g2804), .B(g8386), .Z(g8712) ) ;
AND2    gate7484  (.A(g2777), .B(g8421), .Z(g8713) ) ;
AND2    gate7485  (.A(g2873), .B(g8407), .Z(g8714) ) ;
AND2    gate7486  (.A(g2761), .B(g8386), .Z(g8715) ) ;
AND2    gate7487  (.A(g3506), .B(g8443), .Z(g8716) ) ;
AND2    gate7488  (.A(g2764), .B(g8421), .Z(g8717) ) ;
AND2    gate7489  (.A(g2774), .B(g8386), .Z(g8718) ) ;
AND2    gate7490  (.A(g2821), .B(g8443), .Z(g8719) ) ;
AND2    gate7491  (.A(g3825), .B(g8421), .Z(g8720) ) ;
AND2    gate7492  (.A(g2703), .B(g8464), .Z(g8721) ) ;
AND2    gate7493  (.A(g2787), .B(g8386), .Z(g8722) ) ;
AND2    gate7494  (.A(g2706), .B(g8421), .Z(g8723) ) ;
AND2    gate7495  (.A(g3822), .B(g8464), .Z(g8724) ) ;
AND2    gate7496  (.A(g3008), .B(g8493), .Z(g8725) ) ;
AND2    gate7497  (.A(g2795), .B(g8386), .Z(g8726) ) ;
AND2    gate7498  (.A(g2724), .B(g8421), .Z(g8727) ) ;
AND2    gate7499  (.A(g3815), .B(g8464), .Z(g8728) ) ;
AND2    gate7500  (.A(g2999), .B(g8493), .Z(g8729) ) ;
AND2    gate7501  (.A(g2863), .B(g8407), .Z(g8730) ) ;
AND2    gate7502  (.A(g2743), .B(g8421), .Z(g8731) ) ;
AND2    gate7503  (.A(g3808), .B(g8464), .Z(g8732) ) ;
AND2    gate7504  (.A(g2996), .B(g8493), .Z(g8733) ) ;
AND2    gate7505  (.A(g2807), .B(g8443), .Z(g8735) ) ;
AND2    gate7506  (.A(g3771), .B(g8464), .Z(g8736) ) ;
AND2    gate7507  (.A(g2992), .B(g8493), .Z(g8737) ) ;
AND2    gate7508  (.A(g3780), .B(g8464), .Z(g8739) ) ;
AND2    gate7509  (.A(g2966), .B(g8493), .Z(g8740) ) ;
AND2    gate7510  (.A(g3787), .B(g8464), .Z(g8741) ) ;
AND2    gate7511  (.A(g2973), .B(g8493), .Z(g8742) ) ;
AND2    gate7512  (.A(g3802), .B(g8464), .Z(g8744) ) ;
AND2    gate7513  (.A(g2982), .B(g8493), .Z(g8745) ) ;
AND2    gate7514  (.A(g2721), .B(g8483), .Z(g8748) ) ;
AND2    gate7515  (.A(g2989), .B(g8493), .Z(g8749) ) ;
NAND2   gate7516  (.A(II14473), .B(II14474), .Z(g8231) ) ;
AND2    gate7517  (.A(g8231), .B(g4969), .Z(g8764) ) ;
OR2     gate7518  (.A(g6047), .B(g8060), .Z(g8634) ) ;
OR2     gate7519  (.A(g6057), .B(g8071), .Z(g8637) ) ;
AND2    gate7520  (.A(g255), .B(g8524), .Z(g8813) ) ;
AND2    gate7521  (.A(g3880), .B(g8463), .Z(g8814) ) ;
AND2    gate7522  (.A(g258), .B(g8524), .Z(g8815) ) ;
AND2    gate7523  (.A(g336), .B(g8545), .Z(g8816) ) ;
AND2    gate7524  (.A(g4545), .B(g8482), .Z(g8817) ) ;
AND2    gate7525  (.A(g261), .B(g8524), .Z(g8820) ) ;
AND2    gate7526  (.A(g339), .B(g8545), .Z(g8821) ) ;
AND2    gate7527  (.A(g417), .B(g8564), .Z(g8822) ) ;
AND2    gate7528  (.A(g4561), .B(g8512), .Z(g8823) ) ;
AND2    gate7529  (.A(g264), .B(g8524), .Z(g8824) ) ;
AND2    gate7530  (.A(g342), .B(g8545), .Z(g8825) ) ;
AND2    gate7531  (.A(g420), .B(g8564), .Z(g8826) ) ;
AND2    gate7532  (.A(g498), .B(g8585), .Z(g8827) ) ;
AND2    gate7533  (.A(g4573), .B(g8541), .Z(g8828) ) ;
AND2    gate7534  (.A(g267), .B(g8524), .Z(g8829) ) ;
AND2    gate7535  (.A(g345), .B(g8545), .Z(g8830) ) ;
AND2    gate7536  (.A(g423), .B(g8564), .Z(g8831) ) ;
AND2    gate7537  (.A(g501), .B(g8585), .Z(g8832) ) ;
AND2    gate7538  (.A(g4583), .B(g8562), .Z(g8833) ) ;
AND2    gate7539  (.A(g270), .B(g8524), .Z(g8835) ) ;
AND2    gate7540  (.A(g348), .B(g8545), .Z(g8836) ) ;
AND2    gate7541  (.A(g426), .B(g8564), .Z(g8837) ) ;
AND2    gate7542  (.A(g504), .B(g8585), .Z(g8838) ) ;
AND2    gate7543  (.A(g4050), .B(g8581), .Z(g8839) ) ;
AND2    gate7544  (.A(g4590), .B(g8582), .Z(g8840) ) ;
AND2    gate7545  (.A(g351), .B(g8545), .Z(g8841) ) ;
AND2    gate7546  (.A(g429), .B(g8564), .Z(g8842) ) ;
AND2    gate7547  (.A(g507), .B(g8585), .Z(g8843) ) ;
AND2    gate7548  (.A(g4056), .B(g8602), .Z(g8844) ) ;
AND2    gate7549  (.A(g432), .B(g8564), .Z(g8845) ) ;
AND2    gate7550  (.A(g510), .B(g8585), .Z(g8846) ) ;
AND2    gate7551  (.A(g281), .B(g8524), .Z(g8848) ) ;
AND2    gate7552  (.A(g513), .B(g8585), .Z(g8849) ) ;
AND2    gate7553  (.A(g284), .B(g8524), .Z(g8851) ) ;
AND2    gate7554  (.A(g362), .B(g8545), .Z(g8852) ) ;
AND2    gate7555  (.A(g365), .B(g8545), .Z(g8853) ) ;
AND2    gate7556  (.A(g443), .B(g8564), .Z(g8854) ) ;
AND2    gate7557  (.A(g446), .B(g8564), .Z(g8857) ) ;
AND2    gate7558  (.A(g524), .B(g8585), .Z(g8858) ) ;
AND2    gate7559  (.A(g527), .B(g8585), .Z(g8860) ) ;
OR2     gate7560  (.A(II14951), .B(II14952), .Z(g8769) ) ;
AND2    gate7561  (.A(g8769), .B(g6102), .Z(g8876) ) ;
OR2     gate7562  (.A(II14959), .B(II14960), .Z(g8773) ) ;
AND2    gate7563  (.A(g8773), .B(g6104), .Z(g8877) ) ;
OR2     gate7564  (.A(II14969), .B(II14970), .Z(g8777) ) ;
AND2    gate7565  (.A(g8777), .B(g6106), .Z(g8878) ) ;
OR3     gate7566  (.A(g8624), .B(g8659), .C(II14980), .Z(g8782) ) ;
AND2    gate7567  (.A(g8782), .B(g6108), .Z(g8879) ) ;
NAND2   gate7568  (.A(II14838), .B(II14839), .Z(g8681) ) ;
AND2    gate7569  (.A(g8681), .B(g4969), .Z(g8892) ) ;
OR2     gate7570  (.A(g6060), .B(g8609), .Z(g8804) ) ;
NAND2   gate7571  (.A(g6984), .B(g8644), .Z(g8798) ) ;
OR4     gate7572  (.A(g8150), .B(g8078), .C(g8070), .D(g8360), .Z(g8796) ) ;
NAND2   gate7573  (.A(g8073), .B(g8092), .Z(g8239) ) ;
AND2    gate7574  (.A(g8796), .B(g8239), .Z(g8912) ) ;
OR4     gate7575  (.A(g8151), .B(g8077), .C(g8075), .D(g8279), .Z(g8795) ) ;
AND2    gate7576  (.A(g8795), .B(g8239), .Z(g8914) ) ;
OR4     gate7577  (.A(g8153), .B(g8074), .C(g8069), .D(g8523), .Z(g8794) ) ;
AND2    gate7578  (.A(g8794), .B(g8239), .Z(g8915) ) ;
AND2    gate7579  (.A(g4567), .B(g8743), .Z(g8919) ) ;
AND2    gate7580  (.A(g4578), .B(g8746), .Z(g8920) ) ;
AND2    gate7581  (.A(g4579), .B(g8747), .Z(g8921) ) ;
AND2    gate7582  (.A(g4586), .B(g8750), .Z(g8922) ) ;
AND2    gate7583  (.A(g4587), .B(g8751), .Z(g8923) ) ;
AND2    gate7584  (.A(g4588), .B(g8752), .Z(g8924) ) ;
AND2    gate7585  (.A(g4592), .B(g8754), .Z(g8925) ) ;
AND2    gate7586  (.A(g4593), .B(g8755), .Z(g8926) ) ;
AND2    gate7587  (.A(g4594), .B(g8756), .Z(g8927) ) ;
AND2    gate7588  (.A(g4595), .B(g8757), .Z(g8928) ) ;
AND2    gate7589  (.A(g3865), .B(g8759), .Z(g8929) ) ;
AND2    gate7590  (.A(g3866), .B(g8760), .Z(g8930) ) ;
AND2    gate7591  (.A(g3867), .B(g8761), .Z(g8931) ) ;
AND2    gate7592  (.A(g3868), .B(g8762), .Z(g8932) ) ;
AND2    gate7593  (.A(g4511), .B(g8765), .Z(g8933) ) ;
AND2    gate7594  (.A(g3873), .B(g8766), .Z(g8934) ) ;
AND2    gate7595  (.A(g3874), .B(g8767), .Z(g8935) ) ;
AND2    gate7596  (.A(g3875), .B(g8768), .Z(g8936) ) ;
AND2    gate7597  (.A(g4524), .B(g8770), .Z(g8937) ) ;
AND2    gate7598  (.A(g3878), .B(g8771), .Z(g8938) ) ;
AND2    gate7599  (.A(g3879), .B(g8772), .Z(g8939) ) ;
AND2    gate7600  (.A(g4543), .B(g8775), .Z(g8940) ) ;
AND2    gate7601  (.A(g3882), .B(g8776), .Z(g8941) ) ;
AND2    gate7602  (.A(g4522), .B(g8780), .Z(g8942) ) ;
AND2    gate7603  (.A(g4560), .B(g8781), .Z(g8943) ) ;
AND2    gate7604  (.A(g4539), .B(g8783), .Z(g8944) ) ;
AND2    gate7605  (.A(g4541), .B(g8784), .Z(g8945) ) ;
AND2    gate7606  (.A(g4556), .B(g8786), .Z(g8946) ) ;
AND2    gate7607  (.A(g4558), .B(g8787), .Z(g8947) ) ;
AND2    gate7608  (.A(g4570), .B(g8789), .Z(g8948) ) ;
AND2    gate7609  (.A(g4572), .B(g8790), .Z(g8949) ) ;
AND2    gate7610  (.A(g4582), .B(g8791), .Z(g8950) ) ;
OR3     gate7611  (.A(g8623), .B(g8656), .C(II14985), .Z(g8785) ) ;
AND2    gate7612  (.A(g8785), .B(g6072), .Z(g8951) ) ;
OR3     gate7613  (.A(g8620), .B(g8658), .C(II14990), .Z(g8788) ) ;
AND2    gate7614  (.A(g8788), .B(g6075), .Z(g8952) ) ;
OR3     gate7615  (.A(g8655), .B(II14932), .C(II14933), .Z(g8758) ) ;
AND2    gate7616  (.A(g8758), .B(g6093), .Z(g8953) ) ;
OR3     gate7617  (.A(g8232), .B(II14941), .C(II14942), .Z(g8763) ) ;
AND2    gate7618  (.A(g8763), .B(g6097), .Z(g8954) ) ;
OR3     gate7619  (.A(g8723), .B(g8806), .C(II15243), .Z(g8885) ) ;
AND2    gate7620  (.A(g8885), .B(g5317), .Z(g8961) ) ;
OR3     gate7621  (.A(II15290), .B(II15291), .C(II15292), .Z(g8890) ) ;
AND2    gate7622  (.A(g8890), .B(g5317), .Z(g8962) ) ;
OR4     gate7623  (.A(g8705), .B(g8811), .C(II15297), .D(II15298), .Z(g8891) ) ;
AND2    gate7624  (.A(g8891), .B(g5317), .Z(g8963) ) ;
OR2     gate7625  (.A(g6043), .B(g8764), .Z(g8909) ) ;
OR3     gate7626  (.A(g8079), .B(g8066), .C(g8855), .Z(g8908) ) ;
AND2    gate7627  (.A(g8908), .B(g8239), .Z(g9012) ) ;
OR3     gate7628  (.A(g8081), .B(g8064), .C(g8707), .Z(g8907) ) ;
AND2    gate7629  (.A(g8907), .B(g8239), .Z(g9013) ) ;
OR3     gate7630  (.A(g8088), .B(g8062), .C(g8699), .Z(g8906) ) ;
AND2    gate7631  (.A(g8906), .B(g8239), .Z(g9014) ) ;
OR3     gate7632  (.A(g8089), .B(g8087), .C(g8694), .Z(g8905) ) ;
AND2    gate7633  (.A(g8905), .B(g8239), .Z(g9015) ) ;
OR3     gate7634  (.A(g8090), .B(g8080), .C(g8706), .Z(g8904) ) ;
AND2    gate7635  (.A(g8904), .B(g8239), .Z(g9016) ) ;
OR3     gate7636  (.A(g8727), .B(g8812), .C(II15254), .Z(g8886) ) ;
AND2    gate7637  (.A(g8886), .B(g5317), .Z(g9021) ) ;
OR2     gate7638  (.A(II15265), .B(g8819), .Z(g8887) ) ;
AND2    gate7639  (.A(g8887), .B(g5317), .Z(g9022) ) ;
OR2     gate7640  (.A(II15276), .B(g8807), .Z(g8888) ) ;
AND2    gate7641  (.A(g8888), .B(g5317), .Z(g9023) ) ;
OR3     gate7642  (.A(g8735), .B(g8818), .C(II15232), .Z(g8884) ) ;
AND2    gate7643  (.A(g8884), .B(g5317), .Z(g9024) ) ;
OR3     gate7644  (.A(II15283), .B(II15284), .C(II15285), .Z(g8889) ) ;
AND2    gate7645  (.A(g8889), .B(g5317), .Z(g9025) ) ;
OR4     gate7646  (.A(g8739), .B(g8742), .C(g8914), .D(g8847), .Z(g8965) ) ;
AND2    gate7647  (.A(g8965), .B(g5345), .Z(g9037) ) ;
OR4     gate7648  (.A(g8741), .B(g8745), .C(g8912), .D(g8850), .Z(g8966) ) ;
AND2    gate7649  (.A(g8966), .B(g5345), .Z(g9038) ) ;
OR2     gate7650  (.A(g6046), .B(g8892), .Z(g9011) ) ;
OR3     gate7651  (.A(g8915), .B(g8863), .C(II15400), .Z(g8964) ) ;
AND2    gate7652  (.A(g8964), .B(g5345), .Z(g9084) ) ;
OR4     gate7653  (.A(g8744), .B(g8749), .C(g9016), .D(g8862), .Z(g9046) ) ;
AND2    gate7654  (.A(g9046), .B(g5345), .Z(g9118) ) ;
OR4     gate7655  (.A(g8732), .B(g8737), .C(g9015), .D(g8861), .Z(g9049) ) ;
AND2    gate7656  (.A(g9049), .B(g5345), .Z(g9119) ) ;
OR4     gate7657  (.A(g8728), .B(g8733), .C(g9014), .D(g8679), .Z(g9052) ) ;
AND2    gate7658  (.A(g9052), .B(g5345), .Z(g9120) ) ;
OR4     gate7659  (.A(g8724), .B(g8729), .C(g9013), .D(g8680), .Z(g9054) ) ;
AND2    gate7660  (.A(g9054), .B(g5345), .Z(g9130) ) ;
OR4     gate7661  (.A(g8721), .B(g8725), .C(g9012), .D(g8859), .Z(g9055) ) ;
AND2    gate7662  (.A(g9055), .B(g5345), .Z(g9131) ) ;
OR2     gate7663  (.A(g8876), .B(g9038), .Z(g9124) ) ;
AND2    gate7664  (.A(g9124), .B(g6059), .Z(g9142) ) ;
OR2     gate7665  (.A(g8953), .B(g9084), .Z(g9122) ) ;
AND2    gate7666  (.A(g9122), .B(g6089), .Z(g9143) ) ;
OR2     gate7667  (.A(g8954), .B(g9037), .Z(g9123) ) ;
AND2    gate7668  (.A(g9123), .B(g6096), .Z(g9144) ) ;
OR2     gate7669  (.A(g8951), .B(g9130), .Z(g9135) ) ;
AND2    gate7670  (.A(g9135), .B(g6101), .Z(g9146) ) ;
OR2     gate7671  (.A(g8952), .B(g9131), .Z(g9136) ) ;
AND2    gate7672  (.A(g9136), .B(g6103), .Z(g9147) ) ;
OR2     gate7673  (.A(g8877), .B(g9118), .Z(g9137) ) ;
AND2    gate7674  (.A(g9137), .B(g6070), .Z(g9158) ) ;
OR2     gate7675  (.A(g8878), .B(g9119), .Z(g9138) ) ;
AND2    gate7676  (.A(g9138), .B(g6074), .Z(g9159) ) ;
OR2     gate7677  (.A(g8879), .B(g9120), .Z(g9139) ) ;
AND2    gate7678  (.A(g9139), .B(g6092), .Z(g9160) ) ;
AND2    gate7679  (.A(g9220), .B(g5403), .Z(g9226) ) ;
AND2    gate7680  (.A(g4748), .B(g9223), .Z(g9238) ) ;
AND2    gate7681  (.A(g9223), .B(g5261), .Z(g9240) ) ;
AND2    gate7682  (.A(g4748), .B(g9227), .Z(g9247) ) ;
AND2    gate7683  (.A(g4748), .B(g9230), .Z(g9251) ) ;
AND2    gate7684  (.A(g9227), .B(g5628), .Z(g9258) ) ;
AND2    gate7685  (.A(g9230), .B(g5639), .Z(g9259) ) ;
AND2    gate7686  (.A(g4748), .B(g9241), .Z(g9270) ) ;
AND2    gate7687  (.A(g4748), .B(g9244), .Z(g9271) ) ;
AND2    gate7688  (.A(g4748), .B(g9248), .Z(g9272) ) ;
AND2    gate7689  (.A(g4748), .B(g9252), .Z(g9273) ) ;
AND2    gate7690  (.A(g4748), .B(g9255), .Z(g9274) ) ;
AND2    gate7691  (.A(g9241), .B(g5645), .Z(g9275) ) ;
AND2    gate7692  (.A(g9244), .B(g5649), .Z(g9276) ) ;
AND2    gate7693  (.A(g9248), .B(g5654), .Z(g9277) ) ;
AND2    gate7694  (.A(g9252), .B(g5658), .Z(g9278) ) ;
AND2    gate7695  (.A(g9255), .B(g5665), .Z(g9279) ) ;
AND2    gate7696  (.A(g9316), .B(g5757), .Z(g9327) ) ;
NOR4    gate7697  (.A(g5403), .B(g5802), .C(g5769), .D(g5790), .Z(g6465) ) ;
AND2    gate7698  (.A(g9324), .B(g6465), .Z(g9328) ) ;
AND2    gate7699  (.A(g9318), .B(g6205), .Z(g9334) ) ;
AND2    gate7700  (.A(g9320), .B(g6206), .Z(g9335) ) ;
AND2    gate7701  (.A(g9328), .B(g1738), .Z(g9343) ) ;
AND2    gate7702  (.A(g9329), .B(g6211), .Z(g9344) ) ;
AND2    gate7703  (.A(g9330), .B(g6217), .Z(g9345) ) ;
AND2    gate7704  (.A(g9331), .B(g6222), .Z(g9346) ) ;
AND2    gate7705  (.A(g9332), .B(g6226), .Z(g9347) ) ;
AND2    gate7706  (.A(g9333), .B(g6229), .Z(g9348) ) ;
AND2    gate7707  (.A(g9340), .B(g5690), .Z(g9349) ) ;
AND2    gate7708  (.A(g4748), .B(g9340), .Z(g9359) ) ;
OR2     gate7709  (.A(g9343), .B(g4526), .Z(g9352) ) ;
AND2    gate7710  (.A(g9352), .B(g5917), .Z(g9371) ) ;
AND2    gate7711  (.A(g9383), .B(g6245), .Z(g9384) ) ;
OR4     gate7712  (.A(g969), .B(g970), .C(g966), .D(g963), .Z(II5757) ) ;
OR2     gate7713  (.A(g1263), .B(g1257), .Z(g2043) ) ;
OR4     gate7714  (.A(g1363), .B(g1364), .C(g1365), .D(g1366), .Z(g2206) ) ;
OR4     gate7715  (.A(g1367), .B(g1368), .C(g1369), .D(g1370), .Z(g2213) ) ;
OR4     gate7716  (.A(g1376), .B(g1377), .C(g1378), .D(g1379), .Z(g2214) ) ;
OR4     gate7717  (.A(g1371), .B(g1372), .C(g1373), .D(g1374), .Z(g2229) ) ;
OR4     gate7718  (.A(g1380), .B(g1381), .C(g1382), .D(g1383), .Z(g2230) ) ;
OR4     gate7719  (.A(g1384), .B(g1385), .C(g1386), .D(g1387), .Z(g2262) ) ;
OR4     gate7720  (.A(g891), .B(g896), .C(g901), .D(g906), .Z(II6208) ) ;
OR4     gate7721  (.A(g911), .B(g916), .C(g921), .D(g883), .Z(II6209) ) ;
OR2     gate7722  (.A(II6208), .B(II6209), .Z(g2368) ) ;
NOR2    gate7723  (.A(g1421), .B(g1416), .Z(g2014) ) ;
OR2     gate7724  (.A(g1663), .B(g1421), .Z(g3541) ) ;
NAND2   gate7725  (.A(II6202), .B(II6203), .Z(g2367) ) ;
NAND2   gate7726  (.A(II6171), .B(II6172), .Z(g2352) ) ;
NAND2   gate7727  (.A(II6233), .B(II6234), .Z(g2378) ) ;
NAND2   gate7728  (.A(II6134), .B(II6135), .Z(g2330) ) ;
OR4     gate7729  (.A(g2367), .B(g2352), .C(g2378), .D(g2330), .Z(II7232) ) ;
NAND2   gate7730  (.A(II6103), .B(II6104), .Z(g2315) ) ;
NAND2   gate7731  (.A(II6258), .B(II6259), .Z(g2385) ) ;
NAND2   gate7732  (.A(II6065), .B(II6066), .Z(g2294) ) ;
NAND2   gate7733  (.A(II6274), .B(II6275), .Z(g2395) ) ;
OR4     gate7734  (.A(g2315), .B(g2385), .C(g2294), .D(g2395), .Z(II7233) ) ;
NAND2   gate7735  (.A(II6843), .B(II6844), .Z(g3129) ) ;
NAND2   gate7736  (.A(II6758), .B(II6759), .Z(g3012) ) ;
NAND2   gate7737  (.A(II6740), .B(II6741), .Z(g2995) ) ;
NAND2   gate7738  (.A(II6814), .B(II6815), .Z(g3083) ) ;
NAND2   gate7739  (.A(II6924), .B(II6925), .Z(g3315) ) ;
OR4     gate7740  (.A(g3019), .B(g3029), .C(g3038), .D(g3052), .Z(II8224) ) ;
OR4     gate7741  (.A(g3062), .B(g2712), .C(g2734), .D(g2752), .Z(II8225) ) ;
NAND2   gate7742  (.A(II7069), .B(II7070), .Z(g3602) ) ;
OR3     gate7743  (.A(g2655), .B(g1163), .C(g1160), .Z(II8363) ) ;
OR3     gate7744  (.A(g4504), .B(g4494), .C(g4430), .Z(II9029) ) ;
OR4     gate7745  (.A(g4417), .B(g4172), .C(g4163), .D(II9029), .Z(g4727) ) ;
OR3     gate7746  (.A(g4507), .B(g4497), .C(g4486), .Z(II9038) ) ;
OR3     gate7747  (.A(g4469), .B(g4448), .C(II9038), .Z(g4734) ) ;
OR3     gate7748  (.A(g4483), .B(g4466), .C(g4445), .Z(II9041) ) ;
OR4     gate7749  (.A(g4427), .B(g4414), .C(g4403), .D(II9041), .Z(g4735) ) ;
OR3     gate7750  (.A(g4150), .B(g4142), .C(g4549), .Z(II9044) ) ;
OR3     gate7751  (.A(g4532), .B(g4517), .C(II9044), .Z(g4736) ) ;
OR3     gate7752  (.A(g4155), .B(g4147), .C(g4139), .Z(II9047) ) ;
OR4     gate7753  (.A(g4135), .B(g4529), .C(g4514), .D(II9047), .Z(g4737) ) ;
OR3     gate7754  (.A(g4127), .B(g4123), .C(g4117), .Z(II9099) ) ;
OR4     gate7755  (.A(g4107), .B(g4097), .C(g4124), .D(II9099), .Z(g4786) ) ;
OR4     gate7756  (.A(g4133), .B(g4145), .C(g4138), .D(g4132), .Z(II9107) ) ;
OR4     gate7757  (.A(g4185), .B(g4131), .C(g4129), .D(II9107), .Z(g4790) ) ;
NAND2   gate7758  (.A(II8151), .B(II8152), .Z(g4237) ) ;
NOR2    gate7759  (.A(g3681), .B(g1590), .Z(g4318) ) ;
OR2     gate7760  (.A(g943), .B(g4501), .Z(g5021) ) ;
NAND2   gate7761  (.A(II7486), .B(II7487), .Z(g3900) ) ;
NAND2   gate7762  (.A(II7467), .B(II7468), .Z(g3895) ) ;
NAND2   gate7763  (.A(II7444), .B(II7445), .Z(g3890) ) ;
NAND2   gate7764  (.A(II8339), .B(II8340), .Z(g4363) ) ;
OR4     gate7765  (.A(g3900), .B(g3895), .C(g3890), .D(g4363), .Z(g5040) ) ;
NAND2   gate7766  (.A(II7617), .B(II7618), .Z(g3939) ) ;
NAND2   gate7767  (.A(II7575), .B(II7576), .Z(g3925) ) ;
NAND2   gate7768  (.A(II7539), .B(II7540), .Z(g3915) ) ;
NAND2   gate7769  (.A(II7511), .B(II7512), .Z(g3907) ) ;
OR4     gate7770  (.A(g3939), .B(g3925), .C(g3915), .D(g3907), .Z(g5057) ) ;
NAND2   gate7771  (.A(II9195), .B(II9196), .Z(g4835) ) ;
NAND2   gate7772  (.A(II9182), .B(II9183), .Z(g4824) ) ;
NAND2   gate7773  (.A(II9152), .B(II9153), .Z(g4810) ) ;
NAND2   gate7774  (.A(II10000), .B(II10001), .Z(g5558) ) ;
NAND2   gate7775  (.A(II9964), .B(II9965), .Z(g5546) ) ;
NAND2   gate7776  (.A(II9979), .B(II9980), .Z(g5555) ) ;
NAND2   gate7777  (.A(II9986), .B(II9987), .Z(g5556) ) ;
OR3     gate7778  (.A(g1000), .B(g5335), .C(g1909), .Z(g6270) ) ;
NOR2    gate7779  (.A(g2332), .B(g5305), .Z(g6209) ) ;
NOR2    gate7780  (.A(g875), .B(g5291), .Z(g6184) ) ;
NOR2    gate7781  (.A(g3002), .B(g5312), .Z(g6259) ) ;
NOR2    gate7782  (.A(g1855), .B(g5305), .Z(g6174) ) ;
NOR2    gate7783  (.A(g878), .B(g5284), .Z(g6214) ) ;
NOR2    gate7784  (.A(g1926), .B(g5310), .Z(g6193) ) ;
NOR4    gate7785  (.A(g875), .B(g866), .C(g1590), .D(g5291), .Z(g6197) ) ;
OR3     gate7786  (.A(g6193), .B(g6197), .C(g6175), .Z(II11603) ) ;
NOR2    gate7787  (.A(g5305), .B(g1590), .Z(g6185) ) ;
NAND2   gate7788  (.A(II10744), .B(II10745), .Z(g6119) ) ;
NAND2   gate7789  (.A(II10819), .B(II10820), .Z(g6153) ) ;
OR2     gate7790  (.A(g55), .B(g6264), .Z(g6710) ) ;
OR2     gate7791  (.A(g4048), .B(g6456), .Z(g7062) ) ;
OR3     gate7792  (.A(g5448), .B(g6267), .C(g6710), .Z(g7083) ) ;
OR2     gate7793  (.A(g7071), .B(g6980), .Z(g7191) ) ;
OR3     gate7794  (.A(g58), .B(g6258), .C(g5418), .Z(II13220) ) ;
OR2     gate7795  (.A(g6745), .B(g7202), .Z(g7421) ) ;
OR3     gate7796  (.A(g1166), .B(g1167), .C(g1170), .Z(II13553) ) ;
OR3     gate7797  (.A(g979), .B(g7566), .C(g1865), .Z(II14219) ) ;
OR4     gate7798  (.A(g7406), .B(g6664), .C(g3492), .D(II14219), .Z(g7784) ) ;
OR3     gate7799  (.A(g6664), .B(g3492), .C(g979), .Z(II14302) ) ;
OR4     gate7800  (.A(g3591), .B(g7406), .C(g7566), .D(II14302), .Z(g8009) ) ;
OR3     gate7801  (.A(g7654), .B(g7628), .C(g7611), .Z(g8082) ) ;
OR3     gate7802  (.A(g7566), .B(g1030), .C(g6664), .Z(II14366) ) ;
NOR2    gate7803  (.A(g6270), .B(g2245), .Z(g6452) ) ;
OR3     gate7804  (.A(g7215), .B(g6452), .C(II14366), .Z(g8091) ) ;
NOR4    gate7805  (.A(g1011), .B(g1837), .C(g6559), .D(g1008), .Z(g6910) ) ;
OR3     gate7806  (.A(g7566), .B(g6910), .C(g6452), .Z(g8128) ) ;
OR4     gate7807  (.A(g7566), .B(g1030), .C(g6664), .D(g6452), .Z(g8176) ) ;
OR4     gate7808  (.A(g7993), .B(g7966), .C(g7793), .D(g7811), .Z(II14467) ) ;
OR4     gate7809  (.A(g7937), .B(g7887), .C(g8029), .D(g8018), .Z(II14468) ) ;
OR4     gate7810  (.A(g7993), .B(g7966), .C(g7793), .D(g7811), .Z(II14479) ) ;
OR4     gate7811  (.A(g7937), .B(g7887), .C(g8029), .D(g8018), .Z(II14480) ) ;
OR4     gate7812  (.A(g7993), .B(g7966), .C(g7793), .D(g7811), .Z(II14484) ) ;
OR4     gate7813  (.A(g7937), .B(g7887), .C(g8029), .D(g8018), .Z(II14485) ) ;
OR4     gate7814  (.A(g7993), .B(g7966), .C(g7793), .D(g7811), .Z(II14495) ) ;
OR4     gate7815  (.A(g7937), .B(g7887), .C(g8029), .D(g8018), .Z(II14496) ) ;
OR2     gate7816  (.A(g8082), .B(g7616), .Z(g8613) ) ;
OR4     gate7817  (.A(g7993), .B(g7966), .C(g7793), .D(g7811), .Z(II14753) ) ;
OR4     gate7818  (.A(g7937), .B(g7887), .C(g8029), .D(g8018), .Z(II14754) ) ;
OR4     gate7819  (.A(g7993), .B(g7966), .C(g7793), .D(g7811), .Z(II14758) ) ;
OR4     gate7820  (.A(g7937), .B(g7887), .C(g8029), .D(g8018), .Z(II14759) ) ;
OR4     gate7821  (.A(g7993), .B(g7966), .C(g7793), .D(g7811), .Z(II14766) ) ;
OR4     gate7822  (.A(g7937), .B(g7887), .C(g8029), .D(g8018), .Z(II14767) ) ;
OR4     gate7823  (.A(g7993), .B(g7966), .C(g7793), .D(g7811), .Z(II14771) ) ;
OR4     gate7824  (.A(g7937), .B(g7887), .C(g8029), .D(g8018), .Z(II14772) ) ;
OR3     gate7825  (.A(g8483), .B(g8464), .C(g8514), .Z(II14831) ) ;
OR3     gate7826  (.A(g8483), .B(g8464), .C(g8514), .Z(II14834) ) ;
OR4     gate7827  (.A(g8278), .B(g8329), .C(g8461), .D(g8382), .Z(II14932) ) ;
OR4     gate7828  (.A(g8385), .B(g8404), .C(g8441), .D(g8462), .Z(II14933) ) ;
NOR3    gate7829  (.A(g8199), .B(II14753), .C(II14754), .Z(g8655) ) ;
OR4     gate7830  (.A(g8275), .B(g8323), .C(g8459), .D(g8380), .Z(II14941) ) ;
OR4     gate7831  (.A(g8439), .B(g8440), .C(g8405), .D(g8460), .Z(II14942) ) ;
NOR3    gate7832  (.A(g8199), .B(II14479), .C(II14480), .Z(g8232) ) ;
OR4     gate7833  (.A(g8328), .B(g8316), .C(g8455), .D(g8378), .Z(II14951) ) ;
NOR3    gate7834  (.A(g8199), .B(II14495), .C(II14496), .Z(g8236) ) ;
OR4     gate7835  (.A(g8456), .B(g8513), .C(g8458), .D(g8236), .Z(II14952) ) ;
OR4     gate7836  (.A(g8322), .B(g8308), .C(g8438), .D(g8612), .Z(II14959) ) ;
NOR3    gate7837  (.A(g8199), .B(II14467), .C(II14468), .Z(g8230) ) ;
OR4     gate7838  (.A(g8621), .B(g8622), .C(g8628), .D(g8230), .Z(II14960) ) ;
OR4     gate7839  (.A(g8315), .B(g8377), .C(g8359), .D(g8611), .Z(II14969) ) ;
NOR3    gate7840  (.A(g8199), .B(II14484), .C(II14485), .Z(g8233) ) ;
OR4     gate7841  (.A(g8457), .B(g8383), .C(g8626), .D(g8233), .Z(II14970) ) ;
OR3     gate7842  (.A(g8362), .B(g8403), .C(g8610), .Z(II14980) ) ;
NOR3    gate7843  (.A(g8199), .B(II14771), .C(II14772), .Z(g8659) ) ;
OR3     gate7844  (.A(g8341), .B(g8384), .C(g8542), .Z(II14985) ) ;
NOR3    gate7845  (.A(g8199), .B(II14758), .C(II14759), .Z(g8656) ) ;
OR3     gate7846  (.A(g8337), .B(g8379), .C(g8543), .Z(II14990) ) ;
NOR3    gate7847  (.A(g8199), .B(II14766), .C(II14767), .Z(g8658) ) ;
NOR4    gate7848  (.A(g7658), .B(g7616), .C(g8082), .D(g7634), .Z(g8523) ) ;
NOR4    gate7849  (.A(g7658), .B(g7616), .C(g8082), .D(g7634), .Z(g8279) ) ;
NOR4    gate7850  (.A(g7658), .B(g7616), .C(g8082), .D(g7634), .Z(g8360) ) ;
OR4     gate7851  (.A(g8131), .B(g8111), .C(g8042), .D(g8156), .Z(II15017) ) ;
OR4     gate7852  (.A(g7855), .B(g7838), .C(g7905), .D(g7870), .Z(II15018) ) ;
OR4     gate7853  (.A(g7951), .B(g7920), .C(g7983), .D(g8181), .Z(II15019) ) ;
OR4     gate7854  (.A(g8363), .B(g8342), .C(g8407), .D(g8386), .Z(II15020) ) ;
OR4     gate7855  (.A(II15017), .B(II15018), .C(II15019), .D(II15020), .Z(II15021) ) ;
OR4     gate7856  (.A(g8131), .B(g8111), .C(g8042), .D(g8156), .Z(II15029) ) ;
OR4     gate7857  (.A(g7855), .B(g7838), .C(g7905), .D(g7870), .Z(II15030) ) ;
OR4     gate7858  (.A(g7951), .B(g7920), .C(g7983), .D(g8181), .Z(II15031) ) ;
OR4     gate7859  (.A(g8363), .B(g8342), .C(g8407), .D(g8386), .Z(II15032) ) ;
OR4     gate7860  (.A(II15029), .B(II15030), .C(II15031), .D(II15032), .Z(II15033) ) ;
OR4     gate7861  (.A(g8131), .B(g8111), .C(g8042), .D(g8156), .Z(II15040) ) ;
OR4     gate7862  (.A(g7855), .B(g7838), .C(g7905), .D(g7870), .Z(II15041) ) ;
OR4     gate7863  (.A(g7951), .B(g7920), .C(g7983), .D(g8181), .Z(II15042) ) ;
OR4     gate7864  (.A(g8363), .B(g8342), .C(g8407), .D(g8386), .Z(II15043) ) ;
OR4     gate7865  (.A(II15040), .B(II15041), .C(II15042), .D(II15043), .Z(II15044) ) ;
OR4     gate7866  (.A(g8131), .B(g8111), .C(g8042), .D(g8156), .Z(II15051) ) ;
OR4     gate7867  (.A(g7855), .B(g7838), .C(g7905), .D(g7870), .Z(II15052) ) ;
OR4     gate7868  (.A(g7951), .B(g7920), .C(g7983), .D(g8181), .Z(II15053) ) ;
OR4     gate7869  (.A(g8363), .B(g8342), .C(g8407), .D(g8386), .Z(II15054) ) ;
OR4     gate7870  (.A(II15051), .B(II15052), .C(II15053), .D(II15054), .Z(II15055) ) ;
OR4     gate7871  (.A(g8131), .B(g8111), .C(g8042), .D(g8156), .Z(II15071) ) ;
OR4     gate7872  (.A(g7855), .B(g7838), .C(g7905), .D(g7870), .Z(II15072) ) ;
OR4     gate7873  (.A(g7951), .B(g7920), .C(g7983), .D(g8181), .Z(II15073) ) ;
OR4     gate7874  (.A(g8363), .B(g8342), .C(g8407), .D(g8386), .Z(II15074) ) ;
OR4     gate7875  (.A(II15071), .B(II15072), .C(II15073), .D(II15074), .Z(II15075) ) ;
OR4     gate7876  (.A(g8131), .B(g8111), .C(g8042), .D(g8156), .Z(II15082) ) ;
OR4     gate7877  (.A(g7855), .B(g7838), .C(g7905), .D(g7870), .Z(II15083) ) ;
OR4     gate7878  (.A(g7951), .B(g7920), .C(g7983), .D(g8181), .Z(II15084) ) ;
OR4     gate7879  (.A(g8363), .B(g8342), .C(g8407), .D(g8386), .Z(II15085) ) ;
OR4     gate7880  (.A(II15082), .B(II15083), .C(II15084), .D(II15085), .Z(II15086) ) ;
OR4     gate7881  (.A(g8131), .B(g8111), .C(g8042), .D(g8156), .Z(II15098) ) ;
OR4     gate7882  (.A(g7855), .B(g7838), .C(g7905), .D(g7870), .Z(II15099) ) ;
OR4     gate7883  (.A(g7951), .B(g7920), .C(g7983), .D(g8181), .Z(II15100) ) ;
OR4     gate7884  (.A(g8363), .B(g8342), .C(g8407), .D(g8386), .Z(II15101) ) ;
OR4     gate7885  (.A(II15098), .B(II15099), .C(II15100), .D(II15101), .Z(II15102) ) ;
OR4     gate7886  (.A(g8131), .B(g8111), .C(g8042), .D(g8156), .Z(II15109) ) ;
OR4     gate7887  (.A(g7855), .B(g7838), .C(g7905), .D(g7870), .Z(II15110) ) ;
OR4     gate7888  (.A(g7951), .B(g7920), .C(g7983), .D(g8181), .Z(II15111) ) ;
OR4     gate7889  (.A(g8363), .B(g8342), .C(g8407), .D(g8386), .Z(II15112) ) ;
OR4     gate7890  (.A(II15109), .B(II15110), .C(II15111), .D(II15112), .Z(II15113) ) ;
OR3     gate7891  (.A(g8483), .B(g8464), .C(g8514), .Z(II15147) ) ;
OR3     gate7892  (.A(g8483), .B(g8464), .C(g8514), .Z(II15152) ) ;
OR3     gate7893  (.A(g8483), .B(g8464), .C(g8514), .Z(II15165) ) ;
OR3     gate7894  (.A(g8483), .B(g8464), .C(g8514), .Z(II15169) ) ;
OR3     gate7895  (.A(g8483), .B(g8464), .C(g8514), .Z(II15172) ) ;
OR3     gate7896  (.A(g8483), .B(g8464), .C(g8514), .Z(II15175) ) ;
OR4     gate7897  (.A(g8270), .B(g8258), .C(g8281), .D(g8273), .Z(II15228) ) ;
OR4     gate7898  (.A(g8262), .B(g8303), .C(g8268), .D(g8312), .Z(II15229) ) ;
OR4     gate7899  (.A(g8274), .B(g8321), .C(g8298), .D(g8696), .Z(II15230) ) ;
OR4     gate7900  (.A(g8701), .B(g8715), .C(g8730), .D(g8720), .Z(II15231) ) ;
OR4     gate7901  (.A(II15228), .B(II15229), .C(II15230), .D(II15231), .Z(II15232) ) ;
NOR3    gate7902  (.A(g8443), .B(g8421), .C(II15102), .Z(g8818) ) ;
OR4     gate7903  (.A(g8264), .B(g8260), .C(g8277), .D(g8301), .Z(II15239) ) ;
OR4     gate7904  (.A(g8259), .B(g8294), .C(g8263), .D(g8305), .Z(II15240) ) ;
OR4     gate7905  (.A(g8269), .B(g8314), .C(g8309), .D(g8695), .Z(II15241) ) ;
OR4     gate7906  (.A(g8697), .B(g8714), .C(g8718), .D(g8719), .Z(II15242) ) ;
OR4     gate7907  (.A(II15239), .B(II15240), .C(II15241), .D(II15242), .Z(II15243) ) ;
NOR3    gate7908  (.A(g8443), .B(g8421), .C(II15044), .Z(g8806) ) ;
OR4     gate7909  (.A(g8238), .B(g8265), .C(g8272), .D(g8292), .Z(II15250) ) ;
OR4     gate7910  (.A(g8302), .B(g8288), .C(g8311), .D(g8296), .Z(II15251) ) ;
OR4     gate7911  (.A(g8320), .B(g8307), .C(g8317), .D(g8692), .Z(II15252) ) ;
OR4     gate7912  (.A(g8698), .B(g8711), .C(g8722), .D(g8716), .Z(II15253) ) ;
OR4     gate7913  (.A(II15250), .B(II15251), .C(II15252), .D(II15253), .Z(II15254) ) ;
NOR3    gate7914  (.A(g8443), .B(g8421), .C(II15086), .Z(g8812) ) ;
OR4     gate7915  (.A(g8256), .B(g8271), .C(g8267), .D(g8286), .Z(II15261) ) ;
OR4     gate7916  (.A(g8293), .B(g8283), .C(g8304), .D(g8289), .Z(II15262) ) ;
OR4     gate7917  (.A(g8313), .B(g8297), .C(g8310), .D(g8690), .Z(II15263) ) ;
OR4     gate7918  (.A(g8700), .B(g8708), .C(g8726), .D(g8731), .Z(II15264) ) ;
OR4     gate7919  (.A(II15261), .B(II15262), .C(II15263), .D(II15264), .Z(II15265) ) ;
NOR3    gate7920  (.A(g8443), .B(g8421), .C(II15113), .Z(g8819) ) ;
OR4     gate7921  (.A(g8237), .B(g8300), .C(g8261), .D(g8282), .Z(II15272) ) ;
OR4     gate7922  (.A(g8287), .B(g8334), .C(g8295), .D(g8339), .Z(II15273) ) ;
OR4     gate7923  (.A(g8306), .B(g8361), .C(g8299), .D(g8687), .Z(II15274) ) ;
OR4     gate7924  (.A(g8693), .B(g8703), .C(g8712), .D(g8717), .Z(II15275) ) ;
OR4     gate7925  (.A(II15272), .B(II15273), .C(II15274), .D(II15275), .Z(II15276) ) ;
NOR3    gate7926  (.A(g8443), .B(g8421), .C(II15055), .Z(g8807) ) ;
OR4     gate7927  (.A(g8291), .B(g8276), .C(g8325), .D(g8330), .Z(II15283) ) ;
OR4     gate7928  (.A(g8335), .B(g8340), .C(g8290), .D(g8691), .Z(II15284) ) ;
NOR3    gate7929  (.A(g8443), .B(g8421), .C(II15021), .Z(g8803) ) ;
OR3     gate7930  (.A(g8709), .B(g8713), .C(g8803), .Z(II15285) ) ;
OR4     gate7931  (.A(g8285), .B(g8266), .C(g8318), .D(g8326), .Z(II15290) ) ;
OR4     gate7932  (.A(g8331), .B(g8336), .C(g8338), .D(g8688), .Z(II15291) ) ;
NOR3    gate7933  (.A(g8443), .B(g8421), .C(II15033), .Z(g8805) ) ;
OR3     gate7934  (.A(g8704), .B(g8710), .C(g8805), .Z(II15292) ) ;
OR4     gate7935  (.A(g8280), .B(g8257), .C(g8319), .D(g8327), .Z(II15297) ) ;
OR4     gate7936  (.A(g8332), .B(g8333), .C(g8686), .D(g8702), .Z(II15298) ) ;
NOR3    gate7937  (.A(g8443), .B(g8421), .C(II15075), .Z(g8811) ) ;
NOR3    gate7938  (.A(g7658), .B(g8613), .C(g7634), .Z(g8706) ) ;
NOR3    gate7939  (.A(g7658), .B(g8613), .C(g7634), .Z(g8694) ) ;
NOR3    gate7940  (.A(g7658), .B(g8613), .C(g7634), .Z(g8699) ) ;
NOR3    gate7941  (.A(g7658), .B(g8613), .C(g7634), .Z(g8707) ) ;
NOR3    gate7942  (.A(g7658), .B(g8613), .C(g7634), .Z(g8855) ) ;
OR3     gate7943  (.A(g8736), .B(g8748), .C(g8740), .Z(II15400) ) ;
NOR3    gate7944  (.A(g8493), .B(g8239), .C(II15175), .Z(g8863) ) ;
NOR3    gate7945  (.A(g8493), .B(g8239), .C(II15147), .Z(g8847) ) ;
NOR3    gate7946  (.A(g8493), .B(g8239), .C(II15152), .Z(g8850) ) ;
NOR3    gate7947  (.A(g8493), .B(g8239), .C(II15172), .Z(g8862) ) ;
NOR3    gate7948  (.A(g8493), .B(g8239), .C(II15169), .Z(g8861) ) ;
NOR3    gate7949  (.A(g8493), .B(g8239), .C(II14831), .Z(g8679) ) ;
NOR3    gate7950  (.A(g8493), .B(g8239), .C(II14834), .Z(g8680) ) ;
NOR3    gate7951  (.A(g8493), .B(g8239), .C(II15165), .Z(g8859) ) ;
NAND2   gate7952  (.A(g1532), .B(g1528), .Z(II5505) ) ;
NAND2   gate7953  (.A(g1532), .B(II5505), .Z(II5506) ) ;
NAND2   gate7954  (.A(g1528), .B(II5505), .Z(II5507) ) ;
NAND2   gate7955  (.A(g1087), .B(g1098), .Z(II5519) ) ;
NAND2   gate7956  (.A(g1087), .B(II5519), .Z(II5520) ) ;
NAND2   gate7957  (.A(g1098), .B(II5519), .Z(II5521) ) ;
NAND2   gate7958  (.A(g1481), .B(g1489), .Z(II5598) ) ;
NAND2   gate7959  (.A(g1481), .B(II5598), .Z(II5599) ) ;
NAND2   gate7960  (.A(g1489), .B(II5598), .Z(II5600) ) ;
NAND2   gate7961  (.A(g1092), .B(g1130), .Z(II5619) ) ;
NAND2   gate7962  (.A(g1092), .B(II5619), .Z(II5620) ) ;
NAND2   gate7963  (.A(g1130), .B(II5619), .Z(II5621) ) ;
NAND2   gate7964  (.A(g1513), .B(g1524), .Z(II5695) ) ;
NAND2   gate7965  (.A(g1513), .B(II5695), .Z(II5696) ) ;
NAND2   gate7966  (.A(g1524), .B(II5695), .Z(II5697) ) ;
NAND2   gate7967  (.A(g1435), .B(g1439), .Z(g1910) ) ;
NAND2   gate7968  (.A(g1444), .B(g1450), .Z(g2051) ) ;
NAND2   gate7969  (.A(g852), .B(g883), .Z(II6064) ) ;
NAND2   gate7970  (.A(g852), .B(II6064), .Z(II6065) ) ;
NAND2   gate7971  (.A(g883), .B(II6064), .Z(II6066) ) ;
NAND2   gate7972  (.A(g849), .B(g921), .Z(II6102) ) ;
NAND2   gate7973  (.A(g849), .B(II6102), .Z(II6103) ) ;
NAND2   gate7974  (.A(g921), .B(II6102), .Z(II6104) ) ;
NAND2   gate7975  (.A(g846), .B(g916), .Z(II6133) ) ;
NAND2   gate7976  (.A(g846), .B(II6133), .Z(II6134) ) ;
NAND2   gate7977  (.A(g916), .B(II6133), .Z(II6135) ) ;
NAND2   gate7978  (.A(g985), .B(g990), .Z(g2333) ) ;
NAND2   gate7979  (.A(g843), .B(g911), .Z(II6170) ) ;
NAND2   gate7980  (.A(g843), .B(II6170), .Z(II6171) ) ;
NAND2   gate7981  (.A(g911), .B(II6170), .Z(II6172) ) ;
NAND2   gate7982  (.A(g831), .B(g891), .Z(II6201) ) ;
NAND2   gate7983  (.A(g831), .B(II6201), .Z(II6202) ) ;
NAND2   gate7984  (.A(g891), .B(II6201), .Z(II6203) ) ;
NAND2   gate7985  (.A(g834), .B(g896), .Z(II6232) ) ;
NAND2   gate7986  (.A(g834), .B(II6232), .Z(II6233) ) ;
NAND2   gate7987  (.A(g896), .B(II6232), .Z(II6234) ) ;
NAND2   gate7988  (.A(g837), .B(g901), .Z(II6257) ) ;
NAND2   gate7989  (.A(g837), .B(II6257), .Z(II6258) ) ;
NAND2   gate7990  (.A(g901), .B(II6257), .Z(II6259) ) ;
NAND2   gate7991  (.A(g840), .B(g906), .Z(II6273) ) ;
NAND2   gate7992  (.A(g840), .B(II6273), .Z(II6274) ) ;
NAND2   gate7993  (.A(g906), .B(II6273), .Z(II6275) ) ;
NAND2   gate7994  (.A(g1913), .B(g1537), .Z(II6499) ) ;
NAND2   gate7995  (.A(g1913), .B(II6499), .Z(II6500) ) ;
NAND2   gate7996  (.A(g1537), .B(II6499), .Z(II6501) ) ;
NAND2   gate7997  (.A(g1919), .B(g1102), .Z(II6522) ) ;
NAND2   gate7998  (.A(g1919), .B(II6522), .Z(II6523) ) ;
NAND2   gate7999  (.A(g1102), .B(II6522), .Z(II6524) ) ;
NAND2   gate8000  (.A(g2555), .B(g2557), .Z(II6538) ) ;
NAND2   gate8001  (.A(g2555), .B(II6538), .Z(II6539) ) ;
NAND2   gate8002  (.A(g2557), .B(II6538), .Z(II6540) ) ;
NAND2   gate8003  (.A(g195), .B(g1970), .Z(II6739) ) ;
NAND2   gate8004  (.A(g195), .B(II6739), .Z(II6740) ) ;
NAND2   gate8005  (.A(g1970), .B(II6739), .Z(II6741) ) ;
NAND2   gate8006  (.A(g1733), .B(g1494), .Z(II6750) ) ;
NAND2   gate8007  (.A(g1733), .B(II6750), .Z(II6751) ) ;
NAND2   gate8008  (.A(g1494), .B(II6750), .Z(II6752) ) ;
NAND2   gate8009  (.A(g186), .B(g1983), .Z(II6757) ) ;
NAND2   gate8010  (.A(g186), .B(II6757), .Z(II6758) ) ;
NAND2   gate8011  (.A(g1983), .B(II6757), .Z(II6759) ) ;
NAND2   gate8012  (.A(g2386), .B(g1134), .Z(II6774) ) ;
NAND2   gate8013  (.A(g2386), .B(II6774), .Z(II6775) ) ;
NAND2   gate8014  (.A(g1134), .B(II6774), .Z(II6776) ) ;
NAND2   gate8015  (.A(g210), .B(g2052), .Z(II6813) ) ;
NAND2   gate8016  (.A(g210), .B(II6813), .Z(II6814) ) ;
NAND2   gate8017  (.A(g2052), .B(II6813), .Z(II6815) ) ;
NAND2   gate8018  (.A(g205), .B(g2016), .Z(II6842) ) ;
NAND2   gate8019  (.A(g205), .B(II6842), .Z(II6843) ) ;
NAND2   gate8020  (.A(g2016), .B(II6842), .Z(II6844) ) ;
NAND2   gate8021  (.A(g1967), .B(g1910), .Z(II6876) ) ;
NAND2   gate8022  (.A(g1967), .B(II6876), .Z(II6877) ) ;
NAND2   gate8023  (.A(g1910), .B(II6876), .Z(II6878) ) ;
NAND2   gate8024  (.A(g1889), .B(g1904), .Z(g3231) ) ;
NAND2   gate8025  (.A(g2298), .B(g2276), .Z(g3232) ) ;
NAND2   gate8026  (.A(g2105), .B(g1838), .Z(II6904) ) ;
NAND2   gate8027  (.A(g2105), .B(II6904), .Z(II6905) ) ;
NAND2   gate8028  (.A(g1838), .B(II6904), .Z(II6906) ) ;
NAND2   gate8029  (.A(g2360), .B(g1732), .Z(II6916) ) ;
NAND2   gate8030  (.A(g2360), .B(II6916), .Z(II6917) ) ;
NAND2   gate8031  (.A(g1732), .B(II6916), .Z(II6918) ) ;
NAND2   gate8032  (.A(g1728), .B(g33), .Z(II6923) ) ;
NAND2   gate8033  (.A(g1728), .B(II6923), .Z(II6924) ) ;
NAND2   gate8034  (.A(g33), .B(II6923), .Z(II6925) ) ;
NAND2   gate8035  (.A(g2161), .B(g2051), .Z(II6939) ) ;
NAND2   gate8036  (.A(g2161), .B(II6939), .Z(II6940) ) ;
NAND2   gate8037  (.A(g2051), .B(II6939), .Z(II6941) ) ;
NAND2   gate8038  (.A(g2275), .B(g2242), .Z(II6996) ) ;
NAND2   gate8039  (.A(g2275), .B(II6996), .Z(II6997) ) ;
NAND2   gate8040  (.A(g2242), .B(II6996), .Z(II6998) ) ;
NAND2   gate8041  (.A(g2295), .B(g2333), .Z(II7009) ) ;
NAND2   gate8042  (.A(g2295), .B(II7009), .Z(II7010) ) ;
NAND2   gate8043  (.A(g2333), .B(II7009), .Z(II7011) ) ;
NAND2   gate8044  (.A(g1639), .B(g1643), .Z(II7068) ) ;
NAND2   gate8045  (.A(g1639), .B(II7068), .Z(II7069) ) ;
NAND2   gate8046  (.A(g1643), .B(II7068), .Z(II7070) ) ;
NAND2   gate8047  (.A(g1753), .B(g1918), .Z(II7085) ) ;
NAND2   gate8048  (.A(g1753), .B(II7085), .Z(II7086) ) ;
NAND2   gate8049  (.A(g1918), .B(II7085), .Z(II7087) ) ;
NAND2   gate8050  (.A(g2404), .B(g2397), .Z(II7138) ) ;
NAND2   gate8051  (.A(g2404), .B(II7138), .Z(II7139) ) ;
NAND2   gate8052  (.A(g2397), .B(II7138), .Z(II7140) ) ;
NAND2   gate8053  (.A(g799), .B(g1974), .Z(II7148) ) ;
NAND2   gate8054  (.A(g799), .B(II7148), .Z(II7149) ) ;
NAND2   gate8055  (.A(g1974), .B(II7148), .Z(II7150) ) ;
NAND2   gate8056  (.A(g2331), .B(g929), .Z(II7156) ) ;
NAND2   gate8057  (.A(g2331), .B(II7156), .Z(II7157) ) ;
NAND2   gate8058  (.A(g929), .B(II7156), .Z(II7158) ) ;
NAND2   gate8059  (.A(g1739), .B(g2006), .Z(II7172) ) ;
NAND2   gate8060  (.A(g1739), .B(II7172), .Z(II7173) ) ;
NAND2   gate8061  (.A(g2006), .B(II7172), .Z(II7174) ) ;
NAND2   gate8062  (.A(g2351), .B(g795), .Z(II7179) ) ;
NAND2   gate8063  (.A(g2351), .B(II7179), .Z(II7180) ) ;
NAND2   gate8064  (.A(g795), .B(II7179), .Z(II7181) ) ;
NAND2   gate8065  (.A(g2353), .B(g1834), .Z(II7186) ) ;
NAND2   gate8066  (.A(g2353), .B(II7186), .Z(II7187) ) ;
NAND2   gate8067  (.A(g1834), .B(II7186), .Z(II7188) ) ;
NAND2   gate8068  (.A(g866), .B(g2368), .Z(g3681) ) ;
NAND2   gate8069  (.A(g815), .B(g2091), .Z(II7214) ) ;
NAND2   gate8070  (.A(g815), .B(II7214), .Z(II7215) ) ;
NAND2   gate8071  (.A(g2091), .B(II7214), .Z(II7216) ) ;
NAND2   gate8072  (.A(g1658), .B(g2134), .Z(II7239) ) ;
NAND2   gate8073  (.A(g1658), .B(II7239), .Z(II7240) ) ;
NAND2   gate8074  (.A(g2134), .B(II7239), .Z(II7241) ) ;
NAND2   gate8075  (.A(g2486), .B(g955), .Z(II7268) ) ;
NAND2   gate8076  (.A(g2486), .B(II7268), .Z(II7269) ) ;
NAND2   gate8077  (.A(g955), .B(II7268), .Z(II7270) ) ;
NAND2   gate8078  (.A(g2497), .B(g1898), .Z(II7277) ) ;
NAND2   gate8079  (.A(g2497), .B(II7277), .Z(II7278) ) ;
NAND2   gate8080  (.A(g1898), .B(II7277), .Z(II7279) ) ;
NAND2   gate8081  (.A(g2276), .B(g3188), .Z(g3883) ) ;
NAND2   gate8082  (.A(g2525), .B(g2703), .Z(II7421) ) ;
NAND2   gate8083  (.A(g2525), .B(II7421), .Z(II7422) ) ;
NAND2   gate8084  (.A(g2703), .B(II7421), .Z(II7423) ) ;
NAND2   gate8085  (.A(II7422), .B(II7423), .Z(g3886) ) ;
NAND2   gate8086  (.A(g3222), .B(g1541), .Z(II7428) ) ;
NAND2   gate8087  (.A(g3222), .B(II7428), .Z(II7429) ) ;
NAND2   gate8088  (.A(g1541), .B(II7428), .Z(II7430) ) ;
NAND2   gate8089  (.A(g2517), .B(g3822), .Z(II7436) ) ;
NAND2   gate8090  (.A(g2517), .B(II7436), .Z(II7437) ) ;
NAND2   gate8091  (.A(g3822), .B(II7436), .Z(II7438) ) ;
NAND2   gate8092  (.A(II7437), .B(II7438), .Z(g3889) ) ;
NAND2   gate8093  (.A(g2973), .B(g1701), .Z(II7443) ) ;
NAND2   gate8094  (.A(g2973), .B(II7443), .Z(II7444) ) ;
NAND2   gate8095  (.A(g1701), .B(II7443), .Z(II7445) ) ;
NAND2   gate8096  (.A(g3226), .B(g1106), .Z(II7452) ) ;
NAND2   gate8097  (.A(g3226), .B(II7452), .Z(II7453) ) ;
NAND2   gate8098  (.A(g1106), .B(II7452), .Z(II7454) ) ;
NAND2   gate8099  (.A(g2506), .B(g3815), .Z(II7459) ) ;
NAND2   gate8100  (.A(g2506), .B(II7459), .Z(II7460) ) ;
NAND2   gate8101  (.A(g3815), .B(II7459), .Z(II7461) ) ;
NAND2   gate8102  (.A(II7460), .B(II7461), .Z(g3894) ) ;
NAND2   gate8103  (.A(g2982), .B(g1704), .Z(II7466) ) ;
NAND2   gate8104  (.A(g2982), .B(II7466), .Z(II7467) ) ;
NAND2   gate8105  (.A(g1704), .B(II7466), .Z(II7468) ) ;
NAND2   gate8106  (.A(g2502), .B(g3808), .Z(II7478) ) ;
NAND2   gate8107  (.A(g2502), .B(II7478), .Z(II7479) ) ;
NAND2   gate8108  (.A(g3808), .B(II7478), .Z(II7480) ) ;
NAND2   gate8109  (.A(II7479), .B(II7480), .Z(g3899) ) ;
NAND2   gate8110  (.A(g2989), .B(g1708), .Z(II7485) ) ;
NAND2   gate8111  (.A(g2989), .B(II7485), .Z(II7486) ) ;
NAND2   gate8112  (.A(g1708), .B(II7485), .Z(II7487) ) ;
NAND2   gate8113  (.A(g2498), .B(g3802), .Z(II7503) ) ;
NAND2   gate8114  (.A(g2498), .B(II7503), .Z(II7504) ) ;
NAND2   gate8115  (.A(g3802), .B(II7503), .Z(II7505) ) ;
NAND2   gate8116  (.A(II7504), .B(II7505), .Z(g3906) ) ;
NAND2   gate8117  (.A(g2992), .B(g1711), .Z(II7510) ) ;
NAND2   gate8118  (.A(g2992), .B(II7510), .Z(II7511) ) ;
NAND2   gate8119  (.A(g1711), .B(II7510), .Z(II7512) ) ;
NAND2   gate8120  (.A(g2487), .B(g3787), .Z(II7531) ) ;
NAND2   gate8121  (.A(g2487), .B(II7531), .Z(II7532) ) ;
NAND2   gate8122  (.A(g3787), .B(II7531), .Z(II7533) ) ;
NAND2   gate8123  (.A(II7532), .B(II7533), .Z(g3914) ) ;
NAND2   gate8124  (.A(g2996), .B(g1715), .Z(II7538) ) ;
NAND2   gate8125  (.A(g2996), .B(II7538), .Z(II7539) ) ;
NAND2   gate8126  (.A(g1715), .B(II7538), .Z(II7540) ) ;
NAND2   gate8127  (.A(g2481), .B(g3780), .Z(II7567) ) ;
NAND2   gate8128  (.A(g2481), .B(II7567), .Z(II7568) ) ;
NAND2   gate8129  (.A(g3780), .B(II7567), .Z(II7569) ) ;
NAND2   gate8130  (.A(II7568), .B(II7569), .Z(g3924) ) ;
NAND2   gate8131  (.A(g2999), .B(g1718), .Z(II7574) ) ;
NAND2   gate8132  (.A(g2999), .B(II7574), .Z(II7575) ) ;
NAND2   gate8133  (.A(g1718), .B(II7574), .Z(II7576) ) ;
NAND2   gate8134  (.A(g2471), .B(g3771), .Z(II7609) ) ;
NAND2   gate8135  (.A(g2471), .B(II7609), .Z(II7610) ) ;
NAND2   gate8136  (.A(g3771), .B(II7609), .Z(II7611) ) ;
NAND2   gate8137  (.A(II7610), .B(II7611), .Z(g3938) ) ;
NAND2   gate8138  (.A(g3008), .B(g1721), .Z(II7616) ) ;
NAND2   gate8139  (.A(g3008), .B(II7616), .Z(II7617) ) ;
NAND2   gate8140  (.A(g1721), .B(II7616), .Z(II7618) ) ;
NAND2   gate8141  (.A(g2979), .B(g1499), .Z(II7891) ) ;
NAND2   gate8142  (.A(g2979), .B(II7891), .Z(II7892) ) ;
NAND2   gate8143  (.A(g1499), .B(II7891), .Z(II7893) ) ;
NAND2   gate8144  (.A(g3614), .B(g1138), .Z(II7937) ) ;
NAND2   gate8145  (.A(g3614), .B(II7937), .Z(II7938) ) ;
NAND2   gate8146  (.A(g1138), .B(II7937), .Z(II7939) ) ;
NAND2   gate8147  (.A(g1904), .B(g3220), .Z(II8119) ) ;
NAND2   gate8148  (.A(g1904), .B(II8119), .Z(II8120) ) ;
NAND2   gate8149  (.A(g3220), .B(II8119), .Z(II8121) ) ;
NAND2   gate8150  (.A(g3232), .B(g1646), .Z(II8132) ) ;
NAND2   gate8151  (.A(g3232), .B(II8132), .Z(II8133) ) ;
NAND2   gate8152  (.A(g1646), .B(II8132), .Z(II8134) ) ;
NAND2   gate8153  (.A(g2276), .B(g3258), .Z(g4231) ) ;
NAND2   gate8154  (.A(g3229), .B(g38), .Z(II8150) ) ;
NAND2   gate8155  (.A(g3229), .B(II8150), .Z(II8151) ) ;
NAND2   gate8156  (.A(g38), .B(II8150), .Z(II8152) ) ;
NAND2   gate8157  (.A(g1943), .B(g3231), .Z(II8164) ) ;
NAND2   gate8158  (.A(g1943), .B(II8164), .Z(II8165) ) ;
NAND2   gate8159  (.A(g3231), .B(II8164), .Z(II8166) ) ;
NAND2   gate8160  (.A(g3549), .B(g3533), .Z(g4244) ) ;
NAND2   gate8161  (.A(g2276), .B(g3313), .Z(g4252) ) ;
NAND2   gate8162  (.A(g2011), .B(g3506), .Z(II8243) ) ;
NAND2   gate8163  (.A(g2011), .B(II8243), .Z(II8244) ) ;
NAND2   gate8164  (.A(g3506), .B(II8243), .Z(II8245) ) ;
NAND2   gate8165  (.A(II8244), .B(II8245), .Z(g4294) ) ;
NAND2   gate8166  (.A(g2454), .B(g3825), .Z(II8253) ) ;
NAND2   gate8167  (.A(g2454), .B(II8253), .Z(II8254) ) ;
NAND2   gate8168  (.A(g3825), .B(II8253), .Z(II8255) ) ;
NAND2   gate8169  (.A(II8254), .B(II8255), .Z(g4298) ) ;
NAND3   gate8170  (.A(g3712), .B(g3700), .C(g3732), .Z(g4305) ) ;
NAND2   gate8171  (.A(g3666), .B(g2460), .Z(g4310) ) ;
NAND2   gate8172  (.A(g3712), .B(g3700), .Z(g4313) ) ;
NAND2   gate8173  (.A(g2011), .B(g2721), .Z(II8326) ) ;
NAND2   gate8174  (.A(g2011), .B(II8326), .Z(II8327) ) ;
NAND2   gate8175  (.A(g2721), .B(II8326), .Z(II8328) ) ;
NAND2   gate8176  (.A(II8327), .B(II8328), .Z(g4359) ) ;
NAND2   gate8177  (.A(g2966), .B(g1698), .Z(II8338) ) ;
NAND2   gate8178  (.A(g2966), .B(II8338), .Z(II8339) ) ;
NAND2   gate8179  (.A(g1698), .B(II8338), .Z(II8340) ) ;
NAND2   gate8180  (.A(g2949), .B(g1925), .Z(II8392) ) ;
NAND2   gate8181  (.A(g2949), .B(II8392), .Z(II8393) ) ;
NAND2   gate8182  (.A(g1925), .B(II8392), .Z(II8394) ) ;
NAND2   gate8183  (.A(g2525), .B(g2821), .Z(II8470) ) ;
NAND2   gate8184  (.A(g2525), .B(II8470), .Z(II8471) ) ;
NAND2   gate8185  (.A(g2821), .B(II8470), .Z(II8472) ) ;
NAND2   gate8186  (.A(II8471), .B(II8472), .Z(g4456) ) ;
NAND2   gate8187  (.A(g2986), .B(g2038), .Z(II8502) ) ;
NAND2   gate8188  (.A(g2986), .B(II8502), .Z(II8503) ) ;
NAND2   gate8189  (.A(g2038), .B(II8502), .Z(II8504) ) ;
NAND2   gate8190  (.A(g2517), .B(g2807), .Z(II8510) ) ;
NAND2   gate8191  (.A(g2517), .B(II8510), .Z(II8511) ) ;
NAND2   gate8192  (.A(g2807), .B(II8510), .Z(II8512) ) ;
NAND2   gate8193  (.A(II8511), .B(II8512), .Z(g4476) ) ;
NAND2   gate8194  (.A(g2506), .B(g2798), .Z(II8536) ) ;
NAND2   gate8195  (.A(g2506), .B(II8536), .Z(II8537) ) ;
NAND2   gate8196  (.A(g2798), .B(II8536), .Z(II8538) ) ;
NAND2   gate8197  (.A(II8537), .B(II8538), .Z(g4492) ) ;
NAND2   gate8198  (.A(g2502), .B(g2790), .Z(II8558) ) ;
NAND2   gate8199  (.A(g2502), .B(II8558), .Z(II8559) ) ;
NAND2   gate8200  (.A(g2790), .B(II8558), .Z(II8560) ) ;
NAND2   gate8201  (.A(II8559), .B(II8560), .Z(g4502) ) ;
NAND2   gate8202  (.A(g2498), .B(g2777), .Z(II8581) ) ;
NAND2   gate8203  (.A(g2498), .B(II8581), .Z(II8582) ) ;
NAND2   gate8204  (.A(g2777), .B(II8581), .Z(II8583) ) ;
NAND2   gate8205  (.A(II8582), .B(II8583), .Z(g4513) ) ;
NAND2   gate8206  (.A(g2487), .B(g2764), .Z(II8605) ) ;
NAND2   gate8207  (.A(g2487), .B(II8605), .Z(II8606) ) ;
NAND2   gate8208  (.A(g2764), .B(II8605), .Z(II8607) ) ;
NAND2   gate8209  (.A(II8606), .B(II8607), .Z(g4528) ) ;
NAND2   gate8210  (.A(g2481), .B(g2743), .Z(II8635) ) ;
NAND2   gate8211  (.A(g2481), .B(II8635), .Z(II8636) ) ;
NAND2   gate8212  (.A(g2743), .B(II8635), .Z(II8637) ) ;
NAND2   gate8213  (.A(II8636), .B(II8637), .Z(g4548) ) ;
NAND2   gate8214  (.A(g2471), .B(g2724), .Z(II8658) ) ;
NAND2   gate8215  (.A(g2471), .B(II8658), .Z(II8659) ) ;
NAND2   gate8216  (.A(g2724), .B(II8658), .Z(II8660) ) ;
NAND2   gate8217  (.A(II8659), .B(II8660), .Z(g4563) ) ;
NAND2   gate8218  (.A(g2467), .B(g2706), .Z(II8678) ) ;
NAND2   gate8219  (.A(g2467), .B(II8678), .Z(II8679) ) ;
NAND2   gate8220  (.A(g2706), .B(II8678), .Z(II8680) ) ;
NAND2   gate8221  (.A(II8679), .B(II8680), .Z(g4575) ) ;
NAND2   gate8222  (.A(g4239), .B(g1545), .Z(II8938) ) ;
NAND2   gate8223  (.A(g4239), .B(II8938), .Z(II8939) ) ;
NAND2   gate8224  (.A(g1545), .B(II8938), .Z(II8940) ) ;
NAND2   gate8225  (.A(g4246), .B(g1110), .Z(II8955) ) ;
NAND2   gate8226  (.A(g4246), .B(II8955), .Z(II8956) ) ;
NAND2   gate8227  (.A(g1110), .B(II8955), .Z(II8957) ) ;
NAND2   gate8228  (.A(g2460), .B(g4271), .Z(g4700) ) ;
NAND2   gate8229  (.A(g4059), .B(g1504), .Z(II9057) ) ;
NAND2   gate8230  (.A(g4059), .B(II9057), .Z(II9058) ) ;
NAND2   gate8231  (.A(g1504), .B(II9057), .Z(II9059) ) ;
NAND2   gate8232  (.A(g4400), .B(g1149), .Z(II9069) ) ;
NAND2   gate8233  (.A(g4400), .B(II9069), .Z(II9070) ) ;
NAND2   gate8234  (.A(g1149), .B(II9069), .Z(II9071) ) ;
NAND2   gate8235  (.A(g3883), .B(g1649), .Z(II9151) ) ;
NAND2   gate8236  (.A(g3883), .B(II9151), .Z(II9152) ) ;
NAND2   gate8237  (.A(g1649), .B(II9151), .Z(II9153) ) ;
NAND2   gate8238  (.A(g1935), .B(g4244), .Z(II9169) ) ;
NAND2   gate8239  (.A(g1935), .B(II9169), .Z(II9170) ) ;
NAND2   gate8240  (.A(g4244), .B(II9169), .Z(II9171) ) ;
NAND2   gate8241  (.A(g4220), .B(g3605), .Z(g4821) ) ;
NAND2   gate8242  (.A(g4231), .B(g2007), .Z(II9181) ) ;
NAND2   gate8243  (.A(g4231), .B(II9181), .Z(II9182) ) ;
NAND2   gate8244  (.A(g2007), .B(II9181), .Z(II9183) ) ;
NAND3   gate8245  (.A(g3635), .B(g3605), .C(g4220), .Z(g4831) ) ;
NAND2   gate8246  (.A(g4252), .B(g1652), .Z(II9194) ) ;
NAND2   gate8247  (.A(g4252), .B(II9194), .Z(II9195) ) ;
NAND2   gate8248  (.A(g1652), .B(II9194), .Z(II9196) ) ;
NAND2   gate8249  (.A(g4288), .B(g1879), .Z(g4836) ) ;
NAND2   gate8250  (.A(g1879), .B(g4269), .Z(g4839) ) ;
NAND2   gate8251  (.A(g4254), .B(g3533), .Z(g4869) ) ;
NAND4   gate8252  (.A(g3635), .B(g3605), .C(g4220), .D(g3644), .Z(g4871) ) ;
NAND2   gate8253  (.A(g4287), .B(g1879), .Z(g4880) ) ;
NAND2   gate8254  (.A(g2460), .B(g4315), .Z(g4881) ) ;
NAND2   gate8255  (.A(g4310), .B(g2180), .Z(II9233) ) ;
NAND2   gate8256  (.A(g4310), .B(II9233), .Z(II9234) ) ;
NAND2   gate8257  (.A(g2180), .B(II9233), .Z(II9235) ) ;
NAND2   gate8258  (.A(g2540), .B(g4305), .Z(II9241) ) ;
NAND2   gate8259  (.A(g2540), .B(II9241), .Z(II9242) ) ;
NAND2   gate8260  (.A(g4305), .B(II9241), .Z(II9243) ) ;
NAND2   gate8261  (.A(g2460), .B(g4312), .Z(g4893) ) ;
NAND2   gate8262  (.A(g4282), .B(g3533), .Z(g4905) ) ;
NAND2   gate8263  (.A(g2460), .B(g4314), .Z(g4910) ) ;
NAND2   gate8264  (.A(g4320), .B(g2044), .Z(g4911) ) ;
NAND2   gate8265  (.A(g2533), .B(g4313), .Z(II9276) ) ;
NAND2   gate8266  (.A(g2533), .B(II9276), .Z(II9277) ) ;
NAND2   gate8267  (.A(g4313), .B(II9276), .Z(II9278) ) ;
NAND2   gate8268  (.A(g4319), .B(g2460), .Z(g4954) ) ;
NAND2   gate8269  (.A(g4062), .B(g1908), .Z(II9381) ) ;
NAND2   gate8270  (.A(g4062), .B(II9381), .Z(II9382) ) ;
NAND2   gate8271  (.A(g1908), .B(II9381), .Z(II9383) ) ;
NAND2   gate8272  (.A(g4038), .B(g1942), .Z(II9475) ) ;
NAND2   gate8273  (.A(g4038), .B(II9475), .Z(II9476) ) ;
NAND2   gate8274  (.A(g1942), .B(II9475), .Z(II9477) ) ;
NAND2   gate8275  (.A(g1952), .B(g4307), .Z(II9547) ) ;
NAND2   gate8276  (.A(g1952), .B(II9547), .Z(II9548) ) ;
NAND2   gate8277  (.A(g4307), .B(II9547), .Z(II9549) ) ;
NAND2   gate8278  (.A(g5096), .B(g1037), .Z(II9691) ) ;
NAND2   gate8279  (.A(g5096), .B(II9691), .Z(II9692) ) ;
NAND2   gate8280  (.A(g1037), .B(II9691), .Z(II9693) ) ;
NAND2   gate8281  (.A(g4826), .B(g1549), .Z(II9745) ) ;
NAND2   gate8282  (.A(g4826), .B(II9745), .Z(II9746) ) ;
NAND2   gate8283  (.A(g1549), .B(II9745), .Z(II9747) ) ;
NAND2   gate8284  (.A(g4832), .B(g1114), .Z(II9767) ) ;
NAND2   gate8285  (.A(g4832), .B(II9767), .Z(II9768) ) ;
NAND2   gate8286  (.A(g1114), .B(II9767), .Z(II9769) ) ;
NAND3   gate8287  (.A(g4344), .B(g4335), .C(g4963), .Z(g5284) ) ;
NAND3   gate8288  (.A(g4344), .B(g5002), .C(g4963), .Z(g5291) ) ;
NAND3   gate8289  (.A(g5009), .B(g4335), .C(g4328), .Z(g5305) ) ;
NAND3   gate8290  (.A(g5009), .B(g4335), .C(g4963), .Z(g5310) ) ;
NAND3   gate8291  (.A(g5009), .B(g5002), .C(g4963), .Z(g5312) ) ;
NAND2   gate8292  (.A(g4729), .B(g1509), .Z(II9826) ) ;
NAND2   gate8293  (.A(g4729), .B(II9826), .Z(II9827) ) ;
NAND2   gate8294  (.A(g1509), .B(II9826), .Z(II9828) ) ;
NAND2   gate8295  (.A(g1879), .B(g4877), .Z(g5512) ) ;
NAND2   gate8296  (.A(g2128), .B(g4905), .Z(II9946) ) ;
NAND2   gate8297  (.A(g2128), .B(II9946), .Z(II9947) ) ;
NAND2   gate8298  (.A(g4905), .B(II9946), .Z(II9948) ) ;
NAND2   gate8299  (.A(g2131), .B(g4831), .Z(II9953) ) ;
NAND2   gate8300  (.A(g2131), .B(II9953), .Z(II9954) ) ;
NAND2   gate8301  (.A(g4831), .B(II9953), .Z(II9955) ) ;
NAND2   gate8302  (.A(g1938), .B(g4869), .Z(II9963) ) ;
NAND2   gate8303  (.A(g1938), .B(II9963), .Z(II9964) ) ;
NAND2   gate8304  (.A(g4869), .B(II9963), .Z(II9965) ) ;
NAND2   gate8305  (.A(g1879), .B(g4830), .Z(g5550) ) ;
NAND2   gate8306  (.A(g4880), .B(g2092), .Z(II9978) ) ;
NAND2   gate8307  (.A(g4880), .B(II9978), .Z(II9979) ) ;
NAND2   gate8308  (.A(g2092), .B(II9978), .Z(II9980) ) ;
NAND2   gate8309  (.A(g4836), .B(g2096), .Z(II9985) ) ;
NAND2   gate8310  (.A(g4836), .B(II9985), .Z(II9986) ) ;
NAND2   gate8311  (.A(g2096), .B(II9985), .Z(II9987) ) ;
NAND2   gate8312  (.A(g2145), .B(g4871), .Z(II9992) ) ;
NAND2   gate8313  (.A(g2145), .B(II9992), .Z(II9993) ) ;
NAND2   gate8314  (.A(g4871), .B(II9992), .Z(II9994) ) ;
NAND2   gate8315  (.A(g4839), .B(g1929), .Z(II9999) ) ;
NAND2   gate8316  (.A(g4839), .B(II9999), .Z(II10000) ) ;
NAND2   gate8317  (.A(g1929), .B(II9999), .Z(II10001) ) ;
NAND2   gate8318  (.A(g1949), .B(g4821), .Z(II10009) ) ;
NAND2   gate8319  (.A(g1949), .B(II10009), .Z(II10010) ) ;
NAND2   gate8320  (.A(g4821), .B(II10009), .Z(II10011) ) ;
NAND2   gate8321  (.A(g4700), .B(g2174), .Z(II10017) ) ;
NAND2   gate8322  (.A(g4700), .B(II10017), .Z(II10018) ) ;
NAND2   gate8323  (.A(g2174), .B(II10017), .Z(II10019) ) ;
NAND2   gate8324  (.A(g2044), .B(g4933), .Z(g5565) ) ;
NAND2   gate8325  (.A(g1879), .B(g4883), .Z(g5567) ) ;
NAND3   gate8326  (.A(g2044), .B(g4902), .C(g4320), .Z(g5568) ) ;
NAND2   gate8327  (.A(g4893), .B(g2202), .Z(II10038) ) ;
NAND2   gate8328  (.A(g4893), .B(II10038), .Z(II10039) ) ;
NAND2   gate8329  (.A(g2202), .B(II10038), .Z(II10040) ) ;
NOR3    gate8330  (.A(g4298), .B(g4575), .C(g4563), .Z(g4894) ) ;
NOR4    gate8331  (.A(g4548), .B(g4528), .C(g4513), .D(g4502), .Z(g4888) ) ;
NOR4    gate8332  (.A(g4492), .B(g4476), .C(g4456), .D(g4294), .Z(g4884) ) ;
NAND2   gate8333  (.A(g4910), .B(g2226), .Z(II10060) ) ;
NAND2   gate8334  (.A(g4910), .B(II10060), .Z(II10061) ) ;
NAND2   gate8335  (.A(g2226), .B(II10060), .Z(II10062) ) ;
NAND2   gate8336  (.A(g2044), .B(g4906), .Z(g5590) ) ;
NAND2   gate8337  (.A(g4954), .B(g2253), .Z(II10071) ) ;
NAND2   gate8338  (.A(g4954), .B(II10071), .Z(II10072) ) ;
NAND2   gate8339  (.A(g2253), .B(II10071), .Z(II10073) ) ;
NAND2   gate8340  (.A(g4911), .B(g2256), .Z(II10078) ) ;
NAND2   gate8341  (.A(g4911), .B(II10078), .Z(II10079) ) ;
NAND2   gate8342  (.A(g2256), .B(II10078), .Z(II10080) ) ;
NAND2   gate8343  (.A(g4881), .B(g2177), .Z(II10092) ) ;
NAND2   gate8344  (.A(g4881), .B(II10092), .Z(II10093) ) ;
NAND2   gate8345  (.A(g2177), .B(II10092), .Z(II10094) ) ;
NAND2   gate8346  (.A(g2044), .B(g4957), .Z(g5625) ) ;
NAND2   gate8347  (.A(g2276), .B(g4901), .Z(g5632) ) ;
NAND2   gate8348  (.A(g4707), .B(g1916), .Z(II10142) ) ;
NAND2   gate8349  (.A(g4707), .B(II10142), .Z(II10143) ) ;
NAND2   gate8350  (.A(g1916), .B(II10142), .Z(II10144) ) ;
NOR3    gate8351  (.A(g3556), .B(g2872), .C(g3938), .Z(g5056) ) ;
NOR4    gate8352  (.A(g3924), .B(g3914), .C(g3906), .D(g3899), .Z(g5039) ) ;
NOR4    gate8353  (.A(g3894), .B(g3889), .C(g3886), .D(g4359), .Z(g5023) ) ;
NAND2   gate8354  (.A(g4724), .B(g1958), .Z(II10196) ) ;
NAND2   gate8355  (.A(g4724), .B(II10196), .Z(II10197) ) ;
NAND2   gate8356  (.A(g1958), .B(II10196), .Z(II10198) ) ;
NAND2   gate8357  (.A(g2044), .B(g5005), .Z(g5697) ) ;
NAND2   gate8358  (.A(g2522), .B(g4895), .Z(II10223) ) ;
NAND2   gate8359  (.A(g2522), .B(II10223), .Z(II10224) ) ;
NAND2   gate8360  (.A(g4895), .B(II10223), .Z(II10225) ) ;
NAND2   gate8361  (.A(g5461), .B(g2562), .Z(II10298) ) ;
NAND2   gate8362  (.A(g5461), .B(II10298), .Z(II10299) ) ;
NAND2   gate8363  (.A(g2562), .B(II10298), .Z(II10300) ) ;
NAND2   gate8364  (.A(g5470), .B(g3019), .Z(II10305) ) ;
NAND2   gate8365  (.A(g5470), .B(II10305), .Z(II10306) ) ;
NAND2   gate8366  (.A(g3019), .B(II10305), .Z(II10307) ) ;
NAND2   gate8367  (.A(g5484), .B(g1041), .Z(II10313) ) ;
NAND2   gate8368  (.A(g5484), .B(II10313), .Z(II10314) ) ;
NAND2   gate8369  (.A(g1041), .B(II10313), .Z(II10315) ) ;
NAND2   gate8370  (.A(g5459), .B(g2573), .Z(II10320) ) ;
NAND2   gate8371  (.A(g5459), .B(II10320), .Z(II10321) ) ;
NAND2   gate8372  (.A(g2573), .B(II10320), .Z(II10322) ) ;
NAND2   gate8373  (.A(g5467), .B(g2562), .Z(II10327) ) ;
NAND2   gate8374  (.A(g5467), .B(II10327), .Z(II10328) ) ;
NAND2   gate8375  (.A(g2562), .B(II10327), .Z(II10329) ) ;
NAND2   gate8376  (.A(g5462), .B(g2573), .Z(II10334) ) ;
NAND2   gate8377  (.A(g5462), .B(II10334), .Z(II10335) ) ;
NAND2   gate8378  (.A(g2573), .B(II10334), .Z(II10336) ) ;
NAND2   gate8379  (.A(g5552), .B(g1118), .Z(II10359) ) ;
NAND2   gate8380  (.A(g5552), .B(II10359), .Z(II10360) ) ;
NAND2   gate8381  (.A(g1118), .B(II10359), .Z(II10361) ) ;
NAND2   gate8382  (.A(g5314), .B(g1514), .Z(II10625) ) ;
NAND2   gate8383  (.A(g5314), .B(II10625), .Z(II10626) ) ;
NAND2   gate8384  (.A(g1514), .B(II10625), .Z(II10627) ) ;
NAND2   gate8385  (.A(g5550), .B(g2100), .Z(II10743) ) ;
NAND2   gate8386  (.A(g5550), .B(II10743), .Z(II10744) ) ;
NAND2   gate8387  (.A(g2100), .B(II10743), .Z(II10745) ) ;
NAND2   gate8388  (.A(g5512), .B(g2170), .Z(II10789) ) ;
NAND2   gate8389  (.A(g5512), .B(II10789), .Z(II10790) ) ;
NAND2   gate8390  (.A(g2170), .B(II10789), .Z(II10791) ) ;
NAND2   gate8391  (.A(g5567), .B(g2039), .Z(II10818) ) ;
NAND2   gate8392  (.A(g5567), .B(II10818), .Z(II10819) ) ;
NAND2   gate8393  (.A(g2039), .B(II10818), .Z(II10820) ) ;
NAND4   gate8394  (.A(g3735), .B(g3716), .C(g5633), .D(g3754), .Z(g6158) ) ;
NAND2   gate8395  (.A(g5514), .B(g2584), .Z(II10834) ) ;
NAND2   gate8396  (.A(g5514), .B(II10834), .Z(II10835) ) ;
NAND2   gate8397  (.A(g2584), .B(II10834), .Z(II10836) ) ;
NAND2   gate8398  (.A(g5633), .B(g3716), .Z(g6163) ) ;
NAND2   gate8399  (.A(g5490), .B(g2595), .Z(II10847) ) ;
NAND2   gate8400  (.A(g5490), .B(II10847), .Z(II10848) ) ;
NAND2   gate8401  (.A(g2595), .B(II10847), .Z(II10849) ) ;
NAND2   gate8402  (.A(g5521), .B(g2584), .Z(II10854) ) ;
NAND2   gate8403  (.A(g5521), .B(II10854), .Z(II10855) ) ;
NAND2   gate8404  (.A(g2584), .B(II10854), .Z(II10856) ) ;
NAND2   gate8405  (.A(g5480), .B(g2605), .Z(II10866) ) ;
NAND2   gate8406  (.A(g5480), .B(II10866), .Z(II10867) ) ;
NAND2   gate8407  (.A(g2605), .B(II10866), .Z(II10868) ) ;
NAND2   gate8408  (.A(g5516), .B(g2595), .Z(II10873) ) ;
NAND2   gate8409  (.A(g5516), .B(II10873), .Z(II10874) ) ;
NAND2   gate8410  (.A(g2595), .B(II10873), .Z(II10875) ) ;
NAND2   gate8411  (.A(g5590), .B(g2259), .Z(II10888) ) ;
NAND2   gate8412  (.A(g5590), .B(II10888), .Z(II10889) ) ;
NAND2   gate8413  (.A(g2259), .B(II10888), .Z(II10890) ) ;
NAND2   gate8414  (.A(g5520), .B(g2752), .Z(II10899) ) ;
NAND2   gate8415  (.A(g5520), .B(II10899), .Z(II10900) ) ;
NAND2   gate8416  (.A(g2752), .B(II10899), .Z(II10901) ) ;
NAND2   gate8417  (.A(g5492), .B(g2605), .Z(II10906) ) ;
NAND2   gate8418  (.A(g5492), .B(II10906), .Z(II10907) ) ;
NAND2   gate8419  (.A(g2605), .B(II10906), .Z(II10908) ) ;
NAND3   gate8420  (.A(g5633), .B(g3735), .C(g3716), .Z(g6187) ) ;
NAND2   gate8421  (.A(g5525), .B(g2752), .Z(II10923) ) ;
NAND2   gate8422  (.A(g5525), .B(II10923), .Z(II10924) ) ;
NAND2   gate8423  (.A(g2752), .B(II10923), .Z(II10925) ) ;
NAND2   gate8424  (.A(g5565), .B(g2340), .Z(II10952) ) ;
NAND2   gate8425  (.A(g5565), .B(II10952), .Z(II10953) ) ;
NAND2   gate8426  (.A(g2340), .B(II10952), .Z(II10954) ) ;
NAND2   gate8427  (.A(g5625), .B(g2210), .Z(II10980) ) ;
NAND2   gate8428  (.A(g5625), .B(II10980), .Z(II10981) ) ;
NAND2   gate8429  (.A(g2210), .B(II10980), .Z(II10982) ) ;
NAND2   gate8430  (.A(g5632), .B(g2389), .Z(II10991) ) ;
NAND2   gate8431  (.A(g5632), .B(II10991), .Z(II10992) ) ;
NAND2   gate8432  (.A(g2389), .B(II10991), .Z(II10993) ) ;
NAND2   gate8433  (.A(g5697), .B(g2511), .Z(II11078) ) ;
NAND2   gate8434  (.A(g5697), .B(II11078), .Z(II11079) ) ;
NAND2   gate8435  (.A(g2511), .B(II11078), .Z(II11080) ) ;
NAND2   gate8436  (.A(g5515), .B(g2734), .Z(II11094) ) ;
NAND2   gate8437  (.A(g5515), .B(II11094), .Z(II11095) ) ;
NAND2   gate8438  (.A(g2734), .B(II11094), .Z(II11096) ) ;
NAND2   gate8439  (.A(g5491), .B(g2712), .Z(II11101) ) ;
NAND2   gate8440  (.A(g5491), .B(II11101), .Z(II11102) ) ;
NAND2   gate8441  (.A(g2712), .B(II11101), .Z(II11103) ) ;
NAND2   gate8442  (.A(g5522), .B(g2734), .Z(II11108) ) ;
NAND2   gate8443  (.A(g5522), .B(II11108), .Z(II11109) ) ;
NAND2   gate8444  (.A(g2734), .B(II11108), .Z(II11110) ) ;
NAND2   gate8445  (.A(g5481), .B(g3062), .Z(II11115) ) ;
NAND2   gate8446  (.A(g5481), .B(II11115), .Z(II11116) ) ;
NAND2   gate8447  (.A(g3062), .B(II11115), .Z(II11117) ) ;
NAND2   gate8448  (.A(g5517), .B(g2712), .Z(II11122) ) ;
NAND2   gate8449  (.A(g5517), .B(II11122), .Z(II11123) ) ;
NAND2   gate8450  (.A(g2712), .B(II11122), .Z(II11124) ) ;
NAND2   gate8451  (.A(g5476), .B(g3052), .Z(II11135) ) ;
NAND2   gate8452  (.A(g5476), .B(II11135), .Z(II11136) ) ;
NAND2   gate8453  (.A(g3052), .B(II11135), .Z(II11137) ) ;
NAND2   gate8454  (.A(g5493), .B(g3062), .Z(II11142) ) ;
NAND2   gate8455  (.A(g5493), .B(II11142), .Z(II11143) ) ;
NAND2   gate8456  (.A(g3062), .B(II11142), .Z(II11144) ) ;
NAND2   gate8457  (.A(g5473), .B(g3038), .Z(II11149) ) ;
NAND2   gate8458  (.A(g5473), .B(II11149), .Z(II11150) ) ;
NAND2   gate8459  (.A(g3038), .B(II11149), .Z(II11151) ) ;
NAND2   gate8460  (.A(g5482), .B(g3052), .Z(II11156) ) ;
NAND2   gate8461  (.A(g5482), .B(II11156), .Z(II11157) ) ;
NAND2   gate8462  (.A(g3052), .B(II11156), .Z(II11158) ) ;
NAND2   gate8463  (.A(g5469), .B(g3029), .Z(II11163) ) ;
NAND2   gate8464  (.A(g5469), .B(II11163), .Z(II11164) ) ;
NAND2   gate8465  (.A(g3029), .B(II11163), .Z(II11165) ) ;
NAND2   gate8466  (.A(g5477), .B(g3038), .Z(II11170) ) ;
NAND2   gate8467  (.A(g5477), .B(II11170), .Z(II11171) ) ;
NAND2   gate8468  (.A(g3038), .B(II11170), .Z(II11172) ) ;
NAND2   gate8469  (.A(g5466), .B(g3019), .Z(II11177) ) ;
NAND2   gate8470  (.A(g5466), .B(II11177), .Z(II11178) ) ;
NAND2   gate8471  (.A(g3019), .B(II11177), .Z(II11179) ) ;
NAND2   gate8472  (.A(g5474), .B(g3029), .Z(II11184) ) ;
NAND2   gate8473  (.A(g5474), .B(II11184), .Z(II11185) ) ;
NAND2   gate8474  (.A(g3029), .B(II11184), .Z(II11186) ) ;
NAND2   gate8475  (.A(g5984), .B(g1045), .Z(II11549) ) ;
NAND2   gate8476  (.A(g5984), .B(II11549), .Z(II11550) ) ;
NAND2   gate8477  (.A(g1045), .B(II11549), .Z(II11551) ) ;
NAND2   gate8478  (.A(g5894), .B(g1122), .Z(II11574) ) ;
NAND2   gate8479  (.A(g5894), .B(II11574), .Z(II11575) ) ;
NAND2   gate8480  (.A(g1122), .B(II11574), .Z(II11576) ) ;
NAND2   gate8481  (.A(g6239), .B(g1519), .Z(II11614) ) ;
NAND2   gate8482  (.A(g6239), .B(II11614), .Z(II11615) ) ;
NAND2   gate8483  (.A(g1519), .B(II11614), .Z(II11616) ) ;
NAND2   gate8484  (.A(g5814), .B(g6109), .Z(g6559) ) ;
NAND2   gate8485  (.A(g6112), .B(g1486), .Z(II11750) ) ;
NAND2   gate8486  (.A(g6112), .B(II11750), .Z(II11751) ) ;
NAND2   gate8487  (.A(g1486), .B(II11750), .Z(II11752) ) ;
NAND2   gate8488  (.A(g1758), .B(g6118), .Z(II11757) ) ;
NAND2   gate8489  (.A(g1758), .B(II11757), .Z(II11758) ) ;
NAND2   gate8490  (.A(g6118), .B(II11757), .Z(II11759) ) ;
NAND2   gate8491  (.A(g2548), .B(g6158), .Z(II11841) ) ;
NAND2   gate8492  (.A(g2548), .B(II11841), .Z(II11842) ) ;
NAND2   gate8493  (.A(g6158), .B(II11841), .Z(II11843) ) ;
NAND2   gate8494  (.A(g2543), .B(g6187), .Z(II11873) ) ;
NAND2   gate8495  (.A(g2543), .B(II11873), .Z(II11874) ) ;
NAND2   gate8496  (.A(g6187), .B(II11873), .Z(II11875) ) ;
NAND2   gate8497  (.A(g5403), .B(g6252), .Z(g6680) ) ;
NAND2   gate8498  (.A(g5874), .B(g5847), .Z(II12015) ) ;
NAND2   gate8499  (.A(g5874), .B(II12015), .Z(II12016) ) ;
NAND2   gate8500  (.A(g5847), .B(II12015), .Z(II12017) ) ;
NAND2   gate8501  (.A(II12016), .B(II12017), .Z(g6695) ) ;
NAND2   gate8502  (.A(g5918), .B(g5897), .Z(II12031) ) ;
NAND2   gate8503  (.A(g5918), .B(II12031), .Z(II12032) ) ;
NAND2   gate8504  (.A(g5897), .B(II12031), .Z(II12033) ) ;
NAND2   gate8505  (.A(II12032), .B(II12033), .Z(g6701) ) ;
NAND2   gate8506  (.A(g5956), .B(g5939), .Z(II12051) ) ;
NAND2   gate8507  (.A(g5956), .B(II12051), .Z(II12052) ) ;
NAND2   gate8508  (.A(g5939), .B(II12051), .Z(II12053) ) ;
NAND2   gate8509  (.A(II12052), .B(II12053), .Z(g6709) ) ;
NAND2   gate8510  (.A(g5988), .B(g5971), .Z(II12078) ) ;
NAND2   gate8511  (.A(g5988), .B(II12078), .Z(II12079) ) ;
NAND2   gate8512  (.A(g5971), .B(II12078), .Z(II12080) ) ;
NAND2   gate8513  (.A(II12079), .B(II12080), .Z(g6722) ) ;
NAND2   gate8514  (.A(g1961), .B(g6163), .Z(II12179) ) ;
NAND2   gate8515  (.A(g1961), .B(II12179), .Z(II12180) ) ;
NAND2   gate8516  (.A(g6163), .B(II12179), .Z(II12181) ) ;
NAND2   gate8517  (.A(g6689), .B(g1462), .Z(II12550) ) ;
NAND2   gate8518  (.A(g6689), .B(II12550), .Z(II12551) ) ;
NAND2   gate8519  (.A(g1462), .B(II12550), .Z(II12552) ) ;
NAND2   gate8520  (.A(g6574), .B(g1049), .Z(II12575) ) ;
NAND2   gate8521  (.A(g6574), .B(II12575), .Z(II12576) ) ;
NAND2   gate8522  (.A(g1049), .B(II12575), .Z(II12577) ) ;
NAND2   gate8523  (.A(g6582), .B(g1126), .Z(II12596) ) ;
NAND2   gate8524  (.A(g6582), .B(II12596), .Z(II12597) ) ;
NAND2   gate8525  (.A(g1126), .B(II12596), .Z(II12598) ) ;
NAND2   gate8526  (.A(g6722), .B(g6709), .Z(II12832) ) ;
NAND2   gate8527  (.A(g6722), .B(II12832), .Z(II12833) ) ;
NAND2   gate8528  (.A(g6709), .B(II12832), .Z(II12834) ) ;
NAND2   gate8529  (.A(II12833), .B(II12834), .Z(g7065) ) ;
NAND2   gate8530  (.A(g5435), .B(g6680), .Z(g7069) ) ;
NAND2   gate8531  (.A(g6701), .B(g6695), .Z(II12852) ) ;
NAND2   gate8532  (.A(g6701), .B(II12852), .Z(II12853) ) ;
NAND2   gate8533  (.A(g6695), .B(II12852), .Z(II12854) ) ;
NAND2   gate8534  (.A(II12853), .B(II12854), .Z(g7082) ) ;
NAND2   gate8535  (.A(g2536), .B(g6618), .Z(II12869) ) ;
NAND2   gate8536  (.A(g2536), .B(II12869), .Z(II12870) ) ;
NAND2   gate8537  (.A(g6618), .B(II12869), .Z(II12871) ) ;
NAND2   gate8538  (.A(g7003), .B(g1467), .Z(II12951) ) ;
NAND2   gate8539  (.A(g7003), .B(II12951), .Z(II12952) ) ;
NAND2   gate8540  (.A(g1467), .B(II12951), .Z(II12953) ) ;
NAND2   gate8541  (.A(g7010), .B(g1053), .Z(II13002) ) ;
NAND2   gate8542  (.A(g7010), .B(II13002), .Z(II13003) ) ;
NAND2   gate8543  (.A(g1053), .B(II13002), .Z(II13004) ) ;
NAND2   gate8544  (.A(g6941), .B(g1142), .Z(II13016) ) ;
NAND2   gate8545  (.A(g6941), .B(II13016), .Z(II13017) ) ;
NAND2   gate8546  (.A(g1142), .B(II13016), .Z(II13018) ) ;
NAND4   gate8547  (.A(g3757), .B(g3739), .C(g7050), .D(g3770), .Z(g7234) ) ;
NAND2   gate8548  (.A(g7050), .B(g3739), .Z(g7237) ) ;
NAND3   gate8549  (.A(g7050), .B(g3757), .C(g3739), .Z(g7244) ) ;
NAND2   gate8550  (.A(g7065), .B(g7082), .Z(II13213) ) ;
NAND2   gate8551  (.A(g7065), .B(II13213), .Z(II13214) ) ;
NAND2   gate8552  (.A(g7082), .B(II13213), .Z(II13215) ) ;
NAND2   gate8553  (.A(II13214), .B(II13215), .Z(g7257) ) ;
NAND2   gate8554  (.A(g7199), .B(g1472), .Z(II13376) ) ;
NAND2   gate8555  (.A(g7199), .B(II13376), .Z(II13377) ) ;
NAND2   gate8556  (.A(g1472), .B(II13376), .Z(II13378) ) ;
NAND2   gate8557  (.A(g7212), .B(g1057), .Z(II13395) ) ;
NAND2   gate8558  (.A(g7212), .B(II13395), .Z(II13396) ) ;
NAND2   gate8559  (.A(g1057), .B(II13395), .Z(II13397) ) ;
NAND2   gate8560  (.A(g2556), .B(g7234), .Z(II13587) ) ;
NAND2   gate8561  (.A(g2556), .B(II13587), .Z(II13588) ) ;
NAND2   gate8562  (.A(g7234), .B(II13587), .Z(II13589) ) ;
NAND2   gate8563  (.A(g2551), .B(g7244), .Z(II13598) ) ;
NAND2   gate8564  (.A(g2551), .B(II13598), .Z(II13599) ) ;
NAND2   gate8565  (.A(g7244), .B(II13598), .Z(II13600) ) ;
NAND2   gate8566  (.A(g7257), .B(g7069), .Z(II13638) ) ;
NAND2   gate8567  (.A(g7257), .B(II13638), .Z(II13639) ) ;
NAND2   gate8568  (.A(g7069), .B(II13638), .Z(II13640) ) ;
NAND2   gate8569  (.A(g1977), .B(g7237), .Z(II13685) ) ;
NAND2   gate8570  (.A(g1977), .B(II13685), .Z(II13686) ) ;
NAND2   gate8571  (.A(g7237), .B(II13685), .Z(II13687) ) ;
NAND2   gate8572  (.A(g7427), .B(g1477), .Z(II13785) ) ;
NAND2   gate8573  (.A(g7427), .B(II13785), .Z(II13786) ) ;
NAND2   gate8574  (.A(g1477), .B(II13785), .Z(II13787) ) ;
NAND2   gate8575  (.A(g7429), .B(g1061), .Z(II13800) ) ;
NAND2   gate8576  (.A(g7429), .B(II13800), .Z(II13801) ) ;
NAND2   gate8577  (.A(g1061), .B(II13800), .Z(II13802) ) ;
NAND2   gate8578  (.A(g7683), .B(g1065), .Z(II14244) ) ;
NAND2   gate8579  (.A(g7683), .B(II14244), .Z(II14245) ) ;
NAND2   gate8580  (.A(g1065), .B(II14244), .Z(II14246) ) ;
NAND2   gate8581  (.A(g8147), .B(g1069), .Z(II14472) ) ;
NAND2   gate8582  (.A(g8147), .B(II14472), .Z(II14473) ) ;
NAND2   gate8583  (.A(g1069), .B(II14472), .Z(II14474) ) ;
NOR2    gate8584  (.A(g7658), .B(g7654), .Z(g8073) ) ;
NOR4    gate8585  (.A(g7634), .B(g7628), .C(g7616), .D(g7611), .Z(g8092) ) ;
NAND2   gate8586  (.A(g8660), .B(g1073), .Z(II14837) ) ;
NAND2   gate8587  (.A(g8660), .B(II14837), .Z(II14838) ) ;
NAND2   gate8588  (.A(g1073), .B(II14837), .Z(II14839) ) ;
NOR2    gate8589  (.A(g4146), .B(g8128), .Z(g8644) ) ;
NAND2   gate8590  (.A(g9151), .B(g9148), .Z(II15817) ) ;
NAND2   gate8591  (.A(g9151), .B(II15817), .Z(II15818) ) ;
NAND2   gate8592  (.A(g9148), .B(II15817), .Z(II15819) ) ;
NAND2   gate8593  (.A(II15818), .B(II15819), .Z(g9179) ) ;
NAND2   gate8594  (.A(g9162), .B(g9154), .Z(II15848) ) ;
NAND2   gate8595  (.A(g9162), .B(II15848), .Z(II15849) ) ;
NAND2   gate8596  (.A(g9154), .B(II15848), .Z(II15850) ) ;
NAND2   gate8597  (.A(II15849), .B(II15850), .Z(g9190) ) ;
NAND2   gate8598  (.A(g9168), .B(g9165), .Z(II15855) ) ;
NAND2   gate8599  (.A(g9168), .B(II15855), .Z(II15856) ) ;
NAND2   gate8600  (.A(g9165), .B(II15855), .Z(II15857) ) ;
NAND2   gate8601  (.A(II15856), .B(II15857), .Z(g9191) ) ;
NAND2   gate8602  (.A(g9174), .B(g9171), .Z(II15862) ) ;
NAND2   gate8603  (.A(g9174), .B(II15862), .Z(II15863) ) ;
NAND2   gate8604  (.A(g9171), .B(II15862), .Z(II15864) ) ;
NAND2   gate8605  (.A(II15863), .B(II15864), .Z(g9192) ) ;
NAND2   gate8606  (.A(g9190), .B(g9179), .Z(II15880) ) ;
NAND2   gate8607  (.A(g9190), .B(II15880), .Z(II15881) ) ;
NAND2   gate8608  (.A(g9179), .B(II15880), .Z(II15882) ) ;
NAND2   gate8609  (.A(II15881), .B(II15882), .Z(g9202) ) ;
NAND2   gate8610  (.A(g9192), .B(g9191), .Z(II15887) ) ;
NAND2   gate8611  (.A(g9192), .B(II15887), .Z(II15888) ) ;
NAND2   gate8612  (.A(g9191), .B(II15887), .Z(II15889) ) ;
NAND2   gate8613  (.A(II15888), .B(II15889), .Z(g9203) ) ;
NAND2   gate8614  (.A(g9202), .B(g9203), .Z(II15897) ) ;
NAND2   gate8615  (.A(g9202), .B(II15897), .Z(II15898) ) ;
NAND2   gate8616  (.A(g9203), .B(II15897), .Z(II15899) ) ;
NOR2    gate8617  (.A(g936), .B(g2557), .Z(g3310) ) ;
NOR2    gate8618  (.A(g3310), .B(g3466), .Z(g3885) ) ;
NOR2    gate8619  (.A(g1034), .B(g8128), .Z(g8635) ) ;

endmodule
