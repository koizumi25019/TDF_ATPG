module s5378 (n3065gat, n3066gat, n3067gat, n3068gat, n3069gat
    , n3070gat, n3071gat, n3072gat, n3073gat, n3074gat
    , n3075gat, n3076gat, n3077gat, n3078gat, n3079gat
    , n3080gat, n3081gat, n3082gat, n3083gat, n3084gat
    , n3085gat, n3086gat, n3087gat, n3088gat, n3089gat
    , n3090gat, n3091gat, n3092gat, n3093gat, n3094gat
    , n3095gat, n3097gat, n3098gat, n3099gat, n3100gat
    , CLK
    , n3104gat, n3105gat, n3106gat, n3107gat, n3108gat
    , n3109gat, n3110gat, n3111gat, n3112gat, n3113gat
    , n3114gat, n3115gat, n3116gat, n3117gat, n3118gat
    , n3119gat, n3120gat, n3121gat, n3122gat, n3123gat
    , n3124gat, n3125gat, n3126gat, n3127gat, n3128gat
    , n3129gat, n3130gat, n3131gat, n3132gat, n3133gat
    , n3134gat, n3135gat, n3136gat, n3137gat, n3138gat
    , n3139gat, n3140gat, n3141gat, n3142gat, n3143gat
    , n3144gat, n3145gat, n3146gat, n3147gat, n3148gat
    , n3149gat, n3150gat, n3151gat, n3152gat) ;

input   n3065gat, n3066gat, n3067gat, n3068gat, n3069gat
    , n3070gat, n3071gat, n3072gat, n3073gat, n3074gat
    , n3075gat, n3076gat, n3077gat, n3078gat, n3079gat
    , n3080gat, n3081gat, n3082gat, n3083gat, n3084gat
    , n3085gat, n3086gat, n3087gat, n3088gat, n3089gat
    , n3090gat, n3091gat, n3092gat, n3093gat, n3094gat
    , n3095gat, n3097gat, n3098gat, n3099gat, n3100gat
    , CLK ;

output  n3104gat, n3105gat, n3106gat, n3107gat, n3108gat
    , n3109gat, n3110gat, n3111gat, n3112gat, n3113gat
    , n3114gat, n3115gat, n3116gat, n3117gat, n3118gat
    , n3119gat, n3120gat, n3121gat, n3122gat, n3123gat
    , n3124gat, n3125gat, n3126gat, n3127gat, n3128gat
    , n3129gat, n3130gat, n3131gat, n3132gat, n3133gat
    , n3134gat, n3135gat, n3136gat, n3137gat, n3138gat
    , n3139gat, n3140gat, n3141gat, n3142gat, n3143gat
    , n3144gat, n3145gat, n3146gat, n3147gat, n3148gat
    , n3149gat, n3150gat, n3151gat, n3152gat ;

INV     gate0  (.A(II4654), .Z(n3104gat) ) ;
INV     gate1  (.A(II4657), .Z(n3105gat) ) ;
INV     gate2  (.A(II4660), .Z(n3106gat) ) ;
INV     gate3  (.A(II4663), .Z(n3107gat) ) ;
INV     gate4  (.A(II4666), .Z(n3108gat) ) ;
INV     gate5  (.A(II4669), .Z(n3109gat) ) ;
INV     gate6  (.A(II4672), .Z(n3110gat) ) ;
INV     gate7  (.A(II4675), .Z(n3111gat) ) ;
INV     gate8  (.A(II4678), .Z(n3112gat) ) ;
INV     gate9  (.A(II4681), .Z(n3113gat) ) ;
INV     gate10  (.A(II4684), .Z(n3114gat) ) ;
INV     gate11  (.A(II4687), .Z(n3115gat) ) ;
INV     gate12  (.A(II4690), .Z(n3116gat) ) ;
INV     gate13  (.A(II4693), .Z(n3117gat) ) ;
INV     gate14  (.A(II4696), .Z(n3118gat) ) ;
INV     gate15  (.A(II4699), .Z(n3119gat) ) ;
INV     gate16  (.A(II4702), .Z(n3120gat) ) ;
INV     gate17  (.A(II4705), .Z(n3121gat) ) ;
INV     gate18  (.A(II4708), .Z(n3122gat) ) ;
INV     gate19  (.A(II4711), .Z(n3123gat) ) ;
INV     gate20  (.A(II4714), .Z(n3124gat) ) ;
INV     gate21  (.A(II4717), .Z(n3125gat) ) ;
INV     gate22  (.A(II4720), .Z(n3126gat) ) ;
INV     gate23  (.A(II4723), .Z(n3127gat) ) ;
INV     gate24  (.A(II4726), .Z(n3128gat) ) ;
INV     gate25  (.A(II4729), .Z(n3129gat) ) ;
INV     gate26  (.A(II4732), .Z(n3130gat) ) ;
INV     gate27  (.A(II4735), .Z(n3131gat) ) ;
INV     gate28  (.A(II4738), .Z(n3132gat) ) ;
INV     gate29  (.A(II4741), .Z(n3133gat) ) ;
INV     gate30  (.A(II4744), .Z(n3134gat) ) ;
INV     gate31  (.A(II4747), .Z(n3135gat) ) ;
INV     gate32  (.A(II4750), .Z(n3136gat) ) ;
INV     gate33  (.A(II4753), .Z(n3137gat) ) ;
INV     gate34  (.A(II4756), .Z(n3138gat) ) ;
INV     gate35  (.A(II4759), .Z(n3139gat) ) ;
INV     gate36  (.A(II4762), .Z(n3140gat) ) ;
INV     gate37  (.A(II4765), .Z(n3141gat) ) ;
INV     gate38  (.A(II4768), .Z(n3142gat) ) ;
INV     gate39  (.A(II4771), .Z(n3143gat) ) ;
INV     gate40  (.A(II4774), .Z(n3144gat) ) ;
INV     gate41  (.A(II4777), .Z(n3145gat) ) ;
INV     gate42  (.A(II4780), .Z(n3146gat) ) ;
INV     gate43  (.A(II4783), .Z(n3147gat) ) ;
INV     gate44  (.A(II4786), .Z(n3148gat) ) ;
INV     gate45  (.A(II4789), .Z(n3149gat) ) ;
INV     gate46  (.A(II4792), .Z(n3150gat) ) ;
INV     gate47  (.A(II4795), .Z(n3151gat) ) ;
INV     gate48  (.A(II4798), .Z(n3152gat) ) ;
OR2     gate49  (.A(n648gat), .B(n442gat), .Z(n2897gat) ) ;
DFF     gate50  (.D(n2897gat), .CP(CLK), .Q(n673gat) ) ;
INV     gate51  (.A(II50), .Z(n2782gat) ) ;
DFF     gate52  (.D(n2782gat), .CP(CLK), .Q(n398gat) ) ;
INV     gate53  (.A(II65), .Z(n2790gat) ) ;
DFF     gate54  (.D(n2790gat), .CP(CLK), .Q(n402gat) ) ;
INV     gate55  (.A(II81), .Z(n2670gat) ) ;
DFF     gate56  (.D(n2670gat), .CP(CLK), .Q(n919gat) ) ;
INV     gate57  (.A(II100), .Z(n2793gat) ) ;
DFF     gate58  (.D(n2793gat), .CP(CLK), .Q(n846gat) ) ;
DFF     gate59  (.D(n2782gat), .CP(CLK), .Q(n394gat) ) ;
DFF     gate60  (.D(n2790gat), .CP(CLK), .Q(n703gat) ) ;
DFF     gate61  (.D(n2670gat), .CP(CLK), .Q(n722gat) ) ;
DFF     gate62  (.D(n2793gat), .CP(CLK), .Q(n726gat) ) ;
OR4     gate63  (.A(n749gat), .B(n750gat), .C(n751gat), .D(n752gat), .Z(n748gat) ) ;
DFF     gate64  (.D(n748gat), .CP(CLK), .Q(n2510gat) ) ;
INV     gate65  (.A(II300), .Z(n2732gat) ) ;
DFF     gate66  (.D(n2732gat), .CP(CLK), .Q(n271gat) ) ;
INV     gate67  (.A(II320), .Z(n2776gat) ) ;
DFF     gate68  (.D(n2776gat), .CP(CLK), .Q(n160gat) ) ;
INV     gate69  (.A(II340), .Z(n2735gat) ) ;
DFF     gate70  (.D(n2735gat), .CP(CLK), .Q(n337gat) ) ;
INV     gate71  (.A(II384), .Z(n2673gat) ) ;
DFF     gate72  (.D(n2673gat), .CP(CLK), .Q(n842gat) ) ;
INV     gate73  (.A(II426), .Z(n2779gat) ) ;
DFF     gate74  (.D(n2779gat), .CP(CLK), .Q(n341gat) ) ;
OR4     gate75  (.A(n44gat), .B(n45gat), .C(n46gat), .D(n47gat), .Z(n43gat) ) ;
DFF     gate76  (.D(n43gat), .CP(CLK), .Q(n2522gat) ) ;
NOR2    gate77  (.A(n1448gat), .B(n1446gat), .Z(n1620gat) ) ;
DFF     gate78  (.D(n1620gat), .CP(CLK), .Q(n2472gat) ) ;
INV     gate79  (.A(n2472gat), .Z(n2470gat) ) ;
DFF     gate80  (.D(n2470gat), .CP(CLK), .Q(n2319gat) ) ;
NOR2    gate81  (.A(n2729gat), .B(n2317gat), .Z(n1827gat) ) ;
DFF     gate82  (.D(n1827gat), .CP(CLK), .Q(n1821gat) ) ;
DFF     gate83  (.D(n1827gat), .CP(CLK), .Q(n1825gat) ) ;
INV     gate84  (.A(n1817gat), .Z(n1816gat) ) ;
DFF     gate85  (.D(n1816gat), .CP(CLK), .Q(n2029gat) ) ;
INV     gate86  (.A(n2029gat), .Z(n2027gat) ) ;
DFF     gate87  (.D(n2027gat), .CP(CLK), .Q(n1829gat) ) ;
DFF     gate88  (.D(n2732gat), .CP(CLK), .Q(n283gat) ) ;
DFF     gate89  (.D(n2776gat), .CP(CLK), .Q(n165gat) ) ;
DFF     gate90  (.D(n2735gat), .CP(CLK), .Q(n279gat) ) ;
DFF     gate91  (.D(n2673gat), .CP(CLK), .Q(n1026gat) ) ;
DFF     gate92  (.D(n2779gat), .CP(CLK), .Q(n275gat) ) ;
OR4     gate93  (.A(n56gat), .B(n57gat), .C(n58gat), .D(n59gat), .Z(n55gat) ) ;
DFF     gate94  (.D(n55gat), .CP(CLK), .Q(n2476gat) ) ;
OR2     gate95  (.A(n768gat), .B(n655gat), .Z(n2914gat) ) ;
DFF     gate96  (.D(n2914gat), .CP(CLK), .Q(n1068gat) ) ;
OR2     gate97  (.A(n963gat), .B(n868gat), .Z(n2928gat) ) ;
DFF     gate98  (.D(n2928gat), .CP(CLK), .Q(n957gat) ) ;
OR2     gate99  (.A(n962gat), .B(n959gat), .Z(n2927gat) ) ;
DFF     gate100  (.D(n2927gat), .CP(CLK), .Q(n861gat) ) ;
OR2     gate101  (.A(n647gat), .B(n441gat), .Z(n2896gat) ) ;
DFF     gate102  (.D(n2896gat), .CP(CLK), .Q(n1294gat) ) ;
OR2     gate103  (.A(n967gat), .B(n792gat), .Z(n2922gat) ) ;
DFF     gate104  (.D(n2922gat), .CP(CLK), .Q(n1241gat) ) ;
DFF     gate105  (.D(n2897gat), .CP(CLK), .Q(n1298gat) ) ;
OR2     gate106  (.A(n443gat), .B(n439gat), .Z(n2894gat) ) ;
DFF     gate107  (.D(n2894gat), .CP(CLK), .Q(n865gat) ) ;
OR2     gate108  (.A(n966gat), .B(n790gat), .Z(n2921gat) ) ;
DFF     gate109  (.D(n2921gat), .CP(CLK), .Q(n1080gat) ) ;
OR2     gate110  (.A(n444gat), .B(n440gat), .Z(n2895gat) ) ;
DFF     gate111  (.D(n2895gat), .CP(CLK), .Q(n1148gat) ) ;
OR4     gate112  (.A(n934gat), .B(n935gat), .C(n936gat), .D(n937gat), .Z(n933gat) ) ;
DFF     gate113  (.D(n933gat), .CP(CLK), .Q(n2468gat) ) ;
DFF     gate114  (.D(n2790gat), .CP(CLK), .Q(n618gat) ) ;
DFF     gate115  (.D(n2782gat), .CP(CLK), .Q(n491gat) ) ;
DFF     gate116  (.D(n2793gat), .CP(CLK), .Q(n622gat) ) ;
DFF     gate117  (.D(n2670gat), .CP(CLK), .Q(n626gat) ) ;
INV     gate118  (.A(II3914), .Z(n3064gat) ) ;
DFF     gate119  (.D(n3064gat), .CP(CLK), .Q(n834gat) ) ;
INV     gate120  (.A(II3703), .Z(n3055gat) ) ;
DFF     gate121  (.D(n3055gat), .CP(CLK), .Q(n707gat) ) ;
INV     gate122  (.A(II3891), .Z(n3063gat) ) ;
DFF     gate123  (.D(n3063gat), .CP(CLK), .Q(n838gat) ) ;
INV     gate124  (.A(II3876), .Z(n3062gat) ) ;
DFF     gate125  (.D(n3062gat), .CP(CLK), .Q(n830gat) ) ;
INV     gate126  (.A(II3713), .Z(n3056gat) ) ;
DFF     gate127  (.D(n3056gat), .CP(CLK), .Q(n614gat) ) ;
OR4     gate128  (.A(n505gat), .B(n506gat), .C(n507gat), .D(n508gat), .Z(n504gat) ) ;
DFF     gate129  (.D(n504gat), .CP(CLK), .Q(n2526gat) ) ;
OR2     gate130  (.A(n767gat), .B(n653gat), .Z(n2913gat) ) ;
DFF     gate131  (.D(n2913gat), .CP(CLK), .Q(n680gat) ) ;
OR2     gate132  (.A(n867gat), .B(n771gat), .Z(n2920gat) ) ;
DFF     gate133  (.D(n2920gat), .CP(CLK), .Q(n816gat) ) ;
OR2     gate134  (.A(n964gat), .B(n961gat), .Z(n2905gat) ) ;
DFF     gate135  (.D(n2905gat), .CP(CLK), .Q(n580gat) ) ;
INV     gate136  (.A(II3754), .Z(n3057gat) ) ;
DFF     gate137  (.D(n3057gat), .CP(CLK), .Q(n824gat) ) ;
INV     gate138  (.A(II3801), .Z(n3059gat) ) ;
DFF     gate139  (.D(n3059gat), .CP(CLK), .Q(n820gat) ) ;
INV     gate140  (.A(II3765), .Z(n3058gat) ) ;
DFF     gate141  (.D(n3058gat), .CP(CLK), .Q(n883gat) ) ;
OR2     gate142  (.A(n447gat), .B(n445gat), .Z(n2898gat) ) ;
DFF     gate143  (.D(n2898gat), .CP(CLK), .Q(n584gat) ) ;
INV     gate144  (.A(II3817), .Z(n3060gat) ) ;
DFF     gate145  (.D(n3060gat), .CP(CLK), .Q(n684gat) ) ;
INV     gate146  (.A(II3841), .Z(n3061gat) ) ;
DFF     gate147  (.D(n3061gat), .CP(CLK), .Q(n699gat) ) ;
OR4     gate148  (.A(n568gat), .B(n569gat), .C(n570gat), .D(n571gat), .Z(n567gat) ) ;
DFF     gate149  (.D(n567gat), .CP(CLK), .Q(n2464gat) ) ;
INV     gate150  (.A(II3530), .Z(n3048gat) ) ;
DFF     gate151  (.D(n3048gat), .CP(CLK), .Q(n2399gat) ) ;
INV     gate152  (.A(II3539), .Z(n3049gat) ) ;
DFF     gate153  (.D(n3049gat), .CP(CLK), .Q(n2343gat) ) ;
INV     gate154  (.A(II3558), .Z(n3051gat) ) ;
DFF     gate155  (.D(n3051gat), .CP(CLK), .Q(n2203gat) ) ;
INV     gate156  (.A(II3520), .Z(n3047gat) ) ;
DFF     gate157  (.D(n3047gat), .CP(CLK), .Q(n2562gat) ) ;
INV     gate158  (.A(II3549), .Z(n3050gat) ) ;
DFF     gate159  (.D(n3050gat), .CP(CLK), .Q(n2207gat) ) ;
INV     gate160  (.A(II3472), .Z(n3040gat) ) ;
DFF     gate161  (.D(n3040gat), .CP(CLK), .Q(n2626gat) ) ;
INV     gate162  (.A(II3504), .Z(n3044gat) ) ;
DFF     gate163  (.D(n3044gat), .CP(CLK), .Q(n2490gat) ) ;
INV     gate164  (.A(II3491), .Z(n3042gat) ) ;
DFF     gate165  (.D(n3042gat), .CP(CLK), .Q(n2622gat) ) ;
INV     gate166  (.A(II3457), .Z(n3037gat) ) ;
DFF     gate167  (.D(n3037gat), .CP(CLK), .Q(n2630gat) ) ;
INV     gate168  (.A(II3483), .Z(n3041gat) ) ;
DFF     gate169  (.D(n3041gat), .CP(CLK), .Q(n2543gat) ) ;
NOR2    gate170  (.A(n3020gat), .B(n270gat), .Z(n1606gat) ) ;
DFF     gate171  (.D(n1606gat), .CP(CLK), .Q(n2102gat) ) ;
INV     gate172  (.A(II3610), .Z(n3052gat) ) ;
DFF     gate173  (.D(n3052gat), .CP(CLK), .Q(n1880gat) ) ;
NOR2    gate174  (.A(n1698gat), .B(n1543gat), .Z(n1610gat) ) ;
DFF     gate175  (.D(n1610gat), .CP(CLK), .Q(n1763gat) ) ;
INV     gate176  (.A(n1673gat), .Z(n1858gat) ) ;
DFF     gate177  (.D(n1858gat), .CP(CLK), .Q(n2155gat) ) ;
OR2     gate178  (.A(n769gat), .B(n759gat), .Z(n2918gat) ) ;
DFF     gate179  (.D(n2918gat), .CP(CLK), .Q(n1035gat) ) ;
OR2     gate180  (.A(n1076gat), .B(n1075gat), .Z(n2952gat) ) ;
DFF     gate181  (.D(n2952gat), .CP(CLK), .Q(n1121gat) ) ;
OR2     gate182  (.A(n766gat), .B(n760gat), .Z(n2919gat) ) ;
DFF     gate183  (.D(n2919gat), .CP(CLK), .Q(n1072gat) ) ;
OR2     gate184  (.A(n645gat), .B(n644gat), .Z(n2910gat) ) ;
DFF     gate185  (.D(n2910gat), .CP(CLK), .Q(n1282gat) ) ;
OR2     gate186  (.A(n646gat), .B(n641gat), .Z(n2907gat) ) ;
DFF     gate187  (.D(n2907gat), .CP(CLK), .Q(n1226gat) ) ;
OR2     gate188  (.A(n761gat), .B(n651gat), .Z(n2911gat) ) ;
DFF     gate189  (.D(n2911gat), .CP(CLK), .Q(n931gat) ) ;
OR2     gate190  (.A(n762gat), .B(n652gat), .Z(n2912gat) ) ;
DFF     gate191  (.D(n2912gat), .CP(CLK), .Q(n1135gat) ) ;
OR2     gate192  (.A(n765gat), .B(n643gat), .Z(n2909gat) ) ;
DFF     gate193  (.D(n2909gat), .CP(CLK), .Q(n1045gat) ) ;
OR2     gate194  (.A(n763gat), .B(n642gat), .Z(n2908gat) ) ;
DFF     gate195  (.D(n2908gat), .CP(CLK), .Q(n1197gat) ) ;
OR2     gate196  (.A(n1287gat), .B(n1285gat), .Z(n2971gat) ) ;
DFF     gate197  (.D(n2971gat), .CP(CLK), .Q(n2518gat) ) ;
OR3     gate198  (.A(n793gat), .B(n664gat), .C(n556gat), .Z(n2904gat) ) ;
DFF     gate199  (.D(n2904gat), .CP(CLK), .Q(n667gat) ) ;
OR3     gate200  (.A(n795gat), .B(n656gat), .C(n368gat), .Z(n2891gat) ) ;
DFF     gate201  (.D(n2891gat), .CP(CLK), .Q(n659gat) ) ;
OR3     gate202  (.A(n794gat), .B(n773gat), .C(n662gat), .Z(n2903gat) ) ;
DFF     gate203  (.D(n2903gat), .CP(CLK), .Q(n553gat) ) ;
OR3     gate204  (.A(n965gat), .B(n960gat), .C(n661gat), .Z(n2915gat) ) ;
DFF     gate205  (.D(n2915gat), .CP(CLK), .Q(n777gat) ) ;
OR3     gate206  (.A(n558gat), .B(n555gat), .C(n450gat), .Z(n2901gat) ) ;
DFF     gate207  (.D(n2901gat), .CP(CLK), .Q(n561gat) ) ;
OR3     gate208  (.A(n654gat), .B(n557gat), .C(n371gat), .Z(n2890gat) ) ;
DFF     gate209  (.D(n2890gat), .CP(CLK), .Q(n366gat) ) ;
OR3     gate210  (.A(n663gat), .B(n649gat), .C(n449gat), .Z(n2888gat) ) ;
DFF     gate211  (.D(n2888gat), .CP(CLK), .Q(n322gat) ) ;
OR3     gate212  (.A(n791gat), .B(n650gat), .C(n370gat), .Z(n2887gat) ) ;
DFF     gate213  (.D(n2887gat), .CP(CLK), .Q(n318gat) ) ;
OR3     gate214  (.A(n774gat), .B(n764gat), .C(n369gat), .Z(n2886gat) ) ;
DFF     gate215  (.D(n2886gat), .CP(CLK), .Q(n314gat) ) ;
OR2     gate216  (.A(n2460gat), .B(n2423gat), .Z(n3010gat) ) ;
DFF     gate217  (.D(n3010gat), .CP(CLK), .Q(n2599gat) ) ;
OR2     gate218  (.A(n2596gat), .B(n2595gat), .Z(n3016gat) ) ;
DFF     gate219  (.D(n3016gat), .CP(CLK), .Q(n2588gat) ) ;
INV     gate220  (.A(II3660), .Z(n3054gat) ) ;
DFF     gate221  (.D(n3054gat), .CP(CLK), .Q(n2640gat) ) ;
OR2     gate222  (.A(n2580gat), .B(n2581gat), .Z(n2579gat) ) ;
DFF     gate223  (.D(n2579gat), .CP(CLK), .Q(n2658gat) ) ;
INV     gate224  (.A(II3436), .Z(n3036gat) ) ;
DFF     gate225  (.D(n3036gat), .CP(CLK), .Q(n2495gat) ) ;
INV     gate226  (.A(II3401), .Z(n3034gat) ) ;
DFF     gate227  (.D(n3034gat), .CP(CLK), .Q(n2390gat) ) ;
INV     gate228  (.A(II3387), .Z(n3031gat) ) ;
DFF     gate229  (.D(n3031gat), .CP(CLK), .Q(n2270gat) ) ;
INV     gate230  (.A(II3412), .Z(n3035gat) ) ;
DFF     gate231  (.D(n3035gat), .CP(CLK), .Q(n2339gat) ) ;
OR2     gate232  (.A(n2647gat), .B(n2648gat), .Z(n2646gat) ) ;
DFF     gate233  (.D(n2646gat), .CP(CLK), .Q(n2502gat) ) ;
INV     gate234  (.A(II3635), .Z(n3053gat) ) ;
DFF     gate235  (.D(n3053gat), .CP(CLK), .Q(n2634gat) ) ;
OR2     gate236  (.A(n2614gat), .B(n2615gat), .Z(n2613gat) ) ;
DFF     gate237  (.D(n2613gat), .CP(CLK), .Q(n2506gat) ) ;
NOR2    gate238  (.A(n3021gat), .B(n1628gat), .Z(n1625gat) ) ;
DFF     gate239  (.D(n1625gat), .CP(CLK), .Q(n1834gat) ) ;
NOR2    gate240  (.A(n1627gat), .B(n3022gat), .Z(n1626gat) ) ;
DFF     gate241  (.D(n1626gat), .CP(CLK), .Q(n1767gat) ) ;
INV     gate242  (.A(n1831gat), .Z(n1603gat) ) ;
DFF     gate243  (.D(n1603gat), .CP(CLK), .Q(n2084gat) ) ;
INV     gate244  (.A(n2543gat), .Z(n2541gat) ) ;
DFF     gate245  (.D(n2541gat), .CP(CLK), .Q(n2143gat) ) ;
INV     gate246  (.A(n2621gat), .Z(n2557gat) ) ;
DFF     gate247  (.D(n2557gat), .CP(CLK), .Q(n2061gat) ) ;
INV     gate248  (.A(n2489gat), .Z(n2487gat) ) ;
DFF     gate249  (.D(n2487gat), .CP(CLK), .Q(n2139gat) ) ;
INV     gate250  (.A(n2625gat), .Z(n2532gat) ) ;
DFF     gate251  (.D(n2532gat), .CP(CLK), .Q(n1899gat) ) ;
INV     gate252  (.A(n2630gat), .Z(n2628gat) ) ;
DFF     gate253  (.D(n2628gat), .CP(CLK), .Q(n1850gat) ) ;
INV     gate254  (.A(n2399gat), .Z(n2397gat) ) ;
DFF     gate255  (.D(n2397gat), .CP(CLK), .Q(n2403gat) ) ;
INV     gate256  (.A(n2343gat), .Z(n2341gat) ) ;
DFF     gate257  (.D(n2341gat), .CP(CLK), .Q(n2394gat) ) ;
INV     gate258  (.A(n2562gat), .Z(n2560gat) ) ;
DFF     gate259  (.D(n2560gat), .CP(CLK), .Q(n2440gat) ) ;
INV     gate260  (.A(n2207gat), .Z(n2205gat) ) ;
DFF     gate261  (.D(n2205gat), .CP(CLK), .Q(n2407gat) ) ;
INV     gate262  (.A(n2203gat), .Z(n2201gat) ) ;
DFF     gate263  (.D(n2201gat), .CP(CLK), .Q(n2347gat) ) ;
NOR2    gate264  (.A(n1792gat), .B(n1735gat), .Z(n1793gat) ) ;
DFF     gate265  (.D(n1793gat), .CP(CLK), .Q(n1389gat) ) ;
INV     gate266  (.A(n1780gat), .Z(n1781gat) ) ;
DFF     gate267  (.D(n1781gat), .CP(CLK), .Q(n2021gat) ) ;
NOR2    gate268  (.A(n1551gat), .B(n1517gat), .Z(n1516gat) ) ;
DFF     gate269  (.D(n1516gat), .CP(CLK), .Q(n1394gat) ) ;
INV     gate270  (.A(n1394gat), .Z(n1392gat) ) ;
DFF     gate271  (.D(n1392gat), .CP(CLK), .Q(n1496gat) ) ;
INV     gate272  (.A(n1604gat), .Z(n1685gat) ) ;
DFF     gate273  (.D(n1685gat), .CP(CLK), .Q(n2091gat) ) ;
NOR2    gate274  (.A(n1735gat), .B(n1552gat), .Z(n1565gat) ) ;
DFF     gate275  (.D(n1565gat), .CP(CLK), .Q(n1332gat) ) ;
INV     gate276  (.A(n1332gat), .Z(n1330gat) ) ;
DFF     gate277  (.D(n1330gat), .CP(CLK), .Q(n1740gat) ) ;
INV     gate278  (.A(n1690gat), .Z(n1945gat) ) ;
DFF     gate279  (.D(n1945gat), .CP(CLK), .Q(n2179gat) ) ;
INV     gate280  (.A(n2270gat), .Z(n2268gat) ) ;
DFF     gate281  (.D(n2268gat), .CP(CLK), .Q(n2190gat) ) ;
INV     gate282  (.A(n2339gat), .Z(n2337gat) ) ;
DFF     gate283  (.D(n2337gat), .CP(CLK), .Q(n2135gat) ) ;
INV     gate284  (.A(n2390gat), .Z(n2388gat) ) ;
DFF     gate285  (.D(n2388gat), .CP(CLK), .Q(n2262gat) ) ;
INV     gate286  (.A(n1695gat), .Z(n1836gat) ) ;
DFF     gate287  (.D(n1836gat), .CP(CLK), .Q(n2182gat) ) ;
OR2     gate288  (.A(n2079gat), .B(n2073gat), .Z(n2983gat) ) ;
DFF     gate289  (.D(n2983gat), .CP(CLK), .Q(n1433gat) ) ;
INV     gate290  (.A(n1433gat), .Z(n1431gat) ) ;
DFF     gate291  (.D(n1431gat), .CP(CLK), .Q(n1316gat) ) ;
INV     gate292  (.A(n1316gat), .Z(n1314gat) ) ;
DFF     gate293  (.D(n1314gat), .CP(CLK), .Q(n1363gat) ) ;
INV     gate294  (.A(n1363gat), .Z(n1361gat) ) ;
DFF     gate295  (.D(n1361gat), .CP(CLK), .Q(n1312gat) ) ;
NOR2    gate296  (.A(n1707gat), .B(n1698gat), .Z(n1696gat) ) ;
DFF     gate297  (.D(n1696gat), .CP(CLK), .Q(n1775gat) ) ;
NOR3    gate298  (.A(n2016gat), .B(n2664gat), .C(n2004gat), .Z(n2009gat) ) ;
DFF     gate299  (.D(n2009gat), .CP(CLK), .Q(n1871gat) ) ;
INV     gate300  (.A(n1775gat), .Z(n1773gat) ) ;
DFF     gate301  (.D(n1773gat), .CP(CLK), .Q(n2592gat) ) ;
NOR2    gate302  (.A(n1584gat), .B(n1718gat), .Z(n1636gat) ) ;
DFF     gate303  (.D(n1636gat), .CP(CLK), .Q(n1508gat) ) ;
INV     gate304  (.A(II3179), .Z(n1712gat) ) ;
DFF     gate305  (.D(n1712gat), .CP(CLK), .Q(n1678gat) ) ;
OR2     gate306  (.A(n2000gat), .B(n1999gat), .Z(n3000gat) ) ;
DFF     gate307  (.D(n3000gat), .CP(CLK), .Q(n2309gat) ) ;
INV     gate308  (.A(n2309gat), .Z(n2307gat) ) ;
DFF     gate309  (.D(n2307gat), .CP(CLK), .Q(n2450gat) ) ;
INV     gate310  (.A(n2662gat), .Z(n2661gat) ) ;
DFF     gate311  (.D(n2661gat), .CP(CLK), .Q(n2446gat) ) ;
INV     gate312  (.A(n204gat), .Z(n827gat) ) ;
DFF     gate313  (.D(n827gat), .CP(CLK), .Q(n2095gat) ) ;
INV     gate314  (.A(n2095gat), .Z(n2093gat) ) ;
DFF     gate315  (.D(n2093gat), .CP(CLK), .Q(n2176gat) ) ;
INV     gate316  (.A(n2176gat), .Z(n2174gat) ) ;
DFF     gate317  (.D(n2174gat), .CP(CLK), .Q(n2169gat) ) ;
NOR4    gate318  (.A(n1790gat), .B(n1310gat), .C(n2664gat), .D(n2168gat), .Z(n2163gat) ) ;
DFF     gate319  (.D(n2163gat), .CP(CLK), .Q(n2454gat) ) ;
INV     gate320  (.A(n1694gat), .Z(n1777gat) ) ;
DFF     gate321  (.D(n1777gat), .CP(CLK), .Q(n2040gat) ) ;
NOR3    gate322  (.A(n2039gat), .B(n1774gat), .C(n1315gat), .Z(n2015gat) ) ;
DFF     gate323  (.D(n2015gat), .CP(CLK), .Q(n2044gat) ) ;
INV     gate324  (.A(n2044gat), .Z(n2042gat) ) ;
DFF     gate325  (.D(n2042gat), .CP(CLK), .Q(n2037gat) ) ;
NOR2    gate326  (.A(n1790gat), .B(n2016gat), .Z(n2017gat) ) ;
DFF     gate327  (.D(n2017gat), .CP(CLK), .Q(n2025gat) ) ;
INV     gate328  (.A(n2025gat), .Z(n2023gat) ) ;
DFF     gate329  (.D(n2023gat), .CP(CLK), .Q(n2099gat) ) ;
INV     gate330  (.A(n2495gat), .Z(n2493gat) ) ;
DFF     gate331  (.D(n2493gat), .CP(CLK), .Q(n2266gat) ) ;
INV     gate332  (.A(n2037gat), .Z(n2035gat) ) ;
DFF     gate333  (.D(n2035gat), .CP(CLK), .Q(n2033gat) ) ;
INV     gate334  (.A(n2033gat), .Z(n2031gat) ) ;
DFF     gate335  (.D(n2031gat), .CP(CLK), .Q(n2110gat) ) ;
INV     gate336  (.A(n2110gat), .Z(n2108gat) ) ;
DFF     gate337  (.D(n2108gat), .CP(CLK), .Q(n2125gat) ) ;
INV     gate338  (.A(n2125gat), .Z(n2123gat) ) ;
DFF     gate339  (.D(n2123gat), .CP(CLK), .Q(n2121gat) ) ;
INV     gate340  (.A(n2121gat), .Z(n2119gat) ) ;
DFF     gate341  (.D(n2119gat), .CP(CLK), .Q(n2117gat) ) ;
INV     gate342  (.A(n2634gat), .Z(n2632gat) ) ;
DFF     gate343  (.D(n2632gat), .CP(CLK), .Q(n1975gat) ) ;
INV     gate344  (.A(n2640gat), .Z(n2638gat) ) ;
DFF     gate345  (.D(n2638gat), .CP(CLK), .Q(n2644gat) ) ;
INV     gate346  (.A(n614gat), .Z(n612gat) ) ;
DFF     gate347  (.D(n612gat), .CP(CLK), .Q(n156gat) ) ;
INV     gate348  (.A(n707gat), .Z(n705gat) ) ;
DFF     gate349  (.D(n705gat), .CP(CLK), .Q(n152gat) ) ;
INV     gate350  (.A(n824gat), .Z(n822gat) ) ;
DFF     gate351  (.D(n822gat), .CP(CLK), .Q(n331gat) ) ;
INV     gate352  (.A(n883gat), .Z(n881gat) ) ;
DFF     gate353  (.D(n881gat), .CP(CLK), .Q(n388gat) ) ;
INV     gate354  (.A(n820gat), .Z(n818gat) ) ;
DFF     gate355  (.D(n818gat), .CP(CLK), .Q(n463gat) ) ;
INV     gate356  (.A(n684gat), .Z(n682gat) ) ;
DFF     gate357  (.D(n682gat), .CP(CLK), .Q(n327gat) ) ;
INV     gate358  (.A(n699gat), .Z(n697gat) ) ;
DFF     gate359  (.D(n697gat), .CP(CLK), .Q(n384gat) ) ;
INV     gate360  (.A(n838gat), .Z(n836gat) ) ;
DFF     gate361  (.D(n836gat), .CP(CLK), .Q(n256gat) ) ;
INV     gate362  (.A(n830gat), .Z(n828gat) ) ;
DFF     gate363  (.D(n828gat), .CP(CLK), .Q(n470gat) ) ;
INV     gate364  (.A(n834gat), .Z(n832gat) ) ;
DFF     gate365  (.D(n832gat), .CP(CLK), .Q(n148gat) ) ;
INV     gate366  (.A(n2592gat), .Z(n2590gat) ) ;
DFF     gate367  (.D(n2590gat), .CP(CLK), .Q(n2458gat) ) ;
INV     gate368  (.A(n2458gat), .Z(n2456gat) ) ;
DFF     gate369  (.D(n2456gat), .CP(CLK), .Q(n2514gat) ) ;
NOR2    gate370  (.A(n1544gat), .B(n1698gat), .Z(n1613gat) ) ;
DFF     gate371  (.D(n1613gat), .CP(CLK), .Q(n1771gat) ) ;
NOR2    gate372  (.A(n1513gat), .B(n2442gat), .Z(n1391gat) ) ;
DFF     gate373  (.D(n1391gat), .CP(CLK), .Q(n1336gat) ) ;
NOR2    gate374  (.A(n1790gat), .B(n1635gat), .Z(n1927gat) ) ;
DFF     gate375  (.D(n1927gat), .CP(CLK), .Q(n1748gat) ) ;
INV     gate376  (.A(II2935), .Z(n1713gat) ) ;
DFF     gate377  (.D(n1713gat), .CP(CLK), .Q(n1675gat) ) ;
INV     gate378  (.A(II2926), .Z(n1717gat) ) ;
DFF     gate379  (.D(n1717gat), .CP(CLK), .Q(n1807gat) ) ;
NOR2    gate380  (.A(n1634gat), .B(n1735gat), .Z(n1567gat) ) ;
DFF     gate381  (.D(n1567gat), .CP(CLK), .Q(n1340gat) ) ;
NOR4    gate382  (.A(n1584gat), .B(n1719gat), .C(n1790gat), .D(n1576gat), .Z(n1564gat) ) ;
DFF     gate383  (.D(n1564gat), .CP(CLK), .Q(n1456gat) ) ;
INV     gate384  (.A(II4145), .Z(n1632gat) ) ;
DFF     gate385  (.D(n1632gat), .CP(CLK), .Q(n1525gat) ) ;
NOR2    gate386  (.A(n1859gat), .B(n1919gat), .Z(n1915gat) ) ;
DFF     gate387  (.D(n1915gat), .CP(CLK), .Q(n1462gat) ) ;
NOR2    gate388  (.A(n1635gat), .B(n1919gat), .Z(n1800gat) ) ;
DFF     gate389  (.D(n1800gat), .CP(CLK), .Q(n1596gat) ) ;
NOR2    gate390  (.A(n1551gat), .B(n1310gat), .Z(n1593gat) ) ;
DFF     gate391  (.D(n1593gat), .CP(CLK), .Q(n1588gat) ) ;
INV     gate392  (.A(n3088gat), .Z(II1) ) ;
INV     gate393  (.A(II1), .Z(n2717gat) ) ;
INV     gate394  (.A(n2717gat), .Z(n2715gat) ) ;
INV     gate395  (.A(n3087gat), .Z(II5) ) ;
INV     gate396  (.A(II5), .Z(n2725gat) ) ;
INV     gate397  (.A(n2725gat), .Z(n2723gat) ) ;
NOR2    gate398  (.A(n2715gat), .B(n2723gat), .Z(n421gat) ) ;
INV     gate399  (.A(n421gat), .Z(n296gat) ) ;
INV     gate400  (.A(n3093gat), .Z(II11) ) ;
INV     gate401  (.A(II11), .Z(n2768gat) ) ;
INV     gate402  (.A(n2768gat), .Z(II14) ) ;
INV     gate403  (.A(II14), .Z(n2767gat) ) ;
INV     gate404  (.A(n2767gat), .Z(n373gat) ) ;
INV     gate405  (.A(n3072gat), .Z(II18) ) ;
INV     gate406  (.A(II18), .Z(n2671gat) ) ;
INV     gate407  (.A(n2671gat), .Z(n2669gat) ) ;
INV     gate408  (.A(n3081gat), .Z(II23) ) ;
INV     gate409  (.A(II23), .Z(n2845gat) ) ;
INV     gate410  (.A(n2845gat), .Z(n2844gat) ) ;
INV     gate411  (.A(n3095gat), .Z(II27) ) ;
INV     gate412  (.A(II27), .Z(n2668gat) ) ;
INV     gate413  (.A(n2668gat), .Z(II30) ) ;
INV     gate414  (.A(II30), .Z(n2667gat) ) ;
INV     gate415  (.A(n2667gat), .Z(n856gat) ) ;
INV     gate416  (.A(n673gat), .Z(II44) ) ;
INV     gate417  (.A(II44), .Z(n672gat) ) ;
INV     gate418  (.A(n3069gat), .Z(II47) ) ;
INV     gate419  (.A(II47), .Z(n2783gat) ) ;
INV     gate420  (.A(n2783gat), .Z(II50) ) ;
INV     gate421  (.A(n398gat), .Z(n396gat) ) ;
INV     gate422  (.A(n3070gat), .Z(II62) ) ;
INV     gate423  (.A(II62), .Z(n2791gat) ) ;
INV     gate424  (.A(n2791gat), .Z(II65) ) ;
INV     gate425  (.A(n402gat), .Z(II76) ) ;
INV     gate426  (.A(II76), .Z(n401gat) ) ;
NOR2    gate427  (.A(n396gat), .B(n401gat), .Z(n1499gat) ) ;
INV     gate428  (.A(n1499gat), .Z(n1645gat) ) ;
INV     gate429  (.A(n2671gat), .Z(II81) ) ;
INV     gate430  (.A(n919gat), .Z(II92) ) ;
INV     gate431  (.A(II92), .Z(n918gat) ) ;
NOR2    gate432  (.A(n918gat), .B(n396gat), .Z(n1616gat) ) ;
INV     gate433  (.A(n1616gat), .Z(n1553gat) ) ;
INV     gate434  (.A(n3071gat), .Z(II97) ) ;
INV     gate435  (.A(II97), .Z(n2794gat) ) ;
INV     gate436  (.A(n2794gat), .Z(II100) ) ;
INV     gate437  (.A(n846gat), .Z(II111) ) ;
INV     gate438  (.A(II111), .Z(n845gat) ) ;
NOR2    gate439  (.A(n396gat), .B(n845gat), .Z(n1614gat) ) ;
INV     gate440  (.A(n1614gat), .Z(n1559gat) ) ;
NOR3    gate441  (.A(n1645gat), .B(n1553gat), .C(n1559gat), .Z(n1641gat) ) ;
INV     gate442  (.A(n1641gat), .Z(n1643gat) ) ;
NOR3    gate443  (.A(n1559gat), .B(n1616gat), .C(n1645gat), .Z(n1642gat) ) ;
INV     gate444  (.A(n1642gat), .Z(n1651gat) ) ;
NOR3    gate445  (.A(n1614gat), .B(n1645gat), .C(n1616gat), .Z(n1556gat) ) ;
INV     gate446  (.A(n1556gat), .Z(n1562gat) ) ;
NOR3    gate447  (.A(n1553gat), .B(n1645gat), .C(n1614gat), .Z(n1557gat) ) ;
INV     gate448  (.A(n1557gat), .Z(n1560gat) ) ;
NOR3    gate449  (.A(n1499gat), .B(n1559gat), .C(n1553gat), .Z(n1639gat) ) ;
INV     gate450  (.A(n1639gat), .Z(n1640gat) ) ;
NOR4    gate451  (.A(n1614gat), .B(n1616gat), .C(n1499gat), .D(n396gat), .Z(n1605gat) ) ;
INV     gate452  (.A(n1605gat), .Z(n1566gat) ) ;
NOR3    gate453  (.A(n1616gat), .B(n1559gat), .C(n1499gat), .Z(n1555gat) ) ;
INV     gate454  (.A(n1555gat), .Z(n1554gat) ) ;
NOR3    gate455  (.A(n1614gat), .B(n1553gat), .C(n1499gat), .Z(n1558gat) ) ;
INV     gate456  (.A(n1558gat), .Z(n1722gat) ) ;
INV     gate457  (.A(n394gat), .Z(n392gat) ) ;
INV     gate458  (.A(n703gat), .Z(II149) ) ;
INV     gate459  (.A(II149), .Z(n702gat) ) ;
NOR2    gate460  (.A(n392gat), .B(n702gat), .Z(n1256gat) ) ;
INV     gate461  (.A(n1256gat), .Z(n1319gat) ) ;
INV     gate462  (.A(n722gat), .Z(n720gat) ) ;
INV     gate463  (.A(n726gat), .Z(II171) ) ;
INV     gate464  (.A(II171), .Z(n725gat) ) ;
NOR2    gate465  (.A(n720gat), .B(n725gat), .Z(n1117gat) ) ;
INV     gate466  (.A(n1117gat), .Z(n1447gat) ) ;
NOR2    gate467  (.A(n1319gat), .B(n1447gat), .Z(n1618gat) ) ;
INV     gate468  (.A(n1618gat), .Z(n1627gat) ) ;
INV     gate469  (.A(n722gat), .Z(II178) ) ;
INV     gate470  (.A(II178), .Z(n721gat) ) ;
NOR2    gate471  (.A(n725gat), .B(n721gat), .Z(n1114gat) ) ;
INV     gate472  (.A(n1114gat), .Z(n1380gat) ) ;
NOR2    gate473  (.A(n1319gat), .B(n1380gat), .Z(n1621gat) ) ;
INV     gate474  (.A(n1621gat), .Z(n1628gat) ) ;
INV     gate475  (.A(n703gat), .Z(n701gat) ) ;
NOR2    gate476  (.A(n392gat), .B(n701gat), .Z(n1318gat) ) ;
INV     gate477  (.A(n1318gat), .Z(n1446gat) ) ;
NOR2    gate478  (.A(n1447gat), .B(n1446gat), .Z(n1619gat) ) ;
INV     gate479  (.A(n1619gat), .Z(n1705gat) ) ;
NOR2    gate480  (.A(n1380gat), .B(n1446gat), .Z(n1622gat) ) ;
INV     gate481  (.A(n1622gat), .Z(n1706gat) ) ;
INV     gate482  (.A(n3083gat), .Z(II192) ) ;
INV     gate483  (.A(II192), .Z(n2856gat) ) ;
INV     gate484  (.A(n2856gat), .Z(n2854gat) ) ;
INV     gate485  (.A(n2854gat), .Z(II196) ) ;
INV     gate486  (.A(II196), .Z(n1218gat) ) ;
INV     gate487  (.A(n3085gat), .Z(II199) ) ;
INV     gate488  (.A(II199), .Z(n2861gat) ) ;
INV     gate489  (.A(n2861gat), .Z(n2859gat) ) ;
INV     gate490  (.A(n2859gat), .Z(II203) ) ;
INV     gate491  (.A(II203), .Z(n1219gat) ) ;
INV     gate492  (.A(n3084gat), .Z(II206) ) ;
INV     gate493  (.A(II206), .Z(n2864gat) ) ;
INV     gate494  (.A(n2864gat), .Z(n2862gat) ) ;
INV     gate495  (.A(n2862gat), .Z(II210) ) ;
INV     gate496  (.A(II210), .Z(n1220gat) ) ;
INV     gate497  (.A(n2861gat), .Z(II214) ) ;
INV     gate498  (.A(II214), .Z(n2860gat) ) ;
INV     gate499  (.A(n2860gat), .Z(II217) ) ;
INV     gate500  (.A(II217), .Z(n1221gat) ) ;
INV     gate501  (.A(n2864gat), .Z(II220) ) ;
INV     gate502  (.A(II220), .Z(n2863gat) ) ;
INV     gate503  (.A(n2863gat), .Z(II223) ) ;
INV     gate504  (.A(II223), .Z(n1222gat) ) ;
INV     gate505  (.A(n2856gat), .Z(II227) ) ;
INV     gate506  (.A(II227), .Z(n2855gat) ) ;
INV     gate507  (.A(n2855gat), .Z(II230) ) ;
INV     gate508  (.A(II230), .Z(n1223gat) ) ;
OR4     gate509  (.A(n1214gat), .B(n1215gat), .C(n1216gat), .D(n1217gat), .Z(n1213gat) ) ;
INV     gate510  (.A(n1213gat), .Z(n640gat) ) ;
INV     gate511  (.A(n640gat), .Z(II237) ) ;
INV     gate512  (.A(II237), .Z(n753gat) ) ;
INV     gate513  (.A(n2717gat), .Z(II240) ) ;
INV     gate514  (.A(II240), .Z(n2716gat) ) ;
INV     gate515  (.A(n3089gat), .Z(II243) ) ;
INV     gate516  (.A(II243), .Z(n2869gat) ) ;
INV     gate517  (.A(n2869gat), .Z(n2867gat) ) ;
INV     gate518  (.A(n2869gat), .Z(II248) ) ;
INV     gate519  (.A(II248), .Z(n2868gat) ) ;
OR2     gate520  (.A(n745gat), .B(n638gat), .Z(n2906gat) ) ;
INV     gate521  (.A(n2906gat), .Z(II253) ) ;
INV     gate522  (.A(II253), .Z(n754gat) ) ;
INV     gate523  (.A(n2725gat), .Z(II256) ) ;
INV     gate524  (.A(II256), .Z(n2724gat) ) ;
INV     gate525  (.A(n3086gat), .Z(II259) ) ;
INV     gate526  (.A(II259), .Z(n2728gat) ) ;
INV     gate527  (.A(n2728gat), .Z(n2726gat) ) ;
INV     gate528  (.A(n2728gat), .Z(II264) ) ;
INV     gate529  (.A(II264), .Z(n2727gat) ) ;
OR2     gate530  (.A(n423gat), .B(n362gat), .Z(n2889gat) ) ;
INV     gate531  (.A(n2889gat), .Z(n422gat) ) ;
INV     gate532  (.A(n422gat), .Z(II270) ) ;
INV     gate533  (.A(II270), .Z(n755gat) ) ;
INV     gate534  (.A(n2906gat), .Z(n747gat) ) ;
INV     gate535  (.A(n747gat), .Z(II275) ) ;
INV     gate536  (.A(II275), .Z(n756gat) ) ;
INV     gate537  (.A(n2889gat), .Z(II278) ) ;
INV     gate538  (.A(II278), .Z(n757gat) ) ;
INV     gate539  (.A(n1213gat), .Z(II282) ) ;
INV     gate540  (.A(II282), .Z(n758gat) ) ;
INV     gate541  (.A(n2510gat), .Z(n2508gat) ) ;
INV     gate542  (.A(n3065gat), .Z(II297) ) ;
INV     gate543  (.A(II297), .Z(n2733gat) ) ;
INV     gate544  (.A(n2733gat), .Z(II300) ) ;
INV     gate545  (.A(n271gat), .Z(II311) ) ;
INV     gate546  (.A(II311), .Z(n270gat) ) ;
INV     gate547  (.A(n270gat), .Z(II314) ) ;
INV     gate548  (.A(II314), .Z(n263gat) ) ;
INV     gate549  (.A(n3067gat), .Z(II317) ) ;
INV     gate550  (.A(II317), .Z(n2777gat) ) ;
INV     gate551  (.A(n2777gat), .Z(II320) ) ;
INV     gate552  (.A(n160gat), .Z(II331) ) ;
INV     gate553  (.A(II331), .Z(n159gat) ) ;
INV     gate554  (.A(n159gat), .Z(II334) ) ;
INV     gate555  (.A(II334), .Z(n264gat) ) ;
INV     gate556  (.A(n3066gat), .Z(II337) ) ;
INV     gate557  (.A(II337), .Z(n2736gat) ) ;
INV     gate558  (.A(n2736gat), .Z(II340) ) ;
INV     gate559  (.A(n337gat), .Z(II351) ) ;
INV     gate560  (.A(II351), .Z(n336gat) ) ;
INV     gate561  (.A(n336gat), .Z(II354) ) ;
INV     gate562  (.A(II354), .Z(n265gat) ) ;
INV     gate563  (.A(n160gat), .Z(n158gat) ) ;
INV     gate564  (.A(n158gat), .Z(II359) ) ;
INV     gate565  (.A(II359), .Z(n266gat) ) ;
INV     gate566  (.A(n337gat), .Z(n335gat) ) ;
INV     gate567  (.A(n335gat), .Z(II363) ) ;
INV     gate568  (.A(II363), .Z(n267gat) ) ;
INV     gate569  (.A(n271gat), .Z(n269gat) ) ;
INV     gate570  (.A(n269gat), .Z(II368) ) ;
INV     gate571  (.A(II368), .Z(n268gat) ) ;
OR4     gate572  (.A(n259gat), .B(n260gat), .C(n261gat), .D(n262gat), .Z(n258gat) ) ;
INV     gate573  (.A(n258gat), .Z(n41gat) ) ;
INV     gate574  (.A(n41gat), .Z(II375) ) ;
INV     gate575  (.A(II375), .Z(n48gat) ) ;
INV     gate576  (.A(n725gat), .Z(II378) ) ;
INV     gate577  (.A(II378), .Z(n1018gat) ) ;
INV     gate578  (.A(n3073gat), .Z(II381) ) ;
INV     gate579  (.A(II381), .Z(n2674gat) ) ;
INV     gate580  (.A(n2674gat), .Z(II384) ) ;
INV     gate581  (.A(n842gat), .Z(II395) ) ;
INV     gate582  (.A(II395), .Z(n841gat) ) ;
INV     gate583  (.A(n841gat), .Z(II398) ) ;
INV     gate584  (.A(II398), .Z(n1019gat) ) ;
INV     gate585  (.A(n721gat), .Z(II401) ) ;
INV     gate586  (.A(II401), .Z(n1020gat) ) ;
INV     gate587  (.A(n842gat), .Z(n840gat) ) ;
INV     gate588  (.A(n840gat), .Z(II406) ) ;
INV     gate589  (.A(II406), .Z(n1021gat) ) ;
INV     gate590  (.A(n720gat), .Z(II409) ) ;
INV     gate591  (.A(II409), .Z(n1022gat) ) ;
INV     gate592  (.A(n726gat), .Z(n724gat) ) ;
INV     gate593  (.A(n724gat), .Z(II414) ) ;
INV     gate594  (.A(II414), .Z(n1023gat) ) ;
OR4     gate595  (.A(n1014gat), .B(n1015gat), .C(n1016gat), .D(n1017gat), .Z(n1013gat) ) ;
INV     gate596  (.A(n1013gat), .Z(II420) ) ;
INV     gate597  (.A(II420), .Z(n49gat) ) ;
INV     gate598  (.A(n3068gat), .Z(II423) ) ;
INV     gate599  (.A(II423), .Z(n2780gat) ) ;
INV     gate600  (.A(n2780gat), .Z(II426) ) ;
INV     gate601  (.A(n341gat), .Z(II437) ) ;
INV     gate602  (.A(II437), .Z(n340gat) ) ;
INV     gate603  (.A(n340gat), .Z(II440) ) ;
INV     gate604  (.A(II440), .Z(n480gat) ) ;
INV     gate605  (.A(n702gat), .Z(II443) ) ;
INV     gate606  (.A(II443), .Z(n481gat) ) ;
INV     gate607  (.A(n394gat), .Z(II446) ) ;
INV     gate608  (.A(II446), .Z(n393gat) ) ;
INV     gate609  (.A(n393gat), .Z(II449) ) ;
INV     gate610  (.A(II449), .Z(n482gat) ) ;
INV     gate611  (.A(n701gat), .Z(II453) ) ;
INV     gate612  (.A(II453), .Z(n483gat) ) ;
INV     gate613  (.A(n392gat), .Z(II456) ) ;
INV     gate614  (.A(II456), .Z(n484gat) ) ;
INV     gate615  (.A(n341gat), .Z(n339gat) ) ;
INV     gate616  (.A(n339gat), .Z(II461) ) ;
INV     gate617  (.A(II461), .Z(n485gat) ) ;
OR4     gate618  (.A(n476gat), .B(n477gat), .C(n478gat), .D(n479gat), .Z(n475gat) ) ;
INV     gate619  (.A(n475gat), .Z(n42gat) ) ;
INV     gate620  (.A(n42gat), .Z(II468) ) ;
INV     gate621  (.A(II468), .Z(n50gat) ) ;
INV     gate622  (.A(n1013gat), .Z(n162gat) ) ;
INV     gate623  (.A(n162gat), .Z(II473) ) ;
INV     gate624  (.A(II473), .Z(n51gat) ) ;
INV     gate625  (.A(n475gat), .Z(II476) ) ;
INV     gate626  (.A(II476), .Z(n52gat) ) ;
INV     gate627  (.A(n258gat), .Z(II480) ) ;
INV     gate628  (.A(II480), .Z(n53gat) ) ;
INV     gate629  (.A(n2522gat), .Z(n2520gat) ) ;
NOR2    gate630  (.A(n724gat), .B(n720gat), .Z(n1376gat) ) ;
INV     gate631  (.A(n1376gat), .Z(n1448gat) ) ;
NOR2    gate632  (.A(n1319gat), .B(n1448gat), .Z(n1617gat) ) ;
INV     gate633  (.A(n1617gat), .Z(n1701gat) ) ;
NOR2    gate634  (.A(n724gat), .B(n721gat), .Z(n1377gat) ) ;
INV     gate635  (.A(n1377gat), .Z(n1379gat) ) ;
NOR2    gate636  (.A(n1319gat), .B(n1379gat), .Z(n1624gat) ) ;
INV     gate637  (.A(n1624gat), .Z(n1615gat) ) ;
NOR2    gate638  (.A(n393gat), .B(n701gat), .Z(n1113gat) ) ;
INV     gate639  (.A(n1113gat), .Z(n1500gat) ) ;
NOR2    gate640  (.A(n1448gat), .B(n1500gat), .Z(n1501gat) ) ;
INV     gate641  (.A(n1501gat), .Z(n1503gat) ) ;
NOR2    gate642  (.A(n1379gat), .B(n1446gat), .Z(n1623gat) ) ;
INV     gate643  (.A(n1623gat), .Z(n1779gat) ) ;
INV     gate644  (.A(n3099gat), .Z(II509) ) ;
INV     gate645  (.A(II509), .Z(n2730gat) ) ;
INV     gate646  (.A(n2730gat), .Z(II512) ) ;
INV     gate647  (.A(II512), .Z(n2729gat) ) ;
INV     gate648  (.A(n2319gat), .Z(n2317gat) ) ;
INV     gate649  (.A(n1821gat), .Z(n1819gat) ) ;
INV     gate650  (.A(n1825gat), .Z(n1823gat) ) ;
NOR2    gate651  (.A(n1819gat), .B(n1823gat), .Z(n1817gat) ) ;
INV     gate652  (.A(n1829gat), .Z(II572) ) ;
INV     gate653  (.A(II572), .Z(n1828gat) ) ;
INV     gate654  (.A(n3100gat), .Z(II576) ) ;
INV     gate655  (.A(II576), .Z(n2851gat) ) ;
INV     gate656  (.A(n2851gat), .Z(II579) ) ;
INV     gate657  (.A(II579), .Z(n2850gat) ) ;
OR2     gate658  (.A(n3091gat), .B(n3092gat), .Z(n2786gat) ) ;
INV     gate659  (.A(n2786gat), .Z(II583) ) ;
INV     gate660  (.A(II583), .Z(n2785gat) ) ;
INV     gate661  (.A(n2785gat), .Z(n92gat) ) ;
NOR2    gate662  (.A(n2724gat), .B(n2715gat), .Z(n529gat) ) ;
INV     gate663  (.A(n529gat), .Z(n637gat) ) ;
NOR2    gate664  (.A(n2859gat), .B(n2726gat), .Z(n361gat) ) ;
INV     gate665  (.A(n361gat), .Z(n293gat) ) ;
INV     gate666  (.A(n3094gat), .Z(II591) ) ;
INV     gate667  (.A(II591), .Z(n2722gat) ) ;
INV     gate668  (.A(n2722gat), .Z(II594) ) ;
INV     gate669  (.A(II594), .Z(n2721gat) ) ;
INV     gate670  (.A(n2721gat), .Z(n297gat) ) ;
INV     gate671  (.A(n283gat), .Z(II606) ) ;
INV     gate672  (.A(II606), .Z(n282gat) ) ;
INV     gate673  (.A(n282gat), .Z(II609) ) ;
INV     gate674  (.A(II609), .Z(n172gat) ) ;
INV     gate675  (.A(n165gat), .Z(II620) ) ;
INV     gate676  (.A(II620), .Z(n164gat) ) ;
INV     gate677  (.A(n164gat), .Z(II623) ) ;
INV     gate678  (.A(II623), .Z(n173gat) ) ;
INV     gate679  (.A(n279gat), .Z(II634) ) ;
INV     gate680  (.A(II634), .Z(n278gat) ) ;
INV     gate681  (.A(n278gat), .Z(II637) ) ;
INV     gate682  (.A(II637), .Z(n174gat) ) ;
INV     gate683  (.A(n165gat), .Z(n163gat) ) ;
INV     gate684  (.A(n163gat), .Z(II642) ) ;
INV     gate685  (.A(II642), .Z(n175gat) ) ;
INV     gate686  (.A(n279gat), .Z(n277gat) ) ;
INV     gate687  (.A(n277gat), .Z(II646) ) ;
INV     gate688  (.A(II646), .Z(n176gat) ) ;
INV     gate689  (.A(n283gat), .Z(n281gat) ) ;
INV     gate690  (.A(n281gat), .Z(II651) ) ;
INV     gate691  (.A(II651), .Z(n177gat) ) ;
OR4     gate692  (.A(n168gat), .B(n169gat), .C(n170gat), .D(n171gat), .Z(n167gat) ) ;
INV     gate693  (.A(n167gat), .Z(n54gat) ) ;
INV     gate694  (.A(n54gat), .Z(II658) ) ;
INV     gate695  (.A(II658), .Z(n60gat) ) ;
INV     gate696  (.A(n845gat), .Z(II661) ) ;
INV     gate697  (.A(II661), .Z(n911gat) ) ;
INV     gate698  (.A(n1026gat), .Z(II672) ) ;
INV     gate699  (.A(II672), .Z(n1025gat) ) ;
INV     gate700  (.A(n1025gat), .Z(II675) ) ;
INV     gate701  (.A(II675), .Z(n912gat) ) ;
INV     gate702  (.A(n918gat), .Z(II678) ) ;
INV     gate703  (.A(II678), .Z(n913gat) ) ;
INV     gate704  (.A(n1026gat), .Z(n1024gat) ) ;
INV     gate705  (.A(n1024gat), .Z(II683) ) ;
INV     gate706  (.A(II683), .Z(n914gat) ) ;
INV     gate707  (.A(n919gat), .Z(n917gat) ) ;
INV     gate708  (.A(n917gat), .Z(II687) ) ;
INV     gate709  (.A(II687), .Z(n915gat) ) ;
INV     gate710  (.A(n846gat), .Z(n844gat) ) ;
INV     gate711  (.A(n844gat), .Z(II692) ) ;
INV     gate712  (.A(II692), .Z(n916gat) ) ;
OR4     gate713  (.A(n907gat), .B(n908gat), .C(n909gat), .D(n910gat), .Z(n906gat) ) ;
INV     gate714  (.A(n906gat), .Z(II698) ) ;
INV     gate715  (.A(II698), .Z(n61gat) ) ;
INV     gate716  (.A(n275gat), .Z(II709) ) ;
INV     gate717  (.A(II709), .Z(n274gat) ) ;
INV     gate718  (.A(n274gat), .Z(II712) ) ;
INV     gate719  (.A(II712), .Z(n348gat) ) ;
INV     gate720  (.A(n401gat), .Z(II715) ) ;
INV     gate721  (.A(II715), .Z(n349gat) ) ;
INV     gate722  (.A(n398gat), .Z(II718) ) ;
INV     gate723  (.A(II718), .Z(n397gat) ) ;
INV     gate724  (.A(n397gat), .Z(II721) ) ;
INV     gate725  (.A(II721), .Z(n350gat) ) ;
INV     gate726  (.A(n402gat), .Z(n400gat) ) ;
INV     gate727  (.A(n400gat), .Z(II726) ) ;
INV     gate728  (.A(II726), .Z(n351gat) ) ;
INV     gate729  (.A(n396gat), .Z(II729) ) ;
INV     gate730  (.A(II729), .Z(n352gat) ) ;
INV     gate731  (.A(n275gat), .Z(n273gat) ) ;
INV     gate732  (.A(n273gat), .Z(II734) ) ;
INV     gate733  (.A(II734), .Z(n353gat) ) ;
OR4     gate734  (.A(n344gat), .B(n345gat), .C(n346gat), .D(n347gat), .Z(n343gat) ) ;
INV     gate735  (.A(n343gat), .Z(n178gat) ) ;
INV     gate736  (.A(n178gat), .Z(II741) ) ;
INV     gate737  (.A(II741), .Z(n62gat) ) ;
INV     gate738  (.A(n906gat), .Z(n66gat) ) ;
INV     gate739  (.A(n66gat), .Z(II746) ) ;
INV     gate740  (.A(II746), .Z(n63gat) ) ;
INV     gate741  (.A(n343gat), .Z(II749) ) ;
INV     gate742  (.A(II749), .Z(n64gat) ) ;
INV     gate743  (.A(n167gat), .Z(II753) ) ;
INV     gate744  (.A(II753), .Z(n65gat) ) ;
INV     gate745  (.A(n2476gat), .Z(n2474gat) ) ;
INV     gate746  (.A(n3090gat), .Z(II768) ) ;
INV     gate747  (.A(II768), .Z(n2832gat) ) ;
INV     gate748  (.A(n2832gat), .Z(II771) ) ;
INV     gate749  (.A(II771), .Z(n2831gat) ) ;
INV     gate750  (.A(n2733gat), .Z(n2731gat) ) ;
INV     gate751  (.A(n3074gat), .Z(II776) ) ;
INV     gate752  (.A(II776), .Z(n2719gat) ) ;
INV     gate753  (.A(n2719gat), .Z(n2718gat) ) ;
INV     gate754  (.A(n1068gat), .Z(II790) ) ;
INV     gate755  (.A(II790), .Z(n1067gat) ) ;
INV     gate756  (.A(n1067gat), .Z(II793) ) ;
INV     gate757  (.A(II793), .Z(n949gat) ) ;
INV     gate758  (.A(n3076gat), .Z(II796) ) ;
INV     gate759  (.A(II796), .Z(n2839gat) ) ;
INV     gate760  (.A(n2839gat), .Z(n2838gat) ) ;
INV     gate761  (.A(n2777gat), .Z(n2775gat) ) ;
INV     gate762  (.A(n957gat), .Z(II812) ) ;
INV     gate763  (.A(II812), .Z(n956gat) ) ;
INV     gate764  (.A(n956gat), .Z(II815) ) ;
INV     gate765  (.A(II815), .Z(n950gat) ) ;
INV     gate766  (.A(n3075gat), .Z(II818) ) ;
INV     gate767  (.A(II818), .Z(n2712gat) ) ;
INV     gate768  (.A(n2712gat), .Z(n2711gat) ) ;
INV     gate769  (.A(n2736gat), .Z(n2734gat) ) ;
INV     gate770  (.A(n861gat), .Z(II834) ) ;
INV     gate771  (.A(II834), .Z(n860gat) ) ;
INV     gate772  (.A(n860gat), .Z(II837) ) ;
INV     gate773  (.A(II837), .Z(n951gat) ) ;
INV     gate774  (.A(n957gat), .Z(n955gat) ) ;
INV     gate775  (.A(n955gat), .Z(II842) ) ;
INV     gate776  (.A(II842), .Z(n952gat) ) ;
INV     gate777  (.A(n861gat), .Z(n859gat) ) ;
INV     gate778  (.A(n859gat), .Z(II846) ) ;
INV     gate779  (.A(II846), .Z(n953gat) ) ;
INV     gate780  (.A(n1068gat), .Z(n1066gat) ) ;
INV     gate781  (.A(n1066gat), .Z(II851) ) ;
INV     gate782  (.A(II851), .Z(n954gat) ) ;
OR4     gate783  (.A(n945gat), .B(n946gat), .C(n947gat), .D(n948gat), .Z(n944gat) ) ;
INV     gate784  (.A(n944gat), .Z(n857gat) ) ;
INV     gate785  (.A(n857gat), .Z(II858) ) ;
INV     gate786  (.A(II858), .Z(n938gat) ) ;
INV     gate787  (.A(n2794gat), .Z(n2792gat) ) ;
INV     gate788  (.A(n3080gat), .Z(II863) ) ;
INV     gate789  (.A(II863), .Z(n2847gat) ) ;
INV     gate790  (.A(n2847gat), .Z(n2846gat) ) ;
INV     gate791  (.A(n1294gat), .Z(II877) ) ;
INV     gate792  (.A(II877), .Z(n1293gat) ) ;
INV     gate793  (.A(n1293gat), .Z(II880) ) ;
INV     gate794  (.A(II880), .Z(n1233gat) ) ;
INV     gate795  (.A(n2674gat), .Z(n2672gat) ) ;
INV     gate796  (.A(n3082gat), .Z(II885) ) ;
INV     gate797  (.A(II885), .Z(n2853gat) ) ;
INV     gate798  (.A(n2853gat), .Z(n2852gat) ) ;
INV     gate799  (.A(n1241gat), .Z(II899) ) ;
INV     gate800  (.A(II899), .Z(n1240gat) ) ;
INV     gate801  (.A(n1240gat), .Z(II902) ) ;
INV     gate802  (.A(II902), .Z(n1234gat) ) ;
INV     gate803  (.A(n1298gat), .Z(II913) ) ;
INV     gate804  (.A(II913), .Z(n1297gat) ) ;
INV     gate805  (.A(n1297gat), .Z(II916) ) ;
INV     gate806  (.A(II916), .Z(n1235gat) ) ;
INV     gate807  (.A(n1241gat), .Z(n1239gat) ) ;
INV     gate808  (.A(n1239gat), .Z(II921) ) ;
INV     gate809  (.A(II921), .Z(n1236gat) ) ;
INV     gate810  (.A(n1298gat), .Z(n1296gat) ) ;
INV     gate811  (.A(n1296gat), .Z(II925) ) ;
INV     gate812  (.A(II925), .Z(n1237gat) ) ;
INV     gate813  (.A(n1294gat), .Z(n1292gat) ) ;
INV     gate814  (.A(n1292gat), .Z(II930) ) ;
INV     gate815  (.A(II930), .Z(n1238gat) ) ;
OR4     gate816  (.A(n1229gat), .B(n1230gat), .C(n1231gat), .D(n1232gat), .Z(n1228gat) ) ;
INV     gate817  (.A(n1228gat), .Z(II936) ) ;
INV     gate818  (.A(II936), .Z(n939gat) ) ;
INV     gate819  (.A(n2780gat), .Z(n2778gat) ) ;
INV     gate820  (.A(n3077gat), .Z(II941) ) ;
INV     gate821  (.A(II941), .Z(n2837gat) ) ;
INV     gate822  (.A(n2837gat), .Z(n2836gat) ) ;
INV     gate823  (.A(n865gat), .Z(II955) ) ;
INV     gate824  (.A(II955), .Z(n864gat) ) ;
INV     gate825  (.A(n864gat), .Z(II958) ) ;
INV     gate826  (.A(II958), .Z(n1055gat) ) ;
INV     gate827  (.A(n2791gat), .Z(n2789gat) ) ;
INV     gate828  (.A(n3079gat), .Z(II963) ) ;
INV     gate829  (.A(II963), .Z(n2841gat) ) ;
INV     gate830  (.A(n2841gat), .Z(n2840gat) ) ;
INV     gate831  (.A(n1080gat), .Z(II977) ) ;
INV     gate832  (.A(II977), .Z(n1079gat) ) ;
INV     gate833  (.A(n1079gat), .Z(II980) ) ;
INV     gate834  (.A(II980), .Z(n1056gat) ) ;
INV     gate835  (.A(n2783gat), .Z(n2781gat) ) ;
INV     gate836  (.A(n3078gat), .Z(II985) ) ;
INV     gate837  (.A(II985), .Z(n2843gat) ) ;
INV     gate838  (.A(n2843gat), .Z(n2842gat) ) ;
INV     gate839  (.A(n1148gat), .Z(II999) ) ;
INV     gate840  (.A(II999), .Z(n1147gat) ) ;
INV     gate841  (.A(n1147gat), .Z(II1002) ) ;
INV     gate842  (.A(II1002), .Z(n1057gat) ) ;
INV     gate843  (.A(n1080gat), .Z(n1078gat) ) ;
INV     gate844  (.A(n1078gat), .Z(II1007) ) ;
INV     gate845  (.A(II1007), .Z(n1058gat) ) ;
INV     gate846  (.A(n1148gat), .Z(n1146gat) ) ;
INV     gate847  (.A(n1146gat), .Z(II1011) ) ;
INV     gate848  (.A(II1011), .Z(n1059gat) ) ;
INV     gate849  (.A(n865gat), .Z(n863gat) ) ;
INV     gate850  (.A(n863gat), .Z(II1016) ) ;
INV     gate851  (.A(II1016), .Z(n1060gat) ) ;
OR4     gate852  (.A(n1051gat), .B(n1052gat), .C(n1053gat), .D(n1054gat), .Z(n1050gat) ) ;
INV     gate853  (.A(n1050gat), .Z(n928gat) ) ;
INV     gate854  (.A(n928gat), .Z(II1023) ) ;
INV     gate855  (.A(II1023), .Z(n940gat) ) ;
INV     gate856  (.A(n1228gat), .Z(n858gat) ) ;
INV     gate857  (.A(n858gat), .Z(II1028) ) ;
INV     gate858  (.A(II1028), .Z(n941gat) ) ;
INV     gate859  (.A(n1050gat), .Z(II1031) ) ;
INV     gate860  (.A(II1031), .Z(n942gat) ) ;
INV     gate861  (.A(n944gat), .Z(II1035) ) ;
INV     gate862  (.A(II1035), .Z(n943gat) ) ;
INV     gate863  (.A(n2468gat), .Z(n2466gat) ) ;
INV     gate864  (.A(n2722gat), .Z(n2720gat) ) ;
INV     gate865  (.A(n2667gat), .Z(n740gat) ) ;
INV     gate866  (.A(n2786gat), .Z(n2784gat) ) ;
NOR2    gate867  (.A(n2716gat), .B(n2723gat), .Z(n746gat) ) ;
INV     gate868  (.A(n746gat), .Z(n743gat) ) ;
NOR2    gate869  (.A(n2859gat), .B(n2727gat), .Z(n360gat) ) ;
INV     gate870  (.A(n360gat), .Z(n294gat) ) ;
INV     gate871  (.A(n2767gat), .Z(n374gat) ) ;
INV     gate872  (.A(n618gat), .Z(n616gat) ) ;
INV     gate873  (.A(n616gat), .Z(II1067) ) ;
INV     gate874  (.A(II1067), .Z(n501gat) ) ;
INV     gate875  (.A(n491gat), .Z(n489gat) ) ;
INV     gate876  (.A(n489gat), .Z(II1079) ) ;
INV     gate877  (.A(II1079), .Z(n502gat) ) ;
INV     gate878  (.A(n618gat), .Z(II1082) ) ;
INV     gate879  (.A(II1082), .Z(n617gat) ) ;
INV     gate880  (.A(n617gat), .Z(II1085) ) ;
INV     gate881  (.A(II1085), .Z(n499gat) ) ;
INV     gate882  (.A(n491gat), .Z(II1088) ) ;
INV     gate883  (.A(II1088), .Z(n490gat) ) ;
INV     gate884  (.A(n490gat), .Z(II1091) ) ;
INV     gate885  (.A(II1091), .Z(n500gat) ) ;
INV     gate886  (.A(n622gat), .Z(n620gat) ) ;
INV     gate887  (.A(n620gat), .Z(II1103) ) ;
INV     gate888  (.A(II1103), .Z(n738gat) ) ;
INV     gate889  (.A(n626gat), .Z(n624gat) ) ;
INV     gate890  (.A(n624gat), .Z(II1115) ) ;
INV     gate891  (.A(II1115), .Z(n737gat) ) ;
INV     gate892  (.A(n622gat), .Z(II1118) ) ;
INV     gate893  (.A(II1118), .Z(n621gat) ) ;
INV     gate894  (.A(n621gat), .Z(II1121) ) ;
INV     gate895  (.A(II1121), .Z(n733gat) ) ;
INV     gate896  (.A(n626gat), .Z(II1124) ) ;
INV     gate897  (.A(II1124), .Z(n625gat) ) ;
INV     gate898  (.A(n625gat), .Z(II1127) ) ;
INV     gate899  (.A(II1127), .Z(n735gat) ) ;
INV     gate900  (.A(n834gat), .Z(II1138) ) ;
INV     gate901  (.A(II1138), .Z(n833gat) ) ;
INV     gate902  (.A(n833gat), .Z(II1141) ) ;
INV     gate903  (.A(II1141), .Z(n714gat) ) ;
INV     gate904  (.A(n707gat), .Z(II1152) ) ;
INV     gate905  (.A(II1152), .Z(n706gat) ) ;
INV     gate906  (.A(n706gat), .Z(II1155) ) ;
INV     gate907  (.A(II1155), .Z(n715gat) ) ;
INV     gate908  (.A(n838gat), .Z(II1166) ) ;
INV     gate909  (.A(II1166), .Z(n837gat) ) ;
INV     gate910  (.A(n837gat), .Z(II1169) ) ;
INV     gate911  (.A(II1169), .Z(n716gat) ) ;
INV     gate912  (.A(n705gat), .Z(II1174) ) ;
INV     gate913  (.A(II1174), .Z(n717gat) ) ;
INV     gate914  (.A(n836gat), .Z(II1178) ) ;
INV     gate915  (.A(II1178), .Z(n718gat) ) ;
INV     gate916  (.A(n832gat), .Z(II1183) ) ;
INV     gate917  (.A(II1183), .Z(n719gat) ) ;
OR4     gate918  (.A(n710gat), .B(n711gat), .C(n712gat), .D(n713gat), .Z(n709gat) ) ;
INV     gate919  (.A(n709gat), .Z(n515gat) ) ;
INV     gate920  (.A(n515gat), .Z(II1190) ) ;
INV     gate921  (.A(II1190), .Z(n509gat) ) ;
INV     gate922  (.A(n830gat), .Z(II1201) ) ;
INV     gate923  (.A(II1201), .Z(n829gat) ) ;
INV     gate924  (.A(n829gat), .Z(II1204) ) ;
INV     gate925  (.A(II1204), .Z(n734gat) ) ;
INV     gate926  (.A(n828gat), .Z(II1209) ) ;
INV     gate927  (.A(II1209), .Z(n736gat) ) ;
OR4     gate928  (.A(n729gat), .B(n730gat), .C(n731gat), .D(n732gat), .Z(n728gat) ) ;
INV     gate929  (.A(n728gat), .Z(II1216) ) ;
INV     gate930  (.A(II1216), .Z(n510gat) ) ;
INV     gate931  (.A(n614gat), .Z(II1227) ) ;
INV     gate932  (.A(II1227), .Z(n613gat) ) ;
INV     gate933  (.A(n613gat), .Z(II1230) ) ;
INV     gate934  (.A(II1230), .Z(n498gat) ) ;
INV     gate935  (.A(n612gat), .Z(II1236) ) ;
INV     gate936  (.A(II1236), .Z(n503gat) ) ;
OR4     gate937  (.A(n494gat), .B(n495gat), .C(n496gat), .D(n497gat), .Z(n493gat) ) ;
INV     gate938  (.A(n493gat), .Z(n404gat) ) ;
INV     gate939  (.A(n404gat), .Z(II1243) ) ;
INV     gate940  (.A(II1243), .Z(n511gat) ) ;
INV     gate941  (.A(n728gat), .Z(n405gat) ) ;
INV     gate942  (.A(n405gat), .Z(II1248) ) ;
INV     gate943  (.A(II1248), .Z(n512gat) ) ;
INV     gate944  (.A(n493gat), .Z(II1251) ) ;
INV     gate945  (.A(II1251), .Z(n513gat) ) ;
INV     gate946  (.A(n709gat), .Z(II1255) ) ;
INV     gate947  (.A(II1255), .Z(n514gat) ) ;
INV     gate948  (.A(n2526gat), .Z(n2524gat) ) ;
NOR4    gate949  (.A(n3029gat), .B(n2863gat), .C(n2855gat), .D(n374gat), .Z(n564gat) ) ;
INV     gate950  (.A(n564gat), .Z(n17gat) ) ;
NOR3    gate951  (.A(n743gat), .B(n294gat), .C(n17gat), .Z(n86gat) ) ;
INV     gate952  (.A(n86gat), .Z(n79gat) ) ;
NOR2    gate953  (.A(n2784gat), .B(n79gat), .Z(n78gat) ) ;
INV     gate954  (.A(n78gat), .Z(n219gat) ) ;
OR3     gate955  (.A(n740gat), .B(n3030gat), .C(II1277), .Z(II1278) ) ;
INV     gate956  (.A(II1278), .Z(n563gat) ) ;
INV     gate957  (.A(n563gat), .Z(n289gat) ) ;
NOR2    gate958  (.A(n289gat), .B(n2715gat), .Z(n287gat) ) ;
INV     gate959  (.A(n287gat), .Z(n179gat) ) ;
NOR2    gate960  (.A(n289gat), .B(n2726gat), .Z(n288gat) ) ;
INV     gate961  (.A(n288gat), .Z(n188gat) ) ;
NOR3    gate962  (.A(n286gat), .B(n179gat), .C(n188gat), .Z(n181gat) ) ;
INV     gate963  (.A(n181gat), .Z(n72gat) ) ;
NOR2    gate964  (.A(n72gat), .B(n2720gat), .Z(n182gat) ) ;
INV     gate965  (.A(n182gat), .Z(n111gat) ) ;
INV     gate966  (.A(n680gat), .Z(II1302) ) ;
INV     gate967  (.A(II1302), .Z(n679gat) ) ;
INV     gate968  (.A(n679gat), .Z(II1305) ) ;
INV     gate969  (.A(II1305), .Z(n808gat) ) ;
INV     gate970  (.A(n816gat), .Z(II1319) ) ;
INV     gate971  (.A(II1319), .Z(n815gat) ) ;
INV     gate972  (.A(n815gat), .Z(II1322) ) ;
INV     gate973  (.A(II1322), .Z(n809gat) ) ;
INV     gate974  (.A(n580gat), .Z(II1336) ) ;
INV     gate975  (.A(II1336), .Z(n579gat) ) ;
INV     gate976  (.A(n579gat), .Z(II1339) ) ;
INV     gate977  (.A(II1339), .Z(n810gat) ) ;
INV     gate978  (.A(n816gat), .Z(n814gat) ) ;
INV     gate979  (.A(n814gat), .Z(II1344) ) ;
INV     gate980  (.A(II1344), .Z(n811gat) ) ;
INV     gate981  (.A(n580gat), .Z(n578gat) ) ;
INV     gate982  (.A(n578gat), .Z(II1348) ) ;
INV     gate983  (.A(II1348), .Z(n812gat) ) ;
INV     gate984  (.A(n680gat), .Z(n678gat) ) ;
INV     gate985  (.A(n678gat), .Z(II1353) ) ;
INV     gate986  (.A(II1353), .Z(n813gat) ) ;
OR4     gate987  (.A(n804gat), .B(n805gat), .C(n806gat), .D(n807gat), .Z(n803gat) ) ;
INV     gate988  (.A(n803gat), .Z(n677gat) ) ;
INV     gate989  (.A(n677gat), .Z(II1360) ) ;
INV     gate990  (.A(II1360), .Z(n572gat) ) ;
INV     gate991  (.A(n824gat), .Z(II1371) ) ;
INV     gate992  (.A(II1371), .Z(n823gat) ) ;
INV     gate993  (.A(n823gat), .Z(II1374) ) ;
INV     gate994  (.A(II1374), .Z(n591gat) ) ;
INV     gate995  (.A(n820gat), .Z(II1385) ) ;
INV     gate996  (.A(II1385), .Z(n819gat) ) ;
INV     gate997  (.A(n819gat), .Z(II1388) ) ;
INV     gate998  (.A(II1388), .Z(n592gat) ) ;
INV     gate999  (.A(n883gat), .Z(II1399) ) ;
INV     gate1000  (.A(II1399), .Z(n882gat) ) ;
INV     gate1001  (.A(n882gat), .Z(II1402) ) ;
INV     gate1002  (.A(II1402), .Z(n593gat) ) ;
INV     gate1003  (.A(n818gat), .Z(II1407) ) ;
INV     gate1004  (.A(II1407), .Z(n594gat) ) ;
INV     gate1005  (.A(n881gat), .Z(II1411) ) ;
INV     gate1006  (.A(II1411), .Z(n595gat) ) ;
INV     gate1007  (.A(n822gat), .Z(II1416) ) ;
INV     gate1008  (.A(II1416), .Z(n596gat) ) ;
OR4     gate1009  (.A(n587gat), .B(n588gat), .C(n589gat), .D(n590gat), .Z(n586gat) ) ;
INV     gate1010  (.A(n586gat), .Z(II1422) ) ;
INV     gate1011  (.A(II1422), .Z(n573gat) ) ;
INV     gate1012  (.A(n584gat), .Z(II1436) ) ;
INV     gate1013  (.A(II1436), .Z(n583gat) ) ;
INV     gate1014  (.A(n583gat), .Z(II1439) ) ;
INV     gate1015  (.A(II1439), .Z(n691gat) ) ;
INV     gate1016  (.A(n684gat), .Z(II1450) ) ;
INV     gate1017  (.A(II1450), .Z(n683gat) ) ;
INV     gate1018  (.A(n683gat), .Z(II1453) ) ;
INV     gate1019  (.A(II1453), .Z(n692gat) ) ;
INV     gate1020  (.A(n699gat), .Z(II1464) ) ;
INV     gate1021  (.A(II1464), .Z(n698gat) ) ;
INV     gate1022  (.A(n698gat), .Z(II1467) ) ;
INV     gate1023  (.A(II1467), .Z(n693gat) ) ;
INV     gate1024  (.A(n682gat), .Z(II1472) ) ;
INV     gate1025  (.A(II1472), .Z(n694gat) ) ;
INV     gate1026  (.A(n697gat), .Z(II1476) ) ;
INV     gate1027  (.A(II1476), .Z(n695gat) ) ;
INV     gate1028  (.A(n584gat), .Z(n582gat) ) ;
INV     gate1029  (.A(n582gat), .Z(II1481) ) ;
INV     gate1030  (.A(II1481), .Z(n696gat) ) ;
OR4     gate1031  (.A(n687gat), .B(n688gat), .C(n689gat), .D(n690gat), .Z(n686gat) ) ;
INV     gate1032  (.A(n686gat), .Z(n456gat) ) ;
INV     gate1033  (.A(n456gat), .Z(II1488) ) ;
INV     gate1034  (.A(II1488), .Z(n574gat) ) ;
INV     gate1035  (.A(n586gat), .Z(n565gat) ) ;
INV     gate1036  (.A(n565gat), .Z(II1493) ) ;
INV     gate1037  (.A(II1493), .Z(n575gat) ) ;
INV     gate1038  (.A(n686gat), .Z(II1496) ) ;
INV     gate1039  (.A(II1496), .Z(n576gat) ) ;
INV     gate1040  (.A(n803gat), .Z(II1500) ) ;
INV     gate1041  (.A(II1500), .Z(n577gat) ) ;
INV     gate1042  (.A(n2464gat), .Z(n2462gat) ) ;
OR3     gate1043  (.A(n2466gat), .B(n2462gat), .C(II1515), .Z(II1516) ) ;
INV     gate1044  (.A(II1516), .Z(n2665gat) ) ;
INV     gate1045  (.A(n2665gat), .Z(n2596gat) ) ;
NOR2    gate1046  (.A(n289gat), .B(n2723gat), .Z(n286gat) ) ;
INV     gate1047  (.A(n286gat), .Z(n189gat) ) ;
NOR3    gate1048  (.A(n189gat), .B(n287gat), .C(n188gat), .Z(n187gat) ) ;
INV     gate1049  (.A(n187gat), .Z(n194gat) ) ;
NOR3    gate1050  (.A(n637gat), .B(n17gat), .C(n293gat), .Z(n15gat) ) ;
INV     gate1051  (.A(n15gat), .Z(n21gat) ) ;
INV     gate1052  (.A(n2399gat), .Z(II1538) ) ;
INV     gate1053  (.A(II1538), .Z(n2398gat) ) ;
INV     gate1054  (.A(n2398gat), .Z(n2353gat) ) ;
INV     gate1055  (.A(n2343gat), .Z(II1550) ) ;
INV     gate1056  (.A(II1550), .Z(n2342gat) ) ;
INV     gate1057  (.A(n2342gat), .Z(n2284gat) ) ;
INV     gate1058  (.A(n2201gat), .Z(n2354gat) ) ;
INV     gate1059  (.A(n2560gat), .Z(n2356gat) ) ;
INV     gate1060  (.A(n2205gat), .Z(n2214gat) ) ;
OR3     gate1061  (.A(n2356gat), .B(n2214gat), .C(II1584), .Z(II1585) ) ;
INV     gate1062  (.A(II1585), .Z(n2286gat) ) ;
INV     gate1063  (.A(n2626gat), .Z(n2624gat) ) ;
INV     gate1064  (.A(n2490gat), .Z(II1606) ) ;
INV     gate1065  (.A(II1606), .Z(n2489gat) ) ;
INV     gate1066  (.A(n2622gat), .Z(II1617) ) ;
INV     gate1067  (.A(II1617), .Z(n2621gat) ) ;
NOR3    gate1068  (.A(n2624gat), .B(n2489gat), .C(n2621gat), .Z(n2534gat) ) ;
INV     gate1069  (.A(n2534gat), .Z(n2533gat) ) ;
INV     gate1070  (.A(n2630gat), .Z(II1630) ) ;
INV     gate1071  (.A(II1630), .Z(n2629gat) ) ;
INV     gate1072  (.A(n2629gat), .Z(n2486gat) ) ;
INV     gate1073  (.A(n2541gat), .Z(n2429gat) ) ;
NOR3    gate1074  (.A(n2533gat), .B(n2486gat), .C(n2429gat), .Z(n2430gat) ) ;
INV     gate1075  (.A(n2430gat), .Z(n2432gat) ) ;
INV     gate1076  (.A(n2102gat), .Z(II1655) ) ;
INV     gate1077  (.A(II1655), .Z(n2101gat) ) ;
INV     gate1078  (.A(n2101gat), .Z(n1693gat) ) ;
INV     gate1079  (.A(n1880gat), .Z(II1667) ) ;
INV     gate1080  (.A(II1667), .Z(n1879gat) ) ;
NOR3    gate1081  (.A(n2470gat), .B(n1935gat), .C(n2239gat), .Z(n1934gat) ) ;
INV     gate1082  (.A(n1934gat), .Z(n1698gat) ) ;
INV     gate1083  (.A(n1606gat), .Z(n1543gat) ) ;
INV     gate1084  (.A(n1763gat), .Z(II1683) ) ;
INV     gate1085  (.A(II1683), .Z(n1762gat) ) ;
OR2     gate1086  (.A(n1693gat), .B(n1692gat), .Z(n2989gat) ) ;
INV     gate1087  (.A(n2989gat), .Z(n1673gat) ) ;
INV     gate1088  (.A(n2155gat), .Z(II1698) ) ;
INV     gate1089  (.A(II1698), .Z(n2154gat) ) ;
INV     gate1090  (.A(n2490gat), .Z(n2488gat) ) ;
INV     gate1091  (.A(n2626gat), .Z(II1703) ) ;
INV     gate1092  (.A(II1703), .Z(n2625gat) ) ;
NOR3    gate1093  (.A(n2488gat), .B(n2625gat), .C(n2621gat), .Z(n2531gat) ) ;
INV     gate1094  (.A(n2531gat), .Z(n2530gat) ) ;
INV     gate1095  (.A(n2543gat), .Z(II1708) ) ;
INV     gate1096  (.A(II1708), .Z(n2542gat) ) ;
INV     gate1097  (.A(n2542gat), .Z(n2482gat) ) ;
NOR3    gate1098  (.A(n2530gat), .B(n2482gat), .C(n2486gat), .Z(n2480gat) ) ;
INV     gate1099  (.A(n2480gat), .Z(n2426gat) ) ;
INV     gate1100  (.A(n2155gat), .Z(n2153gat) ) ;
INV     gate1101  (.A(n2341gat), .Z(n2355gat) ) ;
INV     gate1102  (.A(n2562gat), .Z(II1719) ) ;
INV     gate1103  (.A(II1719), .Z(n2561gat) ) ;
INV     gate1104  (.A(n2561gat), .Z(n2443gat) ) ;
OR3     gate1105  (.A(n2355gat), .B(n2443gat), .C(II1723), .Z(II1724) ) ;
INV     gate1106  (.A(II1724), .Z(n2289gat) ) ;
OR3     gate1107  (.A(n1604gat), .B(n2214gat), .C(II1733), .Z(II1734) ) ;
INV     gate1108  (.A(II1734), .Z(n2148gat) ) ;
INV     gate1109  (.A(n2148gat), .Z(n855gat) ) ;
INV     gate1110  (.A(n855gat), .Z(n759gat) ) ;
INV     gate1111  (.A(n1035gat), .Z(II1749) ) ;
INV     gate1112  (.A(II1749), .Z(n1034gat) ) ;
INV     gate1113  (.A(n1034gat), .Z(II1752) ) ;
INV     gate1114  (.A(II1752), .Z(n1189gat) ) ;
INV     gate1115  (.A(n855gat), .Z(n1075gat) ) ;
INV     gate1116  (.A(n1121gat), .Z(II1766) ) ;
INV     gate1117  (.A(II1766), .Z(n1120gat) ) ;
INV     gate1118  (.A(n1120gat), .Z(II1769) ) ;
INV     gate1119  (.A(II1769), .Z(n1190gat) ) ;
INV     gate1120  (.A(n855gat), .Z(n760gat) ) ;
INV     gate1121  (.A(n1072gat), .Z(II1783) ) ;
INV     gate1122  (.A(II1783), .Z(n1071gat) ) ;
INV     gate1123  (.A(n1071gat), .Z(II1786) ) ;
INV     gate1124  (.A(II1786), .Z(n1191gat) ) ;
INV     gate1125  (.A(n1121gat), .Z(n1119gat) ) ;
INV     gate1126  (.A(n1119gat), .Z(II1791) ) ;
INV     gate1127  (.A(II1791), .Z(n1192gat) ) ;
INV     gate1128  (.A(n1072gat), .Z(n1070gat) ) ;
INV     gate1129  (.A(n1070gat), .Z(II1795) ) ;
INV     gate1130  (.A(II1795), .Z(n1193gat) ) ;
INV     gate1131  (.A(n1035gat), .Z(n1033gat) ) ;
INV     gate1132  (.A(n1033gat), .Z(II1800) ) ;
INV     gate1133  (.A(II1800), .Z(n1194gat) ) ;
OR4     gate1134  (.A(n1185gat), .B(n1186gat), .C(n1187gat), .D(n1188gat), .Z(n1184gat) ) ;
INV     gate1135  (.A(n1184gat), .Z(n1183gat) ) ;
INV     gate1136  (.A(n1183gat), .Z(II1807) ) ;
INV     gate1137  (.A(II1807), .Z(n1274gat) ) ;
INV     gate1138  (.A(n855gat), .Z(n644gat) ) ;
INV     gate1139  (.A(n1282gat), .Z(n1280gat) ) ;
INV     gate1140  (.A(n855gat), .Z(n641gat) ) ;
INV     gate1141  (.A(n1226gat), .Z(II1833) ) ;
INV     gate1142  (.A(II1833), .Z(n1225gat) ) ;
INV     gate1143  (.A(n1282gat), .Z(II1837) ) ;
INV     gate1144  (.A(II1837), .Z(n1281gat) ) ;
INV     gate1145  (.A(n1226gat), .Z(n1224gat) ) ;
OR2     gate1146  (.A(n1383gat), .B(n1327gat), .Z(n2970gat) ) ;
INV     gate1147  (.A(n2970gat), .Z(II1843) ) ;
INV     gate1148  (.A(II1843), .Z(n1275gat) ) ;
INV     gate1149  (.A(n855gat), .Z(n761gat) ) ;
INV     gate1150  (.A(n931gat), .Z(II1857) ) ;
INV     gate1151  (.A(II1857), .Z(n930gat) ) ;
INV     gate1152  (.A(n930gat), .Z(II1860) ) ;
INV     gate1153  (.A(II1860), .Z(n1206gat) ) ;
INV     gate1154  (.A(n855gat), .Z(n762gat) ) ;
INV     gate1155  (.A(n1135gat), .Z(II1874) ) ;
INV     gate1156  (.A(II1874), .Z(n1134gat) ) ;
INV     gate1157  (.A(n1134gat), .Z(II1877) ) ;
INV     gate1158  (.A(II1877), .Z(n1207gat) ) ;
INV     gate1159  (.A(n855gat), .Z(n643gat) ) ;
INV     gate1160  (.A(n1045gat), .Z(II1891) ) ;
INV     gate1161  (.A(II1891), .Z(n1044gat) ) ;
INV     gate1162  (.A(n1044gat), .Z(II1894) ) ;
INV     gate1163  (.A(II1894), .Z(n1208gat) ) ;
INV     gate1164  (.A(n1135gat), .Z(n1133gat) ) ;
INV     gate1165  (.A(n1133gat), .Z(II1899) ) ;
INV     gate1166  (.A(II1899), .Z(n1209gat) ) ;
INV     gate1167  (.A(n1045gat), .Z(n1043gat) ) ;
INV     gate1168  (.A(n1043gat), .Z(II1903) ) ;
INV     gate1169  (.A(II1903), .Z(n1210gat) ) ;
INV     gate1170  (.A(n931gat), .Z(n929gat) ) ;
INV     gate1171  (.A(n929gat), .Z(II1908) ) ;
INV     gate1172  (.A(II1908), .Z(n1211gat) ) ;
OR4     gate1173  (.A(n1202gat), .B(n1203gat), .C(n1204gat), .D(n1205gat), .Z(n1201gat) ) ;
INV     gate1174  (.A(n1201gat), .Z(n1268gat) ) ;
INV     gate1175  (.A(n1268gat), .Z(II1915) ) ;
INV     gate1176  (.A(II1915), .Z(n1276gat) ) ;
INV     gate1177  (.A(n2970gat), .Z(n1329gat) ) ;
INV     gate1178  (.A(n1329gat), .Z(II1920) ) ;
INV     gate1179  (.A(II1920), .Z(n1277gat) ) ;
INV     gate1180  (.A(n1201gat), .Z(II1923) ) ;
INV     gate1181  (.A(II1923), .Z(n1278gat) ) ;
INV     gate1182  (.A(n1184gat), .Z(II1927) ) ;
INV     gate1183  (.A(II1927), .Z(n1279gat) ) ;
OR4     gate1184  (.A(n1270gat), .B(n1271gat), .C(n1272gat), .D(n1273gat), .Z(n1269gat) ) ;
INV     gate1185  (.A(n1269gat), .Z(n1284gat) ) ;
INV     gate1186  (.A(n855gat), .Z(n642gat) ) ;
INV     gate1187  (.A(n1197gat), .Z(n1195gat) ) ;
INV     gate1188  (.A(n1197gat), .Z(II1947) ) ;
INV     gate1189  (.A(II1947), .Z(n1196gat) ) ;
INV     gate1190  (.A(n2518gat), .Z(n2516gat) ) ;
INV     gate1191  (.A(n2516gat), .Z(II1961) ) ;
INV     gate1192  (.A(II1961), .Z(n3017gat) ) ;
NOR2    gate1193  (.A(n740gat), .B(n2148gat), .Z(n853gat) ) ;
INV     gate1194  (.A(n853gat), .Z(n851gat) ) ;
INV     gate1195  (.A(n2148gat), .Z(n1725gat) ) ;
INV     gate1196  (.A(n1725gat), .Z(n664gat) ) ;
NOR2    gate1197  (.A(n2148gat), .B(n374gat), .Z(n854gat) ) ;
INV     gate1198  (.A(n854gat), .Z(n852gat) ) ;
INV     gate1199  (.A(n667gat), .Z(II1981) ) ;
INV     gate1200  (.A(II1981), .Z(n666gat) ) ;
INV     gate1201  (.A(n1725gat), .Z(n368gat) ) ;
INV     gate1202  (.A(n659gat), .Z(II1996) ) ;
INV     gate1203  (.A(II1996), .Z(n658gat) ) ;
INV     gate1204  (.A(n658gat), .Z(II1999) ) ;
INV     gate1205  (.A(II1999), .Z(n784gat) ) ;
INV     gate1206  (.A(n1725gat), .Z(n662gat) ) ;
INV     gate1207  (.A(n553gat), .Z(II2014) ) ;
INV     gate1208  (.A(II2014), .Z(n552gat) ) ;
INV     gate1209  (.A(n552gat), .Z(II2017) ) ;
INV     gate1210  (.A(II2017), .Z(n785gat) ) ;
INV     gate1211  (.A(n1725gat), .Z(n661gat) ) ;
INV     gate1212  (.A(n777gat), .Z(II2032) ) ;
INV     gate1213  (.A(II2032), .Z(n776gat) ) ;
INV     gate1214  (.A(n776gat), .Z(II2035) ) ;
INV     gate1215  (.A(II2035), .Z(n786gat) ) ;
INV     gate1216  (.A(n553gat), .Z(n551gat) ) ;
INV     gate1217  (.A(n551gat), .Z(II2040) ) ;
INV     gate1218  (.A(II2040), .Z(n787gat) ) ;
INV     gate1219  (.A(n777gat), .Z(n775gat) ) ;
INV     gate1220  (.A(n775gat), .Z(II2044) ) ;
INV     gate1221  (.A(II2044), .Z(n788gat) ) ;
INV     gate1222  (.A(n659gat), .Z(n657gat) ) ;
INV     gate1223  (.A(n657gat), .Z(II2049) ) ;
INV     gate1224  (.A(II2049), .Z(n789gat) ) ;
OR4     gate1225  (.A(n780gat), .B(n781gat), .C(n782gat), .D(n783gat), .Z(n779gat) ) ;
INV     gate1226  (.A(n779gat), .Z(n35gat) ) ;
INV     gate1227  (.A(n35gat), .Z(II2056) ) ;
INV     gate1228  (.A(II2056), .Z(n125gat) ) ;
INV     gate1229  (.A(n1725gat), .Z(n558gat) ) ;
INV     gate1230  (.A(n561gat), .Z(n559gat) ) ;
INV     gate1231  (.A(n1725gat), .Z(n371gat) ) ;
INV     gate1232  (.A(n366gat), .Z(II2084) ) ;
INV     gate1233  (.A(II2084), .Z(n365gat) ) ;
INV     gate1234  (.A(n561gat), .Z(II2088) ) ;
INV     gate1235  (.A(II2088), .Z(n560gat) ) ;
INV     gate1236  (.A(n366gat), .Z(n364gat) ) ;
OR2     gate1237  (.A(n874gat), .B(n132gat), .Z(n2876gat) ) ;
INV     gate1238  (.A(n2876gat), .Z(II2094) ) ;
INV     gate1239  (.A(II2094), .Z(n126gat) ) ;
INV     gate1240  (.A(n1725gat), .Z(n663gat) ) ;
INV     gate1241  (.A(n322gat), .Z(II2109) ) ;
INV     gate1242  (.A(II2109), .Z(n321gat) ) ;
INV     gate1243  (.A(n321gat), .Z(II2112) ) ;
INV     gate1244  (.A(II2112), .Z(n226gat) ) ;
INV     gate1245  (.A(n1725gat), .Z(n370gat) ) ;
INV     gate1246  (.A(n318gat), .Z(II2127) ) ;
INV     gate1247  (.A(II2127), .Z(n317gat) ) ;
INV     gate1248  (.A(n317gat), .Z(II2130) ) ;
INV     gate1249  (.A(II2130), .Z(n227gat) ) ;
INV     gate1250  (.A(n1725gat), .Z(n369gat) ) ;
INV     gate1251  (.A(n314gat), .Z(II2145) ) ;
INV     gate1252  (.A(II2145), .Z(n313gat) ) ;
INV     gate1253  (.A(n313gat), .Z(II2148) ) ;
INV     gate1254  (.A(II2148), .Z(n228gat) ) ;
INV     gate1255  (.A(n318gat), .Z(n316gat) ) ;
INV     gate1256  (.A(n316gat), .Z(II2153) ) ;
INV     gate1257  (.A(II2153), .Z(n229gat) ) ;
INV     gate1258  (.A(n314gat), .Z(n312gat) ) ;
INV     gate1259  (.A(n312gat), .Z(II2157) ) ;
INV     gate1260  (.A(II2157), .Z(n230gat) ) ;
INV     gate1261  (.A(n322gat), .Z(n320gat) ) ;
INV     gate1262  (.A(n320gat), .Z(II2162) ) ;
INV     gate1263  (.A(II2162), .Z(n231gat) ) ;
OR4     gate1264  (.A(n222gat), .B(n223gat), .C(n224gat), .D(n225gat), .Z(n221gat) ) ;
INV     gate1265  (.A(n221gat), .Z(n34gat) ) ;
INV     gate1266  (.A(n34gat), .Z(II2169) ) ;
INV     gate1267  (.A(II2169), .Z(n127gat) ) ;
INV     gate1268  (.A(n2876gat), .Z(n133gat) ) ;
INV     gate1269  (.A(n133gat), .Z(II2174) ) ;
INV     gate1270  (.A(II2174), .Z(n128gat) ) ;
INV     gate1271  (.A(n221gat), .Z(II2177) ) ;
INV     gate1272  (.A(II2177), .Z(n129gat) ) ;
INV     gate1273  (.A(n779gat), .Z(II2181) ) ;
INV     gate1274  (.A(II2181), .Z(n130gat) ) ;
INV     gate1275  (.A(n667gat), .Z(n665gat) ) ;
OR4     gate1276  (.A(n121gat), .B(n122gat), .C(n123gat), .D(n124gat), .Z(n120gat) ) ;
INV     gate1277  (.A(n120gat), .Z(n1601gat) ) ;
INV     gate1278  (.A(n2599gat), .Z(n2597gat) ) ;
NOR3    gate1279  (.A(n3017gat), .B(n2520gat), .C(n2597gat), .Z(n2594gat) ) ;
INV     gate1280  (.A(n2594gat), .Z(n2595gat) ) ;
INV     gate1281  (.A(n2588gat), .Z(n2586gat) ) ;
INV     gate1282  (.A(n2342gat), .Z(II2213) ) ;
INV     gate1283  (.A(II2213), .Z(n2573gat) ) ;
INV     gate1284  (.A(n2638gat), .Z(II2225) ) ;
INV     gate1285  (.A(II2225), .Z(n2574gat) ) ;
INV     gate1286  (.A(n2561gat), .Z(II2228) ) ;
INV     gate1287  (.A(II2228), .Z(n2575gat) ) ;
INV     gate1288  (.A(n2640gat), .Z(II2232) ) ;
INV     gate1289  (.A(II2232), .Z(n2639gat) ) ;
INV     gate1290  (.A(n2639gat), .Z(II2235) ) ;
INV     gate1291  (.A(II2235), .Z(n2576gat) ) ;
INV     gate1292  (.A(n2560gat), .Z(II2238) ) ;
INV     gate1293  (.A(II2238), .Z(n2577gat) ) ;
INV     gate1294  (.A(n2341gat), .Z(II2242) ) ;
INV     gate1295  (.A(II2242), .Z(n2578gat) ) ;
OR4     gate1296  (.A(n2569gat), .B(n2570gat), .C(n2571gat), .D(n2572gat), .Z(n2568gat) ) ;
INV     gate1297  (.A(n2568gat), .Z(II2248) ) ;
INV     gate1298  (.A(II2248), .Z(n2582gat) ) ;
INV     gate1299  (.A(n2207gat), .Z(II2251) ) ;
INV     gate1300  (.A(II2251), .Z(n2206gat) ) ;
INV     gate1301  (.A(n2206gat), .Z(II2254) ) ;
INV     gate1302  (.A(II2254), .Z(n2414gat) ) ;
INV     gate1303  (.A(n2398gat), .Z(II2257) ) ;
INV     gate1304  (.A(II2257), .Z(n2415gat) ) ;
INV     gate1305  (.A(n2203gat), .Z(II2260) ) ;
INV     gate1306  (.A(II2260), .Z(n2202gat) ) ;
INV     gate1307  (.A(n2202gat), .Z(II2263) ) ;
INV     gate1308  (.A(II2263), .Z(n2416gat) ) ;
INV     gate1309  (.A(n2397gat), .Z(II2268) ) ;
INV     gate1310  (.A(II2268), .Z(n2417gat) ) ;
INV     gate1311  (.A(n2201gat), .Z(II2271) ) ;
INV     gate1312  (.A(II2271), .Z(n2418gat) ) ;
INV     gate1313  (.A(n2205gat), .Z(II2275) ) ;
INV     gate1314  (.A(II2275), .Z(n2419gat) ) ;
OR4     gate1315  (.A(n2410gat), .B(n2411gat), .C(n2412gat), .D(n2413gat), .Z(n2409gat) ) ;
INV     gate1316  (.A(n2409gat), .Z(II2281) ) ;
INV     gate1317  (.A(II2281), .Z(n2585gat) ) ;
INV     gate1318  (.A(n2658gat), .Z(n2656gat) ) ;
INV     gate1319  (.A(n2390gat), .Z(II2316) ) ;
INV     gate1320  (.A(II2316), .Z(n2389gat) ) ;
INV     gate1321  (.A(n2495gat), .Z(II2319) ) ;
INV     gate1322  (.A(II2319), .Z(n2494gat) ) ;
OR2     gate1323  (.A(n2567gat), .B(n2499gat), .Z(n3014gat) ) ;
INV     gate1324  (.A(n3014gat), .Z(II2324) ) ;
INV     gate1325  (.A(II2324), .Z(n2649gat) ) ;
INV     gate1326  (.A(n2339gat), .Z(II2344) ) ;
INV     gate1327  (.A(II2344), .Z(n2338gat) ) ;
INV     gate1328  (.A(n2270gat), .Z(II2349) ) ;
INV     gate1329  (.A(II2349), .Z(n2269gat) ) ;
OR2     gate1330  (.A(n299gat), .B(n207gat), .Z(n2880gat) ) ;
INV     gate1331  (.A(n2880gat), .Z(II2354) ) ;
INV     gate1332  (.A(II2354), .Z(n2652gat) ) ;
INV     gate1333  (.A(n2502gat), .Z(n2500gat) ) ;
INV     gate1334  (.A(n2622gat), .Z(n2620gat) ) ;
INV     gate1335  (.A(n2620gat), .Z(n2612gat) ) ;
INV     gate1336  (.A(n2612gat), .Z(II2372) ) ;
INV     gate1337  (.A(II2372), .Z(n2606gat) ) ;
INV     gate1338  (.A(n2532gat), .Z(II2376) ) ;
INV     gate1339  (.A(II2376), .Z(n2607gat) ) ;
INV     gate1340  (.A(n2488gat), .Z(n2540gat) ) ;
INV     gate1341  (.A(n2540gat), .Z(II2380) ) ;
INV     gate1342  (.A(II2380), .Z(n2608gat) ) ;
INV     gate1343  (.A(n2624gat), .Z(n2536gat) ) ;
INV     gate1344  (.A(n2536gat), .Z(II2385) ) ;
INV     gate1345  (.A(II2385), .Z(n2609gat) ) ;
INV     gate1346  (.A(n2487gat), .Z(II2389) ) ;
INV     gate1347  (.A(II2389), .Z(n2610gat) ) ;
INV     gate1348  (.A(n2557gat), .Z(II2394) ) ;
INV     gate1349  (.A(II2394), .Z(n2611gat) ) ;
OR4     gate1350  (.A(n2602gat), .B(n2603gat), .C(n2604gat), .D(n2605gat), .Z(n2601gat) ) ;
INV     gate1351  (.A(n2601gat), .Z(II2400) ) ;
INV     gate1352  (.A(II2400), .Z(n2616gat) ) ;
INV     gate1353  (.A(n2629gat), .Z(II2403) ) ;
INV     gate1354  (.A(II2403), .Z(n2550gat) ) ;
INV     gate1355  (.A(n2634gat), .Z(II2414) ) ;
INV     gate1356  (.A(II2414), .Z(n2633gat) ) ;
INV     gate1357  (.A(n2633gat), .Z(II2417) ) ;
INV     gate1358  (.A(II2417), .Z(n2551gat) ) ;
INV     gate1359  (.A(n2542gat), .Z(II2420) ) ;
INV     gate1360  (.A(II2420), .Z(n2552gat) ) ;
INV     gate1361  (.A(n2632gat), .Z(II2425) ) ;
INV     gate1362  (.A(II2425), .Z(n2553gat) ) ;
INV     gate1363  (.A(n2541gat), .Z(II2428) ) ;
INV     gate1364  (.A(II2428), .Z(n2554gat) ) ;
INV     gate1365  (.A(n2628gat), .Z(II2433) ) ;
INV     gate1366  (.A(II2433), .Z(n2555gat) ) ;
OR4     gate1367  (.A(n2546gat), .B(n2547gat), .C(n2548gat), .D(n2549gat), .Z(n2545gat) ) ;
INV     gate1368  (.A(n2545gat), .Z(II2439) ) ;
INV     gate1369  (.A(II2439), .Z(n2619gat) ) ;
INV     gate1370  (.A(n2506gat), .Z(n2504gat) ) ;
NOR4    gate1371  (.A(n2508gat), .B(n2656gat), .C(n2500gat), .D(n2504gat), .Z(n2655gat) ) ;
INV     gate1372  (.A(n2655gat), .Z(n2660gat) ) ;
NOR3    gate1373  (.A(n2353gat), .B(n2284gat), .C(n2443gat), .Z(n2293gat) ) ;
INV     gate1374  (.A(n2293gat), .Z(n1528gat) ) ;
NOR2    gate1375  (.A(n2354gat), .B(n2214gat), .Z(n2219gat) ) ;
INV     gate1376  (.A(n2219gat), .Z(n1523gat) ) ;
NOR2    gate1377  (.A(n1528gat), .B(n1523gat), .Z(n1529gat) ) ;
INV     gate1378  (.A(n1529gat), .Z(n1592gat) ) ;
NOR2    gate1379  (.A(n3027gat), .B(n1706gat), .Z(n1704gat) ) ;
INV     gate1380  (.A(n1704gat), .Z(n2666gat) ) ;
OR2     gate1381  (.A(n2461gat), .B(n2421gat), .Z(n3013gat) ) ;
INV     gate1382  (.A(n3013gat), .Z(n2422gat) ) ;
INV     gate1383  (.A(n2202gat), .Z(n2290gat) ) ;
NOR2    gate1384  (.A(n2214gat), .B(n2290gat), .Z(n2218gat) ) ;
INV     gate1385  (.A(n2218gat), .Z(n2081gat) ) ;
INV     gate1386  (.A(n2397gat), .Z(n2285gat) ) ;
NOR3    gate1387  (.A(n2285gat), .B(n2356gat), .C(n2355gat), .Z(n2358gat) ) ;
INV     gate1388  (.A(n2358gat), .Z(n2359gat) ) ;
NOR2    gate1389  (.A(n2081gat), .B(n2359gat), .Z(n1415gat) ) ;
INV     gate1390  (.A(n1415gat), .Z(n1414gat) ) ;
INV     gate1391  (.A(n364gat), .Z(n566gat) ) ;
NOR3    gate1392  (.A(n2443gat), .B(n2284gat), .C(n2285gat), .Z(n2292gat) ) ;
INV     gate1393  (.A(n2292gat), .Z(n1480gat) ) ;
NOR2    gate1394  (.A(n2081gat), .B(n1480gat), .Z(n1416gat) ) ;
INV     gate1395  (.A(n1416gat), .Z(n1301gat) ) ;
INV     gate1396  (.A(n312gat), .Z(n1150gat) ) ;
INV     gate1397  (.A(n316gat), .Z(n873gat) ) ;
NOR3    gate1398  (.A(n2356gat), .B(n2284gat), .C(n2285gat), .Z(n2306gat) ) ;
INV     gate1399  (.A(n2306gat), .Z(n2011gat) ) ;
NOR2    gate1400  (.A(n2081gat), .B(n2011gat), .Z(n1481gat) ) ;
INV     gate1401  (.A(n1481gat), .Z(n1478gat) ) ;
INV     gate1402  (.A(n559gat), .Z(n875gat) ) ;
NOR3    gate1403  (.A(n2285gat), .B(n2355gat), .C(n2443gat), .Z(n2357gat) ) ;
INV     gate1404  (.A(n2357gat), .Z(n1410gat) ) ;
NOR2    gate1405  (.A(n2081gat), .B(n1410gat), .Z(n1347gat) ) ;
INV     gate1406  (.A(n1347gat), .Z(n876gat) ) ;
NOR2    gate1407  (.A(n2081gat), .B(n1528gat), .Z(n1484gat) ) ;
INV     gate1408  (.A(n1484gat), .Z(n1160gat) ) ;
INV     gate1409  (.A(n657gat), .Z(n1084gat) ) ;
INV     gate1410  (.A(n320gat), .Z(n983gat) ) ;
NOR3    gate1411  (.A(n2353gat), .B(n2356gat), .C(n2355gat), .Z(n2363gat) ) ;
INV     gate1412  (.A(n2363gat), .Z(n1482gat) ) ;
NOR2    gate1413  (.A(n2081gat), .B(n1482gat), .Z(n1483gat) ) ;
INV     gate1414  (.A(n1483gat), .Z(n1157gat) ) ;
INV     gate1415  (.A(n775gat), .Z(n985gat) ) ;
NOR3    gate1416  (.A(n2353gat), .B(n2284gat), .C(n2356gat), .Z(n2364gat) ) ;
INV     gate1417  (.A(n2364gat), .Z(n1530gat) ) ;
NOR2    gate1418  (.A(n2081gat), .B(n1530gat), .Z(n1308gat) ) ;
INV     gate1419  (.A(n1308gat), .Z(n1307gat) ) ;
INV     gate1420  (.A(n551gat), .Z(n1085gat) ) ;
NOR3    gate1421  (.A(n2353gat), .B(n2355gat), .C(n2443gat), .Z(n2291gat) ) ;
INV     gate1422  (.A(n2291gat), .Z(n1479gat) ) ;
NOR2    gate1423  (.A(n1479gat), .B(n2081gat), .Z(n1349gat) ) ;
INV     gate1424  (.A(n1349gat), .Z(n1348gat) ) ;
INV     gate1425  (.A(n2206gat), .Z(n2217gat) ) ;
NOR2    gate1426  (.A(n2354gat), .B(n2217gat), .Z(n2223gat) ) ;
INV     gate1427  (.A(n2223gat), .Z(n1591gat) ) ;
NOR2    gate1428  (.A(n1591gat), .B(n1480gat), .Z(n1438gat) ) ;
INV     gate1429  (.A(n1438gat), .Z(n1437gat) ) ;
INV     gate1430  (.A(n1834gat), .Z(n1832gat) ) ;
INV     gate1431  (.A(n1767gat), .Z(n1765gat) ) ;
INV     gate1432  (.A(n1880gat), .Z(n1878gat) ) ;
NOR3    gate1433  (.A(n1832gat), .B(n1765gat), .C(n1878gat), .Z(n1831gat) ) ;
INV     gate1434  (.A(n1831gat), .Z(n1442gat) ) ;
INV     gate1435  (.A(n1442gat), .Z(n1444gat) ) ;
OR2     gate1436  (.A(n1443gat), .B(n1325gat), .Z(n2975gat) ) ;
INV     gate1437  (.A(n2975gat), .Z(n1378gat) ) ;
OR2     gate1438  (.A(n1321gat), .B(n1320gat), .Z(n2974gat) ) ;
INV     gate1439  (.A(n2974gat), .Z(n1322gat) ) ;
NOR2    gate1440  (.A(n1482gat), .B(n1591gat), .Z(n1486gat) ) ;
INV     gate1441  (.A(n1486gat), .Z(n1439gat) ) ;
NOR2    gate1442  (.A(n2011gat), .B(n1591gat), .Z(n1426gat) ) ;
INV     gate1443  (.A(n1426gat), .Z(n1370gat) ) ;
OR2     gate1444  (.A(n1368gat), .B(n1258gat), .Z(n2966gat) ) ;
INV     gate1445  (.A(n2966gat), .Z(n1369gat) ) ;
NOR2    gate1446  (.A(n1479gat), .B(n1591gat), .Z(n1365gat) ) ;
INV     gate1447  (.A(n1365gat), .Z(n1366gat) ) ;
OR2     gate1448  (.A(n1373gat), .B(n1372gat), .Z(n2979gat) ) ;
INV     gate1449  (.A(n2979gat), .Z(n1374gat) ) ;
NOR2    gate1450  (.A(n2290gat), .B(n2217gat), .Z(n2220gat) ) ;
INV     gate1451  (.A(n2220gat), .Z(n2162gat) ) ;
NOR2    gate1452  (.A(n2162gat), .B(n1530gat), .Z(n1423gat) ) ;
INV     gate1453  (.A(n1423gat), .Z(n1450gat) ) ;
NOR2    gate1454  (.A(n1704gat), .B(n1703gat), .Z(n1608gat) ) ;
INV     gate1455  (.A(n1608gat), .Z(n1427gat) ) ;
INV     gate1456  (.A(n2084gat), .Z(n2082gat) ) ;
NOR2    gate1457  (.A(n1528gat), .B(n2162gat), .Z(n1494gat) ) ;
INV     gate1458  (.A(n1494gat), .Z(n1449gat) ) ;
INV     gate1459  (.A(n1603gat), .Z(n1590gat) ) ;
OR2     gate1460  (.A(n1250gat), .B(n1103gat), .Z(n2954gat) ) ;
INV     gate1461  (.A(n2954gat), .Z(n1248gat) ) ;
NOR2    gate1462  (.A(n2162gat), .B(n1480gat), .Z(n1417gat) ) ;
INV     gate1463  (.A(n1417gat), .Z(n1418gat) ) ;
OR2     gate1464  (.A(n1304gat), .B(n1249gat), .Z(n2964gat) ) ;
INV     gate1465  (.A(n2964gat), .Z(n1306gat) ) ;
NOR2    gate1466  (.A(n2162gat), .B(n1479gat), .Z(n1419gat) ) ;
INV     gate1467  (.A(n1419gat), .Z(n1353gat) ) ;
OR2     gate1468  (.A(n1246gat), .B(n1161gat), .Z(n2958gat) ) ;
INV     gate1469  (.A(n2958gat), .Z(n1247gat) ) ;
NOR2    gate1470  (.A(n2011gat), .B(n2162gat), .Z(n1422gat) ) ;
INV     gate1471  (.A(n1422gat), .Z(n1355gat) ) ;
OR2     gate1472  (.A(n1291gat), .B(n1245gat), .Z(n2963gat) ) ;
INV     gate1473  (.A(n2963gat), .Z(n1300gat) ) ;
NOR2    gate1474  (.A(n1482gat), .B(n2162gat), .Z(n1485gat) ) ;
INV     gate1475  (.A(n1485gat), .Z(n1487gat) ) ;
OR2     gate1476  (.A(n1163gat), .B(n1102gat), .Z(n2953gat) ) ;
INV     gate1477  (.A(n2953gat), .Z(n1164gat) ) ;
NOR2    gate1478  (.A(n1591gat), .B(n1530gat), .Z(n1354gat) ) ;
INV     gate1479  (.A(n1354gat), .Z(n1356gat) ) ;
NOR2    gate1480  (.A(n1591gat), .B(n1528gat), .Z(n1435gat) ) ;
INV     gate1481  (.A(n1435gat), .Z(n1436gat) ) ;
OR2     gate1482  (.A(n1101gat), .B(n996gat), .Z(n2949gat) ) ;
INV     gate1483  (.A(n2949gat), .Z(n1106gat) ) ;
NOR2    gate1484  (.A(n2162gat), .B(n2359gat), .Z(n1421gat) ) ;
INV     gate1485  (.A(n1421gat), .Z(n1425gat) ) ;
OR2     gate1486  (.A(n1104gat), .B(n887gat), .Z(n2934gat) ) ;
INV     gate1487  (.A(n2934gat), .Z(n1105gat) ) ;
NOR2    gate1488  (.A(n1410gat), .B(n2162gat), .Z(n1420gat) ) ;
INV     gate1489  (.A(n1420gat), .Z(n1424gat) ) ;
OR2     gate1490  (.A(n1305gat), .B(n1162gat), .Z(n2959gat) ) ;
INV     gate1491  (.A(n2959gat), .Z(n1309gat) ) ;
INV     gate1492  (.A(n2143gat), .Z(II2672) ) ;
INV     gate1493  (.A(II2672), .Z(n2142gat) ) ;
INV     gate1494  (.A(n2142gat), .Z(n1788gat) ) ;
INV     gate1495  (.A(n2061gat), .Z(II2684) ) ;
INV     gate1496  (.A(II2684), .Z(n2060gat) ) ;
INV     gate1497  (.A(n2060gat), .Z(n1786gat) ) ;
INV     gate1498  (.A(n2139gat), .Z(II2696) ) ;
INV     gate1499  (.A(II2696), .Z(n2138gat) ) ;
INV     gate1500  (.A(n2138gat), .Z(n1839gat) ) ;
INV     gate1501  (.A(n1899gat), .Z(n1897gat) ) ;
INV     gate1502  (.A(n1897gat), .Z(n1884gat) ) ;
INV     gate1503  (.A(n1850gat), .Z(n1848gat) ) ;
INV     gate1504  (.A(n1848gat), .Z(n1783gat) ) ;
OR3     gate1505  (.A(n1884gat), .B(n1783gat), .C(II2720), .Z(II2721) ) ;
INV     gate1506  (.A(II2721), .Z(n1548gat) ) ;
INV     gate1507  (.A(n1548gat), .Z(n1719gat) ) ;
INV     gate1508  (.A(n2139gat), .Z(n2137gat) ) ;
INV     gate1509  (.A(n2137gat), .Z(n1633gat) ) ;
INV     gate1510  (.A(n2061gat), .Z(n2059gat) ) ;
INV     gate1511  (.A(n2059gat), .Z(n1785gat) ) ;
INV     gate1512  (.A(n1850gat), .Z(II2731) ) ;
INV     gate1513  (.A(II2731), .Z(n1849gat) ) ;
INV     gate1514  (.A(n1849gat), .Z(n1784gat) ) ;
OR3     gate1515  (.A(n1785gat), .B(n1784gat), .C(II2735), .Z(II2736) ) ;
INV     gate1516  (.A(II2736), .Z(n1716gat) ) ;
INV     gate1517  (.A(n1716gat), .Z(n1635gat) ) ;
INV     gate1518  (.A(n2403gat), .Z(n2401gat) ) ;
INV     gate1519  (.A(n2401gat), .Z(n1989gat) ) ;
INV     gate1520  (.A(n2394gat), .Z(n2392gat) ) ;
INV     gate1521  (.A(n2392gat), .Z(n1918gat) ) ;
INV     gate1522  (.A(n2440gat), .Z(II2771) ) ;
INV     gate1523  (.A(II2771), .Z(n2439gat) ) ;
INV     gate1524  (.A(n2439gat), .Z(n1986gat) ) ;
NOR3    gate1525  (.A(n1989gat), .B(n1918gat), .C(n1986gat), .Z(n1865gat) ) ;
INV     gate1526  (.A(n1865gat), .Z(n1866gat) ) ;
INV     gate1527  (.A(n2407gat), .Z(II2785) ) ;
INV     gate1528  (.A(II2785), .Z(n2406gat) ) ;
INV     gate1529  (.A(n2406gat), .Z(n2216gat) ) ;
INV     gate1530  (.A(n2347gat), .Z(n2345gat) ) ;
INV     gate1531  (.A(n2345gat), .Z(n1988gat) ) ;
NOR3    gate1532  (.A(n1866gat), .B(n2216gat), .C(n1988gat), .Z(n1861gat) ) ;
INV     gate1533  (.A(n1861gat), .Z(n1735gat) ) ;
INV     gate1534  (.A(n1389gat), .Z(n1387gat) ) ;
OR4     gate1535  (.A(n1609gat), .B(n1702gat), .C(n1700gat), .D(II2812), .Z(II2813) ) ;
INV     gate1536  (.A(II2813), .Z(n1694gat) ) ;
NOR3    gate1537  (.A(n1777gat), .B(n1625gat), .C(n1626gat), .Z(n1780gat) ) ;
INV     gate1538  (.A(n2021gat), .Z(n2019gat) ) ;
OR3     gate1539  (.A(n1884gat), .B(n1784gat), .C(II2831), .Z(II2832) ) ;
INV     gate1540  (.A(II2832), .Z(n1549gat) ) ;
INV     gate1541  (.A(n1549gat), .Z(n1551gat) ) ;
INV     gate1542  (.A(n2347gat), .Z(II2837) ) ;
INV     gate1543  (.A(II2837), .Z(n2346gat) ) ;
INV     gate1544  (.A(n2346gat), .Z(n2152gat) ) ;
INV     gate1545  (.A(n2407gat), .Z(n2405gat) ) ;
INV     gate1546  (.A(n2405gat), .Z(n2351gat) ) ;
INV     gate1547  (.A(n2403gat), .Z(II2843) ) ;
INV     gate1548  (.A(II2843), .Z(n2402gat) ) ;
INV     gate1549  (.A(n2402gat), .Z(n2212gat) ) ;
INV     gate1550  (.A(n2394gat), .Z(II2847) ) ;
INV     gate1551  (.A(II2847), .Z(n2393gat) ) ;
INV     gate1552  (.A(n2393gat), .Z(n1991gat) ) ;
NOR3    gate1553  (.A(n1986gat), .B(n2212gat), .C(n1991gat), .Z(n1666gat) ) ;
INV     gate1554  (.A(n1666gat), .Z(n1665gat) ) ;
NOR3    gate1555  (.A(n2152gat), .B(n2351gat), .C(n1665gat), .Z(n1578gat) ) ;
INV     gate1556  (.A(n1578gat), .Z(n1517gat) ) ;
INV     gate1557  (.A(n1496gat), .Z(II2873) ) ;
INV     gate1558  (.A(II2873), .Z(n1495gat) ) ;
NOR4    gate1559  (.A(n1778gat), .B(n1609gat), .C(n1702gat), .D(n1700gat), .Z(n1604gat) ) ;
INV     gate1560  (.A(n2091gat), .Z(II2885) ) ;
INV     gate1561  (.A(II2885), .Z(n2090gat) ) ;
OR3     gate1562  (.A(n1788gat), .B(n1786gat), .C(II2889), .Z(II2890) ) ;
INV     gate1563  (.A(II2890), .Z(n1550gat) ) ;
INV     gate1564  (.A(n1550gat), .Z(n1552gat) ) ;
INV     gate1565  (.A(n1740gat), .Z(n1738gat) ) ;
INV     gate1566  (.A(n1740gat), .Z(II2915) ) ;
INV     gate1567  (.A(II2915), .Z(n1739gat) ) ;
NOR3    gate1568  (.A(n1864gat), .B(n1921gat), .C(n1798gat), .Z(n1920gat) ) ;
INV     gate1569  (.A(n1920gat), .Z(n1925gat) ) ;
NOR2    gate1570  (.A(n1738gat), .B(n1673gat), .Z(n1921gat) ) ;
INV     gate1571  (.A(n1921gat), .Z(n1917gat) ) ;
INV     gate1572  (.A(n2143gat), .Z(n2141gat) ) ;
INV     gate1573  (.A(n2141gat), .Z(n1787gat) ) ;
OR3     gate1574  (.A(n1884gat), .B(n1787gat), .C(II2925), .Z(II2926) ) ;
INV     gate1575  (.A(n1717gat), .Z(n1859gat) ) ;
NOR2    gate1576  (.A(n1739gat), .B(n1673gat), .Z(n1798gat) ) ;
INV     gate1577  (.A(n1798gat), .Z(n1922gat) ) ;
OR3     gate1578  (.A(n1785gat), .B(n1884gat), .C(II2934), .Z(II2935) ) ;
INV     gate1579  (.A(n1713gat), .Z(n1743gat) ) ;
NOR3    gate1580  (.A(n1858gat), .B(n1495gat), .C(n2090gat), .Z(n1864gat) ) ;
INV     gate1581  (.A(n1864gat), .Z(n1923gat) ) ;
NOR2    gate1582  (.A(n1700gat), .B(n1702gat), .Z(n1690gat) ) ;
INV     gate1583  (.A(n2179gat), .Z(II2953) ) ;
INV     gate1584  (.A(II2953), .Z(n2178gat) ) ;
NOR3    gate1585  (.A(n1918gat), .B(n1986gat), .C(n2212gat), .Z(n1660gat) ) ;
INV     gate1586  (.A(n1660gat), .Z(n1661gat) ) ;
NOR3    gate1587  (.A(n2351gat), .B(n1988gat), .C(n1661gat), .Z(n1576gat) ) ;
INV     gate1588  (.A(n1576gat), .Z(n1572gat) ) ;
INV     gate1589  (.A(n2440gat), .Z(n2438gat) ) ;
INV     gate1590  (.A(n2438gat), .Z(n2283gat) ) ;
NOR3    gate1591  (.A(n2283gat), .B(n1991gat), .C(n2212gat), .Z(n1582gat) ) ;
INV     gate1592  (.A(n1582gat), .Z(n1520gat) ) ;
NOR3    gate1593  (.A(n1520gat), .B(n2351gat), .C(n1988gat), .Z(n1577gat) ) ;
INV     gate1594  (.A(n1577gat), .Z(n1580gat) ) ;
OR2     gate1595  (.A(n1733gat), .B(n1581gat), .Z(n2988gat) ) ;
INV     gate1596  (.A(n2988gat), .Z(n1990gat) ) ;
INV     gate1597  (.A(n2190gat), .Z(II2978) ) ;
INV     gate1598  (.A(II2978), .Z(n2189gat) ) ;
INV     gate1599  (.A(n2135gat), .Z(II2989) ) ;
INV     gate1600  (.A(II2989), .Z(n2134gat) ) ;
INV     gate1601  (.A(n2262gat), .Z(II3000) ) ;
INV     gate1602  (.A(II3000), .Z(n2261gat) ) ;
NOR3    gate1603  (.A(n2189gat), .B(n2134gat), .C(n2261gat), .Z(n2129gat) ) ;
INV     gate1604  (.A(n2129gat), .Z(n2128gat) ) ;
NOR4    gate1605  (.A(n1609gat), .B(n1778gat), .C(n1704gat), .D(n1703gat), .Z(n1695gat) ) ;
INV     gate1606  (.A(n2182gat), .Z(II3016) ) ;
INV     gate1607  (.A(II3016), .Z(n2181gat) ) ;
INV     gate1608  (.A(n1312gat), .Z(II3056) ) ;
INV     gate1609  (.A(II3056), .Z(n1311gat) ) ;
INV     gate1610  (.A(n1626gat), .Z(n1707gat) ) ;
OR2     gate1611  (.A(n1574gat), .B(n1573gat), .Z(n2987gat) ) ;
INV     gate1612  (.A(n2987gat), .Z(n1659gat) ) ;
NOR2    gate1613  (.A(n2283gat), .B(n1991gat), .Z(n1521gat) ) ;
INV     gate1614  (.A(n1521gat), .Z(n1515gat) ) ;
NOR2    gate1615  (.A(n2212gat), .B(n2152gat), .Z(n1737gat) ) ;
INV     gate1616  (.A(n1737gat), .Z(n1736gat) ) ;
INV     gate1617  (.A(n2216gat), .Z(n1658gat) ) ;
NOR3    gate1618  (.A(n1515gat), .B(n1736gat), .C(n1658gat), .Z(n1732gat) ) ;
INV     gate1619  (.A(n1732gat), .Z(n1724gat) ) ;
NOR2    gate1620  (.A(n1986gat), .B(n1918gat), .Z(n1663gat) ) ;
INV     gate1621  (.A(n1663gat), .Z(n1662gat) ) ;
NOR3    gate1622  (.A(n1736gat), .B(n1662gat), .C(n1658gat), .Z(n1655gat) ) ;
INV     gate1623  (.A(n1655gat), .Z(n1656gat) ) ;
NOR2    gate1624  (.A(n1991gat), .B(n1986gat), .Z(n1667gat) ) ;
INV     gate1625  (.A(n1667gat), .Z(n1670gat) ) ;
NOR3    gate1626  (.A(n1736gat), .B(n1658gat), .C(n1670gat), .Z(n1570gat) ) ;
INV     gate1627  (.A(n1570gat), .Z(n1569gat) ) ;
NOR2    gate1628  (.A(n1918gat), .B(n2283gat), .Z(n1575gat) ) ;
INV     gate1629  (.A(n1575gat), .Z(n1568gat) ) ;
NOR3    gate1630  (.A(n1568gat), .B(n1736gat), .C(n1658gat), .Z(n1728gat) ) ;
INV     gate1631  (.A(n1728gat), .Z(n1727gat) ) ;
NOR2    gate1632  (.A(n2152gat), .B(n1989gat), .Z(n1801gat) ) ;
INV     gate1633  (.A(n1801gat), .Z(n1797gat) ) ;
NOR3    gate1634  (.A(n1658gat), .B(n1515gat), .C(n1797gat), .Z(n1731gat) ) ;
INV     gate1635  (.A(n1731gat), .Z(n1730gat) ) ;
NOR3    gate1636  (.A(n1670gat), .B(n1658gat), .C(n1797gat), .Z(n1571gat) ) ;
INV     gate1637  (.A(n1571gat), .Z(n1561gat) ) ;
NOR2    gate1638  (.A(n1988gat), .B(n2212gat), .Z(n1734gat) ) ;
INV     gate1639  (.A(n1734gat), .Z(n1668gat) ) ;
INV     gate1640  (.A(n2216gat), .Z(n1742gat) ) ;
NOR3    gate1641  (.A(n1668gat), .B(n1742gat), .C(n1670gat), .Z(n1669gat) ) ;
INV     gate1642  (.A(n1669gat), .Z(n1671gat) ) ;
NOR3    gate1643  (.A(n1662gat), .B(n1797gat), .C(n1658gat), .Z(n1657gat) ) ;
INV     gate1644  (.A(n1657gat), .Z(n1652gat) ) ;
NOR3    gate1645  (.A(n1658gat), .B(n1797gat), .C(n1568gat), .Z(n1729gat) ) ;
INV     gate1646  (.A(n1729gat), .Z(n1648gat) ) ;
NOR3    gate1647  (.A(n2992gat), .B(n2986gat), .C(n2991gat), .Z(n1726gat) ) ;
INV     gate1648  (.A(n1726gat), .Z(n1790gat) ) ;
NOR2    gate1649  (.A(n1758gat), .B(n1790gat), .Z(n1929gat) ) ;
INV     gate1650  (.A(n1929gat), .Z(n2004gat) ) ;
INV     gate1651  (.A(n1871gat), .Z(n1869gat) ) ;
INV     gate1652  (.A(n2592gat), .Z(II3143) ) ;
INV     gate1653  (.A(II3143), .Z(n2591gat) ) ;
INV     gate1654  (.A(n2989gat), .Z(n1584gat) ) ;
OR3     gate1655  (.A(n1786gat), .B(n1787gat), .C(II3148), .Z(II3149) ) ;
INV     gate1656  (.A(II3149), .Z(n1714gat) ) ;
INV     gate1657  (.A(n1714gat), .Z(n1718gat) ) ;
INV     gate1658  (.A(n1508gat), .Z(II3163) ) ;
INV     gate1659  (.A(II3163), .Z(n1507gat) ) ;
NOR2    gate1660  (.A(n1584gat), .B(n1590gat), .Z(n1401gat) ) ;
INV     gate1661  (.A(n1401gat), .Z(n1396gat) ) ;
INV     gate1662  (.A(n1394gat), .Z(II3168) ) ;
INV     gate1663  (.A(II3168), .Z(n1393gat) ) ;
NOR2    gate1664  (.A(n1858gat), .B(n1590gat), .Z(n1476gat) ) ;
INV     gate1665  (.A(n1476gat), .Z(n1409gat) ) ;
INV     gate1666  (.A(n1899gat), .Z(II3174) ) ;
INV     gate1667  (.A(II3174), .Z(n1898gat) ) ;
INV     gate1668  (.A(n1898gat), .Z(n1838gat) ) ;
OR3     gate1669  (.A(n1839gat), .B(n1784gat), .C(II3178), .Z(II3179) ) ;
INV     gate1670  (.A(n1678gat), .Z(II3191) ) ;
INV     gate1671  (.A(II3191), .Z(n1677gat) ) ;
NOR3    gate1672  (.A(n1411gat), .B(n1406gat), .C(n2981gat), .Z(n1412gat) ) ;
INV     gate1673  (.A(n1412gat), .Z(n2000gat) ) ;
INV     gate1674  (.A(n1412gat), .Z(n2001gat) ) ;
INV     gate1675  (.A(n2001gat), .Z(n1999gat) ) ;
NOR3    gate1676  (.A(n2586gat), .B(n2660gat), .C(n2307gat), .Z(n2663gat) ) ;
INV     gate1677  (.A(n2663gat), .Z(II3211) ) ;
INV     gate1678  (.A(II3211), .Z(n3018gat) ) ;
INV     gate1679  (.A(n2450gat), .Z(n2448gat) ) ;
NOR2    gate1680  (.A(n2660gat), .B(n2586gat), .Z(n2662gat) ) ;
INV     gate1681  (.A(n2446gat), .Z(n2444gat) ) ;
NOR2    gate1682  (.A(n2448gat), .B(n2444gat), .Z(n2238gat) ) ;
INV     gate1683  (.A(n2238gat), .Z(II3235) ) ;
INV     gate1684  (.A(II3235), .Z(n3019gat) ) ;
INV     gate1685  (.A(n1312gat), .Z(n1310gat) ) ;
NOR3    gate1686  (.A(n743gat), .B(n17gat), .C(n293gat), .Z(n87gat) ) ;
INV     gate1687  (.A(n87gat), .Z(n199gat) ) ;
NOR3    gate1688  (.A(n189gat), .B(n188gat), .C(n179gat), .Z(n184gat) ) ;
INV     gate1689  (.A(n184gat), .Z(n195gat) ) ;
NOR2    gate1690  (.A(n200gat), .B(n196gat), .Z(n204gat) ) ;
INV     gate1691  (.A(n2169gat), .Z(II3273) ) ;
INV     gate1692  (.A(II3273), .Z(n2168gat) ) ;
INV     gate1693  (.A(n2454gat), .Z(n2452gat) ) ;
INV     gate1694  (.A(n2452gat), .Z(n1691gat) ) ;
INV     gate1695  (.A(n1691gat), .Z(II3287) ) ;
INV     gate1696  (.A(II3287), .Z(n3020gat) ) ;
INV     gate1697  (.A(n1691gat), .Z(II3290) ) ;
INV     gate1698  (.A(II3290), .Z(n3021gat) ) ;
INV     gate1699  (.A(n1691gat), .Z(II3293) ) ;
INV     gate1700  (.A(II3293), .Z(n3022gat) ) ;
INV     gate1701  (.A(n2452gat), .Z(n1699gat) ) ;
INV     gate1702  (.A(n1699gat), .Z(II3297) ) ;
INV     gate1703  (.A(II3297), .Z(n3023gat) ) ;
INV     gate1704  (.A(n1699gat), .Z(II3300) ) ;
INV     gate1705  (.A(II3300), .Z(n3024gat) ) ;
INV     gate1706  (.A(n1691gat), .Z(II3303) ) ;
INV     gate1707  (.A(II3303), .Z(n3025gat) ) ;
INV     gate1708  (.A(n1699gat), .Z(II3306) ) ;
INV     gate1709  (.A(II3306), .Z(n3026gat) ) ;
INV     gate1710  (.A(n1699gat), .Z(II3309) ) ;
INV     gate1711  (.A(II3309), .Z(n3027gat) ) ;
INV     gate1712  (.A(n1699gat), .Z(II3312) ) ;
INV     gate1713  (.A(II3312), .Z(n3028gat) ) ;
INV     gate1714  (.A(n1869gat), .Z(II3315) ) ;
INV     gate1715  (.A(II3315), .Z(n3029gat) ) ;
INV     gate1716  (.A(n1869gat), .Z(II3318) ) ;
INV     gate1717  (.A(II3318), .Z(n3030gat) ) ;
INV     gate1718  (.A(n2262gat), .Z(n2260gat) ) ;
INV     gate1719  (.A(n2189gat), .Z(n2257gat) ) ;
INV     gate1720  (.A(n2190gat), .Z(n2188gat) ) ;
OR3     gate1721  (.A(n2258gat), .B(n2257gat), .C(n2255gat), .Z(n3004gat) ) ;
INV     gate1722  (.A(n3004gat), .Z(n2187gat) ) ;
INV     gate1723  (.A(n2040gat), .Z(II3336) ) ;
INV     gate1724  (.A(II3336), .Z(n2039gat) ) ;
INV     gate1725  (.A(n1775gat), .Z(II3339) ) ;
INV     gate1726  (.A(II3339), .Z(n1774gat) ) ;
INV     gate1727  (.A(n1316gat), .Z(II3342) ) ;
INV     gate1728  (.A(II3342), .Z(n1315gat) ) ;
INV     gate1729  (.A(n2099gat), .Z(n2097gat) ) ;
NOR4    gate1730  (.A(n2035gat), .B(n2093gat), .C(n2018gat), .D(n2664gat), .Z(n2014gat) ) ;
INV     gate1731  (.A(n2014gat), .Z(n1855gat) ) ;
NOR2    gate1732  (.A(n2187gat), .B(n1855gat), .Z(n2194gat) ) ;
INV     gate1733  (.A(n2194gat), .Z(II3387) ) ;
INV     gate1734  (.A(n2261gat), .Z(II3390) ) ;
INV     gate1735  (.A(II3390), .Z(n3032gat) ) ;
INV     gate1736  (.A(n3032gat), .Z(n2256gat) ) ;
INV     gate1737  (.A(n2260gat), .Z(II3394) ) ;
INV     gate1738  (.A(II3394), .Z(n3033gat) ) ;
INV     gate1739  (.A(n3033gat), .Z(n2251gat) ) ;
OR2     gate1740  (.A(n2256gat), .B(n2251gat), .Z(n3003gat) ) ;
INV     gate1741  (.A(n3003gat), .Z(n2184gat) ) ;
NOR2    gate1742  (.A(n2184gat), .B(n1855gat), .Z(n2192gat) ) ;
INV     gate1743  (.A(n2192gat), .Z(II3401) ) ;
INV     gate1744  (.A(n2135gat), .Z(n2133gat) ) ;
NOR2    gate1745  (.A(n2261gat), .B(n2189gat), .Z(n2185gat) ) ;
INV     gate1746  (.A(n2185gat), .Z(n2131gat) ) ;
OR2     gate1747  (.A(n2132gat), .B(n2130gat), .Z(n3001gat) ) ;
INV     gate1748  (.A(n3001gat), .Z(n2049gat) ) ;
NOR2    gate1749  (.A(n2049gat), .B(n1855gat), .Z(n2057gat) ) ;
INV     gate1750  (.A(n2057gat), .Z(II3412) ) ;
INV     gate1751  (.A(n2189gat), .Z(n2253gat) ) ;
INV     gate1752  (.A(n2260gat), .Z(n2252gat) ) ;
OR2     gate1753  (.A(n2253gat), .B(n2252gat), .Z(n3006gat) ) ;
INV     gate1754  (.A(n3006gat), .Z(n2248gat) ) ;
INV     gate1755  (.A(n2266gat), .Z(n2264gat) ) ;
INV     gate1756  (.A(n2266gat), .Z(II3429) ) ;
INV     gate1757  (.A(II3429), .Z(n2265gat) ) ;
NOR2    gate1758  (.A(n1855gat), .B(n3007gat), .Z(n2329gat) ) ;
INV     gate1759  (.A(n2329gat), .Z(n2492gat) ) ;
INV     gate1760  (.A(n2492gat), .Z(II3436) ) ;
INV     gate1761  (.A(n1849gat), .Z(n1709gat) ) ;
INV     gate1762  (.A(n2141gat), .Z(n1845gat) ) ;
INV     gate1763  (.A(n2059gat), .Z(n1891gat) ) ;
INV     gate1764  (.A(n2137gat), .Z(n1963gat) ) ;
INV     gate1765  (.A(n1897gat), .Z(n1886gat) ) ;
NOR2    gate1766  (.A(n1963gat), .B(n1886gat), .Z(n1958gat) ) ;
INV     gate1767  (.A(n1958gat), .Z(n1968gat) ) ;
NOR3    gate1768  (.A(n1845gat), .B(n1891gat), .C(n1968gat), .Z(n1895gat) ) ;
INV     gate1769  (.A(n1895gat), .Z(n1629gat) ) ;
INV     gate1770  (.A(n1848gat), .Z(n1631gat) ) ;
OR2     gate1771  (.A(n1710gat), .B(n1630gat), .Z(n2990gat) ) ;
INV     gate1772  (.A(n2990gat), .Z(n1711gat) ) ;
NOR4    gate1773  (.A(n1926gat), .B(n1916gat), .C(n1994gat), .D(n1924gat), .Z(n2078gat) ) ;
INV     gate1774  (.A(n2078gat), .Z(n2200gat) ) ;
NOR2    gate1775  (.A(n2200gat), .B(n1855gat), .Z(n2195gat) ) ;
INV     gate1776  (.A(n2195gat), .Z(n2437gat) ) ;
NOR2    gate1777  (.A(n1711gat), .B(n2437gat), .Z(n2556gat) ) ;
INV     gate1778  (.A(n2556gat), .Z(II3457) ) ;
INV     gate1779  (.A(n1898gat), .Z(n1956gat) ) ;
INV     gate1780  (.A(n1956gat), .Z(II3461) ) ;
INV     gate1781  (.A(II3461), .Z(n3038gat) ) ;
INV     gate1782  (.A(n3038gat), .Z(n1954gat) ) ;
INV     gate1783  (.A(n1886gat), .Z(II3465) ) ;
INV     gate1784  (.A(II3465), .Z(n3039gat) ) ;
INV     gate1785  (.A(n3039gat), .Z(n1888gat) ) ;
OR2     gate1786  (.A(n1954gat), .B(n1888gat), .Z(n2994gat) ) ;
INV     gate1787  (.A(n2994gat), .Z(n2048gat) ) ;
NOR2    gate1788  (.A(n2048gat), .B(n2437gat), .Z(n2539gat) ) ;
INV     gate1789  (.A(n2539gat), .Z(II3472) ) ;
INV     gate1790  (.A(n2142gat), .Z(n1969gat) ) ;
INV     gate1791  (.A(n2060gat), .Z(n1893gat) ) ;
OR3     gate1792  (.A(n1894gat), .B(n1847gat), .C(n1846gat), .Z(n2993gat) ) ;
INV     gate1793  (.A(n2993gat), .Z(n1892gat) ) ;
NOR2    gate1794  (.A(n2437gat), .B(n1892gat), .Z(n2436gat) ) ;
INV     gate1795  (.A(n2436gat), .Z(II3483) ) ;
OR2     gate1796  (.A(n2055gat), .B(n1967gat), .Z(n2998gat) ) ;
INV     gate1797  (.A(n2998gat), .Z(n2056gat) ) ;
NOR2    gate1798  (.A(n2056gat), .B(n2437gat), .Z(n2387gat) ) ;
INV     gate1799  (.A(n2387gat), .Z(II3491) ) ;
INV     gate1800  (.A(n1963gat), .Z(II3494) ) ;
INV     gate1801  (.A(II3494), .Z(n3043gat) ) ;
INV     gate1802  (.A(n3043gat), .Z(n1960gat) ) ;
INV     gate1803  (.A(n2138gat), .Z(n1887gat) ) ;
OR3     gate1804  (.A(n1960gat), .B(n1959gat), .C(n1957gat), .Z(n2996gat) ) ;
INV     gate1805  (.A(n2996gat), .Z(n1961gat) ) ;
NOR2    gate1806  (.A(n2437gat), .B(n1961gat), .Z(n2330gat) ) ;
INV     gate1807  (.A(n2330gat), .Z(II3504) ) ;
NOR2    gate1808  (.A(n2988gat), .B(n1855gat), .Z(n2147gat) ) ;
INV     gate1809  (.A(n2147gat), .Z(n2199gat) ) ;
INV     gate1810  (.A(n2438gat), .Z(II3509) ) ;
INV     gate1811  (.A(II3509), .Z(n3045gat) ) ;
INV     gate1812  (.A(n3045gat), .Z(n2332gat) ) ;
INV     gate1813  (.A(n2439gat), .Z(II3513) ) ;
INV     gate1814  (.A(II3513), .Z(n3046gat) ) ;
INV     gate1815  (.A(n3046gat), .Z(n2259gat) ) ;
OR2     gate1816  (.A(n2332gat), .B(n2259gat), .Z(n3008gat) ) ;
INV     gate1817  (.A(n3008gat), .Z(n2328gat) ) ;
NOR2    gate1818  (.A(n2199gat), .B(n2328gat), .Z(n2498gat) ) ;
INV     gate1819  (.A(n2498gat), .Z(II3520) ) ;
NOR2    gate1820  (.A(n2393gat), .B(n2439gat), .Z(n2193gat) ) ;
INV     gate1821  (.A(n2193gat), .Z(n2151gat) ) ;
OR2     gate1822  (.A(n2211gat), .B(n2210gat), .Z(n3005gat) ) ;
INV     gate1823  (.A(n3005gat), .Z(n2209gat) ) ;
NOR2    gate1824  (.A(n2199gat), .B(n2209gat), .Z(n2396gat) ) ;
INV     gate1825  (.A(n2396gat), .Z(II3530) ) ;
INV     gate1826  (.A(n2393gat), .Z(n2052gat) ) ;
OR3     gate1827  (.A(n2053gat), .B(n2052gat), .C(n1964gat), .Z(n2997gat) ) ;
INV     gate1828  (.A(n2997gat), .Z(n2058gat) ) ;
NOR2    gate1829  (.A(n2199gat), .B(n2058gat), .Z(n2198gat) ) ;
INV     gate1830  (.A(n2198gat), .Z(II3539) ) ;
NOR3    gate1831  (.A(n2346gat), .B(n2151gat), .C(n2402gat), .Z(n2215gat) ) ;
INV     gate1832  (.A(n2215gat), .Z(n2349gat) ) ;
OR2     gate1833  (.A(n2350gat), .B(n2282gat), .Z(n3009gat) ) ;
INV     gate1834  (.A(n3009gat), .Z(n2281gat) ) ;
NOR2    gate1835  (.A(n2199gat), .B(n2281gat), .Z(n2197gat) ) ;
INV     gate1836  (.A(n2197gat), .Z(II3549) ) ;
OR3     gate1837  (.A(n2213gat), .B(n2150gat), .C(n2149gat), .Z(n3002gat) ) ;
INV     gate1838  (.A(n3002gat), .Z(n2146gat) ) ;
NOR2    gate1839  (.A(n2199gat), .B(n2146gat), .Z(n2196gat) ) ;
INV     gate1840  (.A(n2196gat), .Z(II3558) ) ;
INV     gate1841  (.A(n2125gat), .Z(II3587) ) ;
INV     gate1842  (.A(II3587), .Z(n2124gat) ) ;
INV     gate1843  (.A(n2117gat), .Z(n2115gat) ) ;
NOR3    gate1844  (.A(n2124gat), .B(n2115gat), .C(n2239gat), .Z(n1882gat) ) ;
INV     gate1845  (.A(n1882gat), .Z(II3610) ) ;
INV     gate1846  (.A(n1975gat), .Z(II3621) ) ;
INV     gate1847  (.A(II3621), .Z(n1974gat) ) ;
INV     gate1848  (.A(n1956gat), .Z(n1955gat) ) ;
NOR2    gate1849  (.A(n2995gat), .B(n1895gat), .Z(n1896gat) ) ;
INV     gate1850  (.A(n1896gat), .Z(n1970gat) ) ;
INV     gate1851  (.A(n1975gat), .Z(n1973gat) ) ;
NOR2    gate1852  (.A(n2999gat), .B(n2437gat), .Z(n2559gat) ) ;
INV     gate1853  (.A(n2559gat), .Z(n2558gat) ) ;
INV     gate1854  (.A(n2558gat), .Z(II3635) ) ;
INV     gate1855  (.A(n2644gat), .Z(II3646) ) ;
INV     gate1856  (.A(II3646), .Z(n2643gat) ) ;
INV     gate1857  (.A(n2438gat), .Z(n2333gat) ) ;
NOR2    gate1858  (.A(n3011gat), .B(n2215gat), .Z(n2352gat) ) ;
INV     gate1859  (.A(n2352gat), .Z(n2564gat) ) ;
INV     gate1860  (.A(n2644gat), .Z(n2642gat) ) ;
NOR2    gate1861  (.A(n3015gat), .B(n2199gat), .Z(n2637gat) ) ;
INV     gate1862  (.A(n2637gat), .Z(n2636gat) ) ;
INV     gate1863  (.A(n2636gat), .Z(II3660) ) ;
NOR3    gate1864  (.A(n296gat), .B(n17gat), .C(n294gat), .Z(n84gat) ) ;
INV     gate1865  (.A(n84gat), .Z(n88gat) ) ;
NOR2    gate1866  (.A(n182gat), .B(n89gat), .Z(n110gat) ) ;
INV     gate1867  (.A(n110gat), .Z(n375gat) ) ;
INV     gate1868  (.A(n156gat), .Z(II3677) ) ;
INV     gate1869  (.A(II3677), .Z(n155gat) ) ;
NOR2    gate1870  (.A(n3024gat), .B(n1615gat), .Z(n1702gat) ) ;
INV     gate1871  (.A(n1702gat), .Z(n253gat) ) ;
INV     gate1872  (.A(n152gat), .Z(n150gat) ) ;
INV     gate1873  (.A(n152gat), .Z(II3691) ) ;
INV     gate1874  (.A(II3691), .Z(n151gat) ) ;
INV     gate1875  (.A(n1702gat), .Z(n243gat) ) ;
INV     gate1876  (.A(n243gat), .Z(n233gat) ) ;
INV     gate1877  (.A(n156gat), .Z(n154gat) ) ;
OR3     gate1878  (.A(n141gat), .B(n38gat), .C(n37gat), .Z(n2874gat) ) ;
INV     gate1879  (.A(n2874gat), .Z(n800gat) ) ;
OR2     gate1880  (.A(n1074gat), .B(n872gat), .Z(n2917gat) ) ;
INV     gate1881  (.A(n2917gat), .Z(II3703) ) ;
OR2     gate1882  (.A(n234gat), .B(n137gat), .Z(n2878gat) ) ;
INV     gate1883  (.A(n2878gat), .Z(n235gat) ) ;
OR2     gate1884  (.A(n378gat), .B(n377gat), .Z(n2892gat) ) ;
INV     gate1885  (.A(n2892gat), .Z(II3713) ) ;
NOR2    gate1886  (.A(n182gat), .B(n78gat), .Z(n212gat) ) ;
INV     gate1887  (.A(n212gat), .Z(n372gat) ) ;
INV     gate1888  (.A(n331gat), .Z(n329gat) ) ;
INV     gate1889  (.A(n388gat), .Z(II3736) ) ;
INV     gate1890  (.A(II3736), .Z(n387gat) ) ;
NOR2    gate1891  (.A(n1701gat), .B(n3023gat), .Z(n1700gat) ) ;
INV     gate1892  (.A(n1700gat), .Z(n334gat) ) ;
INV     gate1893  (.A(n388gat), .Z(n386gat) ) ;
INV     gate1894  (.A(n331gat), .Z(II3742) ) ;
INV     gate1895  (.A(II3742), .Z(n330gat) ) ;
INV     gate1896  (.A(n1700gat), .Z(n1430gat) ) ;
INV     gate1897  (.A(n1430gat), .Z(n1490gat) ) ;
OR3     gate1898  (.A(n250gat), .B(n249gat), .C(n248gat), .Z(n2885gat) ) ;
INV     gate1899  (.A(n2885gat), .Z(n452gat) ) ;
OR3     gate1900  (.A(n869gat), .B(n453gat), .C(n448gat), .Z(n2900gat) ) ;
INV     gate1901  (.A(n2900gat), .Z(II3754) ) ;
OR2     gate1902  (.A(n251gat), .B(n244gat), .Z(n2883gat) ) ;
INV     gate1903  (.A(n2883gat), .Z(n333gat) ) ;
OR3     gate1904  (.A(n974gat), .B(n973gat), .C(n870gat), .Z(n2929gat) ) ;
INV     gate1905  (.A(n2929gat), .Z(II3765) ) ;
INV     gate1906  (.A(n463gat), .Z(II3777) ) ;
INV     gate1907  (.A(II3777), .Z(n462gat) ) ;
INV     gate1908  (.A(n327gat), .Z(n325gat) ) ;
OR2     gate1909  (.A(n246gat), .B(n245gat), .Z(n2884gat) ) ;
INV     gate1910  (.A(n2884gat), .Z(n457gat) ) ;
INV     gate1911  (.A(n463gat), .Z(n461gat) ) ;
OR2     gate1912  (.A(n460gat), .B(n459gat), .Z(n2902gat) ) ;
INV     gate1913  (.A(n2902gat), .Z(n458gat) ) ;
OR3     gate1914  (.A(n975gat), .B(n972gat), .C(n969gat), .Z(n2925gat) ) ;
INV     gate1915  (.A(n2925gat), .Z(II3801) ) ;
NOR3    gate1916  (.A(n334gat), .B(n387gat), .C(n330gat), .Z(n247gat) ) ;
INV     gate1917  (.A(n247gat), .Z(n144gat) ) ;
INV     gate1918  (.A(n327gat), .Z(II3808) ) ;
INV     gate1919  (.A(II3808), .Z(n326gat) ) ;
OR2     gate1920  (.A(n145gat), .B(n143gat), .Z(n2879gat) ) ;
INV     gate1921  (.A(n2879gat), .Z(n878gat) ) ;
OR3     gate1922  (.A(n971gat), .B(n970gat), .C(n968gat), .Z(n2916gat) ) ;
INV     gate1923  (.A(n2916gat), .Z(II3817) ) ;
INV     gate1924  (.A(n384gat), .Z(n382gat) ) ;
INV     gate1925  (.A(n384gat), .Z(II3831) ) ;
INV     gate1926  (.A(II3831), .Z(n383gat) ) ;
OR3     gate1927  (.A(n142gat), .B(n40gat), .C(n39gat), .Z(n2875gat) ) ;
INV     gate1928  (.A(n2875gat), .Z(n134gat) ) ;
OR3     gate1929  (.A(n772gat), .B(n451gat), .C(n446gat), .Z(n2899gat) ) ;
INV     gate1930  (.A(n2899gat), .Z(II3841) ) ;
INV     gate1931  (.A(n256gat), .Z(n254gat) ) ;
OR2     gate1932  (.A(n139gat), .B(n136gat), .Z(n2877gat) ) ;
INV     gate1933  (.A(n2877gat), .Z(n252gat) ) ;
INV     gate1934  (.A(n470gat), .Z(n468gat) ) ;
INV     gate1935  (.A(n470gat), .Z(II3867) ) ;
INV     gate1936  (.A(II3867), .Z(n469gat) ) ;
OR2     gate1937  (.A(n391gat), .B(n390gat), .Z(n2893gat) ) ;
INV     gate1938  (.A(n2893gat), .Z(n381gat) ) ;
OR2     gate1939  (.A(n1083gat), .B(n1077gat), .Z(n2926gat) ) ;
INV     gate1940  (.A(n2926gat), .Z(II3876) ) ;
NOR3    gate1941  (.A(n151gat), .B(n253gat), .C(n155gat), .Z(n140gat) ) ;
INV     gate1942  (.A(n140gat), .Z(n241gat) ) ;
INV     gate1943  (.A(n256gat), .Z(II3882) ) ;
INV     gate1944  (.A(II3882), .Z(n255gat) ) ;
OR2     gate1945  (.A(n242gat), .B(n240gat), .Z(n2882gat) ) ;
INV     gate1946  (.A(n2882gat), .Z(n802gat) ) ;
OR2     gate1947  (.A(n871gat), .B(n797gat), .Z(n2924gat) ) ;
INV     gate1948  (.A(n2924gat), .Z(II3891) ) ;
INV     gate1949  (.A(n148gat), .Z(n146gat) ) ;
INV     gate1950  (.A(n148gat), .Z(II3904) ) ;
INV     gate1951  (.A(II3904), .Z(n147gat) ) ;
OR3     gate1952  (.A(n324gat), .B(n238gat), .C(n237gat), .Z(n2881gat) ) ;
INV     gate1953  (.A(n2881gat), .Z(n380gat) ) ;
OR2     gate1954  (.A(n1082gat), .B(n796gat), .Z(n2923gat) ) ;
INV     gate1955  (.A(n2923gat), .Z(II3914) ) ;
NOR2    gate1956  (.A(n85gat), .B(n180gat), .Z(n68gat) ) ;
INV     gate1957  (.A(n68gat), .Z(n69gat) ) ;
INV     gate1958  (.A(n2048gat), .Z(n1885gat) ) ;
OR2     gate1959  (.A(n69gat), .B(n1885gat), .Z(n2710gat) ) ;
INV     gate1960  (.A(n2710gat), .Z(II3923) ) ;
INV     gate1961  (.A(II3923), .Z(n2707gat) ) ;
INV     gate1962  (.A(n564gat), .Z(n16gat) ) ;
NOR2    gate1963  (.A(n2726gat), .B(n2860gat), .Z(n357gat) ) ;
INV     gate1964  (.A(n357gat), .Z(n295gat) ) ;
NOR2    gate1965  (.A(n186gat), .B(n82gat), .Z(n12gat) ) ;
INV     gate1966  (.A(n12gat), .Z(n11gat) ) ;
INV     gate1967  (.A(n1961gat), .Z(n1889gat) ) ;
OR2     gate1968  (.A(n11gat), .B(n1889gat), .Z(n2704gat) ) ;
INV     gate1969  (.A(n2704gat), .Z(II3935) ) ;
INV     gate1970  (.A(II3935), .Z(n2700gat) ) ;
INV     gate1971  (.A(n2056gat), .Z(n2051gat) ) ;
OR2     gate1972  (.A(n1599gat), .B(n2051gat), .Z(n2684gat) ) ;
INV     gate1973  (.A(n2684gat), .Z(II3941) ) ;
INV     gate1974  (.A(II3941), .Z(n2680gat) ) ;
INV     gate1975  (.A(n1831gat), .Z(n1350gat) ) ;
INV     gate1976  (.A(n1350gat), .Z(II3945) ) ;
INV     gate1977  (.A(II3945), .Z(n2696gat) ) ;
INV     gate1978  (.A(n2696gat), .Z(II3948) ) ;
INV     gate1979  (.A(II3948), .Z(n2692gat) ) ;
INV     gate1980  (.A(n2448gat), .Z(II3951) ) ;
INV     gate1981  (.A(II3951), .Z(n2683gat) ) ;
INV     gate1982  (.A(n2683gat), .Z(II3954) ) ;
INV     gate1983  (.A(II3954), .Z(n2679gat) ) ;
INV     gate1984  (.A(n2450gat), .Z(II3957) ) ;
INV     gate1985  (.A(II3957), .Z(n2449gat) ) ;
INV     gate1986  (.A(n2449gat), .Z(n1754gat) ) ;
OR2     gate1987  (.A(n2444gat), .B(n1754gat), .Z(n2830gat) ) ;
INV     gate1988  (.A(n2830gat), .Z(II3962) ) ;
INV     gate1989  (.A(II3962), .Z(n2827gat) ) ;
INV     gate1990  (.A(n2514gat), .Z(n2512gat) ) ;
INV     gate1991  (.A(n1625gat), .Z(n1544gat) ) ;
INV     gate1992  (.A(n1771gat), .Z(n1769gat) ) ;
NOR3    gate1993  (.A(n2512gat), .B(n1769gat), .C(n1773gat), .Z(n1756gat) ) ;
INV     gate1994  (.A(n1756gat), .Z(n1683gat) ) ;
INV     gate1995  (.A(n2169gat), .Z(n2167gat) ) ;
OR4     gate1996  (.A(n2108gat), .B(n2093gat), .C(n2035gat), .D(II3999), .Z(II4000) ) ;
INV     gate1997  (.A(II4000), .Z(n2013gat) ) ;
INV     gate1998  (.A(n2013gat), .Z(n1791gat) ) ;
OR2     gate1999  (.A(n1586gat), .B(n1791gat), .Z(n2695gat) ) ;
INV     gate2000  (.A(n2695gat), .Z(n2691gat) ) ;
INV     gate2001  (.A(n1694gat), .Z(n1518gat) ) ;
OR2     gate2002  (.A(n1755gat), .B(n1518gat), .Z(n2703gat) ) ;
INV     gate2003  (.A(n2703gat), .Z(n2699gat) ) ;
INV     gate2004  (.A(n1412gat), .Z(n2159gat) ) ;
INV     gate2005  (.A(n2579gat), .Z(n2478gat) ) ;
OR2     gate2006  (.A(n2159gat), .B(n2478gat), .Z(n2744gat) ) ;
INV     gate2007  (.A(n2744gat), .Z(II4014) ) ;
INV     gate2008  (.A(II4014), .Z(n2740gat) ) ;
INV     gate2009  (.A(n1412gat), .Z(n2158gat) ) ;
INV     gate2010  (.A(n2613gat), .Z(n2186gat) ) ;
OR2     gate2011  (.A(n2158gat), .B(n2186gat), .Z(n2800gat) ) ;
INV     gate2012  (.A(n2800gat), .Z(II4020) ) ;
INV     gate2013  (.A(II4020), .Z(n2797gat) ) ;
OR3     gate2014  (.A(n2353gat), .B(n2284gat), .C(II4023), .Z(II4024) ) ;
INV     gate2015  (.A(II4024), .Z(n2288gat) ) ;
INV     gate2016  (.A(n2288gat), .Z(n1513gat) ) ;
NOR3    gate2017  (.A(n2620gat), .B(n2625gat), .C(n2488gat), .Z(n2538gat) ) ;
INV     gate2018  (.A(n2538gat), .Z(n2537gat) ) ;
NOR3    gate2019  (.A(n2537gat), .B(n2482gat), .C(n2486gat), .Z(n2483gat) ) ;
INV     gate2020  (.A(n2483gat), .Z(n2442gat) ) ;
INV     gate2021  (.A(n1336gat), .Z(n1334gat) ) ;
INV     gate2022  (.A(n1748gat), .Z(II4055) ) ;
INV     gate2023  (.A(II4055), .Z(n1747gat) ) ;
INV     gate2024  (.A(n1675gat), .Z(II4067) ) ;
INV     gate2025  (.A(II4067), .Z(n1674gat) ) ;
NOR3    gate2026  (.A(n1858gat), .B(n1393gat), .C(n1604gat), .Z(n1402gat) ) ;
INV     gate2027  (.A(n1402gat), .Z(n1403gat) ) ;
INV     gate2028  (.A(n1807gat), .Z(II4081) ) ;
INV     gate2029  (.A(II4081), .Z(n1806gat) ) ;
INV     gate2030  (.A(n1712gat), .Z(n1634gat) ) ;
INV     gate2031  (.A(n1340gat), .Z(n1338gat) ) ;
INV     gate2032  (.A(n1456gat), .Z(II4105) ) ;
INV     gate2033  (.A(II4105), .Z(n1455gat) ) ;
INV     gate2034  (.A(n1340gat), .Z(II4108) ) ;
INV     gate2035  (.A(II4108), .Z(n1339gat) ) ;
OR4     gate2036  (.A(n1470gat), .B(n1400gat), .C(n1399gat), .D(n1398gat), .Z(n2980gat) ) ;
INV     gate2037  (.A(n2980gat), .Z(n1505gat) ) ;
INV     gate2038  (.A(n1505gat), .Z(II4117) ) ;
INV     gate2039  (.A(II4117), .Z(n2758gat) ) ;
INV     gate2040  (.A(n2758gat), .Z(n2755gat) ) ;
INV     gate2041  (.A(n2980gat), .Z(n1546gat) ) ;
INV     gate2042  (.A(n1546gat), .Z(II4122) ) ;
INV     gate2043  (.A(II4122), .Z(n2752gat) ) ;
INV     gate2044  (.A(n2752gat), .Z(n2748gat) ) ;
NOR2    gate2045  (.A(n2019gat), .B(n1878gat), .Z(n2016gat) ) ;
INV     gate2046  (.A(n2016gat), .Z(n2012gat) ) ;
NOR2    gate2047  (.A(n2012gat), .B(n1774gat), .Z(n2008gat) ) ;
INV     gate2048  (.A(n2008gat), .Z(n2002gat) ) ;
INV     gate2049  (.A(n3097gat), .Z(II4129) ) ;
INV     gate2050  (.A(II4129), .Z(n2858gat) ) ;
INV     gate2051  (.A(n2858gat), .Z(n2857gat) ) ;
INV     gate2052  (.A(n3098gat), .Z(II4135) ) ;
INV     gate2053  (.A(II4135), .Z(n2766gat) ) ;
INV     gate2054  (.A(n2766gat), .Z(II4138) ) ;
INV     gate2055  (.A(II4138), .Z(n2765gat) ) ;
NOR3    gate2056  (.A(n1818gat), .B(n1935gat), .C(n2765gat), .Z(n1759gat) ) ;
INV     gate2057  (.A(n1759gat), .Z(n1684gat) ) ;
OR3     gate2058  (.A(n1788gat), .B(n1784gat), .C(II4144), .Z(II4145) ) ;
INV     gate2059  (.A(n1525gat), .Z(II4157) ) ;
INV     gate2060  (.A(II4157), .Z(n1524gat) ) ;
NOR3    gate2061  (.A(n1991gat), .B(n2283gat), .C(n1989gat), .Z(n1863gat) ) ;
INV     gate2062  (.A(n1863gat), .Z(n1862gat) ) ;
NOR3    gate2063  (.A(n1988gat), .B(n2216gat), .C(n1862gat), .Z(n1860gat) ) ;
INV     gate2064  (.A(n1860gat), .Z(n1919gat) ) ;
INV     gate2065  (.A(n1462gat), .Z(n1460gat) ) ;
INV     gate2066  (.A(n1596gat), .Z(II4185) ) ;
INV     gate2067  (.A(II4185), .Z(n1595gat) ) ;
NOR2    gate2068  (.A(n1858gat), .B(n1608gat), .Z(n1469gat) ) ;
INV     gate2069  (.A(n1469gat), .Z(n1454gat) ) ;
NOR3    gate2070  (.A(n1584gat), .B(n1339gat), .C(n1600gat), .Z(n1519gat) ) ;
INV     gate2071  (.A(n1519gat), .Z(n1468gat) ) ;
INV     gate2072  (.A(n1462gat), .Z(II4194) ) ;
INV     gate2073  (.A(II4194), .Z(n1461gat) ) ;
OR2     gate2074  (.A(n1467gat), .B(n1466gat), .Z(n2984gat) ) ;
INV     gate2075  (.A(n2984gat), .Z(n1477gat) ) ;
INV     gate2076  (.A(n1596gat), .Z(n1594gat) ) ;
INV     gate2077  (.A(n1588gat), .Z(II4212) ) ;
INV     gate2078  (.A(II4212), .Z(n1587gat) ) ;
OR3     gate2079  (.A(n1392gat), .B(n2989gat), .C(II4216), .Z(II4217) ) ;
INV     gate2080  (.A(II4217), .Z(n1681gat) ) ;
NOR3    gate2081  (.A(n2985gat), .B(n1602gat), .C(n1681gat), .Z(n1761gat) ) ;
INV     gate2082  (.A(n1761gat), .Z(II4222) ) ;
INV     gate2083  (.A(II4222), .Z(n2751gat) ) ;
INV     gate2084  (.A(n2751gat), .Z(n2747gat) ) ;
NOR3    gate2085  (.A(n1681gat), .B(n1602gat), .C(n2985gat), .Z(n1760gat) ) ;
INV     gate2086  (.A(n1760gat), .Z(II4227) ) ;
INV     gate2087  (.A(II4227), .Z(n2743gat) ) ;
INV     gate2088  (.A(n2743gat), .Z(n2739gat) ) ;
INV     gate2089  (.A(n2286gat), .Z(n1978gat) ) ;
NOR3    gate2090  (.A(n2442gat), .B(n1690gat), .C(n1978gat), .Z(n1721gat) ) ;
INV     gate2091  (.A(n1721gat), .Z(II4233) ) ;
INV     gate2092  (.A(II4233), .Z(n2808gat) ) ;
INV     gate2093  (.A(n2808gat), .Z(II4236) ) ;
INV     gate2094  (.A(II4236), .Z(n2804gat) ) ;
NOR2    gate2095  (.A(n520gat), .B(n519gat), .Z(n518gat) ) ;
INV     gate2096  (.A(n518gat), .Z(n517gat) ) ;
NOR2    gate2097  (.A(n374gat), .B(n2723gat), .Z(n418gat) ) ;
INV     gate2098  (.A(n418gat), .Z(n417gat) ) ;
NOR2    gate2099  (.A(n374gat), .B(n2726gat), .Z(n411gat) ) ;
INV     gate2100  (.A(n411gat), .Z(n413gat) ) ;
NOR2    gate2101  (.A(n374gat), .B(n2859gat), .Z(n522gat) ) ;
INV     gate2102  (.A(n522gat), .Z(n412gat) ) ;
NOR2    gate2103  (.A(n374gat), .B(n2715gat), .Z(n516gat) ) ;
INV     gate2104  (.A(n516gat), .Z(n406gat) ) ;
NOR3    gate2105  (.A(n517gat), .B(n410gat), .C(n354gat), .Z(n355gat) ) ;
INV     gate2106  (.A(n355gat), .Z(n407gat) ) ;
NOR3    gate2107  (.A(n526gat), .B(n531gat), .C(n530gat), .Z(n525gat) ) ;
INV     gate2108  (.A(n525gat), .Z(n290gat) ) ;
NOR2    gate2109  (.A(n2726gat), .B(n740gat), .Z(n356gat) ) ;
INV     gate2110  (.A(n356gat), .Z(n527gat) ) ;
NOR2    gate2111  (.A(n2723gat), .B(n740gat), .Z(n415gat) ) ;
INV     gate2112  (.A(n415gat), .Z(n416gat) ) ;
NOR2    gate2113  (.A(n740gat), .B(n2715gat), .Z(n521gat) ) ;
INV     gate2114  (.A(n521gat), .Z(n528gat) ) ;
NOR3    gate2115  (.A(n527gat), .B(n416gat), .C(n528gat), .Z(n532gat) ) ;
INV     gate2116  (.A(n532gat), .Z(n358gat) ) ;
NOR2    gate2117  (.A(n522gat), .B(n356gat), .Z(n523gat) ) ;
INV     gate2118  (.A(n523gat), .Z(n639gat) ) ;
NOR3    gate2119  (.A(n639gat), .B(n634gat), .C(n414gat), .Z(n635gat) ) ;
INV     gate2120  (.A(n635gat), .Z(n1111gat) ) ;
NOR2    gate2121  (.A(n411gat), .B(n415gat), .Z(n414gat) ) ;
INV     gate2122  (.A(n414gat), .Z(n524gat) ) ;
NOR3    gate2123  (.A(n634gat), .B(n523gat), .C(n524gat), .Z(n630gat) ) ;
INV     gate2124  (.A(n630gat), .Z(n1112gat) ) ;
NOR3    gate2125  (.A(n414gat), .B(n634gat), .C(n523gat), .Z(n629gat) ) ;
INV     gate2126  (.A(n629gat), .Z(n741gat) ) ;
NOR2    gate2127  (.A(n418gat), .B(n521gat), .Z(n634gat) ) ;
INV     gate2128  (.A(n634gat), .Z(n633gat) ) ;
NOR3    gate2129  (.A(n414gat), .B(n523gat), .C(n633gat), .Z(n632gat) ) ;
INV     gate2130  (.A(n632gat), .Z(n926gat) ) ;
NOR3    gate2131  (.A(n414gat), .B(n633gat), .C(n639gat), .Z(n636gat) ) ;
INV     gate2132  (.A(n636gat), .Z(n670gat) ) ;
INV     gate2133  (.A(n632gat), .Z(n1123gat) ) ;
INV     gate2134  (.A(n635gat), .Z(n1007gat) ) ;
INV     gate2135  (.A(n630gat), .Z(n1006gat) ) ;
OR2     gate2136  (.A(n1003gat), .B(n902gat), .Z(n2941gat) ) ;
INV     gate2137  (.A(n2941gat), .Z(II4309) ) ;
INV     gate2138  (.A(II4309), .Z(n2814gat) ) ;
INV     gate2139  (.A(n2814gat), .Z(II4312) ) ;
INV     gate2140  (.A(II4312), .Z(n2811gat) ) ;
OR4     gate2141  (.A(n1099gat), .B(n998gat), .C(n995gat), .D(n980gat), .Z(n2946gat) ) ;
INV     gate2142  (.A(n2946gat), .Z(n1002gat) ) ;
OR2     gate2143  (.A(n1001gat), .B(n999gat), .Z(n2950gat) ) ;
INV     gate2144  (.A(n2950gat), .Z(II4329) ) ;
INV     gate2145  (.A(II4329), .Z(n2813gat) ) ;
INV     gate2146  (.A(n2813gat), .Z(II4332) ) ;
INV     gate2147  (.A(II4332), .Z(n2810gat) ) ;
OR4     gate2148  (.A(n981gat), .B(n890gat), .C(n889gat), .D(n886gat), .Z(n2933gat) ) ;
INV     gate2149  (.A(n2933gat), .Z(n888gat) ) ;
OR2     gate2150  (.A(n892gat), .B(n891gat), .Z(n2935gat) ) ;
INV     gate2151  (.A(n2935gat), .Z(II4349) ) ;
INV     gate2152  (.A(II4349), .Z(n2818gat) ) ;
INV     gate2153  (.A(n2818gat), .Z(II4352) ) ;
INV     gate2154  (.A(II4352), .Z(n2816gat) ) ;
OR4     gate2155  (.A(n1152gat), .B(n1092gat), .C(n997gat), .D(n993gat), .Z(n2940gat) ) ;
INV     gate2156  (.A(n2940gat), .Z(n898gat) ) ;
OR2     gate2157  (.A(n900gat), .B(n895gat), .Z(n2937gat) ) ;
INV     gate2158  (.A(n2937gat), .Z(II4369) ) ;
INV     gate2159  (.A(II4369), .Z(n2817gat) ) ;
INV     gate2160  (.A(n2817gat), .Z(II4372) ) ;
INV     gate2161  (.A(II4372), .Z(n2815gat) ) ;
OR4     gate2162  (.A(n1094gat), .B(n1093gat), .C(n988gat), .D(n984gat), .Z(n2947gat) ) ;
INV     gate2163  (.A(n2947gat), .Z(n1179gat) ) ;
OR2     gate2164  (.A(n1178gat), .B(n1116gat), .Z(n2956gat) ) ;
INV     gate2165  (.A(n2956gat), .Z(II4389) ) ;
INV     gate2166  (.A(II4389), .Z(n2824gat) ) ;
INV     gate2167  (.A(n2824gat), .Z(II4392) ) ;
INV     gate2168  (.A(II4392), .Z(n2821gat) ) ;
OR4     gate2169  (.A(n1091gat), .B(n1088gat), .C(n992gat), .D(n987gat), .Z(n2939gat) ) ;
INV     gate2170  (.A(n2939gat), .Z(n897gat) ) ;
OR2     gate2171  (.A(n899gat), .B(n896gat), .Z(n2938gat) ) ;
INV     gate2172  (.A(n2938gat), .Z(II4409) ) ;
INV     gate2173  (.A(II4409), .Z(n2823gat) ) ;
INV     gate2174  (.A(n2823gat), .Z(II4412) ) ;
INV     gate2175  (.A(II4412), .Z(n2820gat) ) ;
OR4     gate2176  (.A(n1098gat), .B(n1090gat), .C(n986gat), .D(n885gat), .Z(n2932gat) ) ;
INV     gate2177  (.A(n2932gat), .Z(n894gat) ) ;
OR2     gate2178  (.A(n901gat), .B(n893gat), .Z(n2936gat) ) ;
INV     gate2179  (.A(n2936gat), .Z(II4429) ) ;
INV     gate2180  (.A(II4429), .Z(n2829gat) ) ;
INV     gate2181  (.A(n2829gat), .Z(II4432) ) ;
INV     gate2182  (.A(II4432), .Z(n2826gat) ) ;
OR4     gate2183  (.A(n1097gat), .B(n1089gat), .C(n1087gat), .D(n991gat), .Z(n2948gat) ) ;
INV     gate2184  (.A(n2948gat), .Z(n1180gat) ) ;
OR2     gate2185  (.A(n1177gat), .B(n1115gat), .Z(n2955gat) ) ;
INV     gate2186  (.A(n2955gat), .Z(II4449) ) ;
INV     gate2187  (.A(II4449), .Z(n2828gat) ) ;
INV     gate2188  (.A(n2828gat), .Z(II4452) ) ;
INV     gate2189  (.A(II4452), .Z(n2825gat) ) ;
INV     gate2190  (.A(n673gat), .Z(n671gat) ) ;
NOR3    gate2191  (.A(n523gat), .B(n633gat), .C(n524gat), .Z(n631gat) ) ;
INV     gate2192  (.A(n631gat), .Z(n628gat) ) ;
INV     gate2193  (.A(n628gat), .Z(n976gat) ) ;
OR2     gate2194  (.A(n1004gat), .B(n1000gat), .Z(n2951gat) ) ;
INV     gate2195  (.A(n2951gat), .Z(II4475) ) ;
INV     gate2196  (.A(II4475), .Z(n2807gat) ) ;
INV     gate2197  (.A(n2807gat), .Z(II4478) ) ;
INV     gate2198  (.A(II4478), .Z(n2803gat) ) ;
INV     gate2199  (.A(n2389gat), .Z(n2127gat) ) ;
INV     gate2200  (.A(n2127gat), .Z(II4482) ) ;
INV     gate2201  (.A(II4482), .Z(n2682gat) ) ;
INV     gate2202  (.A(n2682gat), .Z(II4485) ) ;
INV     gate2203  (.A(II4485), .Z(n2678gat) ) ;
INV     gate2204  (.A(n2269gat), .Z(n2046gat) ) ;
INV     gate2205  (.A(n2046gat), .Z(II4489) ) ;
INV     gate2206  (.A(II4489), .Z(n2681gat) ) ;
INV     gate2207  (.A(n2681gat), .Z(II4492) ) ;
INV     gate2208  (.A(II4492), .Z(n2677gat) ) ;
INV     gate2209  (.A(n2338gat), .Z(n1708gat) ) ;
INV     gate2210  (.A(n1708gat), .Z(II4496) ) ;
INV     gate2211  (.A(II4496), .Z(n2688gat) ) ;
INV     gate2212  (.A(n2688gat), .Z(II4499) ) ;
INV     gate2213  (.A(II4499), .Z(n2686gat) ) ;
NOR2    gate2214  (.A(n290gat), .B(n292gat), .Z(n291gat) ) ;
INV     gate2215  (.A(n291gat), .Z(n455gat) ) ;
INV     gate2216  (.A(n2646gat), .Z(n2237gat) ) ;
OR2     gate2217  (.A(n1029gat), .B(n2237gat), .Z(n2764gat) ) ;
INV     gate2218  (.A(n2764gat), .Z(II4506) ) ;
INV     gate2219  (.A(II4506), .Z(n2763gat) ) ;
INV     gate2220  (.A(n2971gat), .Z(n1782gat) ) ;
OR2     gate2221  (.A(n1028gat), .B(n1782gat), .Z(n2762gat) ) ;
INV     gate2222  (.A(n2762gat), .Z(II4512) ) ;
INV     gate2223  (.A(II4512), .Z(n2760gat) ) ;
INV     gate2224  (.A(n3010gat), .Z(n2325gat) ) ;
OR2     gate2225  (.A(n1031gat), .B(n2325gat), .Z(n2761gat) ) ;
INV     gate2226  (.A(n2761gat), .Z(II4518) ) ;
INV     gate2227  (.A(II4518), .Z(n2759gat) ) ;
INV     gate2228  (.A(n504gat), .Z(n2245gat) ) ;
OR2     gate2229  (.A(n1030gat), .B(n2245gat), .Z(n2757gat) ) ;
INV     gate2230  (.A(n2757gat), .Z(II4524) ) ;
INV     gate2231  (.A(II4524), .Z(n2754gat) ) ;
INV     gate2232  (.A(n567gat), .Z(n2244gat) ) ;
OR2     gate2233  (.A(n1011gat), .B(n2244gat), .Z(n2756gat) ) ;
INV     gate2234  (.A(n2756gat), .Z(II4530) ) ;
INV     gate2235  (.A(II4530), .Z(n2753gat) ) ;
INV     gate2236  (.A(n55gat), .Z(n2243gat) ) ;
OR2     gate2237  (.A(n1181gat), .B(n2243gat), .Z(n2750gat) ) ;
INV     gate2238  (.A(n2750gat), .Z(II4536) ) ;
INV     gate2239  (.A(II4536), .Z(n2746gat) ) ;
INV     gate2240  (.A(n933gat), .Z(n2246gat) ) ;
OR2     gate2241  (.A(n1010gat), .B(n2246gat), .Z(n2749gat) ) ;
INV     gate2242  (.A(n2749gat), .Z(II4542) ) ;
INV     gate2243  (.A(II4542), .Z(n2745gat) ) ;
INV     gate2244  (.A(n43gat), .Z(n2384gat) ) ;
OR2     gate2245  (.A(n1005gat), .B(n2384gat), .Z(n2742gat) ) ;
INV     gate2246  (.A(n2742gat), .Z(II4548) ) ;
INV     gate2247  (.A(II4548), .Z(n2738gat) ) ;
INV     gate2248  (.A(n748gat), .Z(n2385gat) ) ;
OR2     gate2249  (.A(n1182gat), .B(n2385gat), .Z(n2741gat) ) ;
INV     gate2250  (.A(n2741gat), .Z(II4554) ) ;
INV     gate2251  (.A(II4554), .Z(n2737gat) ) ;
INV     gate2252  (.A(n1269gat), .Z(n1286gat) ) ;
INV     gate2253  (.A(n1286gat), .Z(II4558) ) ;
INV     gate2254  (.A(II4558), .Z(n2687gat) ) ;
INV     gate2255  (.A(n2687gat), .Z(n2685gat) ) ;
INV     gate2256  (.A(n1224gat), .Z(n1328gat) ) ;
INV     gate2257  (.A(n1328gat), .Z(n1381gat) ) ;
INV     gate2258  (.A(n2184gat), .Z(n1384gat) ) ;
OR2     gate2259  (.A(n1381gat), .B(n1384gat), .Z(n2694gat) ) ;
INV     gate2260  (.A(n2694gat), .Z(II4566) ) ;
INV     gate2261  (.A(II4566), .Z(n2690gat) ) ;
INV     gate2262  (.A(n1280gat), .Z(n1382gat) ) ;
INV     gate2263  (.A(n1382gat), .Z(n1451gat) ) ;
INV     gate2264  (.A(n2187gat), .Z(n1453gat) ) ;
OR2     gate2265  (.A(n1451gat), .B(n1453gat), .Z(n2693gat) ) ;
INV     gate2266  (.A(n2693gat), .Z(II4573) ) ;
INV     gate2267  (.A(II4573), .Z(n2689gat) ) ;
INV     gate2268  (.A(n1133gat), .Z(n927gat) ) ;
INV     gate2269  (.A(n927gat), .Z(n925gat) ) ;
INV     gate2270  (.A(n2049gat), .Z(n1452gat) ) ;
OR2     gate2271  (.A(n925gat), .B(n1452gat), .Z(n2702gat) ) ;
INV     gate2272  (.A(n2702gat), .Z(II4580) ) ;
INV     gate2273  (.A(II4580), .Z(n2698gat) ) ;
INV     gate2274  (.A(n1043gat), .Z(n923gat) ) ;
INV     gate2275  (.A(n923gat), .Z(n921gat) ) ;
INV     gate2276  (.A(n2328gat), .Z(n1890gat) ) ;
OR2     gate2277  (.A(n921gat), .B(n1890gat), .Z(n2701gat) ) ;
INV     gate2278  (.A(n2701gat), .Z(II4587) ) ;
INV     gate2279  (.A(II4587), .Z(n2697gat) ) ;
INV     gate2280  (.A(n929gat), .Z(n850gat) ) ;
INV     gate2281  (.A(n850gat), .Z(n739gat) ) ;
INV     gate2282  (.A(n2058gat), .Z(n1841gat) ) ;
OR2     gate2283  (.A(n739gat), .B(n1841gat), .Z(n2709gat) ) ;
INV     gate2284  (.A(n2709gat), .Z(II4594) ) ;
INV     gate2285  (.A(II4594), .Z(n2706gat) ) ;
INV     gate2286  (.A(n1119gat), .Z(n922gat) ) ;
INV     gate2287  (.A(n922gat), .Z(n848gat) ) ;
INV     gate2288  (.A(n2209gat), .Z(n2047gat) ) ;
OR2     gate2289  (.A(n848gat), .B(n2047gat), .Z(n2708gat) ) ;
INV     gate2290  (.A(n2708gat), .Z(II4601) ) ;
INV     gate2291  (.A(II4601), .Z(n2705gat) ) ;
INV     gate2292  (.A(n1070gat), .Z(n924gat) ) ;
INV     gate2293  (.A(n924gat), .Z(n849gat) ) ;
INV     gate2294  (.A(n2146gat), .Z(n2050gat) ) ;
OR2     gate2295  (.A(n849gat), .B(n2050gat), .Z(n2799gat) ) ;
INV     gate2296  (.A(n2799gat), .Z(II4608) ) ;
INV     gate2297  (.A(II4608), .Z(n2796gat) ) ;
INV     gate2298  (.A(n1033gat), .Z(n1118gat) ) ;
INV     gate2299  (.A(n1118gat), .Z(n1032gat) ) ;
INV     gate2300  (.A(n2281gat), .Z(n2054gat) ) ;
OR2     gate2301  (.A(n1032gat), .B(n2054gat), .Z(n2798gat) ) ;
INV     gate2302  (.A(n2798gat), .Z(II4615) ) ;
INV     gate2303  (.A(II4615), .Z(n2795gat) ) ;
NOR2    gate2304  (.A(n1869gat), .B(n1757gat), .Z(n1745gat) ) ;
INV     gate2305  (.A(n1745gat), .Z(II4620) ) ;
INV     gate2306  (.A(II4620), .Z(n2806gat) ) ;
INV     gate2307  (.A(n2806gat), .Z(II4623) ) ;
INV     gate2308  (.A(II4623), .Z(n2802gat) ) ;
INV     gate2309  (.A(n1871gat), .Z(II4626) ) ;
INV     gate2310  (.A(II4626), .Z(n1870gat) ) ;
INV     gate2311  (.A(n1870gat), .Z(n1086gat) ) ;
INV     gate2312  (.A(n1086gat), .Z(II4630) ) ;
INV     gate2313  (.A(II4630), .Z(n2805gat) ) ;
INV     gate2314  (.A(n2805gat), .Z(II4633) ) ;
INV     gate2315  (.A(II4633), .Z(n2801gat) ) ;
NOR3    gate2316  (.A(n17gat), .B(n294gat), .C(n637gat), .Z(n85gat) ) ;
INV     gate2317  (.A(n85gat), .Z(n67gat) ) ;
NOR3    gate2318  (.A(n286gat), .B(n188gat), .C(n287gat), .Z(n180gat) ) ;
INV     gate2319  (.A(n180gat), .Z(n71gat) ) ;
INV     gate2320  (.A(n1892gat), .Z(n1840gat) ) ;
OR3     gate2321  (.A(n73gat), .B(n70gat), .C(n1840gat), .Z(n2812gat) ) ;
INV     gate2322  (.A(n2812gat), .Z(II4642) ) ;
INV     gate2323  (.A(II4642), .Z(n2809gat) ) ;
NOR3    gate2324  (.A(n16gat), .B(n295gat), .C(n637gat), .Z(n82gat) ) ;
INV     gate2325  (.A(n82gat), .Z(n76gat) ) ;
NOR3    gate2326  (.A(n189gat), .B(n287gat), .C(n288gat), .Z(n186gat) ) ;
INV     gate2327  (.A(n186gat), .Z(n14gat) ) ;
INV     gate2328  (.A(n1711gat), .Z(n1842gat) ) ;
OR3     gate2329  (.A(n77gat), .B(n13gat), .C(n1842gat), .Z(n2822gat) ) ;
INV     gate2330  (.A(n2822gat), .Z(II4651) ) ;
INV     gate2331  (.A(II4651), .Z(n2819gat) ) ;
INV     gate2332  (.A(n2819gat), .Z(II4654) ) ;
INV     gate2333  (.A(n2809gat), .Z(II4657) ) ;
INV     gate2334  (.A(n2801gat), .Z(II4660) ) ;
INV     gate2335  (.A(n2802gat), .Z(II4663) ) ;
INV     gate2336  (.A(n2795gat), .Z(II4666) ) ;
INV     gate2337  (.A(n2796gat), .Z(II4669) ) ;
INV     gate2338  (.A(n2705gat), .Z(II4672) ) ;
INV     gate2339  (.A(n2706gat), .Z(II4675) ) ;
INV     gate2340  (.A(n2697gat), .Z(II4678) ) ;
INV     gate2341  (.A(n2698gat), .Z(II4681) ) ;
INV     gate2342  (.A(n2689gat), .Z(II4684) ) ;
INV     gate2343  (.A(n2690gat), .Z(II4687) ) ;
INV     gate2344  (.A(n2685gat), .Z(II4690) ) ;
INV     gate2345  (.A(n2737gat), .Z(II4693) ) ;
INV     gate2346  (.A(n2738gat), .Z(II4696) ) ;
INV     gate2347  (.A(n2745gat), .Z(II4699) ) ;
INV     gate2348  (.A(n2746gat), .Z(II4702) ) ;
INV     gate2349  (.A(n2753gat), .Z(II4705) ) ;
INV     gate2350  (.A(n2754gat), .Z(II4708) ) ;
INV     gate2351  (.A(n2759gat), .Z(II4711) ) ;
INV     gate2352  (.A(n2760gat), .Z(II4714) ) ;
INV     gate2353  (.A(n2763gat), .Z(II4717) ) ;
INV     gate2354  (.A(n2686gat), .Z(II4720) ) ;
INV     gate2355  (.A(n2677gat), .Z(II4723) ) ;
INV     gate2356  (.A(n2678gat), .Z(II4726) ) ;
INV     gate2357  (.A(n2803gat), .Z(II4729) ) ;
INV     gate2358  (.A(n2825gat), .Z(II4732) ) ;
INV     gate2359  (.A(n2826gat), .Z(II4735) ) ;
INV     gate2360  (.A(n2820gat), .Z(II4738) ) ;
INV     gate2361  (.A(n2821gat), .Z(II4741) ) ;
INV     gate2362  (.A(n2815gat), .Z(II4744) ) ;
INV     gate2363  (.A(n2816gat), .Z(II4747) ) ;
INV     gate2364  (.A(n2810gat), .Z(II4750) ) ;
INV     gate2365  (.A(n2811gat), .Z(II4753) ) ;
INV     gate2366  (.A(n2804gat), .Z(II4756) ) ;
INV     gate2367  (.A(n2739gat), .Z(II4759) ) ;
INV     gate2368  (.A(n2747gat), .Z(II4762) ) ;
INV     gate2369  (.A(n2748gat), .Z(II4765) ) ;
INV     gate2370  (.A(n2755gat), .Z(II4768) ) ;
INV     gate2371  (.A(n2797gat), .Z(II4771) ) ;
INV     gate2372  (.A(n2740gat), .Z(II4774) ) ;
INV     gate2373  (.A(n2699gat), .Z(II4777) ) ;
INV     gate2374  (.A(n2691gat), .Z(II4780) ) ;
INV     gate2375  (.A(n2827gat), .Z(II4783) ) ;
INV     gate2376  (.A(n2679gat), .Z(II4786) ) ;
INV     gate2377  (.A(n2692gat), .Z(II4789) ) ;
INV     gate2378  (.A(n2680gat), .Z(II4792) ) ;
INV     gate2379  (.A(n2700gat), .Z(II4795) ) ;
INV     gate2380  (.A(n2707gat), .Z(II4798) ) ;
NOR2    gate2381  (.A(n373gat), .B(n2669gat), .Z(n648gat) ) ;
NOR2    gate2382  (.A(n2844gat), .B(n856gat), .Z(n442gat) ) ;
NOR3    gate2383  (.A(n1218gat), .B(n1219gat), .C(n1220gat), .Z(n1214gat) ) ;
NOR3    gate2384  (.A(n1218gat), .B(n1221gat), .C(n1222gat), .Z(n1215gat) ) ;
NOR3    gate2385  (.A(n1223gat), .B(n1219gat), .C(n1222gat), .Z(n1216gat) ) ;
NOR3    gate2386  (.A(n1223gat), .B(n1221gat), .C(n1220gat), .Z(n1217gat) ) ;
NOR2    gate2387  (.A(n2716gat), .B(n2867gat), .Z(n745gat) ) ;
NOR2    gate2388  (.A(n2715gat), .B(n2868gat), .Z(n638gat) ) ;
NOR2    gate2389  (.A(n2724gat), .B(n2726gat), .Z(n423gat) ) ;
NOR2    gate2390  (.A(n2723gat), .B(n2727gat), .Z(n362gat) ) ;
NOR3    gate2391  (.A(n753gat), .B(n754gat), .C(n755gat), .Z(n749gat) ) ;
NOR3    gate2392  (.A(n753gat), .B(n756gat), .C(n757gat), .Z(n750gat) ) ;
NOR3    gate2393  (.A(n758gat), .B(n754gat), .C(n757gat), .Z(n751gat) ) ;
NOR3    gate2394  (.A(n758gat), .B(n756gat), .C(n755gat), .Z(n752gat) ) ;
NOR3    gate2395  (.A(n263gat), .B(n264gat), .C(n265gat), .Z(n259gat) ) ;
NOR3    gate2396  (.A(n263gat), .B(n266gat), .C(n267gat), .Z(n260gat) ) ;
NOR3    gate2397  (.A(n268gat), .B(n264gat), .C(n267gat), .Z(n261gat) ) ;
NOR3    gate2398  (.A(n268gat), .B(n266gat), .C(n265gat), .Z(n262gat) ) ;
NOR3    gate2399  (.A(n1018gat), .B(n1019gat), .C(n1020gat), .Z(n1014gat) ) ;
NOR3    gate2400  (.A(n1018gat), .B(n1021gat), .C(n1022gat), .Z(n1015gat) ) ;
NOR3    gate2401  (.A(n1023gat), .B(n1019gat), .C(n1022gat), .Z(n1016gat) ) ;
NOR3    gate2402  (.A(n1023gat), .B(n1021gat), .C(n1020gat), .Z(n1017gat) ) ;
NOR3    gate2403  (.A(n480gat), .B(n481gat), .C(n482gat), .Z(n476gat) ) ;
NOR3    gate2404  (.A(n480gat), .B(n483gat), .C(n484gat), .Z(n477gat) ) ;
NOR3    gate2405  (.A(n485gat), .B(n481gat), .C(n484gat), .Z(n478gat) ) ;
NOR3    gate2406  (.A(n485gat), .B(n483gat), .C(n482gat), .Z(n479gat) ) ;
NOR3    gate2407  (.A(n48gat), .B(n49gat), .C(n50gat), .Z(n44gat) ) ;
NOR3    gate2408  (.A(n48gat), .B(n51gat), .C(n52gat), .Z(n45gat) ) ;
NOR3    gate2409  (.A(n53gat), .B(n49gat), .C(n52gat), .Z(n46gat) ) ;
NOR3    gate2410  (.A(n53gat), .B(n51gat), .C(n50gat), .Z(n47gat) ) ;
NOR3    gate2411  (.A(n172gat), .B(n173gat), .C(n174gat), .Z(n168gat) ) ;
NOR3    gate2412  (.A(n172gat), .B(n175gat), .C(n176gat), .Z(n169gat) ) ;
NOR3    gate2413  (.A(n177gat), .B(n173gat), .C(n176gat), .Z(n170gat) ) ;
NOR3    gate2414  (.A(n177gat), .B(n175gat), .C(n174gat), .Z(n171gat) ) ;
NOR3    gate2415  (.A(n911gat), .B(n912gat), .C(n913gat), .Z(n907gat) ) ;
NOR3    gate2416  (.A(n911gat), .B(n914gat), .C(n915gat), .Z(n908gat) ) ;
NOR3    gate2417  (.A(n916gat), .B(n912gat), .C(n915gat), .Z(n909gat) ) ;
NOR3    gate2418  (.A(n916gat), .B(n914gat), .C(n913gat), .Z(n910gat) ) ;
NOR3    gate2419  (.A(n348gat), .B(n349gat), .C(n350gat), .Z(n344gat) ) ;
NOR3    gate2420  (.A(n348gat), .B(n351gat), .C(n352gat), .Z(n345gat) ) ;
NOR3    gate2421  (.A(n353gat), .B(n349gat), .C(n352gat), .Z(n346gat) ) ;
NOR3    gate2422  (.A(n353gat), .B(n351gat), .C(n350gat), .Z(n347gat) ) ;
NOR3    gate2423  (.A(n60gat), .B(n61gat), .C(n62gat), .Z(n56gat) ) ;
NOR3    gate2424  (.A(n60gat), .B(n63gat), .C(n64gat), .Z(n57gat) ) ;
NOR3    gate2425  (.A(n65gat), .B(n61gat), .C(n64gat), .Z(n58gat) ) ;
NOR3    gate2426  (.A(n65gat), .B(n63gat), .C(n62gat), .Z(n59gat) ) ;
NOR2    gate2427  (.A(n373gat), .B(n2731gat), .Z(n768gat) ) ;
NOR2    gate2428  (.A(n856gat), .B(n2718gat), .Z(n655gat) ) ;
NOR2    gate2429  (.A(n856gat), .B(n2838gat), .Z(n963gat) ) ;
NOR2    gate2430  (.A(n2775gat), .B(n373gat), .Z(n868gat) ) ;
NOR2    gate2431  (.A(n856gat), .B(n2711gat), .Z(n962gat) ) ;
NOR2    gate2432  (.A(n373gat), .B(n2734gat), .Z(n959gat) ) ;
NOR3    gate2433  (.A(n949gat), .B(n950gat), .C(n951gat), .Z(n945gat) ) ;
NOR3    gate2434  (.A(n949gat), .B(n952gat), .C(n953gat), .Z(n946gat) ) ;
NOR3    gate2435  (.A(n954gat), .B(n950gat), .C(n953gat), .Z(n947gat) ) ;
NOR3    gate2436  (.A(n954gat), .B(n952gat), .C(n951gat), .Z(n948gat) ) ;
NOR2    gate2437  (.A(n2792gat), .B(n373gat), .Z(n647gat) ) ;
NOR2    gate2438  (.A(n856gat), .B(n2846gat), .Z(n441gat) ) ;
NOR2    gate2439  (.A(n373gat), .B(n2672gat), .Z(n967gat) ) ;
NOR2    gate2440  (.A(n2852gat), .B(n856gat), .Z(n792gat) ) ;
NOR3    gate2441  (.A(n1233gat), .B(n1234gat), .C(n1235gat), .Z(n1229gat) ) ;
NOR3    gate2442  (.A(n1233gat), .B(n1236gat), .C(n1237gat), .Z(n1230gat) ) ;
NOR3    gate2443  (.A(n1238gat), .B(n1234gat), .C(n1237gat), .Z(n1231gat) ) ;
NOR3    gate2444  (.A(n1238gat), .B(n1236gat), .C(n1235gat), .Z(n1232gat) ) ;
NOR2    gate2445  (.A(n2778gat), .B(n373gat), .Z(n443gat) ) ;
NOR2    gate2446  (.A(n856gat), .B(n2836gat), .Z(n439gat) ) ;
NOR2    gate2447  (.A(n2789gat), .B(n373gat), .Z(n966gat) ) ;
NOR2    gate2448  (.A(n856gat), .B(n2840gat), .Z(n790gat) ) ;
NOR2    gate2449  (.A(n373gat), .B(n2781gat), .Z(n444gat) ) ;
NOR2    gate2450  (.A(n856gat), .B(n2842gat), .Z(n440gat) ) ;
NOR3    gate2451  (.A(n1055gat), .B(n1056gat), .C(n1057gat), .Z(n1051gat) ) ;
NOR3    gate2452  (.A(n1055gat), .B(n1058gat), .C(n1059gat), .Z(n1052gat) ) ;
NOR3    gate2453  (.A(n1060gat), .B(n1056gat), .C(n1059gat), .Z(n1053gat) ) ;
NOR3    gate2454  (.A(n1060gat), .B(n1058gat), .C(n1057gat), .Z(n1054gat) ) ;
NOR3    gate2455  (.A(n938gat), .B(n939gat), .C(n940gat), .Z(n934gat) ) ;
NOR3    gate2456  (.A(n938gat), .B(n941gat), .C(n942gat), .Z(n935gat) ) ;
NOR3    gate2457  (.A(n943gat), .B(n939gat), .C(n942gat), .Z(n936gat) ) ;
NOR3    gate2458  (.A(n943gat), .B(n941gat), .C(n940gat), .Z(n937gat) ) ;
NOR3    gate2459  (.A(n714gat), .B(n715gat), .C(n716gat), .Z(n710gat) ) ;
NOR3    gate2460  (.A(n714gat), .B(n717gat), .C(n718gat), .Z(n711gat) ) ;
NOR3    gate2461  (.A(n719gat), .B(n715gat), .C(n718gat), .Z(n712gat) ) ;
NOR3    gate2462  (.A(n719gat), .B(n717gat), .C(n716gat), .Z(n713gat) ) ;
NOR3    gate2463  (.A(n733gat), .B(n734gat), .C(n735gat), .Z(n729gat) ) ;
NOR3    gate2464  (.A(n733gat), .B(n736gat), .C(n737gat), .Z(n730gat) ) ;
NOR3    gate2465  (.A(n738gat), .B(n734gat), .C(n737gat), .Z(n731gat) ) ;
NOR3    gate2466  (.A(n738gat), .B(n736gat), .C(n735gat), .Z(n732gat) ) ;
NOR3    gate2467  (.A(n498gat), .B(n499gat), .C(n500gat), .Z(n494gat) ) ;
NOR3    gate2468  (.A(n498gat), .B(n501gat), .C(n502gat), .Z(n495gat) ) ;
NOR3    gate2469  (.A(n503gat), .B(n499gat), .C(n502gat), .Z(n496gat) ) ;
NOR3    gate2470  (.A(n503gat), .B(n501gat), .C(n500gat), .Z(n497gat) ) ;
NOR3    gate2471  (.A(n509gat), .B(n510gat), .C(n511gat), .Z(n505gat) ) ;
NOR3    gate2472  (.A(n509gat), .B(n512gat), .C(n513gat), .Z(n506gat) ) ;
NOR3    gate2473  (.A(n514gat), .B(n510gat), .C(n513gat), .Z(n507gat) ) ;
NOR3    gate2474  (.A(n514gat), .B(n512gat), .C(n511gat), .Z(n508gat) ) ;
OR3     gate2475  (.A(n2860gat), .B(n2855gat), .C(n2863gat), .Z(II1277) ) ;
NOR2    gate2476  (.A(n219gat), .B(n2731gat), .Z(n767gat) ) ;
NOR2    gate2477  (.A(n2718gat), .B(n111gat), .Z(n653gat) ) ;
NOR2    gate2478  (.A(n219gat), .B(n2775gat), .Z(n867gat) ) ;
NOR2    gate2479  (.A(n2838gat), .B(n111gat), .Z(n771gat) ) ;
NOR2    gate2480  (.A(n111gat), .B(n2711gat), .Z(n964gat) ) ;
NOR2    gate2481  (.A(n219gat), .B(n2734gat), .Z(n961gat) ) ;
NOR3    gate2482  (.A(n808gat), .B(n809gat), .C(n810gat), .Z(n804gat) ) ;
NOR3    gate2483  (.A(n808gat), .B(n811gat), .C(n812gat), .Z(n805gat) ) ;
NOR3    gate2484  (.A(n813gat), .B(n809gat), .C(n812gat), .Z(n806gat) ) ;
NOR3    gate2485  (.A(n813gat), .B(n811gat), .C(n810gat), .Z(n807gat) ) ;
NOR3    gate2486  (.A(n591gat), .B(n592gat), .C(n593gat), .Z(n587gat) ) ;
NOR3    gate2487  (.A(n591gat), .B(n594gat), .C(n595gat), .Z(n588gat) ) ;
NOR3    gate2488  (.A(n596gat), .B(n592gat), .C(n595gat), .Z(n589gat) ) ;
NOR3    gate2489  (.A(n596gat), .B(n594gat), .C(n593gat), .Z(n590gat) ) ;
NOR2    gate2490  (.A(n2836gat), .B(n111gat), .Z(n447gat) ) ;
NOR2    gate2491  (.A(n2778gat), .B(n219gat), .Z(n445gat) ) ;
NOR3    gate2492  (.A(n691gat), .B(n692gat), .C(n693gat), .Z(n687gat) ) ;
NOR3    gate2493  (.A(n691gat), .B(n694gat), .C(n695gat), .Z(n688gat) ) ;
NOR3    gate2494  (.A(n696gat), .B(n692gat), .C(n695gat), .Z(n689gat) ) ;
NOR3    gate2495  (.A(n696gat), .B(n694gat), .C(n693gat), .Z(n690gat) ) ;
NOR3    gate2496  (.A(n572gat), .B(n573gat), .C(n574gat), .Z(n568gat) ) ;
NOR3    gate2497  (.A(n572gat), .B(n575gat), .C(n576gat), .Z(n569gat) ) ;
NOR3    gate2498  (.A(n577gat), .B(n573gat), .C(n576gat), .Z(n570gat) ) ;
NOR3    gate2499  (.A(n577gat), .B(n575gat), .C(n574gat), .Z(n571gat) ) ;
OR3     gate2500  (.A(n2474gat), .B(n2524gat), .C(n2831gat), .Z(II1515) ) ;
OR3     gate2501  (.A(n2353gat), .B(n2284gat), .C(n2354gat), .Z(II1584) ) ;
NOR2    gate2502  (.A(n1879gat), .B(n1762gat), .Z(n1692gat) ) ;
OR3     gate2503  (.A(n2354gat), .B(n2353gat), .C(n2214gat), .Z(II1723) ) ;
NOR2    gate2504  (.A(n2433gat), .B(n2427gat), .Z(n2428gat) ) ;
OR3     gate2505  (.A(n2286gat), .B(n2428gat), .C(n2289gat), .Z(II1733) ) ;
NOR2    gate2506  (.A(n93gat), .B(n2731gat), .Z(n769gat) ) ;
NOR2    gate2507  (.A(n93gat), .B(n2775gat), .Z(n1076gat) ) ;
NOR2    gate2508  (.A(n93gat), .B(n2734gat), .Z(n766gat) ) ;
NOR3    gate2509  (.A(n1189gat), .B(n1190gat), .C(n1191gat), .Z(n1185gat) ) ;
NOR3    gate2510  (.A(n1189gat), .B(n1192gat), .C(n1193gat), .Z(n1186gat) ) ;
NOR3    gate2511  (.A(n1194gat), .B(n1190gat), .C(n1193gat), .Z(n1187gat) ) ;
NOR3    gate2512  (.A(n1194gat), .B(n1192gat), .C(n1191gat), .Z(n1188gat) ) ;
NOR2    gate2513  (.A(n2792gat), .B(n93gat), .Z(n645gat) ) ;
NOR2    gate2514  (.A(n93gat), .B(n2669gat), .Z(n646gat) ) ;
NOR2    gate2515  (.A(n1280gat), .B(n1225gat), .Z(n1383gat) ) ;
NOR2    gate2516  (.A(n1281gat), .B(n1224gat), .Z(n1327gat) ) ;
NOR2    gate2517  (.A(n93gat), .B(n2778gat), .Z(n651gat) ) ;
NOR2    gate2518  (.A(n2789gat), .B(n93gat), .Z(n652gat) ) ;
NOR2    gate2519  (.A(n2781gat), .B(n93gat), .Z(n765gat) ) ;
NOR3    gate2520  (.A(n1206gat), .B(n1207gat), .C(n1208gat), .Z(n1202gat) ) ;
NOR3    gate2521  (.A(n1206gat), .B(n1209gat), .C(n1210gat), .Z(n1203gat) ) ;
NOR3    gate2522  (.A(n1211gat), .B(n1207gat), .C(n1210gat), .Z(n1204gat) ) ;
NOR3    gate2523  (.A(n1211gat), .B(n1209gat), .C(n1208gat), .Z(n1205gat) ) ;
NOR3    gate2524  (.A(n1274gat), .B(n1275gat), .C(n1276gat), .Z(n1270gat) ) ;
NOR3    gate2525  (.A(n1274gat), .B(n1277gat), .C(n1278gat), .Z(n1271gat) ) ;
NOR3    gate2526  (.A(n1279gat), .B(n1275gat), .C(n1278gat), .Z(n1272gat) ) ;
NOR3    gate2527  (.A(n1279gat), .B(n1277gat), .C(n1276gat), .Z(n1273gat) ) ;
NOR2    gate2528  (.A(n2672gat), .B(n93gat), .Z(n763gat) ) ;
NOR2    gate2529  (.A(n1284gat), .B(n1195gat), .Z(n1287gat) ) ;
NOR2    gate2530  (.A(n1196gat), .B(n1269gat), .Z(n1285gat) ) ;
NOR2    gate2531  (.A(n2852gat), .B(n851gat), .Z(n793gat) ) ;
NOR2    gate2532  (.A(n2672gat), .B(n852gat), .Z(n556gat) ) ;
NOR2    gate2533  (.A(n2731gat), .B(n852gat), .Z(n795gat) ) ;
NOR2    gate2534  (.A(n851gat), .B(n2718gat), .Z(n656gat) ) ;
NOR2    gate2535  (.A(n852gat), .B(n2775gat), .Z(n794gat) ) ;
NOR2    gate2536  (.A(n851gat), .B(n2838gat), .Z(n773gat) ) ;
NOR2    gate2537  (.A(n2711gat), .B(n851gat), .Z(n965gat) ) ;
NOR2    gate2538  (.A(n2734gat), .B(n852gat), .Z(n960gat) ) ;
NOR3    gate2539  (.A(n784gat), .B(n785gat), .C(n786gat), .Z(n780gat) ) ;
NOR3    gate2540  (.A(n784gat), .B(n787gat), .C(n788gat), .Z(n781gat) ) ;
NOR3    gate2541  (.A(n789gat), .B(n785gat), .C(n788gat), .Z(n782gat) ) ;
NOR3    gate2542  (.A(n789gat), .B(n787gat), .C(n786gat), .Z(n783gat) ) ;
NOR2    gate2543  (.A(n852gat), .B(n2792gat), .Z(n555gat) ) ;
NOR2    gate2544  (.A(n851gat), .B(n2846gat), .Z(n450gat) ) ;
NOR2    gate2545  (.A(n851gat), .B(n2844gat), .Z(n654gat) ) ;
NOR2    gate2546  (.A(n2669gat), .B(n852gat), .Z(n557gat) ) ;
NOR2    gate2547  (.A(n559gat), .B(n365gat), .Z(n874gat) ) ;
NOR2    gate2548  (.A(n560gat), .B(n364gat), .Z(n132gat) ) ;
NOR2    gate2549  (.A(n2778gat), .B(n852gat), .Z(n649gat) ) ;
NOR2    gate2550  (.A(n2836gat), .B(n851gat), .Z(n449gat) ) ;
NOR2    gate2551  (.A(n851gat), .B(n2840gat), .Z(n791gat) ) ;
NOR2    gate2552  (.A(n852gat), .B(n2789gat), .Z(n650gat) ) ;
NOR2    gate2553  (.A(n2842gat), .B(n851gat), .Z(n774gat) ) ;
NOR2    gate2554  (.A(n852gat), .B(n2781gat), .Z(n764gat) ) ;
NOR3    gate2555  (.A(n226gat), .B(n227gat), .C(n228gat), .Z(n222gat) ) ;
NOR3    gate2556  (.A(n226gat), .B(n229gat), .C(n230gat), .Z(n223gat) ) ;
NOR3    gate2557  (.A(n231gat), .B(n227gat), .C(n230gat), .Z(n224gat) ) ;
NOR3    gate2558  (.A(n231gat), .B(n229gat), .C(n228gat), .Z(n225gat) ) ;
NOR3    gate2559  (.A(n125gat), .B(n126gat), .C(n127gat), .Z(n121gat) ) ;
NOR3    gate2560  (.A(n125gat), .B(n128gat), .C(n129gat), .Z(n122gat) ) ;
NOR3    gate2561  (.A(n130gat), .B(n126gat), .C(n129gat), .Z(n123gat) ) ;
NOR3    gate2562  (.A(n130gat), .B(n128gat), .C(n127gat), .Z(n124gat) ) ;
NOR2    gate2563  (.A(n666gat), .B(n120gat), .Z(n2460gat) ) ;
NOR2    gate2564  (.A(n665gat), .B(n1601gat), .Z(n2423gat) ) ;
NOR3    gate2565  (.A(n2573gat), .B(n2574gat), .C(n2575gat), .Z(n2569gat) ) ;
NOR3    gate2566  (.A(n2573gat), .B(n2576gat), .C(n2577gat), .Z(n2570gat) ) ;
NOR3    gate2567  (.A(n2578gat), .B(n2574gat), .C(n2577gat), .Z(n2571gat) ) ;
NOR3    gate2568  (.A(n2578gat), .B(n2576gat), .C(n2575gat), .Z(n2572gat) ) ;
NOR3    gate2569  (.A(n2414gat), .B(n2415gat), .C(n2416gat), .Z(n2410gat) ) ;
NOR3    gate2570  (.A(n2414gat), .B(n2417gat), .C(n2418gat), .Z(n2411gat) ) ;
NOR3    gate2571  (.A(n2419gat), .B(n2415gat), .C(n2418gat), .Z(n2412gat) ) ;
NOR3    gate2572  (.A(n2419gat), .B(n2417gat), .C(n2416gat), .Z(n2413gat) ) ;
NOR2    gate2573  (.A(n2582gat), .B(n2583gat), .Z(n2580gat) ) ;
NOR2    gate2574  (.A(n2583gat), .B(n2585gat), .Z(n2581gat) ) ;
NOR2    gate2575  (.A(n2493gat), .B(n2388gat), .Z(n2567gat) ) ;
NOR2    gate2576  (.A(n2389gat), .B(n2494gat), .Z(n2499gat) ) ;
NOR2    gate2577  (.A(n2268gat), .B(n2338gat), .Z(n299gat) ) ;
NOR2    gate2578  (.A(n2337gat), .B(n2269gat), .Z(n207gat) ) ;
NOR2    gate2579  (.A(n2649gat), .B(n2650gat), .Z(n2647gat) ) ;
NOR2    gate2580  (.A(n2650gat), .B(n2652gat), .Z(n2648gat) ) ;
NOR3    gate2581  (.A(n2606gat), .B(n2607gat), .C(n2608gat), .Z(n2602gat) ) ;
NOR3    gate2582  (.A(n2606gat), .B(n2609gat), .C(n2610gat), .Z(n2603gat) ) ;
NOR3    gate2583  (.A(n2611gat), .B(n2607gat), .C(n2610gat), .Z(n2604gat) ) ;
NOR3    gate2584  (.A(n2611gat), .B(n2609gat), .C(n2608gat), .Z(n2605gat) ) ;
NOR3    gate2585  (.A(n2550gat), .B(n2551gat), .C(n2552gat), .Z(n2546gat) ) ;
NOR3    gate2586  (.A(n2550gat), .B(n2553gat), .C(n2554gat), .Z(n2547gat) ) ;
NOR3    gate2587  (.A(n2555gat), .B(n2551gat), .C(n2554gat), .Z(n2548gat) ) ;
NOR3    gate2588  (.A(n2555gat), .B(n2553gat), .C(n2552gat), .Z(n2549gat) ) ;
NOR2    gate2589  (.A(n2616gat), .B(n2617gat), .Z(n2614gat) ) ;
NOR2    gate2590  (.A(n2617gat), .B(n2619gat), .Z(n2615gat) ) ;
NOR2    gate2591  (.A(n120gat), .B(n2666gat), .Z(n2461gat) ) ;
NOR2    gate2592  (.A(n1601gat), .B(n1704gat), .Z(n2421gat) ) ;
NOR2    gate2593  (.A(n1414gat), .B(n566gat), .Z(n1153gat) ) ;
NOR2    gate2594  (.A(n1301gat), .B(n1150gat), .Z(n1151gat) ) ;
NOR2    gate2595  (.A(n873gat), .B(n1478gat), .Z(n982gat) ) ;
NOR2    gate2596  (.A(n875gat), .B(n876gat), .Z(n877gat) ) ;
OR4     gate2597  (.A(n1153gat), .B(n1151gat), .C(n982gat), .D(n877gat), .Z(n2930gat) ) ;
NOR2    gate2598  (.A(n1160gat), .B(n1084gat), .Z(n1159gat) ) ;
NOR2    gate2599  (.A(n983gat), .B(n1157gat), .Z(n1158gat) ) ;
NOR2    gate2600  (.A(n985gat), .B(n1307gat), .Z(n1156gat) ) ;
NOR2    gate2601  (.A(n1085gat), .B(n1348gat), .Z(n1155gat) ) ;
OR4     gate2602  (.A(n1159gat), .B(n1158gat), .C(n1156gat), .D(n1155gat), .Z(n2957gat) ) ;
NOR2    gate2603  (.A(n1442gat), .B(n706gat), .Z(n1443gat) ) ;
NOR2    gate2604  (.A(n1444gat), .B(n164gat), .Z(n1325gat) ) ;
NOR2    gate2605  (.A(n1442gat), .B(n837gat), .Z(n1321gat) ) ;
NOR2    gate2606  (.A(n1444gat), .B(n278gat), .Z(n1320gat) ) ;
NOR2    gate2607  (.A(n1442gat), .B(n613gat), .Z(n1368gat) ) ;
NOR2    gate2608  (.A(n274gat), .B(n1444gat), .Z(n1258gat) ) ;
NOR2    gate2609  (.A(n833gat), .B(n1442gat), .Z(n1373gat) ) ;
NOR2    gate2610  (.A(n282gat), .B(n1444gat), .Z(n1372gat) ) ;
NOR2    gate2611  (.A(n1437gat), .B(n1378gat), .Z(n1441gat) ) ;
NOR2    gate2612  (.A(n1322gat), .B(n1439gat), .Z(n1440gat) ) ;
NOR2    gate2613  (.A(n1370gat), .B(n1369gat), .Z(n1371gat) ) ;
NOR2    gate2614  (.A(n1366gat), .B(n1374gat), .Z(n1367gat) ) ;
OR4     gate2615  (.A(n1441gat), .B(n1440gat), .C(n1371gat), .D(n1367gat), .Z(n2978gat) ) ;
NOR2    gate2616  (.A(n1450gat), .B(n1498gat), .Z(n1504gat) ) ;
NOR2    gate2617  (.A(n1607gat), .B(n1449gat), .Z(n1502gat) ) ;
OR2     gate2618  (.A(n1504gat), .B(n1502gat), .Z(n2982gat) ) ;
NOR2    gate2619  (.A(n1603gat), .B(n815gat), .Z(n1250gat) ) ;
NOR2    gate2620  (.A(n956gat), .B(n1590gat), .Z(n1103gat) ) ;
NOR2    gate2621  (.A(n1590gat), .B(n1067gat), .Z(n1304gat) ) ;
NOR2    gate2622  (.A(n679gat), .B(n1603gat), .Z(n1249gat) ) ;
NOR2    gate2623  (.A(n864gat), .B(n1590gat), .Z(n1246gat) ) ;
NOR2    gate2624  (.A(n583gat), .B(n1603gat), .Z(n1161gat) ) ;
NOR2    gate2625  (.A(n1603gat), .B(n579gat), .Z(n1291gat) ) ;
NOR2    gate2626  (.A(n1590gat), .B(n860gat), .Z(n1245gat) ) ;
NOR2    gate2627  (.A(n1248gat), .B(n1418gat), .Z(n1352gat) ) ;
NOR2    gate2628  (.A(n1306gat), .B(n1353gat), .Z(n1351gat) ) ;
NOR2    gate2629  (.A(n1247gat), .B(n1355gat), .Z(n1303gat) ) ;
NOR2    gate2630  (.A(n1300gat), .B(n1487gat), .Z(n1302gat) ) ;
OR4     gate2631  (.A(n1352gat), .B(n1351gat), .C(n1303gat), .D(n1302gat), .Z(n2973gat) ) ;
NOR2    gate2632  (.A(n882gat), .B(n1603gat), .Z(n1163gat) ) ;
NOR2    gate2633  (.A(n1297gat), .B(n1590gat), .Z(n1102gat) ) ;
NOR2    gate2634  (.A(n1590gat), .B(n1293gat), .Z(n1101gat) ) ;
NOR2    gate2635  (.A(n1603gat), .B(n823gat), .Z(n996gat) ) ;
NOR2    gate2636  (.A(n1079gat), .B(n1590gat), .Z(n1104gat) ) ;
NOR2    gate2637  (.A(n1603gat), .B(n683gat), .Z(n887gat) ) ;
NOR2    gate2638  (.A(n1147gat), .B(n1590gat), .Z(n1305gat) ) ;
NOR2    gate2639  (.A(n698gat), .B(n1603gat), .Z(n1162gat) ) ;
NOR2    gate2640  (.A(n1164gat), .B(n1356gat), .Z(n1360gat) ) ;
NOR2    gate2641  (.A(n1436gat), .B(n1106gat), .Z(n1359gat) ) ;
NOR2    gate2642  (.A(n1425gat), .B(n1105gat), .Z(n1358gat) ) ;
NOR2    gate2643  (.A(n1424gat), .B(n1309gat), .Z(n1357gat) ) ;
OR4     gate2644  (.A(n1360gat), .B(n1359gat), .C(n1358gat), .D(n1357gat), .Z(n2977gat) ) ;
OR3     gate2645  (.A(n1788gat), .B(n1786gat), .C(n1839gat), .Z(II2720) ) ;
OR3     gate2646  (.A(n1788gat), .B(n1884gat), .C(n1633gat), .Z(II2735) ) ;
NOR2    gate2647  (.A(n1705gat), .B(n3028gat), .Z(n1703gat) ) ;
NOR2    gate2648  (.A(n3026gat), .B(n1779gat), .Z(n1778gat) ) ;
OR3     gate2649  (.A(n1703gat), .B(n1704gat), .C(n1778gat), .Z(II2812) ) ;
NOR2    gate2650  (.A(n1503gat), .B(n3025gat), .Z(n1609gat) ) ;
OR3     gate2651  (.A(n1839gat), .B(n1786gat), .C(n1788gat), .Z(II2831) ) ;
OR3     gate2652  (.A(n1784gat), .B(n1633gat), .C(n1884gat), .Z(II2889) ) ;
OR3     gate2653  (.A(n1784gat), .B(n1785gat), .C(n1633gat), .Z(II2925) ) ;
OR3     gate2654  (.A(n1784gat), .B(n1839gat), .C(n1788gat), .Z(II2934) ) ;
NOR2    gate2655  (.A(n1673gat), .B(n1572gat), .Z(n1733gat) ) ;
NOR2    gate2656  (.A(n1858gat), .B(n1580gat), .Z(n1581gat) ) ;
NOR4    gate2657  (.A(n2078gat), .B(n2178gat), .C(n1990gat), .D(n2128gat), .Z(n2079gat) ) ;
NOR3    gate2658  (.A(n2078gat), .B(n1990gat), .C(n2181gat), .Z(n2073gat) ) ;
NOR3    gate2659  (.A(n1719gat), .B(n1673gat), .C(n1444gat), .Z(n1574gat) ) ;
NOR3    gate2660  (.A(n1444gat), .B(n1858gat), .C(n1635gat), .Z(n1573gat) ) ;
NOR3    gate2661  (.A(n1659gat), .B(n1722gat), .C(n1724gat), .Z(n1723gat) ) ;
NOR3    gate2662  (.A(n1656gat), .B(n1659gat), .C(n1554gat), .Z(n1647gat) ) ;
NOR3    gate2663  (.A(n1569gat), .B(n1659gat), .C(n1566gat), .Z(n1646gat) ) ;
OR3     gate2664  (.A(n1723gat), .B(n1647gat), .C(n1646gat), .Z(n2992gat) ) ;
NOR3    gate2665  (.A(n1727gat), .B(n1659gat), .C(n1640gat), .Z(n1650gat) ) ;
NOR3    gate2666  (.A(n1560gat), .B(n1659gat), .C(n1730gat), .Z(n1649gat) ) ;
NOR3    gate2667  (.A(n1561gat), .B(n1562gat), .C(n1659gat), .Z(n1563gat) ) ;
OR3     gate2668  (.A(n1650gat), .B(n1649gat), .C(n1563gat), .Z(n2986gat) ) ;
NOR2    gate2669  (.A(n1671gat), .B(n1659gat), .Z(n1654gat) ) ;
NOR3    gate2670  (.A(n1651gat), .B(n1652gat), .C(n1659gat), .Z(n1653gat) ) ;
NOR3    gate2671  (.A(n1643gat), .B(n1648gat), .C(n1659gat), .Z(n1644gat) ) ;
OR3     gate2672  (.A(n1654gat), .B(n1653gat), .C(n1644gat), .Z(n2991gat) ) ;
OR3     gate2673  (.A(n1839gat), .B(n1884gat), .C(n1784gat), .Z(II3148) ) ;
OR3     gate2674  (.A(n1838gat), .B(n1785gat), .C(n1788gat), .Z(II3178) ) ;
NOR3    gate2675  (.A(n1869gat), .B(n672gat), .C(n2591gat), .Z(n1413gat) ) ;
NOR3    gate2676  (.A(n1507gat), .B(n1396gat), .C(n1393gat), .Z(n1408gat) ) ;
NOR3    gate2677  (.A(n1393gat), .B(n1409gat), .C(n1677gat), .Z(n1407gat) ) ;
OR3     gate2678  (.A(n1413gat), .B(n1408gat), .C(n1407gat), .Z(n2981gat) ) ;
NOR2    gate2679  (.A(n2260gat), .B(n2189gat), .Z(n2258gat) ) ;
NOR2    gate2680  (.A(n2261gat), .B(n2188gat), .Z(n2255gat) ) ;
NOR2    gate2681  (.A(n2133gat), .B(n2131gat), .Z(n2132gat) ) ;
NOR2    gate2682  (.A(n2134gat), .B(n2185gat), .Z(n2130gat) ) ;
NOR2    gate2683  (.A(n2248gat), .B(n2264gat), .Z(n2250gat) ) ;
NOR2    gate2684  (.A(n2265gat), .B(n3006gat), .Z(n2249gat) ) ;
OR2     gate2685  (.A(n2250gat), .B(n2249gat), .Z(n3007gat) ) ;
NOR2    gate2686  (.A(n1709gat), .B(n1629gat), .Z(n1710gat) ) ;
NOR2    gate2687  (.A(n1895gat), .B(n1631gat), .Z(n1630gat) ) ;
NOR3    gate2688  (.A(n1968gat), .B(n1891gat), .C(n1969gat), .Z(n1894gat) ) ;
NOR2    gate2689  (.A(n1958gat), .B(n1845gat), .Z(n1847gat) ) ;
NOR2    gate2690  (.A(n1845gat), .B(n1893gat), .Z(n1846gat) ) ;
NOR2    gate2691  (.A(n1891gat), .B(n1958gat), .Z(n2055gat) ) ;
NOR2    gate2692  (.A(n1893gat), .B(n1968gat), .Z(n1967gat) ) ;
NOR2    gate2693  (.A(n1956gat), .B(n1963gat), .Z(n1959gat) ) ;
NOR2    gate2694  (.A(n1886gat), .B(n1887gat), .Z(n1957gat) ) ;
NOR2    gate2695  (.A(n2193gat), .B(n2402gat), .Z(n2211gat) ) ;
NOR2    gate2696  (.A(n2401gat), .B(n2151gat), .Z(n2210gat) ) ;
NOR2    gate2697  (.A(n2393gat), .B(n2438gat), .Z(n2053gat) ) ;
NOR2    gate2698  (.A(n2392gat), .B(n2439gat), .Z(n1964gat) ) ;
NOR2    gate2699  (.A(n2405gat), .B(n2349gat), .Z(n2350gat) ) ;
NOR2    gate2700  (.A(n2406gat), .B(n2215gat), .Z(n2282gat) ) ;
NOR3    gate2701  (.A(n2402gat), .B(n2151gat), .C(n2345gat), .Z(n2213gat) ) ;
NOR2    gate2702  (.A(n2401gat), .B(n2346gat), .Z(n2150gat) ) ;
NOR2    gate2703  (.A(n2193gat), .B(n2346gat), .Z(n2149gat) ) ;
NOR2    gate2704  (.A(n1963gat), .B(n1893gat), .Z(n1962gat) ) ;
OR2     gate2705  (.A(n1962gat), .B(n1955gat), .Z(n2995gat) ) ;
NOR2    gate2706  (.A(n1974gat), .B(n1970gat), .Z(n1972gat) ) ;
NOR2    gate2707  (.A(n1896gat), .B(n1973gat), .Z(n1971gat) ) ;
OR2     gate2708  (.A(n1972gat), .B(n1971gat), .Z(n2999gat) ) ;
NOR2    gate2709  (.A(n2393gat), .B(n2401gat), .Z(n2331gat) ) ;
OR2     gate2710  (.A(n2333gat), .B(n2331gat), .Z(n3011gat) ) ;
NOR2    gate2711  (.A(n2643gat), .B(n2564gat), .Z(n2566gat) ) ;
NOR2    gate2712  (.A(n2352gat), .B(n2642gat), .Z(n2565gat) ) ;
OR2     gate2713  (.A(n2566gat), .B(n2565gat), .Z(n3015gat) ) ;
NOR3    gate2714  (.A(n155gat), .B(n253gat), .C(n150gat), .Z(n141gat) ) ;
NOR2    gate2715  (.A(n151gat), .B(n233gat), .Z(n38gat) ) ;
NOR2    gate2716  (.A(n151gat), .B(n154gat), .Z(n37gat) ) ;
NOR2    gate2717  (.A(n2775gat), .B(n110gat), .Z(n1074gat) ) ;
NOR2    gate2718  (.A(n375gat), .B(n800gat), .Z(n872gat) ) ;
NOR2    gate2719  (.A(n155gat), .B(n233gat), .Z(n234gat) ) ;
NOR2    gate2720  (.A(n154gat), .B(n253gat), .Z(n137gat) ) ;
NOR2    gate2721  (.A(n375gat), .B(n235gat), .Z(n378gat) ) ;
NOR2    gate2722  (.A(n110gat), .B(n2778gat), .Z(n377gat) ) ;
NOR3    gate2723  (.A(n329gat), .B(n387gat), .C(n334gat), .Z(n250gat) ) ;
NOR2    gate2724  (.A(n386gat), .B(n330gat), .Z(n249gat) ) ;
NOR2    gate2725  (.A(n330gat), .B(n1490gat), .Z(n248gat) ) ;
NOR2    gate2726  (.A(n219gat), .B(n2792gat), .Z(n869gat) ) ;
NOR2    gate2727  (.A(n372gat), .B(n452gat), .Z(n453gat) ) ;
NOR2    gate2728  (.A(n111gat), .B(n2846gat), .Z(n448gat) ) ;
NOR2    gate2729  (.A(n1490gat), .B(n387gat), .Z(n251gat) ) ;
NOR2    gate2730  (.A(n334gat), .B(n386gat), .Z(n244gat) ) ;
NOR2    gate2731  (.A(n2844gat), .B(n111gat), .Z(n974gat) ) ;
NOR2    gate2732  (.A(n372gat), .B(n333gat), .Z(n973gat) ) ;
NOR2    gate2733  (.A(n2669gat), .B(n219gat), .Z(n870gat) ) ;
NOR3    gate2734  (.A(n330gat), .B(n325gat), .C(n334gat), .Z(n246gat) ) ;
NOR2    gate2735  (.A(n386gat), .B(n334gat), .Z(n245gat) ) ;
NOR2    gate2736  (.A(n462gat), .B(n2884gat), .Z(n460gat) ) ;
NOR2    gate2737  (.A(n457gat), .B(n461gat), .Z(n459gat) ) ;
NOR2    gate2738  (.A(n111gat), .B(n2852gat), .Z(n975gat) ) ;
NOR2    gate2739  (.A(n372gat), .B(n458gat), .Z(n972gat) ) ;
NOR2    gate2740  (.A(n219gat), .B(n2672gat), .Z(n969gat) ) ;
NOR2    gate2741  (.A(n144gat), .B(n325gat), .Z(n145gat) ) ;
NOR2    gate2742  (.A(n326gat), .B(n247gat), .Z(n143gat) ) ;
NOR2    gate2743  (.A(n111gat), .B(n2840gat), .Z(n971gat) ) ;
NOR2    gate2744  (.A(n372gat), .B(n878gat), .Z(n970gat) ) ;
NOR2    gate2745  (.A(n2789gat), .B(n219gat), .Z(n968gat) ) ;
NOR3    gate2746  (.A(n382gat), .B(n326gat), .C(n144gat), .Z(n142gat) ) ;
NOR2    gate2747  (.A(n325gat), .B(n383gat), .Z(n40gat) ) ;
NOR2    gate2748  (.A(n383gat), .B(n247gat), .Z(n39gat) ) ;
NOR2    gate2749  (.A(n111gat), .B(n2842gat), .Z(n772gat) ) ;
NOR2    gate2750  (.A(n134gat), .B(n372gat), .Z(n451gat) ) ;
NOR2    gate2751  (.A(n219gat), .B(n2781gat), .Z(n446gat) ) ;
NOR3    gate2752  (.A(n253gat), .B(n151gat), .C(n254gat), .Z(n139gat) ) ;
NOR2    gate2753  (.A(n253gat), .B(n154gat), .Z(n136gat) ) ;
NOR2    gate2754  (.A(n252gat), .B(n468gat), .Z(n391gat) ) ;
NOR2    gate2755  (.A(n469gat), .B(n2877gat), .Z(n390gat) ) ;
NOR2    gate2756  (.A(n381gat), .B(n375gat), .Z(n1083gat) ) ;
NOR2    gate2757  (.A(n110gat), .B(n2672gat), .Z(n1077gat) ) ;
NOR2    gate2758  (.A(n254gat), .B(n241gat), .Z(n242gat) ) ;
NOR2    gate2759  (.A(n255gat), .B(n140gat), .Z(n240gat) ) ;
NOR2    gate2760  (.A(n802gat), .B(n375gat), .Z(n871gat) ) ;
NOR2    gate2761  (.A(n110gat), .B(n2734gat), .Z(n797gat) ) ;
NOR3    gate2762  (.A(n255gat), .B(n146gat), .C(n241gat), .Z(n324gat) ) ;
NOR2    gate2763  (.A(n147gat), .B(n254gat), .Z(n238gat) ) ;
NOR2    gate2764  (.A(n140gat), .B(n147gat), .Z(n237gat) ) ;
NOR2    gate2765  (.A(n375gat), .B(n380gat), .Z(n1082gat) ) ;
NOR2    gate2766  (.A(n2731gat), .B(n110gat), .Z(n796gat) ) ;
NOR2    gate2767  (.A(n1691gat), .B(n336gat), .Z(n1599gat) ) ;
OR3     gate2768  (.A(n2167gat), .B(n2031gat), .C(n2174gat), .Z(II3999) ) ;
NOR2    gate2769  (.A(n1869gat), .B(n1683gat), .Z(n1586gat) ) ;
NOR3    gate2770  (.A(n1769gat), .B(n1773gat), .C(n2512gat), .Z(n1755gat) ) ;
OR3     gate2771  (.A(n2443gat), .B(n2290gat), .C(n2214gat), .Z(II4023) ) ;
NOR2    gate2772  (.A(n1472gat), .B(n1747gat), .Z(n1470gat) ) ;
NOR2    gate2773  (.A(n1674gat), .B(n1403gat), .Z(n1400gat) ) ;
NOR3    gate2774  (.A(n1806gat), .B(n1338gat), .C(n1584gat), .Z(n1399gat) ) ;
NOR2    gate2775  (.A(n1455gat), .B(n1397gat), .Z(n1398gat) ) ;
OR3     gate2776  (.A(n1633gat), .B(n1838gat), .C(n1786gat), .Z(II4144) ) ;
NOR2    gate2777  (.A(n2289gat), .B(n1468gat), .Z(n1467gat) ) ;
NOR3    gate2778  (.A(n1392gat), .B(n1461gat), .C(n1396gat), .Z(n1466gat) ) ;
NOR3    gate2779  (.A(n1774gat), .B(n1869gat), .C(n1684gat), .Z(n1686gat) ) ;
NOR2    gate2780  (.A(n1524gat), .B(n1403gat), .Z(n1533gat) ) ;
NOR2    gate2781  (.A(n1677gat), .B(n1458gat), .Z(n1532gat) ) ;
NOR2    gate2782  (.A(n1507gat), .B(n1477gat), .Z(n1531gat) ) ;
OR4     gate2783  (.A(n1686gat), .B(n1533gat), .C(n1532gat), .D(n1531gat), .Z(n2985gat) ) ;
OR3     gate2784  (.A(n1427gat), .B(n1595gat), .C(n1677gat), .Z(II4216) ) ;
NOR2    gate2785  (.A(n1297gat), .B(n1111gat), .Z(n1100gat) ) ;
NOR2    gate2786  (.A(n1112gat), .B(n882gat), .Z(n994gat) ) ;
NOR2    gate2787  (.A(n721gat), .B(n741gat), .Z(n989gat) ) ;
NOR2    gate2788  (.A(n926gat), .B(n566gat), .Z(n880gat) ) ;
OR4     gate2789  (.A(n1100gat), .B(n994gat), .C(n989gat), .D(n880gat), .Z(n2931gat) ) ;
NOR2    gate2790  (.A(n1007gat), .B(n918gat), .Z(n1012gat) ) ;
NOR2    gate2791  (.A(n625gat), .B(n1006gat), .Z(n905gat) ) ;
OR2     gate2792  (.A(n1012gat), .B(n905gat), .Z(n2943gat) ) ;
NOR2    gate2793  (.A(n420gat), .B(n879gat), .Z(n1003gat) ) ;
NOR2    gate2794  (.A(n1009gat), .B(n419gat), .Z(n902gat) ) ;
NOR2    gate2795  (.A(n1111gat), .B(n1293gat), .Z(n1099gat) ) ;
NOR2    gate2796  (.A(n725gat), .B(n741gat), .Z(n998gat) ) ;
NOR2    gate2797  (.A(n823gat), .B(n1112gat), .Z(n995gat) ) ;
NOR2    gate2798  (.A(n875gat), .B(n926gat), .Z(n980gat) ) ;
NOR2    gate2799  (.A(n621gat), .B(n1006gat), .Z(n1175gat) ) ;
NOR2    gate2800  (.A(n845gat), .B(n1007gat), .Z(n1174gat) ) ;
OR2     gate2801  (.A(n1175gat), .B(n1174gat), .Z(n2960gat) ) ;
NOR2    gate2802  (.A(n420gat), .B(n1002gat), .Z(n1001gat) ) ;
NOR2    gate2803  (.A(n419gat), .B(n1171gat), .Z(n999gat) ) ;
NOR2    gate2804  (.A(n1007gat), .B(n401gat), .Z(n1323gat) ) ;
NOR2    gate2805  (.A(n1006gat), .B(n617gat), .Z(n1264gat) ) ;
OR2     gate2806  (.A(n1323gat), .B(n1264gat), .Z(n2969gat) ) ;
NOR2    gate2807  (.A(n926gat), .B(n873gat), .Z(n981gat) ) ;
NOR2    gate2808  (.A(n741gat), .B(n702gat), .Z(n890gat) ) ;
NOR2    gate2809  (.A(n1111gat), .B(n1079gat), .Z(n889gat) ) ;
NOR2    gate2810  (.A(n683gat), .B(n1112gat), .Z(n886gat) ) ;
NOR2    gate2811  (.A(n419gat), .B(n1265gat), .Z(n892gat) ) ;
NOR2    gate2812  (.A(n420gat), .B(n888gat), .Z(n891gat) ) ;
NOR2    gate2813  (.A(n1006gat), .B(n490gat), .Z(n904gat) ) ;
NOR2    gate2814  (.A(n1007gat), .B(n397gat), .Z(n903gat) ) ;
OR2     gate2815  (.A(n904gat), .B(n903gat), .Z(n2942gat) ) ;
NOR2    gate2816  (.A(n926gat), .B(n1150gat), .Z(n1152gat) ) ;
NOR2    gate2817  (.A(n1147gat), .B(n1111gat), .Z(n1092gat) ) ;
NOR2    gate2818  (.A(n741gat), .B(n393gat), .Z(n997gat) ) ;
NOR2    gate2819  (.A(n1112gat), .B(n698gat), .Z(n993gat) ) ;
NOR2    gate2820  (.A(n419gat), .B(n1008gat), .Z(n900gat) ) ;
NOR2    gate2821  (.A(n420gat), .B(n898gat), .Z(n895gat) ) ;
NOR2    gate2822  (.A(n1112gat), .B(n583gat), .Z(n1094gat) ) ;
NOR2    gate2823  (.A(n1111gat), .B(n864gat), .Z(n1093gat) ) ;
NOR2    gate2824  (.A(n340gat), .B(n741gat), .Z(n988gat) ) ;
NOR2    gate2825  (.A(n926gat), .B(n983gat), .Z(n984gat) ) ;
NOR2    gate2826  (.A(n613gat), .B(n1006gat), .Z(n1267gat) ) ;
NOR2    gate2827  (.A(n1007gat), .B(n274gat), .Z(n1257gat) ) ;
OR2     gate2828  (.A(n1267gat), .B(n1257gat), .Z(n2965gat) ) ;
NOR2    gate2829  (.A(n420gat), .B(n1179gat), .Z(n1178gat) ) ;
NOR2    gate2830  (.A(n419gat), .B(n1266gat), .Z(n1116gat) ) ;
NOR2    gate2831  (.A(n1006gat), .B(n706gat), .Z(n1375gat) ) ;
NOR2    gate2832  (.A(n164gat), .B(n1007gat), .Z(n1324gat) ) ;
OR2     gate2833  (.A(n1375gat), .B(n1324gat), .Z(n2961gat) ) ;
NOR2    gate2834  (.A(n1111gat), .B(n956gat), .Z(n1091gat) ) ;
NOR2    gate2835  (.A(n1085gat), .B(n926gat), .Z(n1088gat) ) ;
NOR2    gate2836  (.A(n815gat), .B(n1112gat), .Z(n992gat) ) ;
NOR2    gate2837  (.A(n741gat), .B(n159gat), .Z(n987gat) ) ;
NOR2    gate2838  (.A(n419gat), .B(n1172gat), .Z(n899gat) ) ;
NOR2    gate2839  (.A(n897gat), .B(n420gat), .Z(n896gat) ) ;
NOR2    gate2840  (.A(n837gat), .B(n1006gat), .Z(n1262gat) ) ;
NOR2    gate2841  (.A(n1007gat), .B(n278gat), .Z(n1260gat) ) ;
OR2     gate2842  (.A(n1262gat), .B(n1260gat), .Z(n2967gat) ) ;
NOR2    gate2843  (.A(n336gat), .B(n741gat), .Z(n1098gat) ) ;
NOR2    gate2844  (.A(n1111gat), .B(n860gat), .Z(n1090gat) ) ;
NOR2    gate2845  (.A(n985gat), .B(n926gat), .Z(n986gat) ) ;
NOR2    gate2846  (.A(n579gat), .B(n1112gat), .Z(n885gat) ) ;
NOR2    gate2847  (.A(n419gat), .B(n1259gat), .Z(n901gat) ) ;
NOR2    gate2848  (.A(n894gat), .B(n420gat), .Z(n893gat) ) ;
NOR2    gate2849  (.A(n270gat), .B(n741gat), .Z(n1097gat) ) ;
NOR2    gate2850  (.A(n1067gat), .B(n1111gat), .Z(n1089gat) ) ;
NOR2    gate2851  (.A(n926gat), .B(n1084gat), .Z(n1087gat) ) ;
NOR2    gate2852  (.A(n1112gat), .B(n679gat), .Z(n991gat) ) ;
NOR2    gate2853  (.A(n1007gat), .B(n282gat), .Z(n1326gat) ) ;
NOR2    gate2854  (.A(n833gat), .B(n1006gat), .Z(n1261gat) ) ;
OR2     gate2855  (.A(n1326gat), .B(n1261gat), .Z(n2968gat) ) ;
NOR2    gate2856  (.A(n1180gat), .B(n420gat), .Z(n1177gat) ) ;
NOR2    gate2857  (.A(n1263gat), .B(n419gat), .Z(n1115gat) ) ;
NOR2    gate2858  (.A(n670gat), .B(n671gat), .Z(n977gat) ) ;
OR2     gate2859  (.A(n977gat), .B(n976gat), .Z(n2944gat) ) ;
NOR2    gate2860  (.A(n819gat), .B(n1112gat), .Z(n1096gat) ) ;
NOR2    gate2861  (.A(n1240gat), .B(n1111gat), .Z(n1095gat) ) ;
NOR2    gate2862  (.A(n841gat), .B(n741gat), .Z(n990gat) ) ;
NOR2    gate2863  (.A(n1601gat), .B(n926gat), .Z(n979gat) ) ;
OR4     gate2864  (.A(n1096gat), .B(n1095gat), .C(n990gat), .D(n979gat), .Z(n2945gat) ) ;
NOR2    gate2865  (.A(n829gat), .B(n1006gat), .Z(n1176gat) ) ;
NOR2    gate2866  (.A(n1007gat), .B(n1025gat), .Z(n1173gat) ) ;
OR2     gate2867  (.A(n1176gat), .B(n1173gat), .Z(n2962gat) ) ;
NOR2    gate2868  (.A(n978gat), .B(n420gat), .Z(n1004gat) ) ;
NOR2    gate2869  (.A(n419gat), .B(n1252gat), .Z(n1000gat) ) ;
NOR2    gate2870  (.A(n978gat), .B(n455gat), .Z(n1029gat) ) ;
NOR2    gate2871  (.A(n455gat), .B(n879gat), .Z(n1028gat) ) ;
NOR2    gate2872  (.A(n1002gat), .B(n455gat), .Z(n1031gat) ) ;
NOR2    gate2873  (.A(n455gat), .B(n888gat), .Z(n1030gat) ) ;
NOR2    gate2874  (.A(n455gat), .B(n898gat), .Z(n1011gat) ) ;
NOR2    gate2875  (.A(n455gat), .B(n1179gat), .Z(n1181gat) ) ;
NOR2    gate2876  (.A(n897gat), .B(n455gat), .Z(n1010gat) ) ;
NOR2    gate2877  (.A(n894gat), .B(n455gat), .Z(n1005gat) ) ;
NOR2    gate2878  (.A(n1180gat), .B(n455gat), .Z(n1182gat) ) ;
NOR2    gate2879  (.A(n67gat), .B(n2784gat), .Z(n73gat) ) ;
NOR2    gate2880  (.A(n71gat), .B(n2720gat), .Z(n70gat) ) ;
NOR2    gate2881  (.A(n76gat), .B(n2784gat), .Z(n77gat) ) ;
NOR2    gate2882  (.A(n2720gat), .B(n14gat), .Z(n13gat) ) ;
NOR2    gate2883  (.A(n1816gat), .B(n1828gat), .Z(n1935gat) ) ;
NOR2    gate2884  (.A(n194gat), .B(n297gat), .Z(n197gat) ) ;
NOR2    gate2885  (.A(n92gat), .B(n21gat), .Z(n22gat) ) ;
NOR2    gate2886  (.A(n197gat), .B(n22gat), .Z(n93gat) ) ;
NOR2    gate2887  (.A(n2850gat), .B(n3019gat), .Z(n2239gat) ) ;
NOR2    gate2888  (.A(n2432gat), .B(n2154gat), .Z(n2433gat) ) ;
NOR2    gate2889  (.A(n2426gat), .B(n2153gat), .Z(n2427gat) ) ;
NOR2    gate2890  (.A(n2582gat), .B(n2585gat), .Z(n2583gat) ) ;
NOR2    gate2891  (.A(n2649gat), .B(n2652gat), .Z(n2650gat) ) ;
NOR2    gate2892  (.A(n2616gat), .B(n2619gat), .Z(n2617gat) ) ;
NOR2    gate2893  (.A(n1592gat), .B(n2422gat), .Z(n1598gat) ) ;
NOR3    gate2894  (.A(n1598gat), .B(n2930gat), .C(n2957gat), .Z(n1154gat) ) ;
NOR2    gate2895  (.A(n1154gat), .B(n1608gat), .Z(n1411gat) ) ;
NOR2    gate2896  (.A(n1609gat), .B(n1427gat), .Z(n1498gat) ) ;
NOR2    gate2897  (.A(n2082gat), .B(n1609gat), .Z(n1607gat) ) ;
NOR4    gate2898  (.A(n2978gat), .B(n2982gat), .C(n2973gat), .D(n2977gat), .Z(n1428gat) ) ;
NOR2    gate2899  (.A(n1673gat), .B(n1719gat), .Z(n1794gat) ) ;
NOR2    gate2900  (.A(n1858gat), .B(n1635gat), .Z(n1796gat) ) ;
NOR2    gate2901  (.A(n1794gat), .B(n1796gat), .Z(n1792gat) ) ;
NOR2    gate2902  (.A(n1428gat), .B(n1387gat), .Z(n1406gat) ) ;
NOR2    gate2903  (.A(n2850gat), .B(n3018gat), .Z(n2664gat) ) ;
NOR2    gate2904  (.A(n1925gat), .B(n1635gat), .Z(n1926gat) ) ;
NOR2    gate2905  (.A(n1917gat), .B(n1859gat), .Z(n1916gat) ) ;
NOR2    gate2906  (.A(n1719gat), .B(n1922gat), .Z(n1994gat) ) ;
NOR2    gate2907  (.A(n1743gat), .B(n1923gat), .Z(n1924gat) ) ;
NOR2    gate2908  (.A(n1311gat), .B(n1773gat), .Z(n1758gat) ) ;
NOR2    gate2909  (.A(n199gat), .B(n92gat), .Z(n200gat) ) ;
NOR2    gate2910  (.A(n297gat), .B(n195gat), .Z(n196gat) ) ;
NOR2    gate2911  (.A(n2016gat), .B(n2097gat), .Z(n2018gat) ) ;
NOR2    gate2912  (.A(n88gat), .B(n2784gat), .Z(n89gat) ) ;
NOR3    gate2913  (.A(n1334gat), .B(n1858gat), .C(n1604gat), .Z(n1471gat) ) ;
NOR3    gate2914  (.A(n1476gat), .B(n1471gat), .C(n1469gat), .Z(n1472gat) ) ;
NOR2    gate2915  (.A(n1685gat), .B(n1427gat), .Z(n1600gat) ) ;
NOR2    gate2916  (.A(n1519gat), .B(n1401gat), .Z(n1397gat) ) ;
NOR2    gate2917  (.A(n2002gat), .B(n2857gat), .Z(n2005gat) ) ;
NOR2    gate2918  (.A(n1823gat), .B(n2005gat), .Z(n1818gat) ) ;
NOR2    gate2919  (.A(n1584gat), .B(n1460gat), .Z(n1510gat) ) ;
NOR2    gate2920  (.A(n1595gat), .B(n1454gat), .Z(n1459gat) ) ;
NOR2    gate2921  (.A(n1510gat), .B(n1459gat), .Z(n1458gat) ) ;
NOR3    gate2922  (.A(n1594gat), .B(n1587gat), .C(n2989gat), .Z(n1602gat) ) ;
NOR2    gate2923  (.A(n374gat), .B(n2862gat), .Z(n520gat) ) ;
NOR2    gate2924  (.A(n2854gat), .B(n374gat), .Z(n519gat) ) ;
NOR4    gate2925  (.A(n417gat), .B(n413gat), .C(n412gat), .D(n406gat), .Z(n410gat) ) ;
NOR2    gate2926  (.A(n411gat), .B(n522gat), .Z(n354gat) ) ;
NOR2    gate2927  (.A(n516gat), .B(n407gat), .Z(n408gat) ) ;
NOR2    gate2928  (.A(n2859gat), .B(n740gat), .Z(n526gat) ) ;
NOR2    gate2929  (.A(n740gat), .B(n2854gat), .Z(n531gat) ) ;
NOR2    gate2930  (.A(n2862gat), .B(n740gat), .Z(n530gat) ) ;
NOR2    gate2931  (.A(n290gat), .B(n358gat), .Z(n359gat) ) ;
NOR2    gate2932  (.A(n408gat), .B(n359gat), .Z(n420gat) ) ;
NOR2    gate2933  (.A(n672gat), .B(n670gat), .Z(n801gat) ) ;
NOR2    gate2934  (.A(n2931gat), .B(n801gat), .Z(n879gat) ) ;
NOR2    gate2935  (.A(n1123gat), .B(n1225gat), .Z(n1255gat) ) ;
NOR2    gate2936  (.A(n1255gat), .B(n2943gat), .Z(n1009gat) ) ;
NOR2    gate2937  (.A(n406gat), .B(n407gat), .Z(n409gat) ) ;
NOR2    gate2938  (.A(n415gat), .B(n356gat), .Z(n292gat) ) ;
NOR2    gate2939  (.A(n409gat), .B(n291gat), .Z(n419gat) ) ;
NOR2    gate2940  (.A(n1281gat), .B(n1123gat), .Z(n1243gat) ) ;
NOR2    gate2941  (.A(n2960gat), .B(n1243gat), .Z(n1171gat) ) ;
NOR2    gate2942  (.A(n1123gat), .B(n1134gat), .Z(n1244gat) ) ;
NOR2    gate2943  (.A(n1244gat), .B(n2969gat), .Z(n1265gat) ) ;
NOR2    gate2944  (.A(n1123gat), .B(n1044gat), .Z(n1254gat) ) ;
NOR2    gate2945  (.A(n2942gat), .B(n1254gat), .Z(n1008gat) ) ;
NOR2    gate2946  (.A(n930gat), .B(n1123gat), .Z(n1253gat) ) ;
NOR2    gate2947  (.A(n2965gat), .B(n1253gat), .Z(n1266gat) ) ;
NOR2    gate2948  (.A(n1120gat), .B(n1123gat), .Z(n1200gat) ) ;
NOR2    gate2949  (.A(n2961gat), .B(n1200gat), .Z(n1172gat) ) ;
NOR2    gate2950  (.A(n1123gat), .B(n1071gat), .Z(n1251gat) ) ;
NOR2    gate2951  (.A(n2967gat), .B(n1251gat), .Z(n1259gat) ) ;
NOR2    gate2952  (.A(n1123gat), .B(n1034gat), .Z(n1212gat) ) ;
NOR2    gate2953  (.A(n1212gat), .B(n2968gat), .Z(n1263gat) ) ;
NOR2    gate2954  (.A(n2944gat), .B(n2945gat), .Z(n978gat) ) ;
NOR2    gate2955  (.A(n1123gat), .B(n1284gat), .Z(n1199gat) ) ;
NOR2    gate2956  (.A(n1199gat), .B(n2962gat), .Z(n1252gat) ) ;
NOR2    gate2957  (.A(n1773gat), .B(n1769gat), .Z(n1757gat) ) ;

endmodule
