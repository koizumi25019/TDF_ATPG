module s38417 (g51, g563, g1249, g1943, g2637
    , g3212, g3213, g3214, g3215, g3216
    , g3217, g3218, g3219, g3220, g3221
    , g3222, g3223, g3224, g3225, g3226
    , g3227, g3228, g3229, g3230, g3231
    , g3232, g3233, g3234, CLK
    , g3993, g4088, g4090, g4200, g4321
    , g4323, g4450, g4590, g5388, g5437
    , g5472, g5511, g5549, g5555, g5595
    , g5612, g5629, g5637, g5648, g5657
    , g5686, g5695, g5738, g5747, g5796
    , g6225, g6231, g6313, g6368, g6442
    , g6447, g6485, g6518, g6573, g6642
    , g6677, g6712, g6750, g6782, g6837
    , g6895, g6911, g6944, g6979, g7014
    , g7052, g7084, g7161, g7194, g7229
    , g7264, g7302, g7334, g7357, g7390
    , g7425, g7487, g7519, g7909, g7956
    , g7961, g8007, g8012, g8021, g8023
    , g8030, g8082, g8087, g8096, g8106
    , g8167, g8175, g8249, g8251, g8258
    , g8259, g8260, g8261, g8262, g8263
    , g8264, g8265, g8266, g8267, g8268
    , g8269, g8270, g8271, g8272, g8273
    , g8274, g8275, g16297, g16355, g16399
    , g16437, g16496, g24734, g25420, g25435
    , g25442, g25489, g26104, g26135, g26149
    , g27380) ;

input   g51, g563, g1249, g1943, g2637
    , g3212, g3213, g3214, g3215, g3216
    , g3217, g3218, g3219, g3220, g3221
    , g3222, g3223, g3224, g3225, g3226
    , g3227, g3228, g3229, g3230, g3231
    , g3232, g3233, g3234, CLK ;

output  g3993, g4088, g4090, g4200, g4321
    , g4323, g4450, g4590, g5388, g5437
    , g5472, g5511, g5549, g5555, g5595
    , g5612, g5629, g5637, g5648, g5657
    , g5686, g5695, g5738, g5747, g5796
    , g6225, g6231, g6313, g6368, g6442
    , g6447, g6485, g6518, g6573, g6642
    , g6677, g6712, g6750, g6782, g6837
    , g6895, g6911, g6944, g6979, g7014
    , g7052, g7084, g7161, g7194, g7229
    , g7264, g7302, g7334, g7357, g7390
    , g7425, g7487, g7519, g7909, g7956
    , g7961, g8007, g8012, g8021, g8023
    , g8030, g8082, g8087, g8096, g8106
    , g8167, g8175, g8249, g8251, g8258
    , g8259, g8260, g8261, g8262, g8263
    , g8264, g8265, g8266, g8267, g8268
    , g8269, g8270, g8271, g8272, g8273
    , g8274, g8275, g16297, g16355, g16399
    , g16437, g16496, g24734, g25420, g25435
    , g25442, g25489, g26104, g26135, g26149
    , g27380 ;

INV     gate0  (.A(II13275), .Z(g3993) ) ;
INV     gate1  (.A(II13316), .Z(g4088) ) ;
INV     gate2  (.A(II13320), .Z(g4090) ) ;
INV     gate3  (.A(II13366), .Z(g4200) ) ;
INV     gate4  (.A(II13417), .Z(g4321) ) ;
INV     gate5  (.A(II13421), .Z(g4323) ) ;
INV     gate6  (.A(II13478), .Z(g4450) ) ;
INV     gate7  (.A(II13538), .Z(g4590) ) ;
INV     gate8  (.A(II13892), .Z(g5388) ) ;
INV     gate9  (.A(II13999), .Z(g5437) ) ;
INV     gate10  (.A(II14006), .Z(g5472) ) ;
INV     gate11  (.A(II14017), .Z(g5511) ) ;
INV     gate12  (.A(II14027), .Z(g5549) ) ;
INV     gate13  (.A(II14037), .Z(g5555) ) ;
INV     gate14  (.A(II14049), .Z(g5595) ) ;
INV     gate15  (.A(II14066), .Z(g5612) ) ;
INV     gate16  (.A(II14083), .Z(g5629) ) ;
INV     gate17  (.A(II14091), .Z(g5637) ) ;
INV     gate18  (.A(II14104), .Z(g5648) ) ;
INV     gate19  (.A(II14113), .Z(g5657) ) ;
INV     gate20  (.A(II14134), .Z(g5686) ) ;
INV     gate21  (.A(II14143), .Z(g5695) ) ;
INV     gate22  (.A(II14182), .Z(g5738) ) ;
INV     gate23  (.A(II14191), .Z(g5747) ) ;
INV     gate24  (.A(II14238), .Z(g5796) ) ;
INV     gate25  (.A(II14704), .Z(g6225) ) ;
INV     gate26  (.A(II14712), .Z(g6231) ) ;
INV     gate27  (.A(II14731), .Z(g6313) ) ;
INV     gate28  (.A(II14739), .Z(g6368) ) ;
INV     gate29  (.A(II14755), .Z(g6442) ) ;
INV     gate30  (.A(II14760), .Z(g6447) ) ;
INV     gate31  (.A(II14766), .Z(g6485) ) ;
INV     gate32  (.A(II14775), .Z(g6518) ) ;
INV     gate33  (.A(II14783), .Z(g6573) ) ;
INV     gate34  (.A(II14799), .Z(g6642) ) ;
INV     gate35  (.A(II14808), .Z(g6677) ) ;
INV     gate36  (.A(II14816), .Z(g6712) ) ;
INV     gate37  (.A(II14822), .Z(g6750) ) ;
INV     gate38  (.A(II14831), .Z(g6782) ) ;
INV     gate39  (.A(II14839), .Z(g6837) ) ;
INV     gate40  (.A(II14848), .Z(g6895) ) ;
INV     gate41  (.A(II14857), .Z(g6911) ) ;
INV     gate42  (.A(II14865), .Z(g6944) ) ;
INV     gate43  (.A(II14874), .Z(g6979) ) ;
INV     gate44  (.A(II14882), .Z(g7014) ) ;
INV     gate45  (.A(II14888), .Z(g7052) ) ;
INV     gate46  (.A(II14897), .Z(g7084) ) ;
INV     gate47  (.A(II14917), .Z(g7161) ) ;
INV     gate48  (.A(II14925), .Z(g7194) ) ;
INV     gate49  (.A(II14934), .Z(g7229) ) ;
INV     gate50  (.A(II14942), .Z(g7264) ) ;
INV     gate51  (.A(II14948), .Z(g7302) ) ;
INV     gate52  (.A(II14957), .Z(g7334) ) ;
INV     gate53  (.A(II14973), .Z(g7357) ) ;
INV     gate54  (.A(II14981), .Z(g7390) ) ;
INV     gate55  (.A(II14990), .Z(g7425) ) ;
INV     gate56  (.A(II15012), .Z(g7487) ) ;
INV     gate57  (.A(II15019), .Z(g7519) ) ;
INV     gate58  (.A(II15226), .Z(g7909) ) ;
INV     gate59  (.A(II15262), .Z(g7956) ) ;
INV     gate60  (.A(II15267), .Z(g7961) ) ;
INV     gate61  (.A(II15299), .Z(g8007) ) ;
INV     gate62  (.A(II15304), .Z(g8012) ) ;
INV     gate63  (.A(II15313), .Z(g8021) ) ;
INV     gate64  (.A(II15317), .Z(g8023) ) ;
INV     gate65  (.A(II15326), .Z(g8030) ) ;
INV     gate66  (.A(II15345), .Z(g8082) ) ;
INV     gate67  (.A(II15350), .Z(g8087) ) ;
INV     gate68  (.A(II15359), .Z(g8096) ) ;
INV     gate69  (.A(II15369), .Z(g8106) ) ;
INV     gate70  (.A(II15392), .Z(g8167) ) ;
INV     gate71  (.A(II15398), .Z(g8175) ) ;
INV     gate72  (.A(II15429), .Z(g8249) ) ;
INV     gate73  (.A(II15433), .Z(g8251) ) ;
INV     gate74  (.A(II15442), .Z(g8258) ) ;
INV     gate75  (.A(II15445), .Z(g8259) ) ;
INV     gate76  (.A(II15448), .Z(g8260) ) ;
INV     gate77  (.A(II15451), .Z(g8261) ) ;
INV     gate78  (.A(II15454), .Z(g8262) ) ;
INV     gate79  (.A(II15457), .Z(g8263) ) ;
INV     gate80  (.A(II15460), .Z(g8264) ) ;
INV     gate81  (.A(II15463), .Z(g8265) ) ;
INV     gate82  (.A(II15466), .Z(g8266) ) ;
INV     gate83  (.A(II15469), .Z(g8267) ) ;
INV     gate84  (.A(II15472), .Z(g8268) ) ;
INV     gate85  (.A(II15475), .Z(g8269) ) ;
INV     gate86  (.A(II15478), .Z(g8270) ) ;
INV     gate87  (.A(II15481), .Z(g8271) ) ;
INV     gate88  (.A(II15484), .Z(g8272) ) ;
INV     gate89  (.A(II15487), .Z(g8273) ) ;
INV     gate90  (.A(II15490), .Z(g8274) ) ;
INV     gate91  (.A(II15493), .Z(g8275) ) ;
INV     gate92  (.A(II22382), .Z(g16297) ) ;
INV     gate93  (.A(II22414), .Z(g16355) ) ;
INV     gate94  (.A(II22444), .Z(g16399) ) ;
INV     gate95  (.A(II22475), .Z(g16437) ) ;
INV     gate96  (.A(II22590), .Z(g16496) ) ;
INV     gate97  (.A(II32248), .Z(g24734) ) ;
INV     gate98  (.A(II33246), .Z(g25420) ) ;
INV     gate99  (.A(II33257), .Z(g25435) ) ;
INV     gate100  (.A(II33265), .Z(g25442) ) ;
OR2     gate101  (.A(g24795), .B(g16466), .Z(g25489) ) ;
INV     gate102  (.A(II33999), .Z(g26104) ) ;
INV     gate103  (.A(II34029), .Z(g26135) ) ;
INV     gate104  (.A(II34041), .Z(g26149) ) ;
INV     gate105  (.A(II35708), .Z(g27380) ) ;
INV     gate106  (.A(II22527), .Z(g16475) ) ;
DFF     gate107  (.D(g16475), .CP(CLK), .Q(g2814) ) ;
INV     gate108  (.A(II27038), .Z(g20571) ) ;
DFF     gate109  (.D(g20571), .CP(CLK), .Q(g2817) ) ;
INV     gate110  (.A(II27089), .Z(g20588) ) ;
DFF     gate111  (.D(g20588), .CP(CLK), .Q(g2933) ) ;
INV     gate112  (.A(II28479), .Z(g21951) ) ;
DFF     gate113  (.D(g21951), .CP(CLK), .Q(g2950) ) ;
INV     gate114  (.A(II30398), .Z(g23315) ) ;
DFF     gate115  (.D(g23315), .CP(CLK), .Q(g2883) ) ;
INV     gate116  (.A(II31943), .Z(g24423) ) ;
DFF     gate117  (.D(g24423), .CP(CLK), .Q(g2888) ) ;
INV     gate118  (.A(II33003), .Z(g25175) ) ;
DFF     gate119  (.D(g25175), .CP(CLK), .Q(g2896) ) ;
INV     gate120  (.A(II33909), .Z(g26019) ) ;
DFF     gate121  (.D(g26019), .CP(CLK), .Q(g2892) ) ;
INV     gate122  (.A(II34848), .Z(g26747) ) ;
DFF     gate123  (.D(g26747), .CP(CLK), .Q(g2903) ) ;
INV     gate124  (.A(II35548), .Z(g27237) ) ;
DFF     gate125  (.D(g27237), .CP(CLK), .Q(g2900) ) ;
INV     gate126  (.A(II36156), .Z(g27715) ) ;
DFF     gate127  (.D(g27715), .CP(CLK), .Q(g2908) ) ;
INV     gate128  (.A(II31946), .Z(g24424) ) ;
DFF     gate129  (.D(g24424), .CP(CLK), .Q(g2912) ) ;
INV     gate130  (.A(II33000), .Z(g25174) ) ;
DFF     gate131  (.D(g25174), .CP(CLK), .Q(g2917) ) ;
INV     gate132  (.A(II33912), .Z(g26020) ) ;
DFF     gate133  (.D(g26020), .CP(CLK), .Q(g2924) ) ;
INV     gate134  (.A(II34845), .Z(g26746) ) ;
DFF     gate135  (.D(g26746), .CP(CLK), .Q(g2920) ) ;
INV     gate136  (.A(II25246), .Z(g19061) ) ;
DFF     gate137  (.D(g19061), .CP(CLK), .Q(g2984) ) ;
INV     gate138  (.A(II25243), .Z(g19060) ) ;
DFF     gate139  (.D(g19060), .CP(CLK), .Q(g2985) ) ;
INV     gate140  (.A(II25249), .Z(g19062) ) ;
DFF     gate141  (.D(g19062), .CP(CLK), .Q(g2930) ) ;
DFF     gate142  (.D(g2930), .CP(CLK), .Q(g2929) ) ;
INV     gate143  (.A(II22584), .Z(g16494) ) ;
DFF     gate144  (.D(g16494), .CP(CLK), .Q(g2879) ) ;
INV     gate145  (.A(II22530), .Z(g16476) ) ;
DFF     gate146  (.D(g16476), .CP(CLK), .Q(g2934) ) ;
INV     gate147  (.A(II22533), .Z(g16477) ) ;
DFF     gate148  (.D(g16477), .CP(CLK), .Q(g2935) ) ;
INV     gate149  (.A(II22536), .Z(g16478) ) ;
DFF     gate150  (.D(g16478), .CP(CLK), .Q(g2938) ) ;
INV     gate151  (.A(II22539), .Z(g16479) ) ;
DFF     gate152  (.D(g16479), .CP(CLK), .Q(g2941) ) ;
INV     gate153  (.A(II22542), .Z(g16480) ) ;
DFF     gate154  (.D(g16480), .CP(CLK), .Q(g2944) ) ;
INV     gate155  (.A(II22545), .Z(g16481) ) ;
DFF     gate156  (.D(g16481), .CP(CLK), .Q(g2947) ) ;
INV     gate157  (.A(II22548), .Z(g16482) ) ;
DFF     gate158  (.D(g16482), .CP(CLK), .Q(g2953) ) ;
INV     gate159  (.A(II22551), .Z(g16483) ) ;
DFF     gate160  (.D(g16483), .CP(CLK), .Q(g2956) ) ;
INV     gate161  (.A(II22554), .Z(g16484) ) ;
DFF     gate162  (.D(g16484), .CP(CLK), .Q(g2959) ) ;
INV     gate163  (.A(II22557), .Z(g16485) ) ;
DFF     gate164  (.D(g16485), .CP(CLK), .Q(g2962) ) ;
INV     gate165  (.A(II22560), .Z(g16486) ) ;
DFF     gate166  (.D(g16486), .CP(CLK), .Q(g2963) ) ;
INV     gate167  (.A(II22563), .Z(g16487) ) ;
DFF     gate168  (.D(g16487), .CP(CLK), .Q(g2966) ) ;
INV     gate169  (.A(II22566), .Z(g16488) ) ;
DFF     gate170  (.D(g16488), .CP(CLK), .Q(g2969) ) ;
INV     gate171  (.A(II22569), .Z(g16489) ) ;
DFF     gate172  (.D(g16489), .CP(CLK), .Q(g2972) ) ;
INV     gate173  (.A(II22572), .Z(g16490) ) ;
DFF     gate174  (.D(g16490), .CP(CLK), .Q(g2975) ) ;
INV     gate175  (.A(II22575), .Z(g16491) ) ;
DFF     gate176  (.D(g16491), .CP(CLK), .Q(g2978) ) ;
INV     gate177  (.A(II22578), .Z(g16492) ) ;
DFF     gate178  (.D(g16492), .CP(CLK), .Q(g2981) ) ;
INV     gate179  (.A(II22581), .Z(g16493) ) ;
DFF     gate180  (.D(g16493), .CP(CLK), .Q(g2874) ) ;
INV     gate181  (.A(II27041), .Z(g20572) ) ;
DFF     gate182  (.D(g20572), .CP(CLK), .Q(g1506) ) ;
INV     gate183  (.A(II27044), .Z(g20573) ) ;
DFF     gate184  (.D(g20573), .CP(CLK), .Q(g1501) ) ;
INV     gate185  (.A(II27047), .Z(g20574) ) ;
DFF     gate186  (.D(g20574), .CP(CLK), .Q(g1496) ) ;
INV     gate187  (.A(II27050), .Z(g20575) ) ;
DFF     gate188  (.D(g20575), .CP(CLK), .Q(g1491) ) ;
INV     gate189  (.A(II27053), .Z(g20576) ) ;
DFF     gate190  (.D(g20576), .CP(CLK), .Q(g1486) ) ;
INV     gate191  (.A(II27056), .Z(g20577) ) ;
DFF     gate192  (.D(g20577), .CP(CLK), .Q(g1481) ) ;
INV     gate193  (.A(II27059), .Z(g20578) ) ;
DFF     gate194  (.D(g20578), .CP(CLK), .Q(g1476) ) ;
INV     gate195  (.A(II27062), .Z(g20579) ) ;
DFF     gate196  (.D(g20579), .CP(CLK), .Q(g1471) ) ;
INV     gate197  (.A(II30392), .Z(g23313) ) ;
DFF     gate198  (.D(g23313), .CP(CLK), .Q(g2877) ) ;
INV     gate199  (.A(II28506), .Z(g21960) ) ;
DFF     gate200  (.D(g21960), .CP(CLK), .Q(g2861) ) ;
DFF     gate201  (.D(g2861), .CP(CLK), .Q(g813) ) ;
INV     gate202  (.A(II28509), .Z(g21961) ) ;
DFF     gate203  (.D(g21961), .CP(CLK), .Q(g2864) ) ;
DFF     gate204  (.D(g2864), .CP(CLK), .Q(g809) ) ;
INV     gate205  (.A(II28512), .Z(g21962) ) ;
DFF     gate206  (.D(g21962), .CP(CLK), .Q(g2867) ) ;
DFF     gate207  (.D(g2867), .CP(CLK), .Q(g805) ) ;
INV     gate208  (.A(II28515), .Z(g21963) ) ;
DFF     gate209  (.D(g21963), .CP(CLK), .Q(g2870) ) ;
DFF     gate210  (.D(g2870), .CP(CLK), .Q(g801) ) ;
INV     gate211  (.A(II28467), .Z(g21947) ) ;
DFF     gate212  (.D(g21947), .CP(CLK), .Q(g2818) ) ;
DFF     gate213  (.D(g2818), .CP(CLK), .Q(g797) ) ;
INV     gate214  (.A(II28470), .Z(g21948) ) ;
DFF     gate215  (.D(g21948), .CP(CLK), .Q(g2821) ) ;
DFF     gate216  (.D(g2821), .CP(CLK), .Q(g793) ) ;
INV     gate217  (.A(II28473), .Z(g21949) ) ;
DFF     gate218  (.D(g21949), .CP(CLK), .Q(g2824) ) ;
DFF     gate219  (.D(g2824), .CP(CLK), .Q(g789) ) ;
INV     gate220  (.A(II28476), .Z(g21950) ) ;
DFF     gate221  (.D(g21950), .CP(CLK), .Q(g2827) ) ;
DFF     gate222  (.D(g2827), .CP(CLK), .Q(g785) ) ;
INV     gate223  (.A(II30389), .Z(g23312) ) ;
DFF     gate224  (.D(g23312), .CP(CLK), .Q(g2830) ) ;
DFF     gate225  (.D(g2830), .CP(CLK), .Q(g2873) ) ;
INV     gate226  (.A(II28482), .Z(g21952) ) ;
DFF     gate227  (.D(g21952), .CP(CLK), .Q(g2833) ) ;
DFF     gate228  (.D(g2833), .CP(CLK), .Q(g125) ) ;
INV     gate229  (.A(II28485), .Z(g21953) ) ;
DFF     gate230  (.D(g21953), .CP(CLK), .Q(g2836) ) ;
DFF     gate231  (.D(g2836), .CP(CLK), .Q(g121) ) ;
INV     gate232  (.A(II28488), .Z(g21954) ) ;
DFF     gate233  (.D(g21954), .CP(CLK), .Q(g2839) ) ;
DFF     gate234  (.D(g2839), .CP(CLK), .Q(g117) ) ;
INV     gate235  (.A(II28491), .Z(g21955) ) ;
DFF     gate236  (.D(g21955), .CP(CLK), .Q(g2842) ) ;
DFF     gate237  (.D(g2842), .CP(CLK), .Q(g113) ) ;
INV     gate238  (.A(II28494), .Z(g21956) ) ;
DFF     gate239  (.D(g21956), .CP(CLK), .Q(g2845) ) ;
DFF     gate240  (.D(g2845), .CP(CLK), .Q(g109) ) ;
INV     gate241  (.A(II28497), .Z(g21957) ) ;
DFF     gate242  (.D(g21957), .CP(CLK), .Q(g2848) ) ;
DFF     gate243  (.D(g2848), .CP(CLK), .Q(g105) ) ;
INV     gate244  (.A(II28500), .Z(g21958) ) ;
DFF     gate245  (.D(g21958), .CP(CLK), .Q(g2851) ) ;
DFF     gate246  (.D(g2851), .CP(CLK), .Q(g101) ) ;
INV     gate247  (.A(II28503), .Z(g21959) ) ;
DFF     gate248  (.D(g21959), .CP(CLK), .Q(g2854) ) ;
DFF     gate249  (.D(g2854), .CP(CLK), .Q(g97) ) ;
INV     gate250  (.A(II30401), .Z(g23316) ) ;
DFF     gate251  (.D(g23316), .CP(CLK), .Q(g2858) ) ;
DFF     gate252  (.D(g2858), .CP(CLK), .Q(g2857) ) ;
INV     gate253  (.A(II27086), .Z(g20587) ) ;
DFF     gate254  (.D(g20587), .CP(CLK), .Q(g2200) ) ;
INV     gate255  (.A(II27080), .Z(g20585) ) ;
DFF     gate256  (.D(g20585), .CP(CLK), .Q(g2195) ) ;
INV     gate257  (.A(II27083), .Z(g20586) ) ;
DFF     gate258  (.D(g20586), .CP(CLK), .Q(g2190) ) ;
INV     gate259  (.A(II27077), .Z(g20584) ) ;
DFF     gate260  (.D(g20584), .CP(CLK), .Q(g2185) ) ;
INV     gate261  (.A(II27074), .Z(g20583) ) ;
DFF     gate262  (.D(g20583), .CP(CLK), .Q(g2180) ) ;
INV     gate263  (.A(II27071), .Z(g20582) ) ;
DFF     gate264  (.D(g20582), .CP(CLK), .Q(g2175) ) ;
INV     gate265  (.A(II27068), .Z(g20581) ) ;
DFF     gate266  (.D(g20581), .CP(CLK), .Q(g2170) ) ;
INV     gate267  (.A(II27065), .Z(g20580) ) ;
DFF     gate268  (.D(g20580), .CP(CLK), .Q(g2165) ) ;
INV     gate269  (.A(II30395), .Z(g23314) ) ;
DFF     gate270  (.D(g23314), .CP(CLK), .Q(g2878) ) ;
INV     gate271  (.A(II20709), .Z(g13475) ) ;
DFF     gate272  (.D(g13475), .CP(CLK), .Q(g3129) ) ;
DFF     gate273  (.D(g3129), .CP(CLK), .Q(g3117) ) ;
DFF     gate274  (.D(g3117), .CP(CLK), .Q(g3109) ) ;
INV     gate275  (.A(II27215), .Z(g20630) ) ;
DFF     gate276  (.D(g20630), .CP(CLK), .Q(g3210) ) ;
INV     gate277  (.A(II27218), .Z(g20631) ) ;
DFF     gate278  (.D(g20631), .CP(CLK), .Q(g3211) ) ;
INV     gate279  (.A(II27221), .Z(g20632) ) ;
DFF     gate280  (.D(g20632), .CP(CLK), .Q(g3084) ) ;
INV     gate281  (.A(II27152), .Z(g20609) ) ;
DFF     gate282  (.D(g20609), .CP(CLK), .Q(g3085) ) ;
INV     gate283  (.A(II27155), .Z(g20610) ) ;
DFF     gate284  (.D(g20610), .CP(CLK), .Q(g3086) ) ;
INV     gate285  (.A(II27158), .Z(g20611) ) ;
DFF     gate286  (.D(g20611), .CP(CLK), .Q(g3087) ) ;
INV     gate287  (.A(II27161), .Z(g20612) ) ;
DFF     gate288  (.D(g20612), .CP(CLK), .Q(g3091) ) ;
INV     gate289  (.A(II27164), .Z(g20613) ) ;
DFF     gate290  (.D(g20613), .CP(CLK), .Q(g3092) ) ;
INV     gate291  (.A(II27167), .Z(g20614) ) ;
DFF     gate292  (.D(g20614), .CP(CLK), .Q(g3093) ) ;
INV     gate293  (.A(II27170), .Z(g20615) ) ;
DFF     gate294  (.D(g20615), .CP(CLK), .Q(g3094) ) ;
INV     gate295  (.A(II27173), .Z(g20616) ) ;
DFF     gate296  (.D(g20616), .CP(CLK), .Q(g3095) ) ;
INV     gate297  (.A(II27176), .Z(g20617) ) ;
DFF     gate298  (.D(g20617), .CP(CLK), .Q(g3096) ) ;
INV     gate299  (.A(II34860), .Z(g26751) ) ;
DFF     gate300  (.D(g26751), .CP(CLK), .Q(g3097) ) ;
INV     gate301  (.A(II34863), .Z(g26752) ) ;
DFF     gate302  (.D(g26752), .CP(CLK), .Q(g3098) ) ;
INV     gate303  (.A(II34866), .Z(g26753) ) ;
DFF     gate304  (.D(g26753), .CP(CLK), .Q(g3099) ) ;
INV     gate305  (.A(II38232), .Z(g29163) ) ;
DFF     gate306  (.D(g29163), .CP(CLK), .Q(g3100) ) ;
INV     gate307  (.A(II38235), .Z(g29164) ) ;
DFF     gate308  (.D(g29164), .CP(CLK), .Q(g3101) ) ;
INV     gate309  (.A(II38238), .Z(g29165) ) ;
DFF     gate310  (.D(g29165), .CP(CLK), .Q(g3102) ) ;
INV     gate311  (.A(II39625), .Z(g30120) ) ;
DFF     gate312  (.D(g30120), .CP(CLK), .Q(g3103) ) ;
INV     gate313  (.A(II39628), .Z(g30121) ) ;
DFF     gate314  (.D(g30121), .CP(CLK), .Q(g3104) ) ;
INV     gate315  (.A(II39631), .Z(g30122) ) ;
DFF     gate316  (.D(g30122), .CP(CLK), .Q(g3105) ) ;
INV     gate317  (.A(II41047), .Z(g30941) ) ;
DFF     gate318  (.D(g30941), .CP(CLK), .Q(g3106) ) ;
INV     gate319  (.A(II41050), .Z(g30942) ) ;
DFF     gate320  (.D(g30942), .CP(CLK), .Q(g3107) ) ;
INV     gate321  (.A(II41053), .Z(g30943) ) ;
DFF     gate322  (.D(g30943), .CP(CLK), .Q(g3108) ) ;
INV     gate323  (.A(II27179), .Z(g20618) ) ;
DFF     gate324  (.D(g20618), .CP(CLK), .Q(g3155) ) ;
INV     gate325  (.A(II27182), .Z(g20619) ) ;
DFF     gate326  (.D(g20619), .CP(CLK), .Q(g3158) ) ;
INV     gate327  (.A(II27185), .Z(g20620) ) ;
DFF     gate328  (.D(g20620), .CP(CLK), .Q(g3161) ) ;
INV     gate329  (.A(II27188), .Z(g20621) ) ;
DFF     gate330  (.D(g20621), .CP(CLK), .Q(g3164) ) ;
INV     gate331  (.A(II27191), .Z(g20622) ) ;
DFF     gate332  (.D(g20622), .CP(CLK), .Q(g3167) ) ;
INV     gate333  (.A(II27194), .Z(g20623) ) ;
DFF     gate334  (.D(g20623), .CP(CLK), .Q(g3170) ) ;
INV     gate335  (.A(II27197), .Z(g20624) ) ;
DFF     gate336  (.D(g20624), .CP(CLK), .Q(g3173) ) ;
INV     gate337  (.A(II27200), .Z(g20625) ) ;
DFF     gate338  (.D(g20625), .CP(CLK), .Q(g3176) ) ;
INV     gate339  (.A(II27203), .Z(g20626) ) ;
DFF     gate340  (.D(g20626), .CP(CLK), .Q(g3179) ) ;
INV     gate341  (.A(II27206), .Z(g20627) ) ;
DFF     gate342  (.D(g20627), .CP(CLK), .Q(g3182) ) ;
INV     gate343  (.A(II27209), .Z(g20628) ) ;
DFF     gate344  (.D(g20628), .CP(CLK), .Q(g3185) ) ;
INV     gate345  (.A(II27212), .Z(g20629) ) ;
DFF     gate346  (.D(g20629), .CP(CLK), .Q(g3088) ) ;
INV     gate347  (.A(II36162), .Z(g27717) ) ;
DFF     gate348  (.D(g27717), .CP(CLK), .Q(g3191) ) ;
INV     gate349  (.A(II37197), .Z(g28316) ) ;
DFF     gate350  (.D(g28316), .CP(CLK), .Q(g3194) ) ;
INV     gate351  (.A(II37200), .Z(g28317) ) ;
DFF     gate352  (.D(g28317), .CP(CLK), .Q(g3197) ) ;
INV     gate353  (.A(II37203), .Z(g28318) ) ;
DFF     gate354  (.D(g28318), .CP(CLK), .Q(g3198) ) ;
INV     gate355  (.A(II37659), .Z(g28704) ) ;
DFF     gate356  (.D(g28704), .CP(CLK), .Q(g3201) ) ;
INV     gate357  (.A(II37662), .Z(g28705) ) ;
DFF     gate358  (.D(g28705), .CP(CLK), .Q(g3204) ) ;
INV     gate359  (.A(II37665), .Z(g28706) ) ;
DFF     gate360  (.D(g28706), .CP(CLK), .Q(g3207) ) ;
INV     gate361  (.A(II38770), .Z(g29463) ) ;
DFF     gate362  (.D(g29463), .CP(CLK), .Q(g3188) ) ;
INV     gate363  (.A(II39086), .Z(g29656) ) ;
DFF     gate364  (.D(g29656), .CP(CLK), .Q(g3133) ) ;
INV     gate365  (.A(II37641), .Z(g28698) ) ;
DFF     gate366  (.D(g28698), .CP(CLK), .Q(g3132) ) ;
INV     gate367  (.A(II38241), .Z(g29166) ) ;
DFF     gate368  (.D(g29166), .CP(CLK), .Q(g3128) ) ;
INV     gate369  (.A(II37638), .Z(g28697) ) ;
DFF     gate370  (.D(g28697), .CP(CLK), .Q(g3127) ) ;
INV     gate371  (.A(II37194), .Z(g28315) ) ;
DFF     gate372  (.D(g28315), .CP(CLK), .Q(g3126) ) ;
INV     gate373  (.A(II37635), .Z(g28696) ) ;
DFF     gate374  (.D(g28696), .CP(CLK), .Q(g3125) ) ;
INV     gate375  (.A(II37191), .Z(g28314) ) ;
DFF     gate376  (.D(g28314), .CP(CLK), .Q(g3124) ) ;
INV     gate377  (.A(II37188), .Z(g28313) ) ;
DFF     gate378  (.D(g28313), .CP(CLK), .Q(g3123) ) ;
INV     gate379  (.A(II37632), .Z(g28695) ) ;
DFF     gate380  (.D(g28695), .CP(CLK), .Q(g3120) ) ;
INV     gate381  (.A(II37629), .Z(g28694) ) ;
DFF     gate382  (.D(g28694), .CP(CLK), .Q(g3114) ) ;
INV     gate383  (.A(II37626), .Z(g28693) ) ;
DFF     gate384  (.D(g28693), .CP(CLK), .Q(g3113) ) ;
INV     gate385  (.A(II37185), .Z(g28312) ) ;
DFF     gate386  (.D(g28312), .CP(CLK), .Q(g3112) ) ;
INV     gate387  (.A(II37182), .Z(g28311) ) ;
DFF     gate388  (.D(g28311), .CP(CLK), .Q(g3110) ) ;
INV     gate389  (.A(II37179), .Z(g28310) ) ;
DFF     gate390  (.D(g28310), .CP(CLK), .Q(g3111) ) ;
INV     gate391  (.A(II38764), .Z(g29461) ) ;
DFF     gate392  (.D(g29461), .CP(CLK), .Q(g3139) ) ;
INV     gate393  (.A(II37650), .Z(g28701) ) ;
DFF     gate394  (.D(g28701), .CP(CLK), .Q(g3136) ) ;
INV     gate395  (.A(II37647), .Z(g28700) ) ;
DFF     gate396  (.D(g28700), .CP(CLK), .Q(g3134) ) ;
INV     gate397  (.A(II37644), .Z(g28699) ) ;
DFF     gate398  (.D(g28699), .CP(CLK), .Q(g3135) ) ;
INV     gate399  (.A(II38767), .Z(g29462) ) ;
DFF     gate400  (.D(g29462), .CP(CLK), .Q(g3151) ) ;
INV     gate401  (.A(II37656), .Z(g28703) ) ;
DFF     gate402  (.D(g28703), .CP(CLK), .Q(g3142) ) ;
INV     gate403  (.A(II37653), .Z(g28702) ) ;
DFF     gate404  (.D(g28702), .CP(CLK), .Q(g3147) ) ;
INV     gate405  (.A(II39089), .Z(g29657) ) ;
DFF     gate406  (.D(g29657), .CP(CLK), .Q(g185) ) ;
INV     gate407  (.A(II20514), .Z(g13405) ) ;
DFF     gate408  (.D(g13405), .CP(CLK), .Q(g138) ) ;
DFF     gate409  (.D(g138), .CP(CLK), .Q(g135) ) ;
DFF     gate410  (.D(g135), .CP(CLK), .Q(g165) ) ;
INV     gate411  (.A(II31451), .Z(g24259) ) ;
DFF     gate412  (.D(g24259), .CP(CLK), .Q(g130) ) ;
INV     gate413  (.A(II31454), .Z(g24260) ) ;
DFF     gate414  (.D(g24260), .CP(CLK), .Q(g131) ) ;
INV     gate415  (.A(II31457), .Z(g24261) ) ;
DFF     gate416  (.D(g24261), .CP(CLK), .Q(g129) ) ;
INV     gate417  (.A(II31460), .Z(g24262) ) ;
DFF     gate418  (.D(g24262), .CP(CLK), .Q(g133) ) ;
INV     gate419  (.A(II31463), .Z(g24263) ) ;
DFF     gate420  (.D(g24263), .CP(CLK), .Q(g134) ) ;
INV     gate421  (.A(II31466), .Z(g24264) ) ;
DFF     gate422  (.D(g24264), .CP(CLK), .Q(g132) ) ;
INV     gate423  (.A(II31469), .Z(g24265) ) ;
DFF     gate424  (.D(g24265), .CP(CLK), .Q(g142) ) ;
INV     gate425  (.A(II31472), .Z(g24266) ) ;
DFF     gate426  (.D(g24266), .CP(CLK), .Q(g143) ) ;
INV     gate427  (.A(II31475), .Z(g24267) ) ;
DFF     gate428  (.D(g24267), .CP(CLK), .Q(g141) ) ;
INV     gate429  (.A(II31478), .Z(g24268) ) ;
DFF     gate430  (.D(g24268), .CP(CLK), .Q(g145) ) ;
INV     gate431  (.A(II31481), .Z(g24269) ) ;
DFF     gate432  (.D(g24269), .CP(CLK), .Q(g146) ) ;
INV     gate433  (.A(II31484), .Z(g24270) ) ;
DFF     gate434  (.D(g24270), .CP(CLK), .Q(g144) ) ;
INV     gate435  (.A(II31487), .Z(g24271) ) ;
DFF     gate436  (.D(g24271), .CP(CLK), .Q(g148) ) ;
INV     gate437  (.A(II31490), .Z(g24272) ) ;
DFF     gate438  (.D(g24272), .CP(CLK), .Q(g149) ) ;
INV     gate439  (.A(II31493), .Z(g24273) ) ;
DFF     gate440  (.D(g24273), .CP(CLK), .Q(g147) ) ;
INV     gate441  (.A(II31496), .Z(g24274) ) ;
DFF     gate442  (.D(g24274), .CP(CLK), .Q(g151) ) ;
INV     gate443  (.A(II31499), .Z(g24275) ) ;
DFF     gate444  (.D(g24275), .CP(CLK), .Q(g152) ) ;
INV     gate445  (.A(II31502), .Z(g24276) ) ;
DFF     gate446  (.D(g24276), .CP(CLK), .Q(g150) ) ;
INV     gate447  (.A(II31505), .Z(g24277) ) ;
DFF     gate448  (.D(g24277), .CP(CLK), .Q(g154) ) ;
INV     gate449  (.A(II31508), .Z(g24278) ) ;
DFF     gate450  (.D(g24278), .CP(CLK), .Q(g155) ) ;
INV     gate451  (.A(II31511), .Z(g24279) ) ;
DFF     gate452  (.D(g24279), .CP(CLK), .Q(g153) ) ;
INV     gate453  (.A(II31514), .Z(g24280) ) ;
DFF     gate454  (.D(g24280), .CP(CLK), .Q(g157) ) ;
INV     gate455  (.A(II31517), .Z(g24281) ) ;
DFF     gate456  (.D(g24281), .CP(CLK), .Q(g158) ) ;
INV     gate457  (.A(II31520), .Z(g24282) ) ;
DFF     gate458  (.D(g24282), .CP(CLK), .Q(g156) ) ;
INV     gate459  (.A(II31523), .Z(g24283) ) ;
DFF     gate460  (.D(g24283), .CP(CLK), .Q(g160) ) ;
INV     gate461  (.A(II31526), .Z(g24284) ) ;
DFF     gate462  (.D(g24284), .CP(CLK), .Q(g161) ) ;
INV     gate463  (.A(II31529), .Z(g24285) ) ;
DFF     gate464  (.D(g24285), .CP(CLK), .Q(g159) ) ;
INV     gate465  (.A(II31532), .Z(g24286) ) ;
DFF     gate466  (.D(g24286), .CP(CLK), .Q(g163) ) ;
INV     gate467  (.A(II31535), .Z(g24287) ) ;
DFF     gate468  (.D(g24287), .CP(CLK), .Q(g164) ) ;
INV     gate469  (.A(II31538), .Z(g24288) ) ;
DFF     gate470  (.D(g24288), .CP(CLK), .Q(g162) ) ;
INV     gate471  (.A(II34644), .Z(g26679) ) ;
DFF     gate472  (.D(g26679), .CP(CLK), .Q(g169) ) ;
INV     gate473  (.A(II34647), .Z(g26680) ) ;
DFF     gate474  (.D(g26680), .CP(CLK), .Q(g170) ) ;
INV     gate475  (.A(II34650), .Z(g26681) ) ;
DFF     gate476  (.D(g26681), .CP(CLK), .Q(g168) ) ;
INV     gate477  (.A(II34653), .Z(g26682) ) ;
DFF     gate478  (.D(g26682), .CP(CLK), .Q(g172) ) ;
INV     gate479  (.A(II34656), .Z(g26683) ) ;
DFF     gate480  (.D(g26683), .CP(CLK), .Q(g173) ) ;
INV     gate481  (.A(II34659), .Z(g26684) ) ;
DFF     gate482  (.D(g26684), .CP(CLK), .Q(g171) ) ;
INV     gate483  (.A(II34662), .Z(g26685) ) ;
DFF     gate484  (.D(g26685), .CP(CLK), .Q(g175) ) ;
INV     gate485  (.A(II34665), .Z(g26686) ) ;
DFF     gate486  (.D(g26686), .CP(CLK), .Q(g176) ) ;
INV     gate487  (.A(II34668), .Z(g26687) ) ;
DFF     gate488  (.D(g26687), .CP(CLK), .Q(g174) ) ;
INV     gate489  (.A(II34671), .Z(g26688) ) ;
DFF     gate490  (.D(g26688), .CP(CLK), .Q(g178) ) ;
INV     gate491  (.A(II34674), .Z(g26689) ) ;
DFF     gate492  (.D(g26689), .CP(CLK), .Q(g179) ) ;
INV     gate493  (.A(II34677), .Z(g26690) ) ;
DFF     gate494  (.D(g26690), .CP(CLK), .Q(g177) ) ;
INV     gate495  (.A(II40098), .Z(g30506) ) ;
DFF     gate496  (.D(g30506), .CP(CLK), .Q(g186) ) ;
INV     gate497  (.A(II40101), .Z(g30507) ) ;
DFF     gate498  (.D(g30507), .CP(CLK), .Q(g189) ) ;
INV     gate499  (.A(II40104), .Z(g30508) ) ;
DFF     gate500  (.D(g30508), .CP(CLK), .Q(g192) ) ;
INV     gate501  (.A(II40778), .Z(g30842) ) ;
DFF     gate502  (.D(g30842), .CP(CLK), .Q(g231) ) ;
INV     gate503  (.A(II40781), .Z(g30843) ) ;
DFF     gate504  (.D(g30843), .CP(CLK), .Q(g234) ) ;
INV     gate505  (.A(II40784), .Z(g30844) ) ;
DFF     gate506  (.D(g30844), .CP(CLK), .Q(g237) ) ;
INV     gate507  (.A(II40760), .Z(g30836) ) ;
DFF     gate508  (.D(g30836), .CP(CLK), .Q(g195) ) ;
INV     gate509  (.A(II40763), .Z(g30837) ) ;
DFF     gate510  (.D(g30837), .CP(CLK), .Q(g198) ) ;
INV     gate511  (.A(II40766), .Z(g30838) ) ;
DFF     gate512  (.D(g30838), .CP(CLK), .Q(g201) ) ;
INV     gate513  (.A(II40787), .Z(g30845) ) ;
DFF     gate514  (.D(g30845), .CP(CLK), .Q(g240) ) ;
INV     gate515  (.A(II40790), .Z(g30846) ) ;
DFF     gate516  (.D(g30846), .CP(CLK), .Q(g243) ) ;
INV     gate517  (.A(II40793), .Z(g30847) ) ;
DFF     gate518  (.D(g30847), .CP(CLK), .Q(g246) ) ;
INV     gate519  (.A(II40107), .Z(g30509) ) ;
DFF     gate520  (.D(g30509), .CP(CLK), .Q(g204) ) ;
INV     gate521  (.A(II40110), .Z(g30510) ) ;
DFF     gate522  (.D(g30510), .CP(CLK), .Q(g207) ) ;
INV     gate523  (.A(II40113), .Z(g30511) ) ;
DFF     gate524  (.D(g30511), .CP(CLK), .Q(g210) ) ;
INV     gate525  (.A(II40125), .Z(g30515) ) ;
DFF     gate526  (.D(g30515), .CP(CLK), .Q(g249) ) ;
INV     gate527  (.A(II40128), .Z(g30516) ) ;
DFF     gate528  (.D(g30516), .CP(CLK), .Q(g252) ) ;
INV     gate529  (.A(II40131), .Z(g30517) ) ;
DFF     gate530  (.D(g30517), .CP(CLK), .Q(g255) ) ;
INV     gate531  (.A(II40116), .Z(g30512) ) ;
DFF     gate532  (.D(g30512), .CP(CLK), .Q(g213) ) ;
INV     gate533  (.A(II40119), .Z(g30513) ) ;
DFF     gate534  (.D(g30513), .CP(CLK), .Q(g216) ) ;
INV     gate535  (.A(II40122), .Z(g30514) ) ;
DFF     gate536  (.D(g30514), .CP(CLK), .Q(g219) ) ;
INV     gate537  (.A(II40134), .Z(g30518) ) ;
DFF     gate538  (.D(g30518), .CP(CLK), .Q(g258) ) ;
INV     gate539  (.A(II40137), .Z(g30519) ) ;
DFF     gate540  (.D(g30519), .CP(CLK), .Q(g261) ) ;
INV     gate541  (.A(II40140), .Z(g30520) ) ;
DFF     gate542  (.D(g30520), .CP(CLK), .Q(g264) ) ;
INV     gate543  (.A(II40769), .Z(g30839) ) ;
DFF     gate544  (.D(g30839), .CP(CLK), .Q(g222) ) ;
INV     gate545  (.A(II40772), .Z(g30840) ) ;
DFF     gate546  (.D(g30840), .CP(CLK), .Q(g225) ) ;
INV     gate547  (.A(II40775), .Z(g30841) ) ;
DFF     gate548  (.D(g30841), .CP(CLK), .Q(g228) ) ;
INV     gate549  (.A(II40796), .Z(g30848) ) ;
DFF     gate550  (.D(g30848), .CP(CLK), .Q(g267) ) ;
INV     gate551  (.A(II40799), .Z(g30849) ) ;
DFF     gate552  (.D(g30849), .CP(CLK), .Q(g270) ) ;
INV     gate553  (.A(II40802), .Z(g30850) ) ;
DFF     gate554  (.D(g30850), .CP(CLK), .Q(g273) ) ;
INV     gate555  (.A(II33801), .Z(g25983) ) ;
DFF     gate556  (.D(g25983), .CP(CLK), .Q(g92) ) ;
INV     gate557  (.A(II34641), .Z(g26678) ) ;
DFF     gate558  (.D(g26678), .CP(CLK), .Q(g88) ) ;
INV     gate559  (.A(II35404), .Z(g27189) ) ;
DFF     gate560  (.D(g27189), .CP(CLK), .Q(g83) ) ;
INV     gate561  (.A(II36060), .Z(g27683) ) ;
DFF     gate562  (.D(g27683), .CP(CLK), .Q(g79) ) ;
INV     gate563  (.A(II36867), .Z(g28206) ) ;
DFF     gate564  (.D(g28206), .CP(CLK), .Q(g74) ) ;
INV     gate565  (.A(II37566), .Z(g28673) ) ;
DFF     gate566  (.D(g28673), .CP(CLK), .Q(g70) ) ;
INV     gate567  (.A(II38136), .Z(g29131) ) ;
DFF     gate568  (.D(g29131), .CP(CLK), .Q(g65) ) ;
INV     gate569  (.A(II38620), .Z(g29413) ) ;
DFF     gate570  (.D(g29413), .CP(CLK), .Q(g61) ) ;
INV     gate571  (.A(II38999), .Z(g29627) ) ;
DFF     gate572  (.D(g29627), .CP(CLK), .Q(g56) ) ;
INV     gate573  (.A(II39234), .Z(g29794) ) ;
DFF     gate574  (.D(g29794), .CP(CLK), .Q(g52) ) ;
INV     gate575  (.A(II26990), .Z(g20555) ) ;
DFF     gate576  (.D(g20555), .CP(CLK), .Q(g180) ) ;
DFF     gate577  (.D(g180), .CP(CLK), .Q(g182) ) ;
DFF     gate578  (.D(g182), .CP(CLK), .Q(g181) ) ;
INV     gate579  (.A(II20517), .Z(g13406) ) ;
DFF     gate580  (.D(g13406), .CP(CLK), .Q(g276) ) ;
DFF     gate581  (.D(g276), .CP(CLK), .Q(g405) ) ;
DFF     gate582  (.D(g405), .CP(CLK), .Q(g401) ) ;
INV     gate583  (.A(II18464), .Z(g11496) ) ;
DFF     gate584  (.D(g11496), .CP(CLK), .Q(g309) ) ;
INV     gate585  (.A(II36870), .Z(g28207) ) ;
DFF     gate586  (.D(g28207), .CP(CLK), .Q(g354) ) ;
INV     gate587  (.A(II36873), .Z(g28208) ) ;
DFF     gate588  (.D(g28208), .CP(CLK), .Q(g343) ) ;
INV     gate589  (.A(II36876), .Z(g28209) ) ;
DFF     gate590  (.D(g28209), .CP(CLK), .Q(g346) ) ;
INV     gate591  (.A(II36879), .Z(g28210) ) ;
DFF     gate592  (.D(g28210), .CP(CLK), .Q(g369) ) ;
INV     gate593  (.A(II36882), .Z(g28211) ) ;
DFF     gate594  (.D(g28211), .CP(CLK), .Q(g358) ) ;
INV     gate595  (.A(II36885), .Z(g28212) ) ;
DFF     gate596  (.D(g28212), .CP(CLK), .Q(g361) ) ;
INV     gate597  (.A(II36888), .Z(g28213) ) ;
DFF     gate598  (.D(g28213), .CP(CLK), .Q(g384) ) ;
INV     gate599  (.A(II36891), .Z(g28214) ) ;
DFF     gate600  (.D(g28214), .CP(CLK), .Q(g373) ) ;
INV     gate601  (.A(II36894), .Z(g28215) ) ;
DFF     gate602  (.D(g28215), .CP(CLK), .Q(g376) ) ;
INV     gate603  (.A(II36897), .Z(g28216) ) ;
DFF     gate604  (.D(g28216), .CP(CLK), .Q(g398) ) ;
INV     gate605  (.A(II36900), .Z(g28217) ) ;
DFF     gate606  (.D(g28217), .CP(CLK), .Q(g388) ) ;
INV     gate607  (.A(II36903), .Z(g28218) ) ;
DFF     gate608  (.D(g28218), .CP(CLK), .Q(g391) ) ;
INV     gate609  (.A(II38623), .Z(g29414) ) ;
DFF     gate610  (.D(g29414), .CP(CLK), .Q(g408) ) ;
INV     gate611  (.A(II38626), .Z(g29415) ) ;
DFF     gate612  (.D(g29415), .CP(CLK), .Q(g411) ) ;
INV     gate613  (.A(II38629), .Z(g29416) ) ;
DFF     gate614  (.D(g29416), .CP(CLK), .Q(g414) ) ;
INV     gate615  (.A(II39011), .Z(g29631) ) ;
DFF     gate616  (.D(g29631), .CP(CLK), .Q(g417) ) ;
INV     gate617  (.A(II39014), .Z(g29632) ) ;
DFF     gate618  (.D(g29632), .CP(CLK), .Q(g420) ) ;
INV     gate619  (.A(II39017), .Z(g29633) ) ;
DFF     gate620  (.D(g29633), .CP(CLK), .Q(g423) ) ;
INV     gate621  (.A(II38632), .Z(g29417) ) ;
DFF     gate622  (.D(g29417), .CP(CLK), .Q(g427) ) ;
INV     gate623  (.A(II38635), .Z(g29418) ) ;
DFF     gate624  (.D(g29418), .CP(CLK), .Q(g428) ) ;
INV     gate625  (.A(II38638), .Z(g29419) ) ;
DFF     gate626  (.D(g29419), .CP(CLK), .Q(g426) ) ;
INV     gate627  (.A(II36063), .Z(g27684) ) ;
DFF     gate628  (.D(g27684), .CP(CLK), .Q(g429) ) ;
INV     gate629  (.A(II36066), .Z(g27685) ) ;
DFF     gate630  (.D(g27685), .CP(CLK), .Q(g432) ) ;
INV     gate631  (.A(II36069), .Z(g27686) ) ;
DFF     gate632  (.D(g27686), .CP(CLK), .Q(g435) ) ;
INV     gate633  (.A(II36072), .Z(g27687) ) ;
DFF     gate634  (.D(g27687), .CP(CLK), .Q(g438) ) ;
INV     gate635  (.A(II36075), .Z(g27688) ) ;
DFF     gate636  (.D(g27688), .CP(CLK), .Q(g441) ) ;
INV     gate637  (.A(II36078), .Z(g27689) ) ;
DFF     gate638  (.D(g27689), .CP(CLK), .Q(g444) ) ;
INV     gate639  (.A(II37569), .Z(g28674) ) ;
DFF     gate640  (.D(g28674), .CP(CLK), .Q(g448) ) ;
INV     gate641  (.A(II37572), .Z(g28675) ) ;
DFF     gate642  (.D(g28675), .CP(CLK), .Q(g449) ) ;
INV     gate643  (.A(II37575), .Z(g28676) ) ;
DFF     gate644  (.D(g28676), .CP(CLK), .Q(g447) ) ;
INV     gate645  (.A(II39237), .Z(g29795) ) ;
DFF     gate646  (.D(g29795), .CP(CLK), .Q(g312) ) ;
INV     gate647  (.A(II39240), .Z(g29796) ) ;
DFF     gate648  (.D(g29796), .CP(CLK), .Q(g313) ) ;
INV     gate649  (.A(II39243), .Z(g29797) ) ;
DFF     gate650  (.D(g29797), .CP(CLK), .Q(g314) ) ;
INV     gate651  (.A(II40805), .Z(g30851) ) ;
DFF     gate652  (.D(g30851), .CP(CLK), .Q(g315) ) ;
INV     gate653  (.A(II40808), .Z(g30852) ) ;
DFF     gate654  (.D(g30852), .CP(CLK), .Q(g316) ) ;
INV     gate655  (.A(II40811), .Z(g30853) ) ;
DFF     gate656  (.D(g30853), .CP(CLK), .Q(g317) ) ;
INV     gate657  (.A(II40420), .Z(g30710) ) ;
DFF     gate658  (.D(g30710), .CP(CLK), .Q(g318) ) ;
INV     gate659  (.A(II40423), .Z(g30711) ) ;
DFF     gate660  (.D(g30711), .CP(CLK), .Q(g319) ) ;
INV     gate661  (.A(II40426), .Z(g30712) ) ;
DFF     gate662  (.D(g30712), .CP(CLK), .Q(g320) ) ;
INV     gate663  (.A(II39002), .Z(g29628) ) ;
DFF     gate664  (.D(g29628), .CP(CLK), .Q(g322) ) ;
INV     gate665  (.A(II39005), .Z(g29629) ) ;
DFF     gate666  (.D(g29629), .CP(CLK), .Q(g323) ) ;
INV     gate667  (.A(II39008), .Z(g29630) ) ;
DFF     gate668  (.D(g29630), .CP(CLK), .Q(g321) ) ;
INV     gate669  (.A(II35410), .Z(g27191) ) ;
DFF     gate670  (.D(g27191), .CP(CLK), .Q(g403) ) ;
INV     gate671  (.A(II35413), .Z(g27192) ) ;
DFF     gate672  (.D(g27192), .CP(CLK), .Q(g404) ) ;
INV     gate673  (.A(II35416), .Z(g27193) ) ;
DFF     gate674  (.D(g27193), .CP(CLK), .Q(g402) ) ;
INV     gate675  (.A(II18503), .Z(g11509) ) ;
DFF     gate676  (.D(g11509), .CP(CLK), .Q(g450) ) ;
DFF     gate677  (.D(g450), .CP(CLK), .Q(g451) ) ;
INV     gate678  (.A(II18506), .Z(g11510) ) ;
DFF     gate679  (.D(g11510), .CP(CLK), .Q(g452) ) ;
DFF     gate680  (.D(g452), .CP(CLK), .Q(g453) ) ;
INV     gate681  (.A(II18509), .Z(g11511) ) ;
DFF     gate682  (.D(g11511), .CP(CLK), .Q(g454) ) ;
DFF     gate683  (.D(g454), .CP(CLK), .Q(g279) ) ;
INV     gate684  (.A(II18449), .Z(g11491) ) ;
DFF     gate685  (.D(g11491), .CP(CLK), .Q(g280) ) ;
DFF     gate686  (.D(g280), .CP(CLK), .Q(g281) ) ;
INV     gate687  (.A(II18452), .Z(g11492) ) ;
DFF     gate688  (.D(g11492), .CP(CLK), .Q(g282) ) ;
DFF     gate689  (.D(g282), .CP(CLK), .Q(g283) ) ;
INV     gate690  (.A(II18455), .Z(g11493) ) ;
DFF     gate691  (.D(g11493), .CP(CLK), .Q(g284) ) ;
DFF     gate692  (.D(g284), .CP(CLK), .Q(g285) ) ;
INV     gate693  (.A(II18458), .Z(g11494) ) ;
DFF     gate694  (.D(g11494), .CP(CLK), .Q(g286) ) ;
DFF     gate695  (.D(g286), .CP(CLK), .Q(g287) ) ;
INV     gate696  (.A(II18461), .Z(g11495) ) ;
DFF     gate697  (.D(g11495), .CP(CLK), .Q(g288) ) ;
DFF     gate698  (.D(g288), .CP(CLK), .Q(g289) ) ;
INV     gate699  (.A(II20520), .Z(g13407) ) ;
DFF     gate700  (.D(g13407), .CP(CLK), .Q(g290) ) ;
DFF     gate701  (.D(g290), .CP(CLK), .Q(g291) ) ;
INV     gate702  (.A(II25099), .Z(g19012) ) ;
DFF     gate703  (.D(g19012), .CP(CLK), .Q(g299) ) ;
INV     gate704  (.A(II29897), .Z(g23148) ) ;
DFF     gate705  (.D(g23148), .CP(CLK), .Q(g305) ) ;
INV     gate706  (.A(II29900), .Z(g23149) ) ;
DFF     gate707  (.D(g23149), .CP(CLK), .Q(g308) ) ;
INV     gate708  (.A(II29903), .Z(g23150) ) ;
DFF     gate709  (.D(g23150), .CP(CLK), .Q(g297) ) ;
INV     gate710  (.A(II29906), .Z(g23151) ) ;
DFF     gate711  (.D(g23151), .CP(CLK), .Q(g296) ) ;
INV     gate712  (.A(II29909), .Z(g23152) ) ;
DFF     gate713  (.D(g23152), .CP(CLK), .Q(g295) ) ;
INV     gate714  (.A(II29912), .Z(g23153) ) ;
DFF     gate715  (.D(g23153), .CP(CLK), .Q(g294) ) ;
INV     gate716  (.A(II25111), .Z(g19016) ) ;
DFF     gate717  (.D(g19016), .CP(CLK), .Q(g304) ) ;
INV     gate718  (.A(II25108), .Z(g19015) ) ;
DFF     gate719  (.D(g19015), .CP(CLK), .Q(g303) ) ;
INV     gate720  (.A(II25105), .Z(g19014) ) ;
DFF     gate721  (.D(g19014), .CP(CLK), .Q(g302) ) ;
INV     gate722  (.A(II25102), .Z(g19013) ) ;
DFF     gate723  (.D(g19013), .CP(CLK), .Q(g301) ) ;
INV     gate724  (.A(II32868), .Z(g25130) ) ;
DFF     gate725  (.D(g25130), .CP(CLK), .Q(g300) ) ;
INV     gate726  (.A(II35407), .Z(g27190) ) ;
DFF     gate727  (.D(g27190), .CP(CLK), .Q(g298) ) ;
INV     gate728  (.A(II18467), .Z(g11497) ) ;
DFF     gate729  (.D(g11497), .CP(CLK), .Q(g342) ) ;
DFF     gate730  (.D(g342), .CP(CLK), .Q(g349) ) ;
INV     gate731  (.A(II18470), .Z(g11498) ) ;
DFF     gate732  (.D(g11498), .CP(CLK), .Q(g350) ) ;
DFF     gate733  (.D(g350), .CP(CLK), .Q(g351) ) ;
INV     gate734  (.A(II18473), .Z(g11499) ) ;
DFF     gate735  (.D(g11499), .CP(CLK), .Q(g352) ) ;
DFF     gate736  (.D(g352), .CP(CLK), .Q(g353) ) ;
INV     gate737  (.A(II18476), .Z(g11500) ) ;
DFF     gate738  (.D(g11500), .CP(CLK), .Q(g357) ) ;
DFF     gate739  (.D(g357), .CP(CLK), .Q(g364) ) ;
INV     gate740  (.A(II18479), .Z(g11501) ) ;
DFF     gate741  (.D(g11501), .CP(CLK), .Q(g365) ) ;
DFF     gate742  (.D(g365), .CP(CLK), .Q(g366) ) ;
INV     gate743  (.A(II18482), .Z(g11502) ) ;
DFF     gate744  (.D(g11502), .CP(CLK), .Q(g367) ) ;
DFF     gate745  (.D(g367), .CP(CLK), .Q(g368) ) ;
INV     gate746  (.A(II18485), .Z(g11503) ) ;
DFF     gate747  (.D(g11503), .CP(CLK), .Q(g372) ) ;
DFF     gate748  (.D(g372), .CP(CLK), .Q(g379) ) ;
INV     gate749  (.A(II18488), .Z(g11504) ) ;
DFF     gate750  (.D(g11504), .CP(CLK), .Q(g380) ) ;
DFF     gate751  (.D(g380), .CP(CLK), .Q(g381) ) ;
INV     gate752  (.A(II18491), .Z(g11505) ) ;
DFF     gate753  (.D(g11505), .CP(CLK), .Q(g382) ) ;
DFF     gate754  (.D(g382), .CP(CLK), .Q(g383) ) ;
INV     gate755  (.A(II18494), .Z(g11506) ) ;
DFF     gate756  (.D(g11506), .CP(CLK), .Q(g387) ) ;
DFF     gate757  (.D(g387), .CP(CLK), .Q(g394) ) ;
INV     gate758  (.A(II18497), .Z(g11507) ) ;
DFF     gate759  (.D(g11507), .CP(CLK), .Q(g395) ) ;
DFF     gate760  (.D(g395), .CP(CLK), .Q(g396) ) ;
INV     gate761  (.A(II18500), .Z(g11508) ) ;
DFF     gate762  (.D(g11508), .CP(CLK), .Q(g397) ) ;
DFF     gate763  (.D(g397), .CP(CLK), .Q(g324) ) ;
INV     gate764  (.A(II20523), .Z(g13408) ) ;
DFF     gate765  (.D(g13408), .CP(CLK), .Q(g325) ) ;
DFF     gate766  (.D(g325), .CP(CLK), .Q(g331) ) ;
DFF     gate767  (.D(g331), .CP(CLK), .Q(g337) ) ;
INV     gate768  (.A(II20556), .Z(g13419) ) ;
DFF     gate769  (.D(g13419), .CP(CLK), .Q(g545) ) ;
DFF     gate770  (.D(g545), .CP(CLK), .Q(g551) ) ;
DFF     gate771  (.D(g551), .CP(CLK), .Q(g550) ) ;
INV     gate772  (.A(II29933), .Z(g23160) ) ;
DFF     gate773  (.D(g23160), .CP(CLK), .Q(g554) ) ;
INV     gate774  (.A(II26993), .Z(g20556) ) ;
DFF     gate775  (.D(g20556), .CP(CLK), .Q(g557) ) ;
INV     gate776  (.A(II26996), .Z(g20557) ) ;
DFF     gate777  (.D(g20557), .CP(CLK), .Q(g510) ) ;
INV     gate778  (.A(II22503), .Z(g16467) ) ;
DFF     gate779  (.D(g16467), .CP(CLK), .Q(g513) ) ;
DFF     gate780  (.D(g513), .CP(CLK), .Q(g523) ) ;
DFF     gate781  (.D(g523), .CP(CLK), .Q(g524) ) ;
INV     gate782  (.A(II18512), .Z(g11512) ) ;
DFF     gate783  (.D(g11512), .CP(CLK), .Q(g564) ) ;
DFF     gate784  (.D(g564), .CP(CLK), .Q(g569) ) ;
INV     gate785  (.A(II18521), .Z(g11515) ) ;
DFF     gate786  (.D(g11515), .CP(CLK), .Q(g570) ) ;
DFF     gate787  (.D(g570), .CP(CLK), .Q(g571) ) ;
INV     gate788  (.A(II18524), .Z(g11516) ) ;
DFF     gate789  (.D(g11516), .CP(CLK), .Q(g572) ) ;
DFF     gate790  (.D(g572), .CP(CLK), .Q(g573) ) ;
INV     gate791  (.A(II18527), .Z(g11517) ) ;
DFF     gate792  (.D(g11517), .CP(CLK), .Q(g574) ) ;
DFF     gate793  (.D(g574), .CP(CLK), .Q(g565) ) ;
INV     gate794  (.A(II18515), .Z(g11513) ) ;
DFF     gate795  (.D(g11513), .CP(CLK), .Q(g566) ) ;
DFF     gate796  (.D(g566), .CP(CLK), .Q(g567) ) ;
INV     gate797  (.A(II18518), .Z(g11514) ) ;
DFF     gate798  (.D(g11514), .CP(CLK), .Q(g568) ) ;
DFF     gate799  (.D(g568), .CP(CLK), .Q(g489) ) ;
INV     gate800  (.A(II20526), .Z(g13409) ) ;
DFF     gate801  (.D(g13409), .CP(CLK), .Q(g474) ) ;
DFF     gate802  (.D(g474), .CP(CLK), .Q(g481) ) ;
DFF     gate803  (.D(g481), .CP(CLK), .Q(g485) ) ;
INV     gate804  (.A(II31550), .Z(g24292) ) ;
DFF     gate805  (.D(g24292), .CP(CLK), .Q(g486) ) ;
INV     gate806  (.A(II31553), .Z(g24293) ) ;
DFF     gate807  (.D(g24293), .CP(CLK), .Q(g487) ) ;
INV     gate808  (.A(II31556), .Z(g24294) ) ;
DFF     gate809  (.D(g24294), .CP(CLK), .Q(g488) ) ;
INV     gate810  (.A(II32895), .Z(g25139) ) ;
DFF     gate811  (.D(g25139), .CP(CLK), .Q(g455) ) ;
INV     gate812  (.A(II32871), .Z(g25131) ) ;
DFF     gate813  (.D(g25131), .CP(CLK), .Q(g458) ) ;
INV     gate814  (.A(II32874), .Z(g25132) ) ;
DFF     gate815  (.D(g25132), .CP(CLK), .Q(g461) ) ;
INV     gate816  (.A(II32886), .Z(g25136) ) ;
DFF     gate817  (.D(g25136), .CP(CLK), .Q(g477) ) ;
INV     gate818  (.A(II32889), .Z(g25137) ) ;
DFF     gate819  (.D(g25137), .CP(CLK), .Q(g478) ) ;
INV     gate820  (.A(II32892), .Z(g25138) ) ;
DFF     gate821  (.D(g25138), .CP(CLK), .Q(g479) ) ;
INV     gate822  (.A(II31541), .Z(g24289) ) ;
DFF     gate823  (.D(g24289), .CP(CLK), .Q(g480) ) ;
INV     gate824  (.A(II31544), .Z(g24290) ) ;
DFF     gate825  (.D(g24290), .CP(CLK), .Q(g484) ) ;
INV     gate826  (.A(II31547), .Z(g24291) ) ;
DFF     gate827  (.D(g24291), .CP(CLK), .Q(g464) ) ;
INV     gate828  (.A(II32877), .Z(g25133) ) ;
DFF     gate829  (.D(g25133), .CP(CLK), .Q(g465) ) ;
INV     gate830  (.A(II32880), .Z(g25134) ) ;
DFF     gate831  (.D(g25134), .CP(CLK), .Q(g468) ) ;
INV     gate832  (.A(II32883), .Z(g25135) ) ;
DFF     gate833  (.D(g25135), .CP(CLK), .Q(g471) ) ;
INV     gate834  (.A(II22506), .Z(g16468) ) ;
DFF     gate835  (.D(g16468), .CP(CLK), .Q(g528) ) ;
DFF     gate836  (.D(g528), .CP(CLK), .Q(g535) ) ;
DFF     gate837  (.D(g535), .CP(CLK), .Q(g542) ) ;
INV     gate838  (.A(II25126), .Z(g19021) ) ;
DFF     gate839  (.D(g19021), .CP(CLK), .Q(g543) ) ;
DFF     gate840  (.D(g543), .CP(CLK), .Q(g544) ) ;
INV     gate841  (.A(II29930), .Z(g23159) ) ;
DFF     gate842  (.D(g23159), .CP(CLK), .Q(g548) ) ;
INV     gate843  (.A(II25129), .Z(g19022) ) ;
DFF     gate844  (.D(g19022), .CP(CLK), .Q(g549) ) ;
DFF     gate845  (.D(g549), .CP(CLK), .Q(g499) ) ;
INV     gate846  (.A(II25132), .Z(g19023) ) ;
DFF     gate847  (.D(g19023), .CP(CLK), .Q(g558) ) ;
DFF     gate848  (.D(g558), .CP(CLK), .Q(g559) ) ;
INV     gate849  (.A(II36906), .Z(g28219) ) ;
DFF     gate850  (.D(g28219), .CP(CLK), .Q(g576) ) ;
INV     gate851  (.A(II36909), .Z(g28220) ) ;
DFF     gate852  (.D(g28220), .CP(CLK), .Q(g577) ) ;
INV     gate853  (.A(II36912), .Z(g28221) ) ;
DFF     gate854  (.D(g28221), .CP(CLK), .Q(g575) ) ;
INV     gate855  (.A(II36915), .Z(g28222) ) ;
DFF     gate856  (.D(g28222), .CP(CLK), .Q(g579) ) ;
INV     gate857  (.A(II36918), .Z(g28223) ) ;
DFF     gate858  (.D(g28223), .CP(CLK), .Q(g580) ) ;
INV     gate859  (.A(II36921), .Z(g28224) ) ;
DFF     gate860  (.D(g28224), .CP(CLK), .Q(g578) ) ;
INV     gate861  (.A(II36924), .Z(g28225) ) ;
DFF     gate862  (.D(g28225), .CP(CLK), .Q(g582) ) ;
INV     gate863  (.A(II36927), .Z(g28226) ) ;
DFF     gate864  (.D(g28226), .CP(CLK), .Q(g583) ) ;
INV     gate865  (.A(II36930), .Z(g28227) ) ;
DFF     gate866  (.D(g28227), .CP(CLK), .Q(g581) ) ;
INV     gate867  (.A(II36933), .Z(g28228) ) ;
DFF     gate868  (.D(g28228), .CP(CLK), .Q(g585) ) ;
INV     gate869  (.A(II36936), .Z(g28229) ) ;
DFF     gate870  (.D(g28229), .CP(CLK), .Q(g586) ) ;
INV     gate871  (.A(II36939), .Z(g28230) ) ;
DFF     gate872  (.D(g28230), .CP(CLK), .Q(g584) ) ;
INV     gate873  (.A(II33807), .Z(g25985) ) ;
DFF     gate874  (.D(g25985), .CP(CLK), .Q(g587) ) ;
INV     gate875  (.A(II33810), .Z(g25986) ) ;
DFF     gate876  (.D(g25986), .CP(CLK), .Q(g590) ) ;
INV     gate877  (.A(II33813), .Z(g25987) ) ;
DFF     gate878  (.D(g25987), .CP(CLK), .Q(g593) ) ;
INV     gate879  (.A(II33816), .Z(g25988) ) ;
DFF     gate880  (.D(g25988), .CP(CLK), .Q(g596) ) ;
INV     gate881  (.A(II33819), .Z(g25989) ) ;
DFF     gate882  (.D(g25989), .CP(CLK), .Q(g599) ) ;
INV     gate883  (.A(II33822), .Z(g25990) ) ;
DFF     gate884  (.D(g25990), .CP(CLK), .Q(g602) ) ;
INV     gate885  (.A(II38148), .Z(g29135) ) ;
DFF     gate886  (.D(g29135), .CP(CLK), .Q(g614) ) ;
INV     gate887  (.A(II38151), .Z(g29136) ) ;
DFF     gate888  (.D(g29136), .CP(CLK), .Q(g617) ) ;
INV     gate889  (.A(II38154), .Z(g29137) ) ;
DFF     gate890  (.D(g29137), .CP(CLK), .Q(g620) ) ;
INV     gate891  (.A(II38139), .Z(g29132) ) ;
DFF     gate892  (.D(g29132), .CP(CLK), .Q(g605) ) ;
INV     gate893  (.A(II38142), .Z(g29133) ) ;
DFF     gate894  (.D(g29133), .CP(CLK), .Q(g608) ) ;
INV     gate895  (.A(II38145), .Z(g29134) ) ;
DFF     gate896  (.D(g29134), .CP(CLK), .Q(g611) ) ;
INV     gate897  (.A(II35419), .Z(g27194) ) ;
DFF     gate898  (.D(g27194), .CP(CLK), .Q(g490) ) ;
INV     gate899  (.A(II35422), .Z(g27195) ) ;
DFF     gate900  (.D(g27195), .CP(CLK), .Q(g493) ) ;
INV     gate901  (.A(II35425), .Z(g27196) ) ;
DFF     gate902  (.D(g27196), .CP(CLK), .Q(g496) ) ;
INV     gate903  (.A(II15499), .Z(g8284) ) ;
DFF     gate904  (.D(g8284), .CP(CLK), .Q(g506) ) ;
INV     gate905  (.A(II31559), .Z(g24295) ) ;
DFF     gate906  (.D(g24295), .CP(CLK), .Q(g507) ) ;
INV     gate907  (.A(II25114), .Z(g19017) ) ;
DFF     gate908  (.D(g19017), .CP(CLK), .Q(g508) ) ;
INV     gate909  (.A(II25117), .Z(g19018) ) ;
DFF     gate910  (.D(g19018), .CP(CLK), .Q(g509) ) ;
INV     gate911  (.A(II25120), .Z(g19019) ) ;
DFF     gate912  (.D(g19019), .CP(CLK), .Q(g514) ) ;
INV     gate913  (.A(II25123), .Z(g19020) ) ;
DFF     gate914  (.D(g19020), .CP(CLK), .Q(g515) ) ;
INV     gate915  (.A(II29927), .Z(g23158) ) ;
DFF     gate916  (.D(g23158), .CP(CLK), .Q(g516) ) ;
INV     gate917  (.A(II29924), .Z(g23157) ) ;
DFF     gate918  (.D(g23157), .CP(CLK), .Q(g517) ) ;
INV     gate919  (.A(II29921), .Z(g23156) ) ;
DFF     gate920  (.D(g23156), .CP(CLK), .Q(g518) ) ;
INV     gate921  (.A(II29918), .Z(g23155) ) ;
DFF     gate922  (.D(g23155), .CP(CLK), .Q(g519) ) ;
INV     gate923  (.A(II29915), .Z(g23154) ) ;
DFF     gate924  (.D(g23154), .CP(CLK), .Q(g520) ) ;
DFF     gate925  (.D(g520), .CP(CLK), .Q(g525) ) ;
INV     gate926  (.A(II20529), .Z(g13410) ) ;
DFF     gate927  (.D(g13410), .CP(CLK), .Q(g529) ) ;
INV     gate928  (.A(II20532), .Z(g13411) ) ;
DFF     gate929  (.D(g13411), .CP(CLK), .Q(g530) ) ;
INV     gate930  (.A(II20535), .Z(g13412) ) ;
DFF     gate931  (.D(g13412), .CP(CLK), .Q(g531) ) ;
INV     gate932  (.A(II20538), .Z(g13413) ) ;
DFF     gate933  (.D(g13413), .CP(CLK), .Q(g532) ) ;
INV     gate934  (.A(II20541), .Z(g13414) ) ;
DFF     gate935  (.D(g13414), .CP(CLK), .Q(g533) ) ;
INV     gate936  (.A(II20544), .Z(g13415) ) ;
DFF     gate937  (.D(g13415), .CP(CLK), .Q(g534) ) ;
INV     gate938  (.A(II20547), .Z(g13416) ) ;
DFF     gate939  (.D(g13416), .CP(CLK), .Q(g536) ) ;
INV     gate940  (.A(II20550), .Z(g13417) ) ;
DFF     gate941  (.D(g13417), .CP(CLK), .Q(g537) ) ;
INV     gate942  (.A(II33804), .Z(g25984) ) ;
DFF     gate943  (.D(g25984), .CP(CLK), .Q(g538) ) ;
INV     gate944  (.A(II20553), .Z(g13418) ) ;
DFF     gate945  (.D(g13418), .CP(CLK), .Q(g541) ) ;
INV     gate946  (.A(II20559), .Z(g13420) ) ;
DFF     gate947  (.D(g13420), .CP(CLK), .Q(g623) ) ;
DFF     gate948  (.D(g623), .CP(CLK), .Q(g626) ) ;
DFF     gate949  (.D(g626), .CP(CLK), .Q(g629) ) ;
INV     gate950  (.A(II26999), .Z(g20558) ) ;
DFF     gate951  (.D(g20558), .CP(CLK), .Q(g630) ) ;
INV     gate952  (.A(II28455), .Z(g21943) ) ;
DFF     gate953  (.D(g21943), .CP(CLK), .Q(g659) ) ;
INV     gate954  (.A(II29936), .Z(g23161) ) ;
DFF     gate955  (.D(g23161), .CP(CLK), .Q(g640) ) ;
INV     gate956  (.A(II31562), .Z(g24296) ) ;
DFF     gate957  (.D(g24296), .CP(CLK), .Q(g633) ) ;
INV     gate958  (.A(II32898), .Z(g25140) ) ;
DFF     gate959  (.D(g25140), .CP(CLK), .Q(g653) ) ;
INV     gate960  (.A(II33825), .Z(g25991) ) ;
DFF     gate961  (.D(g25991), .CP(CLK), .Q(g646) ) ;
INV     gate962  (.A(II34680), .Z(g26691) ) ;
DFF     gate963  (.D(g26691), .CP(CLK), .Q(g660) ) ;
INV     gate964  (.A(II35428), .Z(g27197) ) ;
DFF     gate965  (.D(g27197), .CP(CLK), .Q(g672) ) ;
INV     gate966  (.A(II36081), .Z(g27690) ) ;
DFF     gate967  (.D(g27690), .CP(CLK), .Q(g666) ) ;
INV     gate968  (.A(II36942), .Z(g28231) ) ;
DFF     gate969  (.D(g28231), .CP(CLK), .Q(g679) ) ;
INV     gate970  (.A(II37578), .Z(g28677) ) ;
DFF     gate971  (.D(g28677), .CP(CLK), .Q(g686) ) ;
INV     gate972  (.A(II38157), .Z(g29138) ) ;
DFF     gate973  (.D(g29138), .CP(CLK), .Q(g692) ) ;
INV     gate974  (.A(II29939), .Z(g23162) ) ;
DFF     gate975  (.D(g23162), .CP(CLK), .Q(g699) ) ;
INV     gate976  (.A(II29942), .Z(g23163) ) ;
DFF     gate977  (.D(g23163), .CP(CLK), .Q(g700) ) ;
INV     gate978  (.A(II29945), .Z(g23164) ) ;
DFF     gate979  (.D(g23164), .CP(CLK), .Q(g698) ) ;
INV     gate980  (.A(II29948), .Z(g23165) ) ;
DFF     gate981  (.D(g23165), .CP(CLK), .Q(g702) ) ;
INV     gate982  (.A(II29951), .Z(g23166) ) ;
DFF     gate983  (.D(g23166), .CP(CLK), .Q(g703) ) ;
INV     gate984  (.A(II29954), .Z(g23167) ) ;
DFF     gate985  (.D(g23167), .CP(CLK), .Q(g701) ) ;
INV     gate986  (.A(II29957), .Z(g23168) ) ;
DFF     gate987  (.D(g23168), .CP(CLK), .Q(g705) ) ;
INV     gate988  (.A(II29960), .Z(g23169) ) ;
DFF     gate989  (.D(g23169), .CP(CLK), .Q(g706) ) ;
INV     gate990  (.A(II29963), .Z(g23170) ) ;
DFF     gate991  (.D(g23170), .CP(CLK), .Q(g704) ) ;
INV     gate992  (.A(II29966), .Z(g23171) ) ;
DFF     gate993  (.D(g23171), .CP(CLK), .Q(g708) ) ;
INV     gate994  (.A(II29969), .Z(g23172) ) ;
DFF     gate995  (.D(g23172), .CP(CLK), .Q(g709) ) ;
INV     gate996  (.A(II29972), .Z(g23173) ) ;
DFF     gate997  (.D(g23173), .CP(CLK), .Q(g707) ) ;
INV     gate998  (.A(II29975), .Z(g23174) ) ;
DFF     gate999  (.D(g23174), .CP(CLK), .Q(g711) ) ;
INV     gate1000  (.A(II29978), .Z(g23175) ) ;
DFF     gate1001  (.D(g23175), .CP(CLK), .Q(g712) ) ;
INV     gate1002  (.A(II29981), .Z(g23176) ) ;
DFF     gate1003  (.D(g23176), .CP(CLK), .Q(g710) ) ;
INV     gate1004  (.A(II29984), .Z(g23177) ) ;
DFF     gate1005  (.D(g23177), .CP(CLK), .Q(g714) ) ;
INV     gate1006  (.A(II29987), .Z(g23178) ) ;
DFF     gate1007  (.D(g23178), .CP(CLK), .Q(g715) ) ;
INV     gate1008  (.A(II29990), .Z(g23179) ) ;
DFF     gate1009  (.D(g23179), .CP(CLK), .Q(g713) ) ;
INV     gate1010  (.A(II29993), .Z(g23180) ) ;
DFF     gate1011  (.D(g23180), .CP(CLK), .Q(g717) ) ;
INV     gate1012  (.A(II29996), .Z(g23181) ) ;
DFF     gate1013  (.D(g23181), .CP(CLK), .Q(g718) ) ;
INV     gate1014  (.A(II29999), .Z(g23182) ) ;
DFF     gate1015  (.D(g23182), .CP(CLK), .Q(g716) ) ;
INV     gate1016  (.A(II30002), .Z(g23183) ) ;
DFF     gate1017  (.D(g23183), .CP(CLK), .Q(g720) ) ;
INV     gate1018  (.A(II30005), .Z(g23184) ) ;
DFF     gate1019  (.D(g23184), .CP(CLK), .Q(g721) ) ;
INV     gate1020  (.A(II30008), .Z(g23185) ) ;
DFF     gate1021  (.D(g23185), .CP(CLK), .Q(g719) ) ;
INV     gate1022  (.A(II30011), .Z(g23186) ) ;
DFF     gate1023  (.D(g23186), .CP(CLK), .Q(g723) ) ;
INV     gate1024  (.A(II30014), .Z(g23187) ) ;
DFF     gate1025  (.D(g23187), .CP(CLK), .Q(g724) ) ;
INV     gate1026  (.A(II30017), .Z(g23188) ) ;
DFF     gate1027  (.D(g23188), .CP(CLK), .Q(g722) ) ;
INV     gate1028  (.A(II30020), .Z(g23189) ) ;
DFF     gate1029  (.D(g23189), .CP(CLK), .Q(g726) ) ;
INV     gate1030  (.A(II30023), .Z(g23190) ) ;
DFF     gate1031  (.D(g23190), .CP(CLK), .Q(g727) ) ;
INV     gate1032  (.A(II30026), .Z(g23191) ) ;
DFF     gate1033  (.D(g23191), .CP(CLK), .Q(g725) ) ;
INV     gate1034  (.A(II30029), .Z(g23192) ) ;
DFF     gate1035  (.D(g23192), .CP(CLK), .Q(g729) ) ;
INV     gate1036  (.A(II30032), .Z(g23193) ) ;
DFF     gate1037  (.D(g23193), .CP(CLK), .Q(g730) ) ;
INV     gate1038  (.A(II30035), .Z(g23194) ) ;
DFF     gate1039  (.D(g23194), .CP(CLK), .Q(g728) ) ;
INV     gate1040  (.A(II30038), .Z(g23195) ) ;
DFF     gate1041  (.D(g23195), .CP(CLK), .Q(g732) ) ;
INV     gate1042  (.A(II30041), .Z(g23196) ) ;
DFF     gate1043  (.D(g23196), .CP(CLK), .Q(g733) ) ;
INV     gate1044  (.A(II30044), .Z(g23197) ) ;
DFF     gate1045  (.D(g23197), .CP(CLK), .Q(g731) ) ;
INV     gate1046  (.A(II34683), .Z(g26692) ) ;
DFF     gate1047  (.D(g26692), .CP(CLK), .Q(g735) ) ;
INV     gate1048  (.A(II34686), .Z(g26693) ) ;
DFF     gate1049  (.D(g26693), .CP(CLK), .Q(g736) ) ;
INV     gate1050  (.A(II34689), .Z(g26694) ) ;
DFF     gate1051  (.D(g26694), .CP(CLK), .Q(g734) ) ;
INV     gate1052  (.A(II31565), .Z(g24297) ) ;
DFF     gate1053  (.D(g24297), .CP(CLK), .Q(g738) ) ;
INV     gate1054  (.A(II31568), .Z(g24298) ) ;
DFF     gate1055  (.D(g24298), .CP(CLK), .Q(g739) ) ;
INV     gate1056  (.A(II31571), .Z(g24299) ) ;
DFF     gate1057  (.D(g24299), .CP(CLK), .Q(g737) ) ;
INV     gate1058  (.A(II20562), .Z(g13421) ) ;
DFF     gate1059  (.D(g13421), .CP(CLK), .Q(g826) ) ;
DFF     gate1060  (.D(g826), .CP(CLK), .Q(g823) ) ;
DFF     gate1061  (.D(g823), .CP(CLK), .Q(g853) ) ;
INV     gate1062  (.A(II31574), .Z(g24300) ) ;
DFF     gate1063  (.D(g24300), .CP(CLK), .Q(g818) ) ;
INV     gate1064  (.A(II31577), .Z(g24301) ) ;
DFF     gate1065  (.D(g24301), .CP(CLK), .Q(g819) ) ;
INV     gate1066  (.A(II31580), .Z(g24302) ) ;
DFF     gate1067  (.D(g24302), .CP(CLK), .Q(g817) ) ;
INV     gate1068  (.A(II31583), .Z(g24303) ) ;
DFF     gate1069  (.D(g24303), .CP(CLK), .Q(g821) ) ;
INV     gate1070  (.A(II31586), .Z(g24304) ) ;
DFF     gate1071  (.D(g24304), .CP(CLK), .Q(g822) ) ;
INV     gate1072  (.A(II31589), .Z(g24305) ) ;
DFF     gate1073  (.D(g24305), .CP(CLK), .Q(g820) ) ;
INV     gate1074  (.A(II31592), .Z(g24306) ) ;
DFF     gate1075  (.D(g24306), .CP(CLK), .Q(g830) ) ;
INV     gate1076  (.A(II31595), .Z(g24307) ) ;
DFF     gate1077  (.D(g24307), .CP(CLK), .Q(g831) ) ;
INV     gate1078  (.A(II31598), .Z(g24308) ) ;
DFF     gate1079  (.D(g24308), .CP(CLK), .Q(g829) ) ;
INV     gate1080  (.A(II31601), .Z(g24309) ) ;
DFF     gate1081  (.D(g24309), .CP(CLK), .Q(g833) ) ;
INV     gate1082  (.A(II31604), .Z(g24310) ) ;
DFF     gate1083  (.D(g24310), .CP(CLK), .Q(g834) ) ;
INV     gate1084  (.A(II31607), .Z(g24311) ) ;
DFF     gate1085  (.D(g24311), .CP(CLK), .Q(g832) ) ;
INV     gate1086  (.A(II31610), .Z(g24312) ) ;
DFF     gate1087  (.D(g24312), .CP(CLK), .Q(g836) ) ;
INV     gate1088  (.A(II31613), .Z(g24313) ) ;
DFF     gate1089  (.D(g24313), .CP(CLK), .Q(g837) ) ;
INV     gate1090  (.A(II31616), .Z(g24314) ) ;
DFF     gate1091  (.D(g24314), .CP(CLK), .Q(g835) ) ;
INV     gate1092  (.A(II31619), .Z(g24315) ) ;
DFF     gate1093  (.D(g24315), .CP(CLK), .Q(g839) ) ;
INV     gate1094  (.A(II31622), .Z(g24316) ) ;
DFF     gate1095  (.D(g24316), .CP(CLK), .Q(g840) ) ;
INV     gate1096  (.A(II31625), .Z(g24317) ) ;
DFF     gate1097  (.D(g24317), .CP(CLK), .Q(g838) ) ;
INV     gate1098  (.A(II31628), .Z(g24318) ) ;
DFF     gate1099  (.D(g24318), .CP(CLK), .Q(g842) ) ;
INV     gate1100  (.A(II31631), .Z(g24319) ) ;
DFF     gate1101  (.D(g24319), .CP(CLK), .Q(g843) ) ;
INV     gate1102  (.A(II31634), .Z(g24320) ) ;
DFF     gate1103  (.D(g24320), .CP(CLK), .Q(g841) ) ;
INV     gate1104  (.A(II31637), .Z(g24321) ) ;
DFF     gate1105  (.D(g24321), .CP(CLK), .Q(g845) ) ;
INV     gate1106  (.A(II31640), .Z(g24322) ) ;
DFF     gate1107  (.D(g24322), .CP(CLK), .Q(g846) ) ;
INV     gate1108  (.A(II31643), .Z(g24323) ) ;
DFF     gate1109  (.D(g24323), .CP(CLK), .Q(g844) ) ;
INV     gate1110  (.A(II31646), .Z(g24324) ) ;
DFF     gate1111  (.D(g24324), .CP(CLK), .Q(g848) ) ;
INV     gate1112  (.A(II31649), .Z(g24325) ) ;
DFF     gate1113  (.D(g24325), .CP(CLK), .Q(g849) ) ;
INV     gate1114  (.A(II31652), .Z(g24326) ) ;
DFF     gate1115  (.D(g24326), .CP(CLK), .Q(g847) ) ;
INV     gate1116  (.A(II31655), .Z(g24327) ) ;
DFF     gate1117  (.D(g24327), .CP(CLK), .Q(g851) ) ;
INV     gate1118  (.A(II31658), .Z(g24328) ) ;
DFF     gate1119  (.D(g24328), .CP(CLK), .Q(g852) ) ;
INV     gate1120  (.A(II31661), .Z(g24329) ) ;
DFF     gate1121  (.D(g24329), .CP(CLK), .Q(g850) ) ;
INV     gate1122  (.A(II34695), .Z(g26696) ) ;
DFF     gate1123  (.D(g26696), .CP(CLK), .Q(g857) ) ;
INV     gate1124  (.A(II34698), .Z(g26697) ) ;
DFF     gate1125  (.D(g26697), .CP(CLK), .Q(g858) ) ;
INV     gate1126  (.A(II34701), .Z(g26698) ) ;
DFF     gate1127  (.D(g26698), .CP(CLK), .Q(g856) ) ;
INV     gate1128  (.A(II34704), .Z(g26699) ) ;
DFF     gate1129  (.D(g26699), .CP(CLK), .Q(g860) ) ;
INV     gate1130  (.A(II34707), .Z(g26700) ) ;
DFF     gate1131  (.D(g26700), .CP(CLK), .Q(g861) ) ;
INV     gate1132  (.A(II34710), .Z(g26701) ) ;
DFF     gate1133  (.D(g26701), .CP(CLK), .Q(g859) ) ;
INV     gate1134  (.A(II34713), .Z(g26702) ) ;
DFF     gate1135  (.D(g26702), .CP(CLK), .Q(g863) ) ;
INV     gate1136  (.A(II34716), .Z(g26703) ) ;
DFF     gate1137  (.D(g26703), .CP(CLK), .Q(g864) ) ;
INV     gate1138  (.A(II34719), .Z(g26704) ) ;
DFF     gate1139  (.D(g26704), .CP(CLK), .Q(g862) ) ;
INV     gate1140  (.A(II34722), .Z(g26705) ) ;
DFF     gate1141  (.D(g26705), .CP(CLK), .Q(g866) ) ;
INV     gate1142  (.A(II34725), .Z(g26706) ) ;
DFF     gate1143  (.D(g26706), .CP(CLK), .Q(g867) ) ;
INV     gate1144  (.A(II34728), .Z(g26707) ) ;
DFF     gate1145  (.D(g26707), .CP(CLK), .Q(g865) ) ;
INV     gate1146  (.A(II40143), .Z(g30521) ) ;
DFF     gate1147  (.D(g30521), .CP(CLK), .Q(g873) ) ;
INV     gate1148  (.A(II40146), .Z(g30522) ) ;
DFF     gate1149  (.D(g30522), .CP(CLK), .Q(g876) ) ;
INV     gate1150  (.A(II40149), .Z(g30523) ) ;
DFF     gate1151  (.D(g30523), .CP(CLK), .Q(g879) ) ;
INV     gate1152  (.A(II40832), .Z(g30860) ) ;
DFF     gate1153  (.D(g30860), .CP(CLK), .Q(g918) ) ;
INV     gate1154  (.A(II40835), .Z(g30861) ) ;
DFF     gate1155  (.D(g30861), .CP(CLK), .Q(g921) ) ;
INV     gate1156  (.A(II40838), .Z(g30862) ) ;
DFF     gate1157  (.D(g30862), .CP(CLK), .Q(g924) ) ;
INV     gate1158  (.A(II40814), .Z(g30854) ) ;
DFF     gate1159  (.D(g30854), .CP(CLK), .Q(g882) ) ;
INV     gate1160  (.A(II40817), .Z(g30855) ) ;
DFF     gate1161  (.D(g30855), .CP(CLK), .Q(g885) ) ;
INV     gate1162  (.A(II40820), .Z(g30856) ) ;
DFF     gate1163  (.D(g30856), .CP(CLK), .Q(g888) ) ;
INV     gate1164  (.A(II40841), .Z(g30863) ) ;
DFF     gate1165  (.D(g30863), .CP(CLK), .Q(g927) ) ;
INV     gate1166  (.A(II40844), .Z(g30864) ) ;
DFF     gate1167  (.D(g30864), .CP(CLK), .Q(g930) ) ;
INV     gate1168  (.A(II40847), .Z(g30865) ) ;
DFF     gate1169  (.D(g30865), .CP(CLK), .Q(g933) ) ;
INV     gate1170  (.A(II40152), .Z(g30524) ) ;
DFF     gate1171  (.D(g30524), .CP(CLK), .Q(g891) ) ;
INV     gate1172  (.A(II40155), .Z(g30525) ) ;
DFF     gate1173  (.D(g30525), .CP(CLK), .Q(g894) ) ;
INV     gate1174  (.A(II40158), .Z(g30526) ) ;
DFF     gate1175  (.D(g30526), .CP(CLK), .Q(g897) ) ;
INV     gate1176  (.A(II40170), .Z(g30530) ) ;
DFF     gate1177  (.D(g30530), .CP(CLK), .Q(g936) ) ;
INV     gate1178  (.A(II40173), .Z(g30531) ) ;
DFF     gate1179  (.D(g30531), .CP(CLK), .Q(g939) ) ;
INV     gate1180  (.A(II40176), .Z(g30532) ) ;
DFF     gate1181  (.D(g30532), .CP(CLK), .Q(g942) ) ;
INV     gate1182  (.A(II40161), .Z(g30527) ) ;
DFF     gate1183  (.D(g30527), .CP(CLK), .Q(g900) ) ;
INV     gate1184  (.A(II40164), .Z(g30528) ) ;
DFF     gate1185  (.D(g30528), .CP(CLK), .Q(g903) ) ;
INV     gate1186  (.A(II40167), .Z(g30529) ) ;
DFF     gate1187  (.D(g30529), .CP(CLK), .Q(g906) ) ;
INV     gate1188  (.A(II40179), .Z(g30533) ) ;
DFF     gate1189  (.D(g30533), .CP(CLK), .Q(g945) ) ;
INV     gate1190  (.A(II40182), .Z(g30534) ) ;
DFF     gate1191  (.D(g30534), .CP(CLK), .Q(g948) ) ;
INV     gate1192  (.A(II40185), .Z(g30535) ) ;
DFF     gate1193  (.D(g30535), .CP(CLK), .Q(g951) ) ;
INV     gate1194  (.A(II40823), .Z(g30857) ) ;
DFF     gate1195  (.D(g30857), .CP(CLK), .Q(g909) ) ;
INV     gate1196  (.A(II40826), .Z(g30858) ) ;
DFF     gate1197  (.D(g30858), .CP(CLK), .Q(g912) ) ;
INV     gate1198  (.A(II40829), .Z(g30859) ) ;
DFF     gate1199  (.D(g30859), .CP(CLK), .Q(g915) ) ;
INV     gate1200  (.A(II40850), .Z(g30866) ) ;
DFF     gate1201  (.D(g30866), .CP(CLK), .Q(g954) ) ;
INV     gate1202  (.A(II40853), .Z(g30867) ) ;
DFF     gate1203  (.D(g30867), .CP(CLK), .Q(g957) ) ;
INV     gate1204  (.A(II40856), .Z(g30868) ) ;
DFF     gate1205  (.D(g30868), .CP(CLK), .Q(g960) ) ;
INV     gate1206  (.A(II33828), .Z(g25992) ) ;
DFF     gate1207  (.D(g25992), .CP(CLK), .Q(g780) ) ;
INV     gate1208  (.A(II34692), .Z(g26695) ) ;
DFF     gate1209  (.D(g26695), .CP(CLK), .Q(g776) ) ;
INV     gate1210  (.A(II35431), .Z(g27198) ) ;
DFF     gate1211  (.D(g27198), .CP(CLK), .Q(g771) ) ;
INV     gate1212  (.A(II36084), .Z(g27691) ) ;
DFF     gate1213  (.D(g27691), .CP(CLK), .Q(g767) ) ;
INV     gate1214  (.A(II36945), .Z(g28232) ) ;
DFF     gate1215  (.D(g28232), .CP(CLK), .Q(g762) ) ;
INV     gate1216  (.A(II37581), .Z(g28678) ) ;
DFF     gate1217  (.D(g28678), .CP(CLK), .Q(g758) ) ;
INV     gate1218  (.A(II38160), .Z(g29139) ) ;
DFF     gate1219  (.D(g29139), .CP(CLK), .Q(g753) ) ;
INV     gate1220  (.A(II38641), .Z(g29420) ) ;
DFF     gate1221  (.D(g29420), .CP(CLK), .Q(g749) ) ;
INV     gate1222  (.A(II39020), .Z(g29634) ) ;
DFF     gate1223  (.D(g29634), .CP(CLK), .Q(g744) ) ;
INV     gate1224  (.A(II39246), .Z(g29798) ) ;
DFF     gate1225  (.D(g29798), .CP(CLK), .Q(g740) ) ;
INV     gate1226  (.A(II27002), .Z(g20559) ) ;
DFF     gate1227  (.D(g20559), .CP(CLK), .Q(g868) ) ;
DFF     gate1228  (.D(g868), .CP(CLK), .Q(g870) ) ;
DFF     gate1229  (.D(g870), .CP(CLK), .Q(g869) ) ;
INV     gate1230  (.A(II20565), .Z(g13422) ) ;
DFF     gate1231  (.D(g13422), .CP(CLK), .Q(g963) ) ;
DFF     gate1232  (.D(g963), .CP(CLK), .Q(g1092) ) ;
DFF     gate1233  (.D(g1092), .CP(CLK), .Q(g1088) ) ;
INV     gate1234  (.A(II18545), .Z(g11523) ) ;
DFF     gate1235  (.D(g11523), .CP(CLK), .Q(g996) ) ;
INV     gate1236  (.A(II36948), .Z(g28233) ) ;
DFF     gate1237  (.D(g28233), .CP(CLK), .Q(g1041) ) ;
INV     gate1238  (.A(II36951), .Z(g28234) ) ;
DFF     gate1239  (.D(g28234), .CP(CLK), .Q(g1030) ) ;
INV     gate1240  (.A(II36954), .Z(g28235) ) ;
DFF     gate1241  (.D(g28235), .CP(CLK), .Q(g1033) ) ;
INV     gate1242  (.A(II36957), .Z(g28236) ) ;
DFF     gate1243  (.D(g28236), .CP(CLK), .Q(g1056) ) ;
INV     gate1244  (.A(II36960), .Z(g28237) ) ;
DFF     gate1245  (.D(g28237), .CP(CLK), .Q(g1045) ) ;
INV     gate1246  (.A(II36963), .Z(g28238) ) ;
DFF     gate1247  (.D(g28238), .CP(CLK), .Q(g1048) ) ;
INV     gate1248  (.A(II36966), .Z(g28239) ) ;
DFF     gate1249  (.D(g28239), .CP(CLK), .Q(g1071) ) ;
INV     gate1250  (.A(II36969), .Z(g28240) ) ;
DFF     gate1251  (.D(g28240), .CP(CLK), .Q(g1060) ) ;
INV     gate1252  (.A(II36972), .Z(g28241) ) ;
DFF     gate1253  (.D(g28241), .CP(CLK), .Q(g1063) ) ;
INV     gate1254  (.A(II36975), .Z(g28242) ) ;
DFF     gate1255  (.D(g28242), .CP(CLK), .Q(g1085) ) ;
INV     gate1256  (.A(II36978), .Z(g28243) ) ;
DFF     gate1257  (.D(g28243), .CP(CLK), .Q(g1075) ) ;
INV     gate1258  (.A(II36981), .Z(g28244) ) ;
DFF     gate1259  (.D(g28244), .CP(CLK), .Q(g1078) ) ;
INV     gate1260  (.A(II38644), .Z(g29421) ) ;
DFF     gate1261  (.D(g29421), .CP(CLK), .Q(g1095) ) ;
INV     gate1262  (.A(II38647), .Z(g29422) ) ;
DFF     gate1263  (.D(g29422), .CP(CLK), .Q(g1098) ) ;
INV     gate1264  (.A(II38650), .Z(g29423) ) ;
DFF     gate1265  (.D(g29423), .CP(CLK), .Q(g1101) ) ;
INV     gate1266  (.A(II39032), .Z(g29638) ) ;
DFF     gate1267  (.D(g29638), .CP(CLK), .Q(g1104) ) ;
INV     gate1268  (.A(II39035), .Z(g29639) ) ;
DFF     gate1269  (.D(g29639), .CP(CLK), .Q(g1107) ) ;
INV     gate1270  (.A(II39038), .Z(g29640) ) ;
DFF     gate1271  (.D(g29640), .CP(CLK), .Q(g1110) ) ;
INV     gate1272  (.A(II38653), .Z(g29424) ) ;
DFF     gate1273  (.D(g29424), .CP(CLK), .Q(g1114) ) ;
INV     gate1274  (.A(II38656), .Z(g29425) ) ;
DFF     gate1275  (.D(g29425), .CP(CLK), .Q(g1115) ) ;
INV     gate1276  (.A(II38659), .Z(g29426) ) ;
DFF     gate1277  (.D(g29426), .CP(CLK), .Q(g1113) ) ;
INV     gate1278  (.A(II36087), .Z(g27692) ) ;
DFF     gate1279  (.D(g27692), .CP(CLK), .Q(g1116) ) ;
INV     gate1280  (.A(II36090), .Z(g27693) ) ;
DFF     gate1281  (.D(g27693), .CP(CLK), .Q(g1119) ) ;
INV     gate1282  (.A(II36093), .Z(g27694) ) ;
DFF     gate1283  (.D(g27694), .CP(CLK), .Q(g1122) ) ;
INV     gate1284  (.A(II36096), .Z(g27695) ) ;
DFF     gate1285  (.D(g27695), .CP(CLK), .Q(g1125) ) ;
INV     gate1286  (.A(II36099), .Z(g27696) ) ;
DFF     gate1287  (.D(g27696), .CP(CLK), .Q(g1128) ) ;
INV     gate1288  (.A(II36102), .Z(g27697) ) ;
DFF     gate1289  (.D(g27697), .CP(CLK), .Q(g1131) ) ;
INV     gate1290  (.A(II37584), .Z(g28679) ) ;
DFF     gate1291  (.D(g28679), .CP(CLK), .Q(g1135) ) ;
INV     gate1292  (.A(II37587), .Z(g28680) ) ;
DFF     gate1293  (.D(g28680), .CP(CLK), .Q(g1136) ) ;
INV     gate1294  (.A(II37590), .Z(g28681) ) ;
DFF     gate1295  (.D(g28681), .CP(CLK), .Q(g1134) ) ;
INV     gate1296  (.A(II39249), .Z(g29799) ) ;
DFF     gate1297  (.D(g29799), .CP(CLK), .Q(g999) ) ;
INV     gate1298  (.A(II39252), .Z(g29800) ) ;
DFF     gate1299  (.D(g29800), .CP(CLK), .Q(g1000) ) ;
INV     gate1300  (.A(II39255), .Z(g29801) ) ;
DFF     gate1301  (.D(g29801), .CP(CLK), .Q(g1001) ) ;
INV     gate1302  (.A(II40859), .Z(g30869) ) ;
DFF     gate1303  (.D(g30869), .CP(CLK), .Q(g1002) ) ;
INV     gate1304  (.A(II40862), .Z(g30870) ) ;
DFF     gate1305  (.D(g30870), .CP(CLK), .Q(g1003) ) ;
INV     gate1306  (.A(II40865), .Z(g30871) ) ;
DFF     gate1307  (.D(g30871), .CP(CLK), .Q(g1004) ) ;
INV     gate1308  (.A(II40429), .Z(g30713) ) ;
DFF     gate1309  (.D(g30713), .CP(CLK), .Q(g1005) ) ;
INV     gate1310  (.A(II40432), .Z(g30714) ) ;
DFF     gate1311  (.D(g30714), .CP(CLK), .Q(g1006) ) ;
INV     gate1312  (.A(II40435), .Z(g30715) ) ;
DFF     gate1313  (.D(g30715), .CP(CLK), .Q(g1007) ) ;
INV     gate1314  (.A(II39023), .Z(g29635) ) ;
DFF     gate1315  (.D(g29635), .CP(CLK), .Q(g1009) ) ;
INV     gate1316  (.A(II39026), .Z(g29636) ) ;
DFF     gate1317  (.D(g29636), .CP(CLK), .Q(g1010) ) ;
INV     gate1318  (.A(II39029), .Z(g29637) ) ;
DFF     gate1319  (.D(g29637), .CP(CLK), .Q(g1008) ) ;
INV     gate1320  (.A(II35455), .Z(g27206) ) ;
DFF     gate1321  (.D(g27206), .CP(CLK), .Q(g1090) ) ;
INV     gate1322  (.A(II35458), .Z(g27207) ) ;
DFF     gate1323  (.D(g27207), .CP(CLK), .Q(g1091) ) ;
INV     gate1324  (.A(II35461), .Z(g27208) ) ;
DFF     gate1325  (.D(g27208), .CP(CLK), .Q(g1089) ) ;
INV     gate1326  (.A(II18584), .Z(g11536) ) ;
DFF     gate1327  (.D(g11536), .CP(CLK), .Q(g1137) ) ;
DFF     gate1328  (.D(g1137), .CP(CLK), .Q(g1138) ) ;
INV     gate1329  (.A(II18587), .Z(g11537) ) ;
DFF     gate1330  (.D(g11537), .CP(CLK), .Q(g1139) ) ;
DFF     gate1331  (.D(g1139), .CP(CLK), .Q(g1140) ) ;
INV     gate1332  (.A(II18590), .Z(g11538) ) ;
DFF     gate1333  (.D(g11538), .CP(CLK), .Q(g1141) ) ;
DFF     gate1334  (.D(g1141), .CP(CLK), .Q(g966) ) ;
INV     gate1335  (.A(II18530), .Z(g11518) ) ;
DFF     gate1336  (.D(g11518), .CP(CLK), .Q(g967) ) ;
DFF     gate1337  (.D(g967), .CP(CLK), .Q(g968) ) ;
INV     gate1338  (.A(II18533), .Z(g11519) ) ;
DFF     gate1339  (.D(g11519), .CP(CLK), .Q(g969) ) ;
DFF     gate1340  (.D(g969), .CP(CLK), .Q(g970) ) ;
INV     gate1341  (.A(II18536), .Z(g11520) ) ;
DFF     gate1342  (.D(g11520), .CP(CLK), .Q(g971) ) ;
DFF     gate1343  (.D(g971), .CP(CLK), .Q(g972) ) ;
INV     gate1344  (.A(II18539), .Z(g11521) ) ;
DFF     gate1345  (.D(g11521), .CP(CLK), .Q(g973) ) ;
DFF     gate1346  (.D(g973), .CP(CLK), .Q(g974) ) ;
INV     gate1347  (.A(II18542), .Z(g11522) ) ;
DFF     gate1348  (.D(g11522), .CP(CLK), .Q(g975) ) ;
DFF     gate1349  (.D(g975), .CP(CLK), .Q(g976) ) ;
INV     gate1350  (.A(II20568), .Z(g13423) ) ;
DFF     gate1351  (.D(g13423), .CP(CLK), .Q(g977) ) ;
DFF     gate1352  (.D(g977), .CP(CLK), .Q(g978) ) ;
INV     gate1353  (.A(II25135), .Z(g19024) ) ;
DFF     gate1354  (.D(g19024), .CP(CLK), .Q(g986) ) ;
INV     gate1355  (.A(II35437), .Z(g27200) ) ;
DFF     gate1356  (.D(g27200), .CP(CLK), .Q(g992) ) ;
INV     gate1357  (.A(II35440), .Z(g27201) ) ;
DFF     gate1358  (.D(g27201), .CP(CLK), .Q(g995) ) ;
INV     gate1359  (.A(II35443), .Z(g27202) ) ;
DFF     gate1360  (.D(g27202), .CP(CLK), .Q(g984) ) ;
INV     gate1361  (.A(II35446), .Z(g27203) ) ;
DFF     gate1362  (.D(g27203), .CP(CLK), .Q(g983) ) ;
INV     gate1363  (.A(II35449), .Z(g27204) ) ;
DFF     gate1364  (.D(g27204), .CP(CLK), .Q(g982) ) ;
INV     gate1365  (.A(II35452), .Z(g27205) ) ;
DFF     gate1366  (.D(g27205), .CP(CLK), .Q(g981) ) ;
INV     gate1367  (.A(II25147), .Z(g19028) ) ;
DFF     gate1368  (.D(g19028), .CP(CLK), .Q(g991) ) ;
INV     gate1369  (.A(II25144), .Z(g19027) ) ;
DFF     gate1370  (.D(g19027), .CP(CLK), .Q(g990) ) ;
INV     gate1371  (.A(II25141), .Z(g19026) ) ;
DFF     gate1372  (.D(g19026), .CP(CLK), .Q(g989) ) ;
INV     gate1373  (.A(II25138), .Z(g19025) ) ;
DFF     gate1374  (.D(g19025), .CP(CLK), .Q(g988) ) ;
INV     gate1375  (.A(II32901), .Z(g25141) ) ;
DFF     gate1376  (.D(g25141), .CP(CLK), .Q(g987) ) ;
INV     gate1377  (.A(II35434), .Z(g27199) ) ;
DFF     gate1378  (.D(g27199), .CP(CLK), .Q(g985) ) ;
INV     gate1379  (.A(II18548), .Z(g11524) ) ;
DFF     gate1380  (.D(g11524), .CP(CLK), .Q(g1029) ) ;
DFF     gate1381  (.D(g1029), .CP(CLK), .Q(g1036) ) ;
INV     gate1382  (.A(II18551), .Z(g11525) ) ;
DFF     gate1383  (.D(g11525), .CP(CLK), .Q(g1037) ) ;
DFF     gate1384  (.D(g1037), .CP(CLK), .Q(g1038) ) ;
INV     gate1385  (.A(II18554), .Z(g11526) ) ;
DFF     gate1386  (.D(g11526), .CP(CLK), .Q(g1039) ) ;
DFF     gate1387  (.D(g1039), .CP(CLK), .Q(g1040) ) ;
INV     gate1388  (.A(II18557), .Z(g11527) ) ;
DFF     gate1389  (.D(g11527), .CP(CLK), .Q(g1044) ) ;
DFF     gate1390  (.D(g1044), .CP(CLK), .Q(g1051) ) ;
INV     gate1391  (.A(II18560), .Z(g11528) ) ;
DFF     gate1392  (.D(g11528), .CP(CLK), .Q(g1052) ) ;
DFF     gate1393  (.D(g1052), .CP(CLK), .Q(g1053) ) ;
INV     gate1394  (.A(II18563), .Z(g11529) ) ;
DFF     gate1395  (.D(g11529), .CP(CLK), .Q(g1054) ) ;
DFF     gate1396  (.D(g1054), .CP(CLK), .Q(g1055) ) ;
INV     gate1397  (.A(II18566), .Z(g11530) ) ;
DFF     gate1398  (.D(g11530), .CP(CLK), .Q(g1059) ) ;
DFF     gate1399  (.D(g1059), .CP(CLK), .Q(g1066) ) ;
INV     gate1400  (.A(II18569), .Z(g11531) ) ;
DFF     gate1401  (.D(g11531), .CP(CLK), .Q(g1067) ) ;
DFF     gate1402  (.D(g1067), .CP(CLK), .Q(g1068) ) ;
INV     gate1403  (.A(II18572), .Z(g11532) ) ;
DFF     gate1404  (.D(g11532), .CP(CLK), .Q(g1069) ) ;
DFF     gate1405  (.D(g1069), .CP(CLK), .Q(g1070) ) ;
INV     gate1406  (.A(II18575), .Z(g11533) ) ;
DFF     gate1407  (.D(g11533), .CP(CLK), .Q(g1074) ) ;
DFF     gate1408  (.D(g1074), .CP(CLK), .Q(g1081) ) ;
INV     gate1409  (.A(II18578), .Z(g11534) ) ;
DFF     gate1410  (.D(g11534), .CP(CLK), .Q(g1082) ) ;
DFF     gate1411  (.D(g1082), .CP(CLK), .Q(g1083) ) ;
INV     gate1412  (.A(II18581), .Z(g11535) ) ;
DFF     gate1413  (.D(g11535), .CP(CLK), .Q(g1084) ) ;
DFF     gate1414  (.D(g1084), .CP(CLK), .Q(g1011) ) ;
INV     gate1415  (.A(II20571), .Z(g13424) ) ;
DFF     gate1416  (.D(g13424), .CP(CLK), .Q(g1012) ) ;
DFF     gate1417  (.D(g1012), .CP(CLK), .Q(g1018) ) ;
DFF     gate1418  (.D(g1018), .CP(CLK), .Q(g1024) ) ;
INV     gate1419  (.A(II20604), .Z(g13435) ) ;
DFF     gate1420  (.D(g13435), .CP(CLK), .Q(g1231) ) ;
DFF     gate1421  (.D(g1231), .CP(CLK), .Q(g1237) ) ;
DFF     gate1422  (.D(g1237), .CP(CLK), .Q(g1236) ) ;
INV     gate1423  (.A(II30047), .Z(g23198) ) ;
DFF     gate1424  (.D(g23198), .CP(CLK), .Q(g1240) ) ;
INV     gate1425  (.A(II27005), .Z(g20560) ) ;
DFF     gate1426  (.D(g20560), .CP(CLK), .Q(g1243) ) ;
INV     gate1427  (.A(II27008), .Z(g20561) ) ;
DFF     gate1428  (.D(g20561), .CP(CLK), .Q(g1196) ) ;
INV     gate1429  (.A(II22509), .Z(g16469) ) ;
DFF     gate1430  (.D(g16469), .CP(CLK), .Q(g1199) ) ;
DFF     gate1431  (.D(g1199), .CP(CLK), .Q(g1209) ) ;
DFF     gate1432  (.D(g1209), .CP(CLK), .Q(g1210) ) ;
INV     gate1433  (.A(II18593), .Z(g11539) ) ;
DFF     gate1434  (.D(g11539), .CP(CLK), .Q(g1250) ) ;
DFF     gate1435  (.D(g1250), .CP(CLK), .Q(g1255) ) ;
INV     gate1436  (.A(II18602), .Z(g11542) ) ;
DFF     gate1437  (.D(g11542), .CP(CLK), .Q(g1256) ) ;
DFF     gate1438  (.D(g1256), .CP(CLK), .Q(g1257) ) ;
INV     gate1439  (.A(II18605), .Z(g11543) ) ;
DFF     gate1440  (.D(g11543), .CP(CLK), .Q(g1258) ) ;
DFF     gate1441  (.D(g1258), .CP(CLK), .Q(g1259) ) ;
INV     gate1442  (.A(II18608), .Z(g11544) ) ;
DFF     gate1443  (.D(g11544), .CP(CLK), .Q(g1260) ) ;
DFF     gate1444  (.D(g1260), .CP(CLK), .Q(g1251) ) ;
INV     gate1445  (.A(II18596), .Z(g11540) ) ;
DFF     gate1446  (.D(g11540), .CP(CLK), .Q(g1252) ) ;
DFF     gate1447  (.D(g1252), .CP(CLK), .Q(g1253) ) ;
INV     gate1448  (.A(II18599), .Z(g11541) ) ;
DFF     gate1449  (.D(g11541), .CP(CLK), .Q(g1254) ) ;
DFF     gate1450  (.D(g1254), .CP(CLK), .Q(g1176) ) ;
INV     gate1451  (.A(II20574), .Z(g13425) ) ;
DFF     gate1452  (.D(g13425), .CP(CLK), .Q(g1161) ) ;
DFF     gate1453  (.D(g1161), .CP(CLK), .Q(g1168) ) ;
DFF     gate1454  (.D(g1168), .CP(CLK), .Q(g1172) ) ;
INV     gate1455  (.A(II31673), .Z(g24333) ) ;
DFF     gate1456  (.D(g24333), .CP(CLK), .Q(g1173) ) ;
INV     gate1457  (.A(II31676), .Z(g24334) ) ;
DFF     gate1458  (.D(g24334), .CP(CLK), .Q(g1174) ) ;
INV     gate1459  (.A(II31679), .Z(g24335) ) ;
DFF     gate1460  (.D(g24335), .CP(CLK), .Q(g1175) ) ;
INV     gate1461  (.A(II32928), .Z(g25150) ) ;
DFF     gate1462  (.D(g25150), .CP(CLK), .Q(g1142) ) ;
INV     gate1463  (.A(II32904), .Z(g25142) ) ;
DFF     gate1464  (.D(g25142), .CP(CLK), .Q(g1145) ) ;
INV     gate1465  (.A(II32907), .Z(g25143) ) ;
DFF     gate1466  (.D(g25143), .CP(CLK), .Q(g1148) ) ;
INV     gate1467  (.A(II32919), .Z(g25147) ) ;
DFF     gate1468  (.D(g25147), .CP(CLK), .Q(g1164) ) ;
INV     gate1469  (.A(II32922), .Z(g25148) ) ;
DFF     gate1470  (.D(g25148), .CP(CLK), .Q(g1165) ) ;
INV     gate1471  (.A(II32925), .Z(g25149) ) ;
DFF     gate1472  (.D(g25149), .CP(CLK), .Q(g1166) ) ;
INV     gate1473  (.A(II31664), .Z(g24330) ) ;
DFF     gate1474  (.D(g24330), .CP(CLK), .Q(g1167) ) ;
INV     gate1475  (.A(II31667), .Z(g24331) ) ;
DFF     gate1476  (.D(g24331), .CP(CLK), .Q(g1171) ) ;
INV     gate1477  (.A(II31670), .Z(g24332) ) ;
DFF     gate1478  (.D(g24332), .CP(CLK), .Q(g1151) ) ;
INV     gate1479  (.A(II32910), .Z(g25144) ) ;
DFF     gate1480  (.D(g25144), .CP(CLK), .Q(g1152) ) ;
INV     gate1481  (.A(II32913), .Z(g25145) ) ;
DFF     gate1482  (.D(g25145), .CP(CLK), .Q(g1155) ) ;
INV     gate1483  (.A(II32916), .Z(g25146) ) ;
DFF     gate1484  (.D(g25146), .CP(CLK), .Q(g1158) ) ;
INV     gate1485  (.A(II22512), .Z(g16470) ) ;
DFF     gate1486  (.D(g16470), .CP(CLK), .Q(g1214) ) ;
DFF     gate1487  (.D(g1214), .CP(CLK), .Q(g1221) ) ;
DFF     gate1488  (.D(g1221), .CP(CLK), .Q(g1228) ) ;
INV     gate1489  (.A(II25162), .Z(g19033) ) ;
DFF     gate1490  (.D(g19033), .CP(CLK), .Q(g1229) ) ;
DFF     gate1491  (.D(g1229), .CP(CLK), .Q(g1230) ) ;
INV     gate1492  (.A(II35488), .Z(g27217) ) ;
DFF     gate1493  (.D(g27217), .CP(CLK), .Q(g1234) ) ;
INV     gate1494  (.A(II25165), .Z(g19034) ) ;
DFF     gate1495  (.D(g19034), .CP(CLK), .Q(g1235) ) ;
DFF     gate1496  (.D(g1235), .CP(CLK), .Q(g1186) ) ;
INV     gate1497  (.A(II25168), .Z(g19035) ) ;
DFF     gate1498  (.D(g19035), .CP(CLK), .Q(g1244) ) ;
DFF     gate1499  (.D(g1244), .CP(CLK), .Q(g1245) ) ;
INV     gate1500  (.A(II36984), .Z(g28245) ) ;
DFF     gate1501  (.D(g28245), .CP(CLK), .Q(g1262) ) ;
INV     gate1502  (.A(II36987), .Z(g28246) ) ;
DFF     gate1503  (.D(g28246), .CP(CLK), .Q(g1263) ) ;
INV     gate1504  (.A(II36990), .Z(g28247) ) ;
DFF     gate1505  (.D(g28247), .CP(CLK), .Q(g1261) ) ;
INV     gate1506  (.A(II36993), .Z(g28248) ) ;
DFF     gate1507  (.D(g28248), .CP(CLK), .Q(g1265) ) ;
INV     gate1508  (.A(II36996), .Z(g28249) ) ;
DFF     gate1509  (.D(g28249), .CP(CLK), .Q(g1266) ) ;
INV     gate1510  (.A(II36999), .Z(g28250) ) ;
DFF     gate1511  (.D(g28250), .CP(CLK), .Q(g1264) ) ;
INV     gate1512  (.A(II37002), .Z(g28251) ) ;
DFF     gate1513  (.D(g28251), .CP(CLK), .Q(g1268) ) ;
INV     gate1514  (.A(II37005), .Z(g28252) ) ;
DFF     gate1515  (.D(g28252), .CP(CLK), .Q(g1269) ) ;
INV     gate1516  (.A(II37008), .Z(g28253) ) ;
DFF     gate1517  (.D(g28253), .CP(CLK), .Q(g1267) ) ;
INV     gate1518  (.A(II37011), .Z(g28254) ) ;
DFF     gate1519  (.D(g28254), .CP(CLK), .Q(g1271) ) ;
INV     gate1520  (.A(II37014), .Z(g28255) ) ;
DFF     gate1521  (.D(g28255), .CP(CLK), .Q(g1272) ) ;
INV     gate1522  (.A(II37017), .Z(g28256) ) ;
DFF     gate1523  (.D(g28256), .CP(CLK), .Q(g1270) ) ;
INV     gate1524  (.A(II33834), .Z(g25994) ) ;
DFF     gate1525  (.D(g25994), .CP(CLK), .Q(g1273) ) ;
INV     gate1526  (.A(II33837), .Z(g25995) ) ;
DFF     gate1527  (.D(g25995), .CP(CLK), .Q(g1276) ) ;
INV     gate1528  (.A(II33840), .Z(g25996) ) ;
DFF     gate1529  (.D(g25996), .CP(CLK), .Q(g1279) ) ;
INV     gate1530  (.A(II33843), .Z(g25997) ) ;
DFF     gate1531  (.D(g25997), .CP(CLK), .Q(g1282) ) ;
INV     gate1532  (.A(II33846), .Z(g25998) ) ;
DFF     gate1533  (.D(g25998), .CP(CLK), .Q(g1285) ) ;
INV     gate1534  (.A(II33849), .Z(g25999) ) ;
DFF     gate1535  (.D(g25999), .CP(CLK), .Q(g1288) ) ;
INV     gate1536  (.A(II38172), .Z(g29143) ) ;
DFF     gate1537  (.D(g29143), .CP(CLK), .Q(g1300) ) ;
INV     gate1538  (.A(II38175), .Z(g29144) ) ;
DFF     gate1539  (.D(g29144), .CP(CLK), .Q(g1303) ) ;
INV     gate1540  (.A(II38178), .Z(g29145) ) ;
DFF     gate1541  (.D(g29145), .CP(CLK), .Q(g1306) ) ;
INV     gate1542  (.A(II38163), .Z(g29140) ) ;
DFF     gate1543  (.D(g29140), .CP(CLK), .Q(g1291) ) ;
INV     gate1544  (.A(II38166), .Z(g29141) ) ;
DFF     gate1545  (.D(g29141), .CP(CLK), .Q(g1294) ) ;
INV     gate1546  (.A(II38169), .Z(g29142) ) ;
DFF     gate1547  (.D(g29142), .CP(CLK), .Q(g1297) ) ;
INV     gate1548  (.A(II35464), .Z(g27209) ) ;
DFF     gate1549  (.D(g27209), .CP(CLK), .Q(g1177) ) ;
INV     gate1550  (.A(II35467), .Z(g27210) ) ;
DFF     gate1551  (.D(g27210), .CP(CLK), .Q(g1180) ) ;
INV     gate1552  (.A(II35470), .Z(g27211) ) ;
DFF     gate1553  (.D(g27211), .CP(CLK), .Q(g1183) ) ;
INV     gate1554  (.A(II15505), .Z(g8293) ) ;
DFF     gate1555  (.D(g8293), .CP(CLK), .Q(g1192) ) ;
INV     gate1556  (.A(II31682), .Z(g24336) ) ;
DFF     gate1557  (.D(g24336), .CP(CLK), .Q(g1193) ) ;
INV     gate1558  (.A(II25150), .Z(g19029) ) ;
DFF     gate1559  (.D(g19029), .CP(CLK), .Q(g1194) ) ;
INV     gate1560  (.A(II25153), .Z(g19030) ) ;
DFF     gate1561  (.D(g19030), .CP(CLK), .Q(g1195) ) ;
INV     gate1562  (.A(II25156), .Z(g19031) ) ;
DFF     gate1563  (.D(g19031), .CP(CLK), .Q(g1200) ) ;
INV     gate1564  (.A(II25159), .Z(g19032) ) ;
DFF     gate1565  (.D(g19032), .CP(CLK), .Q(g1201) ) ;
INV     gate1566  (.A(II35485), .Z(g27216) ) ;
DFF     gate1567  (.D(g27216), .CP(CLK), .Q(g1202) ) ;
INV     gate1568  (.A(II35482), .Z(g27215) ) ;
DFF     gate1569  (.D(g27215), .CP(CLK), .Q(g1203) ) ;
INV     gate1570  (.A(II35479), .Z(g27214) ) ;
DFF     gate1571  (.D(g27214), .CP(CLK), .Q(g1204) ) ;
INV     gate1572  (.A(II35476), .Z(g27213) ) ;
DFF     gate1573  (.D(g27213), .CP(CLK), .Q(g1205) ) ;
INV     gate1574  (.A(II35473), .Z(g27212) ) ;
DFF     gate1575  (.D(g27212), .CP(CLK), .Q(g1206) ) ;
DFF     gate1576  (.D(g1206), .CP(CLK), .Q(g1211) ) ;
INV     gate1577  (.A(II20577), .Z(g13426) ) ;
DFF     gate1578  (.D(g13426), .CP(CLK), .Q(g1215) ) ;
INV     gate1579  (.A(II20580), .Z(g13427) ) ;
DFF     gate1580  (.D(g13427), .CP(CLK), .Q(g1216) ) ;
INV     gate1581  (.A(II20583), .Z(g13428) ) ;
DFF     gate1582  (.D(g13428), .CP(CLK), .Q(g1217) ) ;
INV     gate1583  (.A(II20586), .Z(g13429) ) ;
DFF     gate1584  (.D(g13429), .CP(CLK), .Q(g1218) ) ;
INV     gate1585  (.A(II20589), .Z(g13430) ) ;
DFF     gate1586  (.D(g13430), .CP(CLK), .Q(g1219) ) ;
INV     gate1587  (.A(II20592), .Z(g13431) ) ;
DFF     gate1588  (.D(g13431), .CP(CLK), .Q(g1220) ) ;
INV     gate1589  (.A(II20595), .Z(g13432) ) ;
DFF     gate1590  (.D(g13432), .CP(CLK), .Q(g1222) ) ;
INV     gate1591  (.A(II20598), .Z(g13433) ) ;
DFF     gate1592  (.D(g13433), .CP(CLK), .Q(g1223) ) ;
INV     gate1593  (.A(II33831), .Z(g25993) ) ;
DFF     gate1594  (.D(g25993), .CP(CLK), .Q(g1224) ) ;
INV     gate1595  (.A(II20601), .Z(g13434) ) ;
DFF     gate1596  (.D(g13434), .CP(CLK), .Q(g1227) ) ;
INV     gate1597  (.A(II20607), .Z(g13436) ) ;
DFF     gate1598  (.D(g13436), .CP(CLK), .Q(g1309) ) ;
DFF     gate1599  (.D(g1309), .CP(CLK), .Q(g1312) ) ;
DFF     gate1600  (.D(g1312), .CP(CLK), .Q(g1315) ) ;
INV     gate1601  (.A(II27011), .Z(g20562) ) ;
DFF     gate1602  (.D(g20562), .CP(CLK), .Q(g1316) ) ;
INV     gate1603  (.A(II28458), .Z(g21944) ) ;
DFF     gate1604  (.D(g21944), .CP(CLK), .Q(g1345) ) ;
INV     gate1605  (.A(II30050), .Z(g23199) ) ;
DFF     gate1606  (.D(g23199), .CP(CLK), .Q(g1326) ) ;
INV     gate1607  (.A(II31685), .Z(g24337) ) ;
DFF     gate1608  (.D(g24337), .CP(CLK), .Q(g1319) ) ;
INV     gate1609  (.A(II32931), .Z(g25151) ) ;
DFF     gate1610  (.D(g25151), .CP(CLK), .Q(g1339) ) ;
INV     gate1611  (.A(II33852), .Z(g26000) ) ;
DFF     gate1612  (.D(g26000), .CP(CLK), .Q(g1332) ) ;
INV     gate1613  (.A(II34731), .Z(g26708) ) ;
DFF     gate1614  (.D(g26708), .CP(CLK), .Q(g1346) ) ;
INV     gate1615  (.A(II35491), .Z(g27218) ) ;
DFF     gate1616  (.D(g27218), .CP(CLK), .Q(g1358) ) ;
INV     gate1617  (.A(II36105), .Z(g27698) ) ;
DFF     gate1618  (.D(g27698), .CP(CLK), .Q(g1352) ) ;
INV     gate1619  (.A(II37020), .Z(g28257) ) ;
DFF     gate1620  (.D(g28257), .CP(CLK), .Q(g1365) ) ;
INV     gate1621  (.A(II37593), .Z(g28682) ) ;
DFF     gate1622  (.D(g28682), .CP(CLK), .Q(g1372) ) ;
INV     gate1623  (.A(II38181), .Z(g29146) ) ;
DFF     gate1624  (.D(g29146), .CP(CLK), .Q(g1378) ) ;
INV     gate1625  (.A(II30053), .Z(g23200) ) ;
DFF     gate1626  (.D(g23200), .CP(CLK), .Q(g1385) ) ;
INV     gate1627  (.A(II30056), .Z(g23201) ) ;
DFF     gate1628  (.D(g23201), .CP(CLK), .Q(g1386) ) ;
INV     gate1629  (.A(II30059), .Z(g23202) ) ;
DFF     gate1630  (.D(g23202), .CP(CLK), .Q(g1384) ) ;
INV     gate1631  (.A(II30062), .Z(g23203) ) ;
DFF     gate1632  (.D(g23203), .CP(CLK), .Q(g1388) ) ;
INV     gate1633  (.A(II30065), .Z(g23204) ) ;
DFF     gate1634  (.D(g23204), .CP(CLK), .Q(g1389) ) ;
INV     gate1635  (.A(II30068), .Z(g23205) ) ;
DFF     gate1636  (.D(g23205), .CP(CLK), .Q(g1387) ) ;
INV     gate1637  (.A(II30071), .Z(g23206) ) ;
DFF     gate1638  (.D(g23206), .CP(CLK), .Q(g1391) ) ;
INV     gate1639  (.A(II30074), .Z(g23207) ) ;
DFF     gate1640  (.D(g23207), .CP(CLK), .Q(g1392) ) ;
INV     gate1641  (.A(II30077), .Z(g23208) ) ;
DFF     gate1642  (.D(g23208), .CP(CLK), .Q(g1390) ) ;
INV     gate1643  (.A(II30080), .Z(g23209) ) ;
DFF     gate1644  (.D(g23209), .CP(CLK), .Q(g1394) ) ;
INV     gate1645  (.A(II30083), .Z(g23210) ) ;
DFF     gate1646  (.D(g23210), .CP(CLK), .Q(g1395) ) ;
INV     gate1647  (.A(II30086), .Z(g23211) ) ;
DFF     gate1648  (.D(g23211), .CP(CLK), .Q(g1393) ) ;
INV     gate1649  (.A(II30089), .Z(g23212) ) ;
DFF     gate1650  (.D(g23212), .CP(CLK), .Q(g1397) ) ;
INV     gate1651  (.A(II30092), .Z(g23213) ) ;
DFF     gate1652  (.D(g23213), .CP(CLK), .Q(g1398) ) ;
INV     gate1653  (.A(II30095), .Z(g23214) ) ;
DFF     gate1654  (.D(g23214), .CP(CLK), .Q(g1396) ) ;
INV     gate1655  (.A(II30098), .Z(g23215) ) ;
DFF     gate1656  (.D(g23215), .CP(CLK), .Q(g1400) ) ;
INV     gate1657  (.A(II30101), .Z(g23216) ) ;
DFF     gate1658  (.D(g23216), .CP(CLK), .Q(g1401) ) ;
INV     gate1659  (.A(II30104), .Z(g23217) ) ;
DFF     gate1660  (.D(g23217), .CP(CLK), .Q(g1399) ) ;
INV     gate1661  (.A(II30107), .Z(g23218) ) ;
DFF     gate1662  (.D(g23218), .CP(CLK), .Q(g1403) ) ;
INV     gate1663  (.A(II30110), .Z(g23219) ) ;
DFF     gate1664  (.D(g23219), .CP(CLK), .Q(g1404) ) ;
INV     gate1665  (.A(II30113), .Z(g23220) ) ;
DFF     gate1666  (.D(g23220), .CP(CLK), .Q(g1402) ) ;
INV     gate1667  (.A(II30116), .Z(g23221) ) ;
DFF     gate1668  (.D(g23221), .CP(CLK), .Q(g1406) ) ;
INV     gate1669  (.A(II30119), .Z(g23222) ) ;
DFF     gate1670  (.D(g23222), .CP(CLK), .Q(g1407) ) ;
INV     gate1671  (.A(II30122), .Z(g23223) ) ;
DFF     gate1672  (.D(g23223), .CP(CLK), .Q(g1405) ) ;
INV     gate1673  (.A(II30125), .Z(g23224) ) ;
DFF     gate1674  (.D(g23224), .CP(CLK), .Q(g1409) ) ;
INV     gate1675  (.A(II30128), .Z(g23225) ) ;
DFF     gate1676  (.D(g23225), .CP(CLK), .Q(g1410) ) ;
INV     gate1677  (.A(II30131), .Z(g23226) ) ;
DFF     gate1678  (.D(g23226), .CP(CLK), .Q(g1408) ) ;
INV     gate1679  (.A(II30134), .Z(g23227) ) ;
DFF     gate1680  (.D(g23227), .CP(CLK), .Q(g1412) ) ;
INV     gate1681  (.A(II30137), .Z(g23228) ) ;
DFF     gate1682  (.D(g23228), .CP(CLK), .Q(g1413) ) ;
INV     gate1683  (.A(II30140), .Z(g23229) ) ;
DFF     gate1684  (.D(g23229), .CP(CLK), .Q(g1411) ) ;
INV     gate1685  (.A(II30143), .Z(g23230) ) ;
DFF     gate1686  (.D(g23230), .CP(CLK), .Q(g1415) ) ;
INV     gate1687  (.A(II30146), .Z(g23231) ) ;
DFF     gate1688  (.D(g23231), .CP(CLK), .Q(g1416) ) ;
INV     gate1689  (.A(II30149), .Z(g23232) ) ;
DFF     gate1690  (.D(g23232), .CP(CLK), .Q(g1414) ) ;
INV     gate1691  (.A(II30152), .Z(g23233) ) ;
DFF     gate1692  (.D(g23233), .CP(CLK), .Q(g1418) ) ;
INV     gate1693  (.A(II30155), .Z(g23234) ) ;
DFF     gate1694  (.D(g23234), .CP(CLK), .Q(g1419) ) ;
INV     gate1695  (.A(II30158), .Z(g23235) ) ;
DFF     gate1696  (.D(g23235), .CP(CLK), .Q(g1417) ) ;
INV     gate1697  (.A(II34734), .Z(g26709) ) ;
DFF     gate1698  (.D(g26709), .CP(CLK), .Q(g1421) ) ;
INV     gate1699  (.A(II34737), .Z(g26710) ) ;
DFF     gate1700  (.D(g26710), .CP(CLK), .Q(g1422) ) ;
INV     gate1701  (.A(II34740), .Z(g26711) ) ;
DFF     gate1702  (.D(g26711), .CP(CLK), .Q(g1420) ) ;
INV     gate1703  (.A(II31688), .Z(g24338) ) ;
DFF     gate1704  (.D(g24338), .CP(CLK), .Q(g1424) ) ;
INV     gate1705  (.A(II31691), .Z(g24339) ) ;
DFF     gate1706  (.D(g24339), .CP(CLK), .Q(g1425) ) ;
INV     gate1707  (.A(II31694), .Z(g24340) ) ;
DFF     gate1708  (.D(g24340), .CP(CLK), .Q(g1423) ) ;
INV     gate1709  (.A(II20610), .Z(g13437) ) ;
DFF     gate1710  (.D(g13437), .CP(CLK), .Q(g1520) ) ;
DFF     gate1711  (.D(g1520), .CP(CLK), .Q(g1517) ) ;
DFF     gate1712  (.D(g1517), .CP(CLK), .Q(g1547) ) ;
INV     gate1713  (.A(II31697), .Z(g24341) ) ;
DFF     gate1714  (.D(g24341), .CP(CLK), .Q(g1512) ) ;
INV     gate1715  (.A(II31700), .Z(g24342) ) ;
DFF     gate1716  (.D(g24342), .CP(CLK), .Q(g1513) ) ;
INV     gate1717  (.A(II31703), .Z(g24343) ) ;
DFF     gate1718  (.D(g24343), .CP(CLK), .Q(g1511) ) ;
INV     gate1719  (.A(II31706), .Z(g24344) ) ;
DFF     gate1720  (.D(g24344), .CP(CLK), .Q(g1515) ) ;
INV     gate1721  (.A(II31709), .Z(g24345) ) ;
DFF     gate1722  (.D(g24345), .CP(CLK), .Q(g1516) ) ;
INV     gate1723  (.A(II31712), .Z(g24346) ) ;
DFF     gate1724  (.D(g24346), .CP(CLK), .Q(g1514) ) ;
INV     gate1725  (.A(II31715), .Z(g24347) ) ;
DFF     gate1726  (.D(g24347), .CP(CLK), .Q(g1524) ) ;
INV     gate1727  (.A(II31718), .Z(g24348) ) ;
DFF     gate1728  (.D(g24348), .CP(CLK), .Q(g1525) ) ;
INV     gate1729  (.A(II31721), .Z(g24349) ) ;
DFF     gate1730  (.D(g24349), .CP(CLK), .Q(g1523) ) ;
INV     gate1731  (.A(II31724), .Z(g24350) ) ;
DFF     gate1732  (.D(g24350), .CP(CLK), .Q(g1527) ) ;
INV     gate1733  (.A(II31727), .Z(g24351) ) ;
DFF     gate1734  (.D(g24351), .CP(CLK), .Q(g1528) ) ;
INV     gate1735  (.A(II31730), .Z(g24352) ) ;
DFF     gate1736  (.D(g24352), .CP(CLK), .Q(g1526) ) ;
INV     gate1737  (.A(II31733), .Z(g24353) ) ;
DFF     gate1738  (.D(g24353), .CP(CLK), .Q(g1530) ) ;
INV     gate1739  (.A(II31736), .Z(g24354) ) ;
DFF     gate1740  (.D(g24354), .CP(CLK), .Q(g1531) ) ;
INV     gate1741  (.A(II31739), .Z(g24355) ) ;
DFF     gate1742  (.D(g24355), .CP(CLK), .Q(g1529) ) ;
INV     gate1743  (.A(II31742), .Z(g24356) ) ;
DFF     gate1744  (.D(g24356), .CP(CLK), .Q(g1533) ) ;
INV     gate1745  (.A(II31745), .Z(g24357) ) ;
DFF     gate1746  (.D(g24357), .CP(CLK), .Q(g1534) ) ;
INV     gate1747  (.A(II31748), .Z(g24358) ) ;
DFF     gate1748  (.D(g24358), .CP(CLK), .Q(g1532) ) ;
INV     gate1749  (.A(II31751), .Z(g24359) ) ;
DFF     gate1750  (.D(g24359), .CP(CLK), .Q(g1536) ) ;
INV     gate1751  (.A(II31754), .Z(g24360) ) ;
DFF     gate1752  (.D(g24360), .CP(CLK), .Q(g1537) ) ;
INV     gate1753  (.A(II31757), .Z(g24361) ) ;
DFF     gate1754  (.D(g24361), .CP(CLK), .Q(g1535) ) ;
INV     gate1755  (.A(II31760), .Z(g24362) ) ;
DFF     gate1756  (.D(g24362), .CP(CLK), .Q(g1539) ) ;
INV     gate1757  (.A(II31763), .Z(g24363) ) ;
DFF     gate1758  (.D(g24363), .CP(CLK), .Q(g1540) ) ;
INV     gate1759  (.A(II31766), .Z(g24364) ) ;
DFF     gate1760  (.D(g24364), .CP(CLK), .Q(g1538) ) ;
INV     gate1761  (.A(II31769), .Z(g24365) ) ;
DFF     gate1762  (.D(g24365), .CP(CLK), .Q(g1542) ) ;
INV     gate1763  (.A(II31772), .Z(g24366) ) ;
DFF     gate1764  (.D(g24366), .CP(CLK), .Q(g1543) ) ;
INV     gate1765  (.A(II31775), .Z(g24367) ) ;
DFF     gate1766  (.D(g24367), .CP(CLK), .Q(g1541) ) ;
INV     gate1767  (.A(II31778), .Z(g24368) ) ;
DFF     gate1768  (.D(g24368), .CP(CLK), .Q(g1545) ) ;
INV     gate1769  (.A(II31781), .Z(g24369) ) ;
DFF     gate1770  (.D(g24369), .CP(CLK), .Q(g1546) ) ;
INV     gate1771  (.A(II31784), .Z(g24370) ) ;
DFF     gate1772  (.D(g24370), .CP(CLK), .Q(g1544) ) ;
INV     gate1773  (.A(II34746), .Z(g26713) ) ;
DFF     gate1774  (.D(g26713), .CP(CLK), .Q(g1551) ) ;
INV     gate1775  (.A(II34749), .Z(g26714) ) ;
DFF     gate1776  (.D(g26714), .CP(CLK), .Q(g1552) ) ;
INV     gate1777  (.A(II34752), .Z(g26715) ) ;
DFF     gate1778  (.D(g26715), .CP(CLK), .Q(g1550) ) ;
INV     gate1779  (.A(II34755), .Z(g26716) ) ;
DFF     gate1780  (.D(g26716), .CP(CLK), .Q(g1554) ) ;
INV     gate1781  (.A(II34758), .Z(g26717) ) ;
DFF     gate1782  (.D(g26717), .CP(CLK), .Q(g1555) ) ;
INV     gate1783  (.A(II34761), .Z(g26718) ) ;
DFF     gate1784  (.D(g26718), .CP(CLK), .Q(g1553) ) ;
INV     gate1785  (.A(II34764), .Z(g26719) ) ;
DFF     gate1786  (.D(g26719), .CP(CLK), .Q(g1557) ) ;
INV     gate1787  (.A(II34767), .Z(g26720) ) ;
DFF     gate1788  (.D(g26720), .CP(CLK), .Q(g1558) ) ;
INV     gate1789  (.A(II34770), .Z(g26721) ) ;
DFF     gate1790  (.D(g26721), .CP(CLK), .Q(g1556) ) ;
INV     gate1791  (.A(II34773), .Z(g26722) ) ;
DFF     gate1792  (.D(g26722), .CP(CLK), .Q(g1560) ) ;
INV     gate1793  (.A(II34776), .Z(g26723) ) ;
DFF     gate1794  (.D(g26723), .CP(CLK), .Q(g1561) ) ;
INV     gate1795  (.A(II34779), .Z(g26724) ) ;
DFF     gate1796  (.D(g26724), .CP(CLK), .Q(g1559) ) ;
INV     gate1797  (.A(II40188), .Z(g30536) ) ;
DFF     gate1798  (.D(g30536), .CP(CLK), .Q(g1567) ) ;
INV     gate1799  (.A(II40191), .Z(g30537) ) ;
DFF     gate1800  (.D(g30537), .CP(CLK), .Q(g1570) ) ;
INV     gate1801  (.A(II40194), .Z(g30538) ) ;
DFF     gate1802  (.D(g30538), .CP(CLK), .Q(g1573) ) ;
INV     gate1803  (.A(II40886), .Z(g30878) ) ;
DFF     gate1804  (.D(g30878), .CP(CLK), .Q(g1612) ) ;
INV     gate1805  (.A(II40889), .Z(g30879) ) ;
DFF     gate1806  (.D(g30879), .CP(CLK), .Q(g1615) ) ;
INV     gate1807  (.A(II40892), .Z(g30880) ) ;
DFF     gate1808  (.D(g30880), .CP(CLK), .Q(g1618) ) ;
INV     gate1809  (.A(II40868), .Z(g30872) ) ;
DFF     gate1810  (.D(g30872), .CP(CLK), .Q(g1576) ) ;
INV     gate1811  (.A(II40871), .Z(g30873) ) ;
DFF     gate1812  (.D(g30873), .CP(CLK), .Q(g1579) ) ;
INV     gate1813  (.A(II40874), .Z(g30874) ) ;
DFF     gate1814  (.D(g30874), .CP(CLK), .Q(g1582) ) ;
INV     gate1815  (.A(II40895), .Z(g30881) ) ;
DFF     gate1816  (.D(g30881), .CP(CLK), .Q(g1621) ) ;
INV     gate1817  (.A(II40898), .Z(g30882) ) ;
DFF     gate1818  (.D(g30882), .CP(CLK), .Q(g1624) ) ;
INV     gate1819  (.A(II40901), .Z(g30883) ) ;
DFF     gate1820  (.D(g30883), .CP(CLK), .Q(g1627) ) ;
INV     gate1821  (.A(II40197), .Z(g30539) ) ;
DFF     gate1822  (.D(g30539), .CP(CLK), .Q(g1585) ) ;
INV     gate1823  (.A(II40200), .Z(g30540) ) ;
DFF     gate1824  (.D(g30540), .CP(CLK), .Q(g1588) ) ;
INV     gate1825  (.A(II40203), .Z(g30541) ) ;
DFF     gate1826  (.D(g30541), .CP(CLK), .Q(g1591) ) ;
INV     gate1827  (.A(II40215), .Z(g30545) ) ;
DFF     gate1828  (.D(g30545), .CP(CLK), .Q(g1630) ) ;
INV     gate1829  (.A(II40218), .Z(g30546) ) ;
DFF     gate1830  (.D(g30546), .CP(CLK), .Q(g1633) ) ;
INV     gate1831  (.A(II40221), .Z(g30547) ) ;
DFF     gate1832  (.D(g30547), .CP(CLK), .Q(g1636) ) ;
INV     gate1833  (.A(II40206), .Z(g30542) ) ;
DFF     gate1834  (.D(g30542), .CP(CLK), .Q(g1594) ) ;
INV     gate1835  (.A(II40209), .Z(g30543) ) ;
DFF     gate1836  (.D(g30543), .CP(CLK), .Q(g1597) ) ;
INV     gate1837  (.A(II40212), .Z(g30544) ) ;
DFF     gate1838  (.D(g30544), .CP(CLK), .Q(g1600) ) ;
INV     gate1839  (.A(II40224), .Z(g30548) ) ;
DFF     gate1840  (.D(g30548), .CP(CLK), .Q(g1639) ) ;
INV     gate1841  (.A(II40227), .Z(g30549) ) ;
DFF     gate1842  (.D(g30549), .CP(CLK), .Q(g1642) ) ;
INV     gate1843  (.A(II40230), .Z(g30550) ) ;
DFF     gate1844  (.D(g30550), .CP(CLK), .Q(g1645) ) ;
INV     gate1845  (.A(II40877), .Z(g30875) ) ;
DFF     gate1846  (.D(g30875), .CP(CLK), .Q(g1603) ) ;
INV     gate1847  (.A(II40880), .Z(g30876) ) ;
DFF     gate1848  (.D(g30876), .CP(CLK), .Q(g1606) ) ;
INV     gate1849  (.A(II40883), .Z(g30877) ) ;
DFF     gate1850  (.D(g30877), .CP(CLK), .Q(g1609) ) ;
INV     gate1851  (.A(II40904), .Z(g30884) ) ;
DFF     gate1852  (.D(g30884), .CP(CLK), .Q(g1648) ) ;
INV     gate1853  (.A(II40907), .Z(g30885) ) ;
DFF     gate1854  (.D(g30885), .CP(CLK), .Q(g1651) ) ;
INV     gate1855  (.A(II40910), .Z(g30886) ) ;
DFF     gate1856  (.D(g30886), .CP(CLK), .Q(g1654) ) ;
INV     gate1857  (.A(II33855), .Z(g26001) ) ;
DFF     gate1858  (.D(g26001), .CP(CLK), .Q(g1466) ) ;
INV     gate1859  (.A(II34743), .Z(g26712) ) ;
DFF     gate1860  (.D(g26712), .CP(CLK), .Q(g1462) ) ;
INV     gate1861  (.A(II35494), .Z(g27219) ) ;
DFF     gate1862  (.D(g27219), .CP(CLK), .Q(g1457) ) ;
INV     gate1863  (.A(II36108), .Z(g27699) ) ;
DFF     gate1864  (.D(g27699), .CP(CLK), .Q(g1453) ) ;
INV     gate1865  (.A(II37023), .Z(g28258) ) ;
DFF     gate1866  (.D(g28258), .CP(CLK), .Q(g1448) ) ;
INV     gate1867  (.A(II37596), .Z(g28683) ) ;
DFF     gate1868  (.D(g28683), .CP(CLK), .Q(g1444) ) ;
INV     gate1869  (.A(II38184), .Z(g29147) ) ;
DFF     gate1870  (.D(g29147), .CP(CLK), .Q(g1439) ) ;
INV     gate1871  (.A(II38662), .Z(g29427) ) ;
DFF     gate1872  (.D(g29427), .CP(CLK), .Q(g1435) ) ;
INV     gate1873  (.A(II39041), .Z(g29641) ) ;
DFF     gate1874  (.D(g29641), .CP(CLK), .Q(g1430) ) ;
INV     gate1875  (.A(II39258), .Z(g29802) ) ;
DFF     gate1876  (.D(g29802), .CP(CLK), .Q(g1426) ) ;
INV     gate1877  (.A(II27014), .Z(g20563) ) ;
DFF     gate1878  (.D(g20563), .CP(CLK), .Q(g1562) ) ;
DFF     gate1879  (.D(g1562), .CP(CLK), .Q(g1564) ) ;
DFF     gate1880  (.D(g1564), .CP(CLK), .Q(g1563) ) ;
INV     gate1881  (.A(II20613), .Z(g13438) ) ;
DFF     gate1882  (.D(g13438), .CP(CLK), .Q(g1657) ) ;
DFF     gate1883  (.D(g1657), .CP(CLK), .Q(g1786) ) ;
DFF     gate1884  (.D(g1786), .CP(CLK), .Q(g1782) ) ;
INV     gate1885  (.A(II18626), .Z(g11550) ) ;
DFF     gate1886  (.D(g11550), .CP(CLK), .Q(g1690) ) ;
INV     gate1887  (.A(II37026), .Z(g28259) ) ;
DFF     gate1888  (.D(g28259), .CP(CLK), .Q(g1735) ) ;
INV     gate1889  (.A(II37029), .Z(g28260) ) ;
DFF     gate1890  (.D(g28260), .CP(CLK), .Q(g1724) ) ;
INV     gate1891  (.A(II37032), .Z(g28261) ) ;
DFF     gate1892  (.D(g28261), .CP(CLK), .Q(g1727) ) ;
INV     gate1893  (.A(II37035), .Z(g28262) ) ;
DFF     gate1894  (.D(g28262), .CP(CLK), .Q(g1750) ) ;
INV     gate1895  (.A(II37038), .Z(g28263) ) ;
DFF     gate1896  (.D(g28263), .CP(CLK), .Q(g1739) ) ;
INV     gate1897  (.A(II37041), .Z(g28264) ) ;
DFF     gate1898  (.D(g28264), .CP(CLK), .Q(g1742) ) ;
INV     gate1899  (.A(II37044), .Z(g28265) ) ;
DFF     gate1900  (.D(g28265), .CP(CLK), .Q(g1765) ) ;
INV     gate1901  (.A(II37047), .Z(g28266) ) ;
DFF     gate1902  (.D(g28266), .CP(CLK), .Q(g1754) ) ;
INV     gate1903  (.A(II37050), .Z(g28267) ) ;
DFF     gate1904  (.D(g28267), .CP(CLK), .Q(g1757) ) ;
INV     gate1905  (.A(II37053), .Z(g28268) ) ;
DFF     gate1906  (.D(g28268), .CP(CLK), .Q(g1779) ) ;
INV     gate1907  (.A(II37056), .Z(g28269) ) ;
DFF     gate1908  (.D(g28269), .CP(CLK), .Q(g1769) ) ;
INV     gate1909  (.A(II37059), .Z(g28270) ) ;
DFF     gate1910  (.D(g28270), .CP(CLK), .Q(g1772) ) ;
INV     gate1911  (.A(II38683), .Z(g29434) ) ;
DFF     gate1912  (.D(g29434), .CP(CLK), .Q(g1789) ) ;
INV     gate1913  (.A(II38686), .Z(g29435) ) ;
DFF     gate1914  (.D(g29435), .CP(CLK), .Q(g1792) ) ;
INV     gate1915  (.A(II38689), .Z(g29436) ) ;
DFF     gate1916  (.D(g29436), .CP(CLK), .Q(g1795) ) ;
INV     gate1917  (.A(II39053), .Z(g29645) ) ;
DFF     gate1918  (.D(g29645), .CP(CLK), .Q(g1798) ) ;
INV     gate1919  (.A(II39056), .Z(g29646) ) ;
DFF     gate1920  (.D(g29646), .CP(CLK), .Q(g1801) ) ;
INV     gate1921  (.A(II39059), .Z(g29647) ) ;
DFF     gate1922  (.D(g29647), .CP(CLK), .Q(g1804) ) ;
INV     gate1923  (.A(II38692), .Z(g29437) ) ;
DFF     gate1924  (.D(g29437), .CP(CLK), .Q(g1808) ) ;
INV     gate1925  (.A(II38695), .Z(g29438) ) ;
DFF     gate1926  (.D(g29438), .CP(CLK), .Q(g1809) ) ;
INV     gate1927  (.A(II38698), .Z(g29439) ) ;
DFF     gate1928  (.D(g29439), .CP(CLK), .Q(g1807) ) ;
INV     gate1929  (.A(II36111), .Z(g27700) ) ;
DFF     gate1930  (.D(g27700), .CP(CLK), .Q(g1810) ) ;
INV     gate1931  (.A(II36114), .Z(g27701) ) ;
DFF     gate1932  (.D(g27701), .CP(CLK), .Q(g1813) ) ;
INV     gate1933  (.A(II36117), .Z(g27702) ) ;
DFF     gate1934  (.D(g27702), .CP(CLK), .Q(g1816) ) ;
INV     gate1935  (.A(II36120), .Z(g27703) ) ;
DFF     gate1936  (.D(g27703), .CP(CLK), .Q(g1819) ) ;
INV     gate1937  (.A(II36123), .Z(g27704) ) ;
DFF     gate1938  (.D(g27704), .CP(CLK), .Q(g1822) ) ;
INV     gate1939  (.A(II36126), .Z(g27705) ) ;
DFF     gate1940  (.D(g27705), .CP(CLK), .Q(g1825) ) ;
INV     gate1941  (.A(II37599), .Z(g28684) ) ;
DFF     gate1942  (.D(g28684), .CP(CLK), .Q(g1829) ) ;
INV     gate1943  (.A(II37602), .Z(g28685) ) ;
DFF     gate1944  (.D(g28685), .CP(CLK), .Q(g1830) ) ;
INV     gate1945  (.A(II37605), .Z(g28686) ) ;
DFF     gate1946  (.D(g28686), .CP(CLK), .Q(g1828) ) ;
INV     gate1947  (.A(II39261), .Z(g29803) ) ;
DFF     gate1948  (.D(g29803), .CP(CLK), .Q(g1693) ) ;
INV     gate1949  (.A(II39264), .Z(g29804) ) ;
DFF     gate1950  (.D(g29804), .CP(CLK), .Q(g1694) ) ;
INV     gate1951  (.A(II39267), .Z(g29805) ) ;
DFF     gate1952  (.D(g29805), .CP(CLK), .Q(g1695) ) ;
INV     gate1953  (.A(II40913), .Z(g30887) ) ;
DFF     gate1954  (.D(g30887), .CP(CLK), .Q(g1696) ) ;
INV     gate1955  (.A(II40916), .Z(g30888) ) ;
DFF     gate1956  (.D(g30888), .CP(CLK), .Q(g1697) ) ;
INV     gate1957  (.A(II40919), .Z(g30889) ) ;
DFF     gate1958  (.D(g30889), .CP(CLK), .Q(g1698) ) ;
INV     gate1959  (.A(II40438), .Z(g30716) ) ;
DFF     gate1960  (.D(g30716), .CP(CLK), .Q(g1699) ) ;
INV     gate1961  (.A(II40441), .Z(g30717) ) ;
DFF     gate1962  (.D(g30717), .CP(CLK), .Q(g1700) ) ;
INV     gate1963  (.A(II40444), .Z(g30718) ) ;
DFF     gate1964  (.D(g30718), .CP(CLK), .Q(g1701) ) ;
INV     gate1965  (.A(II39044), .Z(g29642) ) ;
DFF     gate1966  (.D(g29642), .CP(CLK), .Q(g1703) ) ;
INV     gate1967  (.A(II39047), .Z(g29643) ) ;
DFF     gate1968  (.D(g29643), .CP(CLK), .Q(g1704) ) ;
INV     gate1969  (.A(II39050), .Z(g29644) ) ;
DFF     gate1970  (.D(g29644), .CP(CLK), .Q(g1702) ) ;
INV     gate1971  (.A(II35500), .Z(g27221) ) ;
DFF     gate1972  (.D(g27221), .CP(CLK), .Q(g1784) ) ;
INV     gate1973  (.A(II35503), .Z(g27222) ) ;
DFF     gate1974  (.D(g27222), .CP(CLK), .Q(g1785) ) ;
INV     gate1975  (.A(II35506), .Z(g27223) ) ;
DFF     gate1976  (.D(g27223), .CP(CLK), .Q(g1783) ) ;
INV     gate1977  (.A(II18665), .Z(g11563) ) ;
DFF     gate1978  (.D(g11563), .CP(CLK), .Q(g1831) ) ;
DFF     gate1979  (.D(g1831), .CP(CLK), .Q(g1832) ) ;
INV     gate1980  (.A(II18668), .Z(g11564) ) ;
DFF     gate1981  (.D(g11564), .CP(CLK), .Q(g1833) ) ;
DFF     gate1982  (.D(g1833), .CP(CLK), .Q(g1834) ) ;
INV     gate1983  (.A(II18671), .Z(g11565) ) ;
DFF     gate1984  (.D(g11565), .CP(CLK), .Q(g1835) ) ;
DFF     gate1985  (.D(g1835), .CP(CLK), .Q(g1660) ) ;
INV     gate1986  (.A(II18611), .Z(g11545) ) ;
DFF     gate1987  (.D(g11545), .CP(CLK), .Q(g1661) ) ;
DFF     gate1988  (.D(g1661), .CP(CLK), .Q(g1662) ) ;
INV     gate1989  (.A(II18614), .Z(g11546) ) ;
DFF     gate1990  (.D(g11546), .CP(CLK), .Q(g1663) ) ;
DFF     gate1991  (.D(g1663), .CP(CLK), .Q(g1664) ) ;
INV     gate1992  (.A(II18617), .Z(g11547) ) ;
DFF     gate1993  (.D(g11547), .CP(CLK), .Q(g1665) ) ;
DFF     gate1994  (.D(g1665), .CP(CLK), .Q(g1666) ) ;
INV     gate1995  (.A(II18620), .Z(g11548) ) ;
DFF     gate1996  (.D(g11548), .CP(CLK), .Q(g1667) ) ;
DFF     gate1997  (.D(g1667), .CP(CLK), .Q(g1668) ) ;
INV     gate1998  (.A(II18623), .Z(g11549) ) ;
DFF     gate1999  (.D(g11549), .CP(CLK), .Q(g1669) ) ;
DFF     gate2000  (.D(g1669), .CP(CLK), .Q(g1670) ) ;
INV     gate2001  (.A(II20616), .Z(g13439) ) ;
DFF     gate2002  (.D(g13439), .CP(CLK), .Q(g1671) ) ;
DFF     gate2003  (.D(g1671), .CP(CLK), .Q(g1672) ) ;
INV     gate2004  (.A(II25171), .Z(g19036) ) ;
DFF     gate2005  (.D(g19036), .CP(CLK), .Q(g1680) ) ;
INV     gate2006  (.A(II38665), .Z(g29428) ) ;
DFF     gate2007  (.D(g29428), .CP(CLK), .Q(g1686) ) ;
INV     gate2008  (.A(II38668), .Z(g29429) ) ;
DFF     gate2009  (.D(g29429), .CP(CLK), .Q(g1689) ) ;
INV     gate2010  (.A(II38671), .Z(g29430) ) ;
DFF     gate2011  (.D(g29430), .CP(CLK), .Q(g1678) ) ;
INV     gate2012  (.A(II38674), .Z(g29431) ) ;
DFF     gate2013  (.D(g29431), .CP(CLK), .Q(g1677) ) ;
INV     gate2014  (.A(II38677), .Z(g29432) ) ;
DFF     gate2015  (.D(g29432), .CP(CLK), .Q(g1676) ) ;
INV     gate2016  (.A(II38680), .Z(g29433) ) ;
DFF     gate2017  (.D(g29433), .CP(CLK), .Q(g1675) ) ;
INV     gate2018  (.A(II25183), .Z(g19040) ) ;
DFF     gate2019  (.D(g19040), .CP(CLK), .Q(g1685) ) ;
INV     gate2020  (.A(II25180), .Z(g19039) ) ;
DFF     gate2021  (.D(g19039), .CP(CLK), .Q(g1684) ) ;
INV     gate2022  (.A(II25177), .Z(g19038) ) ;
DFF     gate2023  (.D(g19038), .CP(CLK), .Q(g1683) ) ;
INV     gate2024  (.A(II25174), .Z(g19037) ) ;
DFF     gate2025  (.D(g19037), .CP(CLK), .Q(g1682) ) ;
INV     gate2026  (.A(II32934), .Z(g25152) ) ;
DFF     gate2027  (.D(g25152), .CP(CLK), .Q(g1681) ) ;
INV     gate2028  (.A(II35497), .Z(g27220) ) ;
DFF     gate2029  (.D(g27220), .CP(CLK), .Q(g1679) ) ;
INV     gate2030  (.A(II18629), .Z(g11551) ) ;
DFF     gate2031  (.D(g11551), .CP(CLK), .Q(g1723) ) ;
DFF     gate2032  (.D(g1723), .CP(CLK), .Q(g1730) ) ;
INV     gate2033  (.A(II18632), .Z(g11552) ) ;
DFF     gate2034  (.D(g11552), .CP(CLK), .Q(g1731) ) ;
DFF     gate2035  (.D(g1731), .CP(CLK), .Q(g1732) ) ;
INV     gate2036  (.A(II18635), .Z(g11553) ) ;
DFF     gate2037  (.D(g11553), .CP(CLK), .Q(g1733) ) ;
DFF     gate2038  (.D(g1733), .CP(CLK), .Q(g1734) ) ;
INV     gate2039  (.A(II18638), .Z(g11554) ) ;
DFF     gate2040  (.D(g11554), .CP(CLK), .Q(g1738) ) ;
DFF     gate2041  (.D(g1738), .CP(CLK), .Q(g1745) ) ;
INV     gate2042  (.A(II18641), .Z(g11555) ) ;
DFF     gate2043  (.D(g11555), .CP(CLK), .Q(g1746) ) ;
DFF     gate2044  (.D(g1746), .CP(CLK), .Q(g1747) ) ;
INV     gate2045  (.A(II18644), .Z(g11556) ) ;
DFF     gate2046  (.D(g11556), .CP(CLK), .Q(g1748) ) ;
DFF     gate2047  (.D(g1748), .CP(CLK), .Q(g1749) ) ;
INV     gate2048  (.A(II18647), .Z(g11557) ) ;
DFF     gate2049  (.D(g11557), .CP(CLK), .Q(g1753) ) ;
DFF     gate2050  (.D(g1753), .CP(CLK), .Q(g1760) ) ;
INV     gate2051  (.A(II18650), .Z(g11558) ) ;
DFF     gate2052  (.D(g11558), .CP(CLK), .Q(g1761) ) ;
DFF     gate2053  (.D(g1761), .CP(CLK), .Q(g1762) ) ;
INV     gate2054  (.A(II18653), .Z(g11559) ) ;
DFF     gate2055  (.D(g11559), .CP(CLK), .Q(g1763) ) ;
DFF     gate2056  (.D(g1763), .CP(CLK), .Q(g1764) ) ;
INV     gate2057  (.A(II18656), .Z(g11560) ) ;
DFF     gate2058  (.D(g11560), .CP(CLK), .Q(g1768) ) ;
DFF     gate2059  (.D(g1768), .CP(CLK), .Q(g1775) ) ;
INV     gate2060  (.A(II18659), .Z(g11561) ) ;
DFF     gate2061  (.D(g11561), .CP(CLK), .Q(g1776) ) ;
DFF     gate2062  (.D(g1776), .CP(CLK), .Q(g1777) ) ;
INV     gate2063  (.A(II18662), .Z(g11562) ) ;
DFF     gate2064  (.D(g11562), .CP(CLK), .Q(g1778) ) ;
DFF     gate2065  (.D(g1778), .CP(CLK), .Q(g1705) ) ;
INV     gate2066  (.A(II20619), .Z(g13440) ) ;
DFF     gate2067  (.D(g13440), .CP(CLK), .Q(g1706) ) ;
DFF     gate2068  (.D(g1706), .CP(CLK), .Q(g1712) ) ;
DFF     gate2069  (.D(g1712), .CP(CLK), .Q(g1718) ) ;
INV     gate2070  (.A(II20652), .Z(g13451) ) ;
DFF     gate2071  (.D(g13451), .CP(CLK), .Q(g1925) ) ;
DFF     gate2072  (.D(g1925), .CP(CLK), .Q(g1931) ) ;
DFF     gate2073  (.D(g1931), .CP(CLK), .Q(g1930) ) ;
INV     gate2074  (.A(II30161), .Z(g23236) ) ;
DFF     gate2075  (.D(g23236), .CP(CLK), .Q(g1934) ) ;
INV     gate2076  (.A(II27017), .Z(g20564) ) ;
DFF     gate2077  (.D(g20564), .CP(CLK), .Q(g1937) ) ;
INV     gate2078  (.A(II27020), .Z(g20565) ) ;
DFF     gate2079  (.D(g20565), .CP(CLK), .Q(g1890) ) ;
INV     gate2080  (.A(II22515), .Z(g16471) ) ;
DFF     gate2081  (.D(g16471), .CP(CLK), .Q(g1893) ) ;
DFF     gate2082  (.D(g1893), .CP(CLK), .Q(g1903) ) ;
DFF     gate2083  (.D(g1903), .CP(CLK), .Q(g1904) ) ;
INV     gate2084  (.A(II18674), .Z(g11566) ) ;
DFF     gate2085  (.D(g11566), .CP(CLK), .Q(g1944) ) ;
DFF     gate2086  (.D(g1944), .CP(CLK), .Q(g1949) ) ;
INV     gate2087  (.A(II18683), .Z(g11569) ) ;
DFF     gate2088  (.D(g11569), .CP(CLK), .Q(g1950) ) ;
DFF     gate2089  (.D(g1950), .CP(CLK), .Q(g1951) ) ;
INV     gate2090  (.A(II18686), .Z(g11570) ) ;
DFF     gate2091  (.D(g11570), .CP(CLK), .Q(g1952) ) ;
DFF     gate2092  (.D(g1952), .CP(CLK), .Q(g1953) ) ;
INV     gate2093  (.A(II18689), .Z(g11571) ) ;
DFF     gate2094  (.D(g11571), .CP(CLK), .Q(g1954) ) ;
DFF     gate2095  (.D(g1954), .CP(CLK), .Q(g1945) ) ;
INV     gate2096  (.A(II18677), .Z(g11567) ) ;
DFF     gate2097  (.D(g11567), .CP(CLK), .Q(g1946) ) ;
DFF     gate2098  (.D(g1946), .CP(CLK), .Q(g1947) ) ;
INV     gate2099  (.A(II18680), .Z(g11568) ) ;
DFF     gate2100  (.D(g11568), .CP(CLK), .Q(g1948) ) ;
DFF     gate2101  (.D(g1948), .CP(CLK), .Q(g1870) ) ;
INV     gate2102  (.A(II20622), .Z(g13441) ) ;
DFF     gate2103  (.D(g13441), .CP(CLK), .Q(g1855) ) ;
DFF     gate2104  (.D(g1855), .CP(CLK), .Q(g1862) ) ;
DFF     gate2105  (.D(g1862), .CP(CLK), .Q(g1866) ) ;
INV     gate2106  (.A(II31796), .Z(g24374) ) ;
DFF     gate2107  (.D(g24374), .CP(CLK), .Q(g1867) ) ;
INV     gate2108  (.A(II31799), .Z(g24375) ) ;
DFF     gate2109  (.D(g24375), .CP(CLK), .Q(g1868) ) ;
INV     gate2110  (.A(II31802), .Z(g24376) ) ;
DFF     gate2111  (.D(g24376), .CP(CLK), .Q(g1869) ) ;
INV     gate2112  (.A(II32961), .Z(g25161) ) ;
DFF     gate2113  (.D(g25161), .CP(CLK), .Q(g1836) ) ;
INV     gate2114  (.A(II32937), .Z(g25153) ) ;
DFF     gate2115  (.D(g25153), .CP(CLK), .Q(g1839) ) ;
INV     gate2116  (.A(II32940), .Z(g25154) ) ;
DFF     gate2117  (.D(g25154), .CP(CLK), .Q(g1842) ) ;
INV     gate2118  (.A(II32952), .Z(g25158) ) ;
DFF     gate2119  (.D(g25158), .CP(CLK), .Q(g1858) ) ;
INV     gate2120  (.A(II32955), .Z(g25159) ) ;
DFF     gate2121  (.D(g25159), .CP(CLK), .Q(g1859) ) ;
INV     gate2122  (.A(II32958), .Z(g25160) ) ;
DFF     gate2123  (.D(g25160), .CP(CLK), .Q(g1860) ) ;
INV     gate2124  (.A(II31787), .Z(g24371) ) ;
DFF     gate2125  (.D(g24371), .CP(CLK), .Q(g1861) ) ;
INV     gate2126  (.A(II31790), .Z(g24372) ) ;
DFF     gate2127  (.D(g24372), .CP(CLK), .Q(g1865) ) ;
INV     gate2128  (.A(II31793), .Z(g24373) ) ;
DFF     gate2129  (.D(g24373), .CP(CLK), .Q(g1845) ) ;
INV     gate2130  (.A(II32943), .Z(g25155) ) ;
DFF     gate2131  (.D(g25155), .CP(CLK), .Q(g1846) ) ;
INV     gate2132  (.A(II32946), .Z(g25156) ) ;
DFF     gate2133  (.D(g25156), .CP(CLK), .Q(g1849) ) ;
INV     gate2134  (.A(II32949), .Z(g25157) ) ;
DFF     gate2135  (.D(g25157), .CP(CLK), .Q(g1852) ) ;
INV     gate2136  (.A(II22518), .Z(g16472) ) ;
DFF     gate2137  (.D(g16472), .CP(CLK), .Q(g1908) ) ;
DFF     gate2138  (.D(g1908), .CP(CLK), .Q(g1915) ) ;
DFF     gate2139  (.D(g1915), .CP(CLK), .Q(g1922) ) ;
INV     gate2140  (.A(II25198), .Z(g19045) ) ;
DFF     gate2141  (.D(g19045), .CP(CLK), .Q(g1923) ) ;
DFF     gate2142  (.D(g1923), .CP(CLK), .Q(g1924) ) ;
INV     gate2143  (.A(II38716), .Z(g29445) ) ;
DFF     gate2144  (.D(g29445), .CP(CLK), .Q(g1928) ) ;
INV     gate2145  (.A(II25201), .Z(g19046) ) ;
DFF     gate2146  (.D(g19046), .CP(CLK), .Q(g1929) ) ;
DFF     gate2147  (.D(g1929), .CP(CLK), .Q(g1880) ) ;
INV     gate2148  (.A(II25204), .Z(g19047) ) ;
DFF     gate2149  (.D(g19047), .CP(CLK), .Q(g1938) ) ;
DFF     gate2150  (.D(g1938), .CP(CLK), .Q(g1939) ) ;
INV     gate2151  (.A(II37062), .Z(g28271) ) ;
DFF     gate2152  (.D(g28271), .CP(CLK), .Q(g1956) ) ;
INV     gate2153  (.A(II37065), .Z(g28272) ) ;
DFF     gate2154  (.D(g28272), .CP(CLK), .Q(g1957) ) ;
INV     gate2155  (.A(II37068), .Z(g28273) ) ;
DFF     gate2156  (.D(g28273), .CP(CLK), .Q(g1955) ) ;
INV     gate2157  (.A(II37071), .Z(g28274) ) ;
DFF     gate2158  (.D(g28274), .CP(CLK), .Q(g1959) ) ;
INV     gate2159  (.A(II37074), .Z(g28275) ) ;
DFF     gate2160  (.D(g28275), .CP(CLK), .Q(g1960) ) ;
INV     gate2161  (.A(II37077), .Z(g28276) ) ;
DFF     gate2162  (.D(g28276), .CP(CLK), .Q(g1958) ) ;
INV     gate2163  (.A(II37080), .Z(g28277) ) ;
DFF     gate2164  (.D(g28277), .CP(CLK), .Q(g1962) ) ;
INV     gate2165  (.A(II37083), .Z(g28278) ) ;
DFF     gate2166  (.D(g28278), .CP(CLK), .Q(g1963) ) ;
INV     gate2167  (.A(II37086), .Z(g28279) ) ;
DFF     gate2168  (.D(g28279), .CP(CLK), .Q(g1961) ) ;
INV     gate2169  (.A(II37089), .Z(g28280) ) ;
DFF     gate2170  (.D(g28280), .CP(CLK), .Q(g1965) ) ;
INV     gate2171  (.A(II37092), .Z(g28281) ) ;
DFF     gate2172  (.D(g28281), .CP(CLK), .Q(g1966) ) ;
INV     gate2173  (.A(II37095), .Z(g28282) ) ;
DFF     gate2174  (.D(g28282), .CP(CLK), .Q(g1964) ) ;
INV     gate2175  (.A(II33861), .Z(g26003) ) ;
DFF     gate2176  (.D(g26003), .CP(CLK), .Q(g1967) ) ;
INV     gate2177  (.A(II33864), .Z(g26004) ) ;
DFF     gate2178  (.D(g26004), .CP(CLK), .Q(g1970) ) ;
INV     gate2179  (.A(II33867), .Z(g26005) ) ;
DFF     gate2180  (.D(g26005), .CP(CLK), .Q(g1973) ) ;
INV     gate2181  (.A(II33870), .Z(g26006) ) ;
DFF     gate2182  (.D(g26006), .CP(CLK), .Q(g1976) ) ;
INV     gate2183  (.A(II33873), .Z(g26007) ) ;
DFF     gate2184  (.D(g26007), .CP(CLK), .Q(g1979) ) ;
INV     gate2185  (.A(II33876), .Z(g26008) ) ;
DFF     gate2186  (.D(g26008), .CP(CLK), .Q(g1982) ) ;
INV     gate2187  (.A(II38196), .Z(g29151) ) ;
DFF     gate2188  (.D(g29151), .CP(CLK), .Q(g1994) ) ;
INV     gate2189  (.A(II38199), .Z(g29152) ) ;
DFF     gate2190  (.D(g29152), .CP(CLK), .Q(g1997) ) ;
INV     gate2191  (.A(II38202), .Z(g29153) ) ;
DFF     gate2192  (.D(g29153), .CP(CLK), .Q(g2000) ) ;
INV     gate2193  (.A(II38187), .Z(g29148) ) ;
DFF     gate2194  (.D(g29148), .CP(CLK), .Q(g1985) ) ;
INV     gate2195  (.A(II38190), .Z(g29149) ) ;
DFF     gate2196  (.D(g29149), .CP(CLK), .Q(g1988) ) ;
INV     gate2197  (.A(II38193), .Z(g29150) ) ;
DFF     gate2198  (.D(g29150), .CP(CLK), .Q(g1991) ) ;
INV     gate2199  (.A(II35509), .Z(g27224) ) ;
DFF     gate2200  (.D(g27224), .CP(CLK), .Q(g1871) ) ;
INV     gate2201  (.A(II35512), .Z(g27225) ) ;
DFF     gate2202  (.D(g27225), .CP(CLK), .Q(g1874) ) ;
INV     gate2203  (.A(II35515), .Z(g27226) ) ;
DFF     gate2204  (.D(g27226), .CP(CLK), .Q(g1877) ) ;
INV     gate2205  (.A(II15511), .Z(g8302) ) ;
DFF     gate2206  (.D(g8302), .CP(CLK), .Q(g1886) ) ;
INV     gate2207  (.A(II31805), .Z(g24377) ) ;
DFF     gate2208  (.D(g24377), .CP(CLK), .Q(g1887) ) ;
INV     gate2209  (.A(II25186), .Z(g19041) ) ;
DFF     gate2210  (.D(g19041), .CP(CLK), .Q(g1888) ) ;
INV     gate2211  (.A(II25189), .Z(g19042) ) ;
DFF     gate2212  (.D(g19042), .CP(CLK), .Q(g1889) ) ;
INV     gate2213  (.A(II25192), .Z(g19043) ) ;
DFF     gate2214  (.D(g19043), .CP(CLK), .Q(g1894) ) ;
INV     gate2215  (.A(II25195), .Z(g19044) ) ;
DFF     gate2216  (.D(g19044), .CP(CLK), .Q(g1895) ) ;
INV     gate2217  (.A(II38713), .Z(g29444) ) ;
DFF     gate2218  (.D(g29444), .CP(CLK), .Q(g1896) ) ;
INV     gate2219  (.A(II38710), .Z(g29443) ) ;
DFF     gate2220  (.D(g29443), .CP(CLK), .Q(g1897) ) ;
INV     gate2221  (.A(II38707), .Z(g29442) ) ;
DFF     gate2222  (.D(g29442), .CP(CLK), .Q(g1898) ) ;
INV     gate2223  (.A(II38704), .Z(g29441) ) ;
DFF     gate2224  (.D(g29441), .CP(CLK), .Q(g1899) ) ;
INV     gate2225  (.A(II38701), .Z(g29440) ) ;
DFF     gate2226  (.D(g29440), .CP(CLK), .Q(g1900) ) ;
DFF     gate2227  (.D(g1900), .CP(CLK), .Q(g1905) ) ;
INV     gate2228  (.A(II20625), .Z(g13442) ) ;
DFF     gate2229  (.D(g13442), .CP(CLK), .Q(g1909) ) ;
INV     gate2230  (.A(II20628), .Z(g13443) ) ;
DFF     gate2231  (.D(g13443), .CP(CLK), .Q(g1910) ) ;
INV     gate2232  (.A(II20631), .Z(g13444) ) ;
DFF     gate2233  (.D(g13444), .CP(CLK), .Q(g1911) ) ;
INV     gate2234  (.A(II20634), .Z(g13445) ) ;
DFF     gate2235  (.D(g13445), .CP(CLK), .Q(g1912) ) ;
INV     gate2236  (.A(II20637), .Z(g13446) ) ;
DFF     gate2237  (.D(g13446), .CP(CLK), .Q(g1913) ) ;
INV     gate2238  (.A(II20640), .Z(g13447) ) ;
DFF     gate2239  (.D(g13447), .CP(CLK), .Q(g1914) ) ;
INV     gate2240  (.A(II20643), .Z(g13448) ) ;
DFF     gate2241  (.D(g13448), .CP(CLK), .Q(g1916) ) ;
INV     gate2242  (.A(II20646), .Z(g13449) ) ;
DFF     gate2243  (.D(g13449), .CP(CLK), .Q(g1917) ) ;
INV     gate2244  (.A(II33858), .Z(g26002) ) ;
DFF     gate2245  (.D(g26002), .CP(CLK), .Q(g1918) ) ;
INV     gate2246  (.A(II20649), .Z(g13450) ) ;
DFF     gate2247  (.D(g13450), .CP(CLK), .Q(g1921) ) ;
INV     gate2248  (.A(II20655), .Z(g13452) ) ;
DFF     gate2249  (.D(g13452), .CP(CLK), .Q(g2003) ) ;
DFF     gate2250  (.D(g2003), .CP(CLK), .Q(g2006) ) ;
DFF     gate2251  (.D(g2006), .CP(CLK), .Q(g2009) ) ;
INV     gate2252  (.A(II27023), .Z(g20566) ) ;
DFF     gate2253  (.D(g20566), .CP(CLK), .Q(g2010) ) ;
INV     gate2254  (.A(II28461), .Z(g21945) ) ;
DFF     gate2255  (.D(g21945), .CP(CLK), .Q(g2039) ) ;
INV     gate2256  (.A(II30164), .Z(g23237) ) ;
DFF     gate2257  (.D(g23237), .CP(CLK), .Q(g2020) ) ;
INV     gate2258  (.A(II31808), .Z(g24378) ) ;
DFF     gate2259  (.D(g24378), .CP(CLK), .Q(g2013) ) ;
INV     gate2260  (.A(II32964), .Z(g25162) ) ;
DFF     gate2261  (.D(g25162), .CP(CLK), .Q(g2033) ) ;
INV     gate2262  (.A(II33879), .Z(g26009) ) ;
DFF     gate2263  (.D(g26009), .CP(CLK), .Q(g2026) ) ;
INV     gate2264  (.A(II34782), .Z(g26725) ) ;
DFF     gate2265  (.D(g26725), .CP(CLK), .Q(g2040) ) ;
INV     gate2266  (.A(II35518), .Z(g27227) ) ;
DFF     gate2267  (.D(g27227), .CP(CLK), .Q(g2052) ) ;
INV     gate2268  (.A(II36129), .Z(g27706) ) ;
DFF     gate2269  (.D(g27706), .CP(CLK), .Q(g2046) ) ;
INV     gate2270  (.A(II37098), .Z(g28283) ) ;
DFF     gate2271  (.D(g28283), .CP(CLK), .Q(g2059) ) ;
INV     gate2272  (.A(II37608), .Z(g28687) ) ;
DFF     gate2273  (.D(g28687), .CP(CLK), .Q(g2066) ) ;
INV     gate2274  (.A(II38205), .Z(g29154) ) ;
DFF     gate2275  (.D(g29154), .CP(CLK), .Q(g2072) ) ;
INV     gate2276  (.A(II30167), .Z(g23238) ) ;
DFF     gate2277  (.D(g23238), .CP(CLK), .Q(g2079) ) ;
INV     gate2278  (.A(II30170), .Z(g23239) ) ;
DFF     gate2279  (.D(g23239), .CP(CLK), .Q(g2080) ) ;
INV     gate2280  (.A(II30173), .Z(g23240) ) ;
DFF     gate2281  (.D(g23240), .CP(CLK), .Q(g2078) ) ;
INV     gate2282  (.A(II30176), .Z(g23241) ) ;
DFF     gate2283  (.D(g23241), .CP(CLK), .Q(g2082) ) ;
INV     gate2284  (.A(II30179), .Z(g23242) ) ;
DFF     gate2285  (.D(g23242), .CP(CLK), .Q(g2083) ) ;
INV     gate2286  (.A(II30182), .Z(g23243) ) ;
DFF     gate2287  (.D(g23243), .CP(CLK), .Q(g2081) ) ;
INV     gate2288  (.A(II30185), .Z(g23244) ) ;
DFF     gate2289  (.D(g23244), .CP(CLK), .Q(g2085) ) ;
INV     gate2290  (.A(II30188), .Z(g23245) ) ;
DFF     gate2291  (.D(g23245), .CP(CLK), .Q(g2086) ) ;
INV     gate2292  (.A(II30191), .Z(g23246) ) ;
DFF     gate2293  (.D(g23246), .CP(CLK), .Q(g2084) ) ;
INV     gate2294  (.A(II30194), .Z(g23247) ) ;
DFF     gate2295  (.D(g23247), .CP(CLK), .Q(g2088) ) ;
INV     gate2296  (.A(II30197), .Z(g23248) ) ;
DFF     gate2297  (.D(g23248), .CP(CLK), .Q(g2089) ) ;
INV     gate2298  (.A(II30200), .Z(g23249) ) ;
DFF     gate2299  (.D(g23249), .CP(CLK), .Q(g2087) ) ;
INV     gate2300  (.A(II30203), .Z(g23250) ) ;
DFF     gate2301  (.D(g23250), .CP(CLK), .Q(g2091) ) ;
INV     gate2302  (.A(II30206), .Z(g23251) ) ;
DFF     gate2303  (.D(g23251), .CP(CLK), .Q(g2092) ) ;
INV     gate2304  (.A(II30209), .Z(g23252) ) ;
DFF     gate2305  (.D(g23252), .CP(CLK), .Q(g2090) ) ;
INV     gate2306  (.A(II30212), .Z(g23253) ) ;
DFF     gate2307  (.D(g23253), .CP(CLK), .Q(g2094) ) ;
INV     gate2308  (.A(II30215), .Z(g23254) ) ;
DFF     gate2309  (.D(g23254), .CP(CLK), .Q(g2095) ) ;
INV     gate2310  (.A(II30218), .Z(g23255) ) ;
DFF     gate2311  (.D(g23255), .CP(CLK), .Q(g2093) ) ;
INV     gate2312  (.A(II30221), .Z(g23256) ) ;
DFF     gate2313  (.D(g23256), .CP(CLK), .Q(g2097) ) ;
INV     gate2314  (.A(II30224), .Z(g23257) ) ;
DFF     gate2315  (.D(g23257), .CP(CLK), .Q(g2098) ) ;
INV     gate2316  (.A(II30227), .Z(g23258) ) ;
DFF     gate2317  (.D(g23258), .CP(CLK), .Q(g2096) ) ;
INV     gate2318  (.A(II30230), .Z(g23259) ) ;
DFF     gate2319  (.D(g23259), .CP(CLK), .Q(g2100) ) ;
INV     gate2320  (.A(II30233), .Z(g23260) ) ;
DFF     gate2321  (.D(g23260), .CP(CLK), .Q(g2101) ) ;
INV     gate2322  (.A(II30236), .Z(g23261) ) ;
DFF     gate2323  (.D(g23261), .CP(CLK), .Q(g2099) ) ;
INV     gate2324  (.A(II30239), .Z(g23262) ) ;
DFF     gate2325  (.D(g23262), .CP(CLK), .Q(g2103) ) ;
INV     gate2326  (.A(II30242), .Z(g23263) ) ;
DFF     gate2327  (.D(g23263), .CP(CLK), .Q(g2104) ) ;
INV     gate2328  (.A(II30245), .Z(g23264) ) ;
DFF     gate2329  (.D(g23264), .CP(CLK), .Q(g2102) ) ;
INV     gate2330  (.A(II30248), .Z(g23265) ) ;
DFF     gate2331  (.D(g23265), .CP(CLK), .Q(g2106) ) ;
INV     gate2332  (.A(II30251), .Z(g23266) ) ;
DFF     gate2333  (.D(g23266), .CP(CLK), .Q(g2107) ) ;
INV     gate2334  (.A(II30254), .Z(g23267) ) ;
DFF     gate2335  (.D(g23267), .CP(CLK), .Q(g2105) ) ;
INV     gate2336  (.A(II30257), .Z(g23268) ) ;
DFF     gate2337  (.D(g23268), .CP(CLK), .Q(g2109) ) ;
INV     gate2338  (.A(II30260), .Z(g23269) ) ;
DFF     gate2339  (.D(g23269), .CP(CLK), .Q(g2110) ) ;
INV     gate2340  (.A(II30263), .Z(g23270) ) ;
DFF     gate2341  (.D(g23270), .CP(CLK), .Q(g2108) ) ;
INV     gate2342  (.A(II30266), .Z(g23271) ) ;
DFF     gate2343  (.D(g23271), .CP(CLK), .Q(g2112) ) ;
INV     gate2344  (.A(II30269), .Z(g23272) ) ;
DFF     gate2345  (.D(g23272), .CP(CLK), .Q(g2113) ) ;
INV     gate2346  (.A(II30272), .Z(g23273) ) ;
DFF     gate2347  (.D(g23273), .CP(CLK), .Q(g2111) ) ;
INV     gate2348  (.A(II34785), .Z(g26726) ) ;
DFF     gate2349  (.D(g26726), .CP(CLK), .Q(g2115) ) ;
INV     gate2350  (.A(II34788), .Z(g26727) ) ;
DFF     gate2351  (.D(g26727), .CP(CLK), .Q(g2116) ) ;
INV     gate2352  (.A(II34791), .Z(g26728) ) ;
DFF     gate2353  (.D(g26728), .CP(CLK), .Q(g2114) ) ;
INV     gate2354  (.A(II31811), .Z(g24379) ) ;
DFF     gate2355  (.D(g24379), .CP(CLK), .Q(g2118) ) ;
INV     gate2356  (.A(II31814), .Z(g24380) ) ;
DFF     gate2357  (.D(g24380), .CP(CLK), .Q(g2119) ) ;
INV     gate2358  (.A(II31817), .Z(g24381) ) ;
DFF     gate2359  (.D(g24381), .CP(CLK), .Q(g2117) ) ;
INV     gate2360  (.A(II20658), .Z(g13453) ) ;
DFF     gate2361  (.D(g13453), .CP(CLK), .Q(g2214) ) ;
DFF     gate2362  (.D(g2214), .CP(CLK), .Q(g2211) ) ;
DFF     gate2363  (.D(g2211), .CP(CLK), .Q(g2241) ) ;
INV     gate2364  (.A(II31820), .Z(g24382) ) ;
DFF     gate2365  (.D(g24382), .CP(CLK), .Q(g2206) ) ;
INV     gate2366  (.A(II31823), .Z(g24383) ) ;
DFF     gate2367  (.D(g24383), .CP(CLK), .Q(g2207) ) ;
INV     gate2368  (.A(II31826), .Z(g24384) ) ;
DFF     gate2369  (.D(g24384), .CP(CLK), .Q(g2205) ) ;
INV     gate2370  (.A(II31829), .Z(g24385) ) ;
DFF     gate2371  (.D(g24385), .CP(CLK), .Q(g2209) ) ;
INV     gate2372  (.A(II31832), .Z(g24386) ) ;
DFF     gate2373  (.D(g24386), .CP(CLK), .Q(g2210) ) ;
INV     gate2374  (.A(II31835), .Z(g24387) ) ;
DFF     gate2375  (.D(g24387), .CP(CLK), .Q(g2208) ) ;
INV     gate2376  (.A(II31838), .Z(g24388) ) ;
DFF     gate2377  (.D(g24388), .CP(CLK), .Q(g2218) ) ;
INV     gate2378  (.A(II31841), .Z(g24389) ) ;
DFF     gate2379  (.D(g24389), .CP(CLK), .Q(g2219) ) ;
INV     gate2380  (.A(II31844), .Z(g24390) ) ;
DFF     gate2381  (.D(g24390), .CP(CLK), .Q(g2217) ) ;
INV     gate2382  (.A(II31847), .Z(g24391) ) ;
DFF     gate2383  (.D(g24391), .CP(CLK), .Q(g2221) ) ;
INV     gate2384  (.A(II31850), .Z(g24392) ) ;
DFF     gate2385  (.D(g24392), .CP(CLK), .Q(g2222) ) ;
INV     gate2386  (.A(II31853), .Z(g24393) ) ;
DFF     gate2387  (.D(g24393), .CP(CLK), .Q(g2220) ) ;
INV     gate2388  (.A(II31856), .Z(g24394) ) ;
DFF     gate2389  (.D(g24394), .CP(CLK), .Q(g2224) ) ;
INV     gate2390  (.A(II31859), .Z(g24395) ) ;
DFF     gate2391  (.D(g24395), .CP(CLK), .Q(g2225) ) ;
INV     gate2392  (.A(II31862), .Z(g24396) ) ;
DFF     gate2393  (.D(g24396), .CP(CLK), .Q(g2223) ) ;
INV     gate2394  (.A(II31865), .Z(g24397) ) ;
DFF     gate2395  (.D(g24397), .CP(CLK), .Q(g2227) ) ;
INV     gate2396  (.A(II31868), .Z(g24398) ) ;
DFF     gate2397  (.D(g24398), .CP(CLK), .Q(g2228) ) ;
INV     gate2398  (.A(II31871), .Z(g24399) ) ;
DFF     gate2399  (.D(g24399), .CP(CLK), .Q(g2226) ) ;
INV     gate2400  (.A(II31874), .Z(g24400) ) ;
DFF     gate2401  (.D(g24400), .CP(CLK), .Q(g2230) ) ;
INV     gate2402  (.A(II31877), .Z(g24401) ) ;
DFF     gate2403  (.D(g24401), .CP(CLK), .Q(g2231) ) ;
INV     gate2404  (.A(II31880), .Z(g24402) ) ;
DFF     gate2405  (.D(g24402), .CP(CLK), .Q(g2229) ) ;
INV     gate2406  (.A(II31883), .Z(g24403) ) ;
DFF     gate2407  (.D(g24403), .CP(CLK), .Q(g2233) ) ;
INV     gate2408  (.A(II31886), .Z(g24404) ) ;
DFF     gate2409  (.D(g24404), .CP(CLK), .Q(g2234) ) ;
INV     gate2410  (.A(II31889), .Z(g24405) ) ;
DFF     gate2411  (.D(g24405), .CP(CLK), .Q(g2232) ) ;
INV     gate2412  (.A(II31892), .Z(g24406) ) ;
DFF     gate2413  (.D(g24406), .CP(CLK), .Q(g2236) ) ;
INV     gate2414  (.A(II31895), .Z(g24407) ) ;
DFF     gate2415  (.D(g24407), .CP(CLK), .Q(g2237) ) ;
INV     gate2416  (.A(II31898), .Z(g24408) ) ;
DFF     gate2417  (.D(g24408), .CP(CLK), .Q(g2235) ) ;
INV     gate2418  (.A(II31901), .Z(g24409) ) ;
DFF     gate2419  (.D(g24409), .CP(CLK), .Q(g2239) ) ;
INV     gate2420  (.A(II31904), .Z(g24410) ) ;
DFF     gate2421  (.D(g24410), .CP(CLK), .Q(g2240) ) ;
INV     gate2422  (.A(II31907), .Z(g24411) ) ;
DFF     gate2423  (.D(g24411), .CP(CLK), .Q(g2238) ) ;
INV     gate2424  (.A(II34797), .Z(g26730) ) ;
DFF     gate2425  (.D(g26730), .CP(CLK), .Q(g2245) ) ;
INV     gate2426  (.A(II34800), .Z(g26731) ) ;
DFF     gate2427  (.D(g26731), .CP(CLK), .Q(g2246) ) ;
INV     gate2428  (.A(II34803), .Z(g26732) ) ;
DFF     gate2429  (.D(g26732), .CP(CLK), .Q(g2244) ) ;
INV     gate2430  (.A(II34806), .Z(g26733) ) ;
DFF     gate2431  (.D(g26733), .CP(CLK), .Q(g2248) ) ;
INV     gate2432  (.A(II34809), .Z(g26734) ) ;
DFF     gate2433  (.D(g26734), .CP(CLK), .Q(g2249) ) ;
INV     gate2434  (.A(II34812), .Z(g26735) ) ;
DFF     gate2435  (.D(g26735), .CP(CLK), .Q(g2247) ) ;
INV     gate2436  (.A(II34815), .Z(g26736) ) ;
DFF     gate2437  (.D(g26736), .CP(CLK), .Q(g2251) ) ;
INV     gate2438  (.A(II34818), .Z(g26737) ) ;
DFF     gate2439  (.D(g26737), .CP(CLK), .Q(g2252) ) ;
INV     gate2440  (.A(II34821), .Z(g26738) ) ;
DFF     gate2441  (.D(g26738), .CP(CLK), .Q(g2250) ) ;
INV     gate2442  (.A(II34824), .Z(g26739) ) ;
DFF     gate2443  (.D(g26739), .CP(CLK), .Q(g2254) ) ;
INV     gate2444  (.A(II34827), .Z(g26740) ) ;
DFF     gate2445  (.D(g26740), .CP(CLK), .Q(g2255) ) ;
INV     gate2446  (.A(II34830), .Z(g26741) ) ;
DFF     gate2447  (.D(g26741), .CP(CLK), .Q(g2253) ) ;
INV     gate2448  (.A(II40233), .Z(g30551) ) ;
DFF     gate2449  (.D(g30551), .CP(CLK), .Q(g2261) ) ;
INV     gate2450  (.A(II40236), .Z(g30552) ) ;
DFF     gate2451  (.D(g30552), .CP(CLK), .Q(g2264) ) ;
INV     gate2452  (.A(II40239), .Z(g30553) ) ;
DFF     gate2453  (.D(g30553), .CP(CLK), .Q(g2267) ) ;
INV     gate2454  (.A(II40940), .Z(g30896) ) ;
DFF     gate2455  (.D(g30896), .CP(CLK), .Q(g2306) ) ;
INV     gate2456  (.A(II40943), .Z(g30897) ) ;
DFF     gate2457  (.D(g30897), .CP(CLK), .Q(g2309) ) ;
INV     gate2458  (.A(II40946), .Z(g30898) ) ;
DFF     gate2459  (.D(g30898), .CP(CLK), .Q(g2312) ) ;
INV     gate2460  (.A(II40922), .Z(g30890) ) ;
DFF     gate2461  (.D(g30890), .CP(CLK), .Q(g2270) ) ;
INV     gate2462  (.A(II40925), .Z(g30891) ) ;
DFF     gate2463  (.D(g30891), .CP(CLK), .Q(g2273) ) ;
INV     gate2464  (.A(II40928), .Z(g30892) ) ;
DFF     gate2465  (.D(g30892), .CP(CLK), .Q(g2276) ) ;
INV     gate2466  (.A(II40949), .Z(g30899) ) ;
DFF     gate2467  (.D(g30899), .CP(CLK), .Q(g2315) ) ;
INV     gate2468  (.A(II40952), .Z(g30900) ) ;
DFF     gate2469  (.D(g30900), .CP(CLK), .Q(g2318) ) ;
INV     gate2470  (.A(II40955), .Z(g30901) ) ;
DFF     gate2471  (.D(g30901), .CP(CLK), .Q(g2321) ) ;
INV     gate2472  (.A(II40242), .Z(g30554) ) ;
DFF     gate2473  (.D(g30554), .CP(CLK), .Q(g2279) ) ;
INV     gate2474  (.A(II40245), .Z(g30555) ) ;
DFF     gate2475  (.D(g30555), .CP(CLK), .Q(g2282) ) ;
INV     gate2476  (.A(II40248), .Z(g30556) ) ;
DFF     gate2477  (.D(g30556), .CP(CLK), .Q(g2285) ) ;
INV     gate2478  (.A(II40260), .Z(g30560) ) ;
DFF     gate2479  (.D(g30560), .CP(CLK), .Q(g2324) ) ;
INV     gate2480  (.A(II40263), .Z(g30561) ) ;
DFF     gate2481  (.D(g30561), .CP(CLK), .Q(g2327) ) ;
INV     gate2482  (.A(II40266), .Z(g30562) ) ;
DFF     gate2483  (.D(g30562), .CP(CLK), .Q(g2330) ) ;
INV     gate2484  (.A(II40251), .Z(g30557) ) ;
DFF     gate2485  (.D(g30557), .CP(CLK), .Q(g2288) ) ;
INV     gate2486  (.A(II40254), .Z(g30558) ) ;
DFF     gate2487  (.D(g30558), .CP(CLK), .Q(g2291) ) ;
INV     gate2488  (.A(II40257), .Z(g30559) ) ;
DFF     gate2489  (.D(g30559), .CP(CLK), .Q(g2294) ) ;
INV     gate2490  (.A(II40269), .Z(g30563) ) ;
DFF     gate2491  (.D(g30563), .CP(CLK), .Q(g2333) ) ;
INV     gate2492  (.A(II40272), .Z(g30564) ) ;
DFF     gate2493  (.D(g30564), .CP(CLK), .Q(g2336) ) ;
INV     gate2494  (.A(II40275), .Z(g30565) ) ;
DFF     gate2495  (.D(g30565), .CP(CLK), .Q(g2339) ) ;
INV     gate2496  (.A(II40931), .Z(g30893) ) ;
DFF     gate2497  (.D(g30893), .CP(CLK), .Q(g2297) ) ;
INV     gate2498  (.A(II40934), .Z(g30894) ) ;
DFF     gate2499  (.D(g30894), .CP(CLK), .Q(g2300) ) ;
INV     gate2500  (.A(II40937), .Z(g30895) ) ;
DFF     gate2501  (.D(g30895), .CP(CLK), .Q(g2303) ) ;
INV     gate2502  (.A(II40958), .Z(g30902) ) ;
DFF     gate2503  (.D(g30902), .CP(CLK), .Q(g2342) ) ;
INV     gate2504  (.A(II40961), .Z(g30903) ) ;
DFF     gate2505  (.D(g30903), .CP(CLK), .Q(g2345) ) ;
INV     gate2506  (.A(II40964), .Z(g30904) ) ;
DFF     gate2507  (.D(g30904), .CP(CLK), .Q(g2348) ) ;
INV     gate2508  (.A(II33882), .Z(g26010) ) ;
DFF     gate2509  (.D(g26010), .CP(CLK), .Q(g2160) ) ;
INV     gate2510  (.A(II34794), .Z(g26729) ) ;
DFF     gate2511  (.D(g26729), .CP(CLK), .Q(g2156) ) ;
INV     gate2512  (.A(II35521), .Z(g27228) ) ;
DFF     gate2513  (.D(g27228), .CP(CLK), .Q(g2151) ) ;
INV     gate2514  (.A(II36132), .Z(g27707) ) ;
DFF     gate2515  (.D(g27707), .CP(CLK), .Q(g2147) ) ;
INV     gate2516  (.A(II37101), .Z(g28284) ) ;
DFF     gate2517  (.D(g28284), .CP(CLK), .Q(g2142) ) ;
INV     gate2518  (.A(II37611), .Z(g28688) ) ;
DFF     gate2519  (.D(g28688), .CP(CLK), .Q(g2138) ) ;
INV     gate2520  (.A(II38208), .Z(g29155) ) ;
DFF     gate2521  (.D(g29155), .CP(CLK), .Q(g2133) ) ;
INV     gate2522  (.A(II38719), .Z(g29446) ) ;
DFF     gate2523  (.D(g29446), .CP(CLK), .Q(g2129) ) ;
INV     gate2524  (.A(II39062), .Z(g29648) ) ;
DFF     gate2525  (.D(g29648), .CP(CLK), .Q(g2124) ) ;
INV     gate2526  (.A(II39270), .Z(g29806) ) ;
DFF     gate2527  (.D(g29806), .CP(CLK), .Q(g2120) ) ;
INV     gate2528  (.A(II27026), .Z(g20567) ) ;
DFF     gate2529  (.D(g20567), .CP(CLK), .Q(g2256) ) ;
DFF     gate2530  (.D(g2256), .CP(CLK), .Q(g2258) ) ;
DFF     gate2531  (.D(g2258), .CP(CLK), .Q(g2257) ) ;
INV     gate2532  (.A(II20661), .Z(g13454) ) ;
DFF     gate2533  (.D(g13454), .CP(CLK), .Q(g2351) ) ;
DFF     gate2534  (.D(g2351), .CP(CLK), .Q(g2480) ) ;
DFF     gate2535  (.D(g2480), .CP(CLK), .Q(g2476) ) ;
INV     gate2536  (.A(II18707), .Z(g11577) ) ;
DFF     gate2537  (.D(g11577), .CP(CLK), .Q(g2384) ) ;
INV     gate2538  (.A(II37104), .Z(g28285) ) ;
DFF     gate2539  (.D(g28285), .CP(CLK), .Q(g2429) ) ;
INV     gate2540  (.A(II37107), .Z(g28286) ) ;
DFF     gate2541  (.D(g28286), .CP(CLK), .Q(g2418) ) ;
INV     gate2542  (.A(II37110), .Z(g28287) ) ;
DFF     gate2543  (.D(g28287), .CP(CLK), .Q(g2421) ) ;
INV     gate2544  (.A(II37113), .Z(g28288) ) ;
DFF     gate2545  (.D(g28288), .CP(CLK), .Q(g2444) ) ;
INV     gate2546  (.A(II37116), .Z(g28289) ) ;
DFF     gate2547  (.D(g28289), .CP(CLK), .Q(g2433) ) ;
INV     gate2548  (.A(II37119), .Z(g28290) ) ;
DFF     gate2549  (.D(g28290), .CP(CLK), .Q(g2436) ) ;
INV     gate2550  (.A(II37122), .Z(g28291) ) ;
DFF     gate2551  (.D(g28291), .CP(CLK), .Q(g2459) ) ;
INV     gate2552  (.A(II37125), .Z(g28292) ) ;
DFF     gate2553  (.D(g28292), .CP(CLK), .Q(g2448) ) ;
INV     gate2554  (.A(II37128), .Z(g28293) ) ;
DFF     gate2555  (.D(g28293), .CP(CLK), .Q(g2451) ) ;
INV     gate2556  (.A(II37131), .Z(g28294) ) ;
DFF     gate2557  (.D(g28294), .CP(CLK), .Q(g2473) ) ;
INV     gate2558  (.A(II37134), .Z(g28295) ) ;
DFF     gate2559  (.D(g28295), .CP(CLK), .Q(g2463) ) ;
INV     gate2560  (.A(II37137), .Z(g28296) ) ;
DFF     gate2561  (.D(g28296), .CP(CLK), .Q(g2466) ) ;
INV     gate2562  (.A(II38722), .Z(g29447) ) ;
DFF     gate2563  (.D(g29447), .CP(CLK), .Q(g2483) ) ;
INV     gate2564  (.A(II38725), .Z(g29448) ) ;
DFF     gate2565  (.D(g29448), .CP(CLK), .Q(g2486) ) ;
INV     gate2566  (.A(II38728), .Z(g29449) ) ;
DFF     gate2567  (.D(g29449), .CP(CLK), .Q(g2489) ) ;
INV     gate2568  (.A(II39074), .Z(g29652) ) ;
DFF     gate2569  (.D(g29652), .CP(CLK), .Q(g2492) ) ;
INV     gate2570  (.A(II39077), .Z(g29653) ) ;
DFF     gate2571  (.D(g29653), .CP(CLK), .Q(g2495) ) ;
INV     gate2572  (.A(II39080), .Z(g29654) ) ;
DFF     gate2573  (.D(g29654), .CP(CLK), .Q(g2498) ) ;
INV     gate2574  (.A(II38731), .Z(g29450) ) ;
DFF     gate2575  (.D(g29450), .CP(CLK), .Q(g2502) ) ;
INV     gate2576  (.A(II38734), .Z(g29451) ) ;
DFF     gate2577  (.D(g29451), .CP(CLK), .Q(g2503) ) ;
INV     gate2578  (.A(II38737), .Z(g29452) ) ;
DFF     gate2579  (.D(g29452), .CP(CLK), .Q(g2501) ) ;
INV     gate2580  (.A(II36135), .Z(g27708) ) ;
DFF     gate2581  (.D(g27708), .CP(CLK), .Q(g2504) ) ;
INV     gate2582  (.A(II36138), .Z(g27709) ) ;
DFF     gate2583  (.D(g27709), .CP(CLK), .Q(g2507) ) ;
INV     gate2584  (.A(II36141), .Z(g27710) ) ;
DFF     gate2585  (.D(g27710), .CP(CLK), .Q(g2510) ) ;
INV     gate2586  (.A(II36144), .Z(g27711) ) ;
DFF     gate2587  (.D(g27711), .CP(CLK), .Q(g2513) ) ;
INV     gate2588  (.A(II36147), .Z(g27712) ) ;
DFF     gate2589  (.D(g27712), .CP(CLK), .Q(g2516) ) ;
INV     gate2590  (.A(II36150), .Z(g27713) ) ;
DFF     gate2591  (.D(g27713), .CP(CLK), .Q(g2519) ) ;
INV     gate2592  (.A(II37614), .Z(g28689) ) ;
DFF     gate2593  (.D(g28689), .CP(CLK), .Q(g2523) ) ;
INV     gate2594  (.A(II37617), .Z(g28690) ) ;
DFF     gate2595  (.D(g28690), .CP(CLK), .Q(g2524) ) ;
INV     gate2596  (.A(II37620), .Z(g28691) ) ;
DFF     gate2597  (.D(g28691), .CP(CLK), .Q(g2522) ) ;
INV     gate2598  (.A(II39273), .Z(g29807) ) ;
DFF     gate2599  (.D(g29807), .CP(CLK), .Q(g2387) ) ;
INV     gate2600  (.A(II39276), .Z(g29808) ) ;
DFF     gate2601  (.D(g29808), .CP(CLK), .Q(g2388) ) ;
INV     gate2602  (.A(II39279), .Z(g29809) ) ;
DFF     gate2603  (.D(g29809), .CP(CLK), .Q(g2389) ) ;
INV     gate2604  (.A(II40967), .Z(g30905) ) ;
DFF     gate2605  (.D(g30905), .CP(CLK), .Q(g2390) ) ;
INV     gate2606  (.A(II40970), .Z(g30906) ) ;
DFF     gate2607  (.D(g30906), .CP(CLK), .Q(g2391) ) ;
INV     gate2608  (.A(II40973), .Z(g30907) ) ;
DFF     gate2609  (.D(g30907), .CP(CLK), .Q(g2392) ) ;
INV     gate2610  (.A(II40447), .Z(g30719) ) ;
DFF     gate2611  (.D(g30719), .CP(CLK), .Q(g2393) ) ;
INV     gate2612  (.A(II40450), .Z(g30720) ) ;
DFF     gate2613  (.D(g30720), .CP(CLK), .Q(g2394) ) ;
INV     gate2614  (.A(II40453), .Z(g30721) ) ;
DFF     gate2615  (.D(g30721), .CP(CLK), .Q(g2395) ) ;
INV     gate2616  (.A(II39065), .Z(g29649) ) ;
DFF     gate2617  (.D(g29649), .CP(CLK), .Q(g2397) ) ;
INV     gate2618  (.A(II39068), .Z(g29650) ) ;
DFF     gate2619  (.D(g29650), .CP(CLK), .Q(g2398) ) ;
INV     gate2620  (.A(II39071), .Z(g29651) ) ;
DFF     gate2621  (.D(g29651), .CP(CLK), .Q(g2396) ) ;
INV     gate2622  (.A(II35527), .Z(g27230) ) ;
DFF     gate2623  (.D(g27230), .CP(CLK), .Q(g2478) ) ;
INV     gate2624  (.A(II35530), .Z(g27231) ) ;
DFF     gate2625  (.D(g27231), .CP(CLK), .Q(g2479) ) ;
INV     gate2626  (.A(II35533), .Z(g27232) ) ;
DFF     gate2627  (.D(g27232), .CP(CLK), .Q(g2477) ) ;
INV     gate2628  (.A(II18746), .Z(g11590) ) ;
DFF     gate2629  (.D(g11590), .CP(CLK), .Q(g2525) ) ;
DFF     gate2630  (.D(g2525), .CP(CLK), .Q(g2526) ) ;
INV     gate2631  (.A(II18749), .Z(g11591) ) ;
DFF     gate2632  (.D(g11591), .CP(CLK), .Q(g2527) ) ;
DFF     gate2633  (.D(g2527), .CP(CLK), .Q(g2528) ) ;
INV     gate2634  (.A(II18752), .Z(g11592) ) ;
DFF     gate2635  (.D(g11592), .CP(CLK), .Q(g2529) ) ;
DFF     gate2636  (.D(g2529), .CP(CLK), .Q(g2354) ) ;
INV     gate2637  (.A(II18692), .Z(g11572) ) ;
DFF     gate2638  (.D(g11572), .CP(CLK), .Q(g2355) ) ;
DFF     gate2639  (.D(g2355), .CP(CLK), .Q(g2356) ) ;
INV     gate2640  (.A(II18695), .Z(g11573) ) ;
DFF     gate2641  (.D(g11573), .CP(CLK), .Q(g2357) ) ;
DFF     gate2642  (.D(g2357), .CP(CLK), .Q(g2358) ) ;
INV     gate2643  (.A(II18698), .Z(g11574) ) ;
DFF     gate2644  (.D(g11574), .CP(CLK), .Q(g2359) ) ;
DFF     gate2645  (.D(g2359), .CP(CLK), .Q(g2360) ) ;
INV     gate2646  (.A(II18701), .Z(g11575) ) ;
DFF     gate2647  (.D(g11575), .CP(CLK), .Q(g2361) ) ;
DFF     gate2648  (.D(g2361), .CP(CLK), .Q(g2362) ) ;
INV     gate2649  (.A(II18704), .Z(g11576) ) ;
DFF     gate2650  (.D(g11576), .CP(CLK), .Q(g2363) ) ;
DFF     gate2651  (.D(g2363), .CP(CLK), .Q(g2364) ) ;
INV     gate2652  (.A(II20664), .Z(g13455) ) ;
DFF     gate2653  (.D(g13455), .CP(CLK), .Q(g2365) ) ;
DFF     gate2654  (.D(g2365), .CP(CLK), .Q(g2366) ) ;
INV     gate2655  (.A(II25207), .Z(g19048) ) ;
DFF     gate2656  (.D(g19048), .CP(CLK), .Q(g2374) ) ;
INV     gate2657  (.A(II39785), .Z(g30314) ) ;
DFF     gate2658  (.D(g30314), .CP(CLK), .Q(g2380) ) ;
INV     gate2659  (.A(II39788), .Z(g30315) ) ;
DFF     gate2660  (.D(g30315), .CP(CLK), .Q(g2383) ) ;
INV     gate2661  (.A(II39791), .Z(g30316) ) ;
DFF     gate2662  (.D(g30316), .CP(CLK), .Q(g2372) ) ;
INV     gate2663  (.A(II39794), .Z(g30317) ) ;
DFF     gate2664  (.D(g30317), .CP(CLK), .Q(g2371) ) ;
INV     gate2665  (.A(II39797), .Z(g30318) ) ;
DFF     gate2666  (.D(g30318), .CP(CLK), .Q(g2370) ) ;
INV     gate2667  (.A(II39800), .Z(g30319) ) ;
DFF     gate2668  (.D(g30319), .CP(CLK), .Q(g2369) ) ;
INV     gate2669  (.A(II25219), .Z(g19052) ) ;
DFF     gate2670  (.D(g19052), .CP(CLK), .Q(g2379) ) ;
INV     gate2671  (.A(II25216), .Z(g19051) ) ;
DFF     gate2672  (.D(g19051), .CP(CLK), .Q(g2378) ) ;
INV     gate2673  (.A(II25213), .Z(g19050) ) ;
DFF     gate2674  (.D(g19050), .CP(CLK), .Q(g2377) ) ;
INV     gate2675  (.A(II25210), .Z(g19049) ) ;
DFF     gate2676  (.D(g19049), .CP(CLK), .Q(g2376) ) ;
INV     gate2677  (.A(II32967), .Z(g25163) ) ;
DFF     gate2678  (.D(g25163), .CP(CLK), .Q(g2375) ) ;
INV     gate2679  (.A(II35524), .Z(g27229) ) ;
DFF     gate2680  (.D(g27229), .CP(CLK), .Q(g2373) ) ;
INV     gate2681  (.A(II18710), .Z(g11578) ) ;
DFF     gate2682  (.D(g11578), .CP(CLK), .Q(g2417) ) ;
DFF     gate2683  (.D(g2417), .CP(CLK), .Q(g2424) ) ;
INV     gate2684  (.A(II18713), .Z(g11579) ) ;
DFF     gate2685  (.D(g11579), .CP(CLK), .Q(g2425) ) ;
DFF     gate2686  (.D(g2425), .CP(CLK), .Q(g2426) ) ;
INV     gate2687  (.A(II18716), .Z(g11580) ) ;
DFF     gate2688  (.D(g11580), .CP(CLK), .Q(g2427) ) ;
DFF     gate2689  (.D(g2427), .CP(CLK), .Q(g2428) ) ;
INV     gate2690  (.A(II18719), .Z(g11581) ) ;
DFF     gate2691  (.D(g11581), .CP(CLK), .Q(g2432) ) ;
DFF     gate2692  (.D(g2432), .CP(CLK), .Q(g2439) ) ;
INV     gate2693  (.A(II18722), .Z(g11582) ) ;
DFF     gate2694  (.D(g11582), .CP(CLK), .Q(g2440) ) ;
DFF     gate2695  (.D(g2440), .CP(CLK), .Q(g2441) ) ;
INV     gate2696  (.A(II18725), .Z(g11583) ) ;
DFF     gate2697  (.D(g11583), .CP(CLK), .Q(g2442) ) ;
DFF     gate2698  (.D(g2442), .CP(CLK), .Q(g2443) ) ;
INV     gate2699  (.A(II18728), .Z(g11584) ) ;
DFF     gate2700  (.D(g11584), .CP(CLK), .Q(g2447) ) ;
DFF     gate2701  (.D(g2447), .CP(CLK), .Q(g2454) ) ;
INV     gate2702  (.A(II18731), .Z(g11585) ) ;
DFF     gate2703  (.D(g11585), .CP(CLK), .Q(g2455) ) ;
DFF     gate2704  (.D(g2455), .CP(CLK), .Q(g2456) ) ;
INV     gate2705  (.A(II18734), .Z(g11586) ) ;
DFF     gate2706  (.D(g11586), .CP(CLK), .Q(g2457) ) ;
DFF     gate2707  (.D(g2457), .CP(CLK), .Q(g2458) ) ;
INV     gate2708  (.A(II18737), .Z(g11587) ) ;
DFF     gate2709  (.D(g11587), .CP(CLK), .Q(g2462) ) ;
DFF     gate2710  (.D(g2462), .CP(CLK), .Q(g2469) ) ;
INV     gate2711  (.A(II18740), .Z(g11588) ) ;
DFF     gate2712  (.D(g11588), .CP(CLK), .Q(g2470) ) ;
DFF     gate2713  (.D(g2470), .CP(CLK), .Q(g2471) ) ;
INV     gate2714  (.A(II18743), .Z(g11589) ) ;
DFF     gate2715  (.D(g11589), .CP(CLK), .Q(g2472) ) ;
DFF     gate2716  (.D(g2472), .CP(CLK), .Q(g2399) ) ;
INV     gate2717  (.A(II20667), .Z(g13456) ) ;
DFF     gate2718  (.D(g13456), .CP(CLK), .Q(g2400) ) ;
DFF     gate2719  (.D(g2400), .CP(CLK), .Q(g2406) ) ;
DFF     gate2720  (.D(g2406), .CP(CLK), .Q(g2412) ) ;
INV     gate2721  (.A(II20700), .Z(g13467) ) ;
DFF     gate2722  (.D(g13467), .CP(CLK), .Q(g2619) ) ;
DFF     gate2723  (.D(g2619), .CP(CLK), .Q(g2625) ) ;
DFF     gate2724  (.D(g2625), .CP(CLK), .Q(g2624) ) ;
INV     gate2725  (.A(II30275), .Z(g23274) ) ;
DFF     gate2726  (.D(g23274), .CP(CLK), .Q(g2628) ) ;
INV     gate2727  (.A(II27029), .Z(g20568) ) ;
DFF     gate2728  (.D(g20568), .CP(CLK), .Q(g2631) ) ;
INV     gate2729  (.A(II27032), .Z(g20569) ) ;
DFF     gate2730  (.D(g20569), .CP(CLK), .Q(g2584) ) ;
INV     gate2731  (.A(II22521), .Z(g16473) ) ;
DFF     gate2732  (.D(g16473), .CP(CLK), .Q(g2587) ) ;
DFF     gate2733  (.D(g2587), .CP(CLK), .Q(g2597) ) ;
DFF     gate2734  (.D(g2597), .CP(CLK), .Q(g2598) ) ;
INV     gate2735  (.A(II18755), .Z(g11593) ) ;
DFF     gate2736  (.D(g11593), .CP(CLK), .Q(g2638) ) ;
DFF     gate2737  (.D(g2638), .CP(CLK), .Q(g2643) ) ;
INV     gate2738  (.A(II18764), .Z(g11596) ) ;
DFF     gate2739  (.D(g11596), .CP(CLK), .Q(g2644) ) ;
DFF     gate2740  (.D(g2644), .CP(CLK), .Q(g2645) ) ;
INV     gate2741  (.A(II18767), .Z(g11597) ) ;
DFF     gate2742  (.D(g11597), .CP(CLK), .Q(g2646) ) ;
DFF     gate2743  (.D(g2646), .CP(CLK), .Q(g2647) ) ;
INV     gate2744  (.A(II18770), .Z(g11598) ) ;
DFF     gate2745  (.D(g11598), .CP(CLK), .Q(g2648) ) ;
DFF     gate2746  (.D(g2648), .CP(CLK), .Q(g2639) ) ;
INV     gate2747  (.A(II18758), .Z(g11594) ) ;
DFF     gate2748  (.D(g11594), .CP(CLK), .Q(g2640) ) ;
DFF     gate2749  (.D(g2640), .CP(CLK), .Q(g2641) ) ;
INV     gate2750  (.A(II18761), .Z(g11595) ) ;
DFF     gate2751  (.D(g11595), .CP(CLK), .Q(g2642) ) ;
DFF     gate2752  (.D(g2642), .CP(CLK), .Q(g2564) ) ;
INV     gate2753  (.A(II20670), .Z(g13457) ) ;
DFF     gate2754  (.D(g13457), .CP(CLK), .Q(g2549) ) ;
DFF     gate2755  (.D(g2549), .CP(CLK), .Q(g2556) ) ;
DFF     gate2756  (.D(g2556), .CP(CLK), .Q(g2560) ) ;
INV     gate2757  (.A(II31919), .Z(g24415) ) ;
DFF     gate2758  (.D(g24415), .CP(CLK), .Q(g2561) ) ;
INV     gate2759  (.A(II31922), .Z(g24416) ) ;
DFF     gate2760  (.D(g24416), .CP(CLK), .Q(g2562) ) ;
INV     gate2761  (.A(II31925), .Z(g24417) ) ;
DFF     gate2762  (.D(g24417), .CP(CLK), .Q(g2563) ) ;
INV     gate2763  (.A(II32994), .Z(g25172) ) ;
DFF     gate2764  (.D(g25172), .CP(CLK), .Q(g2530) ) ;
INV     gate2765  (.A(II32970), .Z(g25164) ) ;
DFF     gate2766  (.D(g25164), .CP(CLK), .Q(g2533) ) ;
INV     gate2767  (.A(II32973), .Z(g25165) ) ;
DFF     gate2768  (.D(g25165), .CP(CLK), .Q(g2536) ) ;
INV     gate2769  (.A(II32985), .Z(g25169) ) ;
DFF     gate2770  (.D(g25169), .CP(CLK), .Q(g2552) ) ;
INV     gate2771  (.A(II32988), .Z(g25170) ) ;
DFF     gate2772  (.D(g25170), .CP(CLK), .Q(g2553) ) ;
INV     gate2773  (.A(II32991), .Z(g25171) ) ;
DFF     gate2774  (.D(g25171), .CP(CLK), .Q(g2554) ) ;
INV     gate2775  (.A(II31910), .Z(g24412) ) ;
DFF     gate2776  (.D(g24412), .CP(CLK), .Q(g2555) ) ;
INV     gate2777  (.A(II31913), .Z(g24413) ) ;
DFF     gate2778  (.D(g24413), .CP(CLK), .Q(g2559) ) ;
INV     gate2779  (.A(II31916), .Z(g24414) ) ;
DFF     gate2780  (.D(g24414), .CP(CLK), .Q(g2539) ) ;
INV     gate2781  (.A(II32976), .Z(g25166) ) ;
DFF     gate2782  (.D(g25166), .CP(CLK), .Q(g2540) ) ;
INV     gate2783  (.A(II32979), .Z(g25167) ) ;
DFF     gate2784  (.D(g25167), .CP(CLK), .Q(g2543) ) ;
INV     gate2785  (.A(II32982), .Z(g25168) ) ;
DFF     gate2786  (.D(g25168), .CP(CLK), .Q(g2546) ) ;
INV     gate2787  (.A(II22524), .Z(g16474) ) ;
DFF     gate2788  (.D(g16474), .CP(CLK), .Q(g2602) ) ;
DFF     gate2789  (.D(g2602), .CP(CLK), .Q(g2609) ) ;
DFF     gate2790  (.D(g2609), .CP(CLK), .Q(g2616) ) ;
INV     gate2791  (.A(II25234), .Z(g19057) ) ;
DFF     gate2792  (.D(g19057), .CP(CLK), .Q(g2617) ) ;
DFF     gate2793  (.D(g2617), .CP(CLK), .Q(g2618) ) ;
INV     gate2794  (.A(II39818), .Z(g30325) ) ;
DFF     gate2795  (.D(g30325), .CP(CLK), .Q(g2622) ) ;
INV     gate2796  (.A(II25237), .Z(g19058) ) ;
DFF     gate2797  (.D(g19058), .CP(CLK), .Q(g2623) ) ;
DFF     gate2798  (.D(g2623), .CP(CLK), .Q(g2574) ) ;
INV     gate2799  (.A(II25240), .Z(g19059) ) ;
DFF     gate2800  (.D(g19059), .CP(CLK), .Q(g2632) ) ;
DFF     gate2801  (.D(g2632), .CP(CLK), .Q(g2633) ) ;
INV     gate2802  (.A(II37140), .Z(g28297) ) ;
DFF     gate2803  (.D(g28297), .CP(CLK), .Q(g2650) ) ;
INV     gate2804  (.A(II37143), .Z(g28298) ) ;
DFF     gate2805  (.D(g28298), .CP(CLK), .Q(g2651) ) ;
INV     gate2806  (.A(II37146), .Z(g28299) ) ;
DFF     gate2807  (.D(g28299), .CP(CLK), .Q(g2649) ) ;
INV     gate2808  (.A(II37149), .Z(g28300) ) ;
DFF     gate2809  (.D(g28300), .CP(CLK), .Q(g2653) ) ;
INV     gate2810  (.A(II37152), .Z(g28301) ) ;
DFF     gate2811  (.D(g28301), .CP(CLK), .Q(g2654) ) ;
INV     gate2812  (.A(II37155), .Z(g28302) ) ;
DFF     gate2813  (.D(g28302), .CP(CLK), .Q(g2652) ) ;
INV     gate2814  (.A(II37158), .Z(g28303) ) ;
DFF     gate2815  (.D(g28303), .CP(CLK), .Q(g2656) ) ;
INV     gate2816  (.A(II37161), .Z(g28304) ) ;
DFF     gate2817  (.D(g28304), .CP(CLK), .Q(g2657) ) ;
INV     gate2818  (.A(II37164), .Z(g28305) ) ;
DFF     gate2819  (.D(g28305), .CP(CLK), .Q(g2655) ) ;
INV     gate2820  (.A(II37167), .Z(g28306) ) ;
DFF     gate2821  (.D(g28306), .CP(CLK), .Q(g2659) ) ;
INV     gate2822  (.A(II37170), .Z(g28307) ) ;
DFF     gate2823  (.D(g28307), .CP(CLK), .Q(g2660) ) ;
INV     gate2824  (.A(II37173), .Z(g28308) ) ;
DFF     gate2825  (.D(g28308), .CP(CLK), .Q(g2658) ) ;
INV     gate2826  (.A(II33888), .Z(g26012) ) ;
DFF     gate2827  (.D(g26012), .CP(CLK), .Q(g2661) ) ;
INV     gate2828  (.A(II33891), .Z(g26013) ) ;
DFF     gate2829  (.D(g26013), .CP(CLK), .Q(g2664) ) ;
INV     gate2830  (.A(II33894), .Z(g26014) ) ;
DFF     gate2831  (.D(g26014), .CP(CLK), .Q(g2667) ) ;
INV     gate2832  (.A(II33897), .Z(g26015) ) ;
DFF     gate2833  (.D(g26015), .CP(CLK), .Q(g2670) ) ;
INV     gate2834  (.A(II33900), .Z(g26016) ) ;
DFF     gate2835  (.D(g26016), .CP(CLK), .Q(g2673) ) ;
INV     gate2836  (.A(II33903), .Z(g26017) ) ;
DFF     gate2837  (.D(g26017), .CP(CLK), .Q(g2676) ) ;
INV     gate2838  (.A(II38220), .Z(g29159) ) ;
DFF     gate2839  (.D(g29159), .CP(CLK), .Q(g2688) ) ;
INV     gate2840  (.A(II38223), .Z(g29160) ) ;
DFF     gate2841  (.D(g29160), .CP(CLK), .Q(g2691) ) ;
INV     gate2842  (.A(II38226), .Z(g29161) ) ;
DFF     gate2843  (.D(g29161), .CP(CLK), .Q(g2694) ) ;
INV     gate2844  (.A(II38211), .Z(g29156) ) ;
DFF     gate2845  (.D(g29156), .CP(CLK), .Q(g2679) ) ;
INV     gate2846  (.A(II38214), .Z(g29157) ) ;
DFF     gate2847  (.D(g29157), .CP(CLK), .Q(g2682) ) ;
INV     gate2848  (.A(II38217), .Z(g29158) ) ;
DFF     gate2849  (.D(g29158), .CP(CLK), .Q(g2685) ) ;
INV     gate2850  (.A(II35536), .Z(g27233) ) ;
DFF     gate2851  (.D(g27233), .CP(CLK), .Q(g2565) ) ;
INV     gate2852  (.A(II35539), .Z(g27234) ) ;
DFF     gate2853  (.D(g27234), .CP(CLK), .Q(g2568) ) ;
INV     gate2854  (.A(II35542), .Z(g27235) ) ;
DFF     gate2855  (.D(g27235), .CP(CLK), .Q(g2571) ) ;
INV     gate2856  (.A(II15517), .Z(g8311) ) ;
DFF     gate2857  (.D(g8311), .CP(CLK), .Q(g2580) ) ;
INV     gate2858  (.A(II31928), .Z(g24418) ) ;
DFF     gate2859  (.D(g24418), .CP(CLK), .Q(g2581) ) ;
INV     gate2860  (.A(II25222), .Z(g19053) ) ;
DFF     gate2861  (.D(g19053), .CP(CLK), .Q(g2582) ) ;
INV     gate2862  (.A(II25225), .Z(g19054) ) ;
DFF     gate2863  (.D(g19054), .CP(CLK), .Q(g2583) ) ;
INV     gate2864  (.A(II25228), .Z(g19055) ) ;
DFF     gate2865  (.D(g19055), .CP(CLK), .Q(g2588) ) ;
INV     gate2866  (.A(II25231), .Z(g19056) ) ;
DFF     gate2867  (.D(g19056), .CP(CLK), .Q(g2589) ) ;
INV     gate2868  (.A(II39815), .Z(g30324) ) ;
DFF     gate2869  (.D(g30324), .CP(CLK), .Q(g2590) ) ;
INV     gate2870  (.A(II39812), .Z(g30323) ) ;
DFF     gate2871  (.D(g30323), .CP(CLK), .Q(g2591) ) ;
INV     gate2872  (.A(II39809), .Z(g30322) ) ;
DFF     gate2873  (.D(g30322), .CP(CLK), .Q(g2592) ) ;
INV     gate2874  (.A(II39806), .Z(g30321) ) ;
DFF     gate2875  (.D(g30321), .CP(CLK), .Q(g2593) ) ;
INV     gate2876  (.A(II39803), .Z(g30320) ) ;
DFF     gate2877  (.D(g30320), .CP(CLK), .Q(g2594) ) ;
DFF     gate2878  (.D(g2594), .CP(CLK), .Q(g2599) ) ;
INV     gate2879  (.A(II20673), .Z(g13458) ) ;
DFF     gate2880  (.D(g13458), .CP(CLK), .Q(g2603) ) ;
INV     gate2881  (.A(II20676), .Z(g13459) ) ;
DFF     gate2882  (.D(g13459), .CP(CLK), .Q(g2604) ) ;
INV     gate2883  (.A(II20679), .Z(g13460) ) ;
DFF     gate2884  (.D(g13460), .CP(CLK), .Q(g2605) ) ;
INV     gate2885  (.A(II20682), .Z(g13461) ) ;
DFF     gate2886  (.D(g13461), .CP(CLK), .Q(g2606) ) ;
INV     gate2887  (.A(II20685), .Z(g13462) ) ;
DFF     gate2888  (.D(g13462), .CP(CLK), .Q(g2607) ) ;
INV     gate2889  (.A(II20688), .Z(g13463) ) ;
DFF     gate2890  (.D(g13463), .CP(CLK), .Q(g2608) ) ;
INV     gate2891  (.A(II20691), .Z(g13464) ) ;
DFF     gate2892  (.D(g13464), .CP(CLK), .Q(g2610) ) ;
INV     gate2893  (.A(II20694), .Z(g13465) ) ;
DFF     gate2894  (.D(g13465), .CP(CLK), .Q(g2611) ) ;
INV     gate2895  (.A(II33885), .Z(g26011) ) ;
DFF     gate2896  (.D(g26011), .CP(CLK), .Q(g2612) ) ;
INV     gate2897  (.A(II20697), .Z(g13466) ) ;
DFF     gate2898  (.D(g13466), .CP(CLK), .Q(g2615) ) ;
INV     gate2899  (.A(II20703), .Z(g13468) ) ;
DFF     gate2900  (.D(g13468), .CP(CLK), .Q(g2697) ) ;
DFF     gate2901  (.D(g2697), .CP(CLK), .Q(g2700) ) ;
DFF     gate2902  (.D(g2700), .CP(CLK), .Q(g2703) ) ;
INV     gate2903  (.A(II27035), .Z(g20570) ) ;
DFF     gate2904  (.D(g20570), .CP(CLK), .Q(g2704) ) ;
INV     gate2905  (.A(II28464), .Z(g21946) ) ;
DFF     gate2906  (.D(g21946), .CP(CLK), .Q(g2733) ) ;
INV     gate2907  (.A(II30278), .Z(g23275) ) ;
DFF     gate2908  (.D(g23275), .CP(CLK), .Q(g2714) ) ;
INV     gate2909  (.A(II31931), .Z(g24419) ) ;
DFF     gate2910  (.D(g24419), .CP(CLK), .Q(g2707) ) ;
INV     gate2911  (.A(II32997), .Z(g25173) ) ;
DFF     gate2912  (.D(g25173), .CP(CLK), .Q(g2727) ) ;
INV     gate2913  (.A(II33906), .Z(g26018) ) ;
DFF     gate2914  (.D(g26018), .CP(CLK), .Q(g2720) ) ;
INV     gate2915  (.A(II34833), .Z(g26742) ) ;
DFF     gate2916  (.D(g26742), .CP(CLK), .Q(g2734) ) ;
INV     gate2917  (.A(II35545), .Z(g27236) ) ;
DFF     gate2918  (.D(g27236), .CP(CLK), .Q(g2746) ) ;
INV     gate2919  (.A(II36153), .Z(g27714) ) ;
DFF     gate2920  (.D(g27714), .CP(CLK), .Q(g2740) ) ;
INV     gate2921  (.A(II37176), .Z(g28309) ) ;
DFF     gate2922  (.D(g28309), .CP(CLK), .Q(g2753) ) ;
INV     gate2923  (.A(II37623), .Z(g28692) ) ;
DFF     gate2924  (.D(g28692), .CP(CLK), .Q(g2760) ) ;
INV     gate2925  (.A(II38229), .Z(g29162) ) ;
DFF     gate2926  (.D(g29162), .CP(CLK), .Q(g2766) ) ;
INV     gate2927  (.A(II30281), .Z(g23276) ) ;
DFF     gate2928  (.D(g23276), .CP(CLK), .Q(g2773) ) ;
INV     gate2929  (.A(II30284), .Z(g23277) ) ;
DFF     gate2930  (.D(g23277), .CP(CLK), .Q(g2774) ) ;
INV     gate2931  (.A(II30287), .Z(g23278) ) ;
DFF     gate2932  (.D(g23278), .CP(CLK), .Q(g2772) ) ;
INV     gate2933  (.A(II30290), .Z(g23279) ) ;
DFF     gate2934  (.D(g23279), .CP(CLK), .Q(g2776) ) ;
INV     gate2935  (.A(II30293), .Z(g23280) ) ;
DFF     gate2936  (.D(g23280), .CP(CLK), .Q(g2777) ) ;
INV     gate2937  (.A(II30296), .Z(g23281) ) ;
DFF     gate2938  (.D(g23281), .CP(CLK), .Q(g2775) ) ;
INV     gate2939  (.A(II30299), .Z(g23282) ) ;
DFF     gate2940  (.D(g23282), .CP(CLK), .Q(g2779) ) ;
INV     gate2941  (.A(II30302), .Z(g23283) ) ;
DFF     gate2942  (.D(g23283), .CP(CLK), .Q(g2780) ) ;
INV     gate2943  (.A(II30305), .Z(g23284) ) ;
DFF     gate2944  (.D(g23284), .CP(CLK), .Q(g2778) ) ;
INV     gate2945  (.A(II30308), .Z(g23285) ) ;
DFF     gate2946  (.D(g23285), .CP(CLK), .Q(g2782) ) ;
INV     gate2947  (.A(II30311), .Z(g23286) ) ;
DFF     gate2948  (.D(g23286), .CP(CLK), .Q(g2783) ) ;
INV     gate2949  (.A(II30314), .Z(g23287) ) ;
DFF     gate2950  (.D(g23287), .CP(CLK), .Q(g2781) ) ;
INV     gate2951  (.A(II30317), .Z(g23288) ) ;
DFF     gate2952  (.D(g23288), .CP(CLK), .Q(g2785) ) ;
INV     gate2953  (.A(II30320), .Z(g23289) ) ;
DFF     gate2954  (.D(g23289), .CP(CLK), .Q(g2786) ) ;
INV     gate2955  (.A(II30323), .Z(g23290) ) ;
DFF     gate2956  (.D(g23290), .CP(CLK), .Q(g2784) ) ;
INV     gate2957  (.A(II30326), .Z(g23291) ) ;
DFF     gate2958  (.D(g23291), .CP(CLK), .Q(g2788) ) ;
INV     gate2959  (.A(II30329), .Z(g23292) ) ;
DFF     gate2960  (.D(g23292), .CP(CLK), .Q(g2789) ) ;
INV     gate2961  (.A(II30332), .Z(g23293) ) ;
DFF     gate2962  (.D(g23293), .CP(CLK), .Q(g2787) ) ;
INV     gate2963  (.A(II30335), .Z(g23294) ) ;
DFF     gate2964  (.D(g23294), .CP(CLK), .Q(g2791) ) ;
INV     gate2965  (.A(II30338), .Z(g23295) ) ;
DFF     gate2966  (.D(g23295), .CP(CLK), .Q(g2792) ) ;
INV     gate2967  (.A(II30341), .Z(g23296) ) ;
DFF     gate2968  (.D(g23296), .CP(CLK), .Q(g2790) ) ;
INV     gate2969  (.A(II30344), .Z(g23297) ) ;
DFF     gate2970  (.D(g23297), .CP(CLK), .Q(g2794) ) ;
INV     gate2971  (.A(II30347), .Z(g23298) ) ;
DFF     gate2972  (.D(g23298), .CP(CLK), .Q(g2795) ) ;
INV     gate2973  (.A(II30350), .Z(g23299) ) ;
DFF     gate2974  (.D(g23299), .CP(CLK), .Q(g2793) ) ;
INV     gate2975  (.A(II30353), .Z(g23300) ) ;
DFF     gate2976  (.D(g23300), .CP(CLK), .Q(g2797) ) ;
INV     gate2977  (.A(II30356), .Z(g23301) ) ;
DFF     gate2978  (.D(g23301), .CP(CLK), .Q(g2798) ) ;
INV     gate2979  (.A(II30359), .Z(g23302) ) ;
DFF     gate2980  (.D(g23302), .CP(CLK), .Q(g2796) ) ;
INV     gate2981  (.A(II30362), .Z(g23303) ) ;
DFF     gate2982  (.D(g23303), .CP(CLK), .Q(g2800) ) ;
INV     gate2983  (.A(II30365), .Z(g23304) ) ;
DFF     gate2984  (.D(g23304), .CP(CLK), .Q(g2801) ) ;
INV     gate2985  (.A(II30368), .Z(g23305) ) ;
DFF     gate2986  (.D(g23305), .CP(CLK), .Q(g2799) ) ;
INV     gate2987  (.A(II30371), .Z(g23306) ) ;
DFF     gate2988  (.D(g23306), .CP(CLK), .Q(g2803) ) ;
INV     gate2989  (.A(II30374), .Z(g23307) ) ;
DFF     gate2990  (.D(g23307), .CP(CLK), .Q(g2804) ) ;
INV     gate2991  (.A(II30377), .Z(g23308) ) ;
DFF     gate2992  (.D(g23308), .CP(CLK), .Q(g2802) ) ;
INV     gate2993  (.A(II30380), .Z(g23309) ) ;
DFF     gate2994  (.D(g23309), .CP(CLK), .Q(g2806) ) ;
INV     gate2995  (.A(II30383), .Z(g23310) ) ;
DFF     gate2996  (.D(g23310), .CP(CLK), .Q(g2807) ) ;
INV     gate2997  (.A(II30386), .Z(g23311) ) ;
DFF     gate2998  (.D(g23311), .CP(CLK), .Q(g2805) ) ;
INV     gate2999  (.A(II34836), .Z(g26743) ) ;
DFF     gate3000  (.D(g26743), .CP(CLK), .Q(g2809) ) ;
INV     gate3001  (.A(II34839), .Z(g26744) ) ;
DFF     gate3002  (.D(g26744), .CP(CLK), .Q(g2810) ) ;
INV     gate3003  (.A(II34842), .Z(g26745) ) ;
DFF     gate3004  (.D(g26745), .CP(CLK), .Q(g2808) ) ;
INV     gate3005  (.A(II31934), .Z(g24420) ) ;
DFF     gate3006  (.D(g24420), .CP(CLK), .Q(g2812) ) ;
INV     gate3007  (.A(II31937), .Z(g24421) ) ;
DFF     gate3008  (.D(g24421), .CP(CLK), .Q(g2813) ) ;
INV     gate3009  (.A(II31940), .Z(g24422) ) ;
DFF     gate3010  (.D(g24422), .CP(CLK), .Q(g2811) ) ;
INV     gate3011  (.A(II30404), .Z(g23317) ) ;
DFF     gate3012  (.D(g23317), .CP(CLK), .Q(g3054) ) ;
INV     gate3013  (.A(II30407), .Z(g23318) ) ;
DFF     gate3014  (.D(g23318), .CP(CLK), .Q(g3079) ) ;
INV     gate3015  (.A(II28521), .Z(g21965) ) ;
DFF     gate3016  (.D(g21965), .CP(CLK), .Q(g3080) ) ;
INV     gate3017  (.A(II38740), .Z(g29453) ) ;
DFF     gate3018  (.D(g29453), .CP(CLK), .Q(g3043) ) ;
INV     gate3019  (.A(II38743), .Z(g29454) ) ;
DFF     gate3020  (.D(g29454), .CP(CLK), .Q(g3044) ) ;
INV     gate3021  (.A(II38746), .Z(g29455) ) ;
DFF     gate3022  (.D(g29455), .CP(CLK), .Q(g3045) ) ;
INV     gate3023  (.A(II38749), .Z(g29456) ) ;
DFF     gate3024  (.D(g29456), .CP(CLK), .Q(g3046) ) ;
INV     gate3025  (.A(II38752), .Z(g29457) ) ;
DFF     gate3026  (.D(g29457), .CP(CLK), .Q(g3047) ) ;
INV     gate3027  (.A(II38755), .Z(g29458) ) ;
DFF     gate3028  (.D(g29458), .CP(CLK), .Q(g3048) ) ;
INV     gate3029  (.A(II38758), .Z(g29459) ) ;
DFF     gate3030  (.D(g29459), .CP(CLK), .Q(g3049) ) ;
INV     gate3031  (.A(II38761), .Z(g29460) ) ;
DFF     gate3032  (.D(g29460), .CP(CLK), .Q(g3050) ) ;
INV     gate3033  (.A(II39083), .Z(g29655) ) ;
DFF     gate3034  (.D(g29655), .CP(CLK), .Q(g3051) ) ;
INV     gate3035  (.A(II39454), .Z(g29972) ) ;
DFF     gate3036  (.D(g29972), .CP(CLK), .Q(g3052) ) ;
INV     gate3037  (.A(II39457), .Z(g29973) ) ;
DFF     gate3038  (.D(g29973), .CP(CLK), .Q(g3053) ) ;
INV     gate3039  (.A(II39460), .Z(g29974) ) ;
DFF     gate3040  (.D(g29974), .CP(CLK), .Q(g3055) ) ;
INV     gate3041  (.A(II39463), .Z(g29975) ) ;
DFF     gate3042  (.D(g29975), .CP(CLK), .Q(g3056) ) ;
INV     gate3043  (.A(II39466), .Z(g29976) ) ;
DFF     gate3044  (.D(g29976), .CP(CLK), .Q(g3057) ) ;
INV     gate3045  (.A(II39469), .Z(g29977) ) ;
DFF     gate3046  (.D(g29977), .CP(CLK), .Q(g3058) ) ;
INV     gate3047  (.A(II39472), .Z(g29978) ) ;
DFF     gate3048  (.D(g29978), .CP(CLK), .Q(g3059) ) ;
INV     gate3049  (.A(II39475), .Z(g29979) ) ;
DFF     gate3050  (.D(g29979), .CP(CLK), .Q(g3060) ) ;
INV     gate3051  (.A(II39622), .Z(g30119) ) ;
DFF     gate3052  (.D(g30119), .CP(CLK), .Q(g3061) ) ;
INV     gate3053  (.A(II40976), .Z(g30908) ) ;
DFF     gate3054  (.D(g30908), .CP(CLK), .Q(g3062) ) ;
INV     gate3055  (.A(II40979), .Z(g30909) ) ;
DFF     gate3056  (.D(g30909), .CP(CLK), .Q(g3063) ) ;
INV     gate3057  (.A(II40982), .Z(g30910) ) ;
DFF     gate3058  (.D(g30910), .CP(CLK), .Q(g3064) ) ;
INV     gate3059  (.A(II40985), .Z(g30911) ) ;
DFF     gate3060  (.D(g30911), .CP(CLK), .Q(g3065) ) ;
INV     gate3061  (.A(II40988), .Z(g30912) ) ;
DFF     gate3062  (.D(g30912), .CP(CLK), .Q(g3066) ) ;
INV     gate3063  (.A(II40991), .Z(g30913) ) ;
DFF     gate3064  (.D(g30913), .CP(CLK), .Q(g3067) ) ;
INV     gate3065  (.A(II40994), .Z(g30914) ) ;
DFF     gate3066  (.D(g30914), .CP(CLK), .Q(g3068) ) ;
INV     gate3067  (.A(II40997), .Z(g30915) ) ;
DFF     gate3068  (.D(g30915), .CP(CLK), .Q(g3069) ) ;
INV     gate3069  (.A(II41044), .Z(g30940) ) ;
DFF     gate3070  (.D(g30940), .CP(CLK), .Q(g3070) ) ;
INV     gate3071  (.A(II41114), .Z(g30980) ) ;
DFF     gate3072  (.D(g30980), .CP(CLK), .Q(g3071) ) ;
INV     gate3073  (.A(II41117), .Z(g30981) ) ;
DFF     gate3074  (.D(g30981), .CP(CLK), .Q(g3072) ) ;
INV     gate3075  (.A(II41120), .Z(g30982) ) ;
DFF     gate3076  (.D(g30982), .CP(CLK), .Q(g3073) ) ;
INV     gate3077  (.A(II41123), .Z(g30983) ) ;
DFF     gate3078  (.D(g30983), .CP(CLK), .Q(g3074) ) ;
INV     gate3079  (.A(II41126), .Z(g30984) ) ;
DFF     gate3080  (.D(g30984), .CP(CLK), .Q(g3075) ) ;
INV     gate3081  (.A(II41129), .Z(g30985) ) ;
DFF     gate3082  (.D(g30985), .CP(CLK), .Q(g3076) ) ;
INV     gate3083  (.A(II41132), .Z(g30986) ) ;
DFF     gate3084  (.D(g30986), .CP(CLK), .Q(g3077) ) ;
INV     gate3085  (.A(II41135), .Z(g30987) ) ;
DFF     gate3086  (.D(g30987), .CP(CLK), .Q(g3078) ) ;
INV     gate3087  (.A(II41141), .Z(g30989) ) ;
DFF     gate3088  (.D(g30989), .CP(CLK), .Q(g2997) ) ;
INV     gate3089  (.A(II34851), .Z(g26748) ) ;
DFF     gate3090  (.D(g26748), .CP(CLK), .Q(g2993) ) ;
INV     gate3091  (.A(II35551), .Z(g27238) ) ;
DFF     gate3092  (.D(g27238), .CP(CLK), .Q(g2998) ) ;
INV     gate3093  (.A(II33009), .Z(g25177) ) ;
DFF     gate3094  (.D(g25177), .CP(CLK), .Q(g3006) ) ;
INV     gate3095  (.A(II33915), .Z(g26021) ) ;
DFF     gate3096  (.D(g26021), .CP(CLK), .Q(g3002) ) ;
INV     gate3097  (.A(II34857), .Z(g26750) ) ;
DFF     gate3098  (.D(g26750), .CP(CLK), .Q(g3013) ) ;
INV     gate3099  (.A(II35554), .Z(g27239) ) ;
DFF     gate3100  (.D(g27239), .CP(CLK), .Q(g3010) ) ;
INV     gate3101  (.A(II36159), .Z(g27716) ) ;
DFF     gate3102  (.D(g27716), .CP(CLK), .Q(g3024) ) ;
INV     gate3103  (.A(II31949), .Z(g24425) ) ;
DFF     gate3104  (.D(g24425), .CP(CLK), .Q(g3018) ) ;
INV     gate3105  (.A(II33006), .Z(g25176) ) ;
DFF     gate3106  (.D(g25176), .CP(CLK), .Q(g3028) ) ;
INV     gate3107  (.A(II33918), .Z(g26022) ) ;
DFF     gate3108  (.D(g26022), .CP(CLK), .Q(g3036) ) ;
INV     gate3109  (.A(II34854), .Z(g26749) ) ;
DFF     gate3110  (.D(g26749), .CP(CLK), .Q(g3032) ) ;
INV     gate3111  (.A(II22593), .Z(g16497) ) ;
DFF     gate3112  (.D(g16497), .CP(CLK), .Q(g3040) ) ;
DFF     gate3113  (.D(g3040), .CP(CLK), .Q(g2986) ) ;
INV     gate3114  (.A(II22587), .Z(g16495) ) ;
DFF     gate3115  (.D(g16495), .CP(CLK), .Q(g2987) ) ;
INV     gate3116  (.A(II27110), .Z(g20595) ) ;
DFF     gate3117  (.D(g20595), .CP(CLK), .Q(g48) ) ;
INV     gate3118  (.A(II27113), .Z(g20596) ) ;
DFF     gate3119  (.D(g20596), .CP(CLK), .Q(g45) ) ;
INV     gate3120  (.A(II27116), .Z(g20597) ) ;
DFF     gate3121  (.D(g20597), .CP(CLK), .Q(g42) ) ;
INV     gate3122  (.A(II27119), .Z(g20598) ) ;
DFF     gate3123  (.D(g20598), .CP(CLK), .Q(g39) ) ;
INV     gate3124  (.A(II27122), .Z(g20599) ) ;
DFF     gate3125  (.D(g20599), .CP(CLK), .Q(g27) ) ;
INV     gate3126  (.A(II27125), .Z(g20600) ) ;
DFF     gate3127  (.D(g20600), .CP(CLK), .Q(g30) ) ;
INV     gate3128  (.A(II27128), .Z(g20601) ) ;
DFF     gate3129  (.D(g20601), .CP(CLK), .Q(g33) ) ;
INV     gate3130  (.A(II27131), .Z(g20602) ) ;
DFF     gate3131  (.D(g20602), .CP(CLK), .Q(g36) ) ;
INV     gate3132  (.A(II27134), .Z(g20603) ) ;
DFF     gate3133  (.D(g20603), .CP(CLK), .Q(g3083) ) ;
INV     gate3134  (.A(II27137), .Z(g20604) ) ;
DFF     gate3135  (.D(g20604), .CP(CLK), .Q(g26) ) ;
INV     gate3136  (.A(II28524), .Z(g21966) ) ;
DFF     gate3137  (.D(g21966), .CP(CLK), .Q(g2992) ) ;
INV     gate3138  (.A(II27140), .Z(g20605) ) ;
DFF     gate3139  (.D(g20605), .CP(CLK), .Q(g23) ) ;
INV     gate3140  (.A(II27143), .Z(g20606) ) ;
DFF     gate3141  (.D(g20606), .CP(CLK), .Q(g20) ) ;
INV     gate3142  (.A(II27146), .Z(g20607) ) ;
DFF     gate3143  (.D(g20607), .CP(CLK), .Q(g17) ) ;
INV     gate3144  (.A(II27149), .Z(g20608) ) ;
DFF     gate3145  (.D(g20608), .CP(CLK), .Q(g11) ) ;
INV     gate3146  (.A(II27092), .Z(g20589) ) ;
DFF     gate3147  (.D(g20589), .CP(CLK), .Q(g14) ) ;
INV     gate3148  (.A(II27095), .Z(g20590) ) ;
DFF     gate3149  (.D(g20590), .CP(CLK), .Q(g5) ) ;
INV     gate3150  (.A(II27098), .Z(g20591) ) ;
DFF     gate3151  (.D(g20591), .CP(CLK), .Q(g8) ) ;
INV     gate3152  (.A(II27101), .Z(g20592) ) ;
DFF     gate3153  (.D(g20592), .CP(CLK), .Q(g2) ) ;
INV     gate3154  (.A(II27104), .Z(g20593) ) ;
DFF     gate3155  (.D(g20593), .CP(CLK), .Q(g2990) ) ;
INV     gate3156  (.A(II28518), .Z(g21964) ) ;
DFF     gate3157  (.D(g21964), .CP(CLK), .Q(g2991) ) ;
INV     gate3158  (.A(II27107), .Z(g20594) ) ;
DFF     gate3159  (.D(g20594), .CP(CLK), .Q(g1) ) ;
INV     gate3160  (.A(g563), .Z(II13089) ) ;
INV     gate3161  (.A(II13089), .Z(g562) ) ;
INV     gate3162  (.A(g1249), .Z(II13092) ) ;
INV     gate3163  (.A(II13092), .Z(g1248) ) ;
INV     gate3164  (.A(g1943), .Z(II13095) ) ;
INV     gate3165  (.A(II13095), .Z(g1942) ) ;
INV     gate3166  (.A(g2637), .Z(II13098) ) ;
INV     gate3167  (.A(II13098), .Z(g2636) ) ;
INV     gate3168  (.A(g1), .Z(II13101) ) ;
INV     gate3169  (.A(II13101), .Z(g3235) ) ;
INV     gate3170  (.A(g2), .Z(II13104) ) ;
INV     gate3171  (.A(II13104), .Z(g3236) ) ;
INV     gate3172  (.A(g5), .Z(II13107) ) ;
INV     gate3173  (.A(II13107), .Z(g3237) ) ;
INV     gate3174  (.A(g8), .Z(II13110) ) ;
INV     gate3175  (.A(II13110), .Z(g3238) ) ;
INV     gate3176  (.A(g11), .Z(II13113) ) ;
INV     gate3177  (.A(II13113), .Z(g3239) ) ;
INV     gate3178  (.A(g14), .Z(II13116) ) ;
INV     gate3179  (.A(II13116), .Z(g3240) ) ;
INV     gate3180  (.A(g17), .Z(II13119) ) ;
INV     gate3181  (.A(II13119), .Z(g3241) ) ;
INV     gate3182  (.A(g20), .Z(II13122) ) ;
INV     gate3183  (.A(II13122), .Z(g3242) ) ;
INV     gate3184  (.A(g23), .Z(II13125) ) ;
INV     gate3185  (.A(II13125), .Z(g3243) ) ;
INV     gate3186  (.A(g26), .Z(II13128) ) ;
INV     gate3187  (.A(II13128), .Z(g3244) ) ;
INV     gate3188  (.A(g27), .Z(II13131) ) ;
INV     gate3189  (.A(II13131), .Z(g3245) ) ;
INV     gate3190  (.A(g30), .Z(II13134) ) ;
INV     gate3191  (.A(II13134), .Z(g3246) ) ;
INV     gate3192  (.A(g33), .Z(II13137) ) ;
INV     gate3193  (.A(II13137), .Z(g3247) ) ;
INV     gate3194  (.A(g36), .Z(II13140) ) ;
INV     gate3195  (.A(II13140), .Z(g3248) ) ;
INV     gate3196  (.A(g39), .Z(II13143) ) ;
INV     gate3197  (.A(II13143), .Z(g3249) ) ;
INV     gate3198  (.A(g42), .Z(II13146) ) ;
INV     gate3199  (.A(II13146), .Z(g3250) ) ;
INV     gate3200  (.A(g45), .Z(II13149) ) ;
INV     gate3201  (.A(II13149), .Z(g3251) ) ;
INV     gate3202  (.A(g48), .Z(II13152) ) ;
INV     gate3203  (.A(II13152), .Z(g3252) ) ;
INV     gate3204  (.A(g51), .Z(II13155) ) ;
INV     gate3205  (.A(II13155), .Z(g3253) ) ;
INV     gate3206  (.A(g165), .Z(II13158) ) ;
INV     gate3207  (.A(II13158), .Z(g3254) ) ;
INV     gate3208  (.A(g308), .Z(II13161) ) ;
INV     gate3209  (.A(II13161), .Z(g3304) ) ;
INV     gate3210  (.A(g305), .Z(g3305) ) ;
INV     gate3211  (.A(g401), .Z(II13165) ) ;
INV     gate3212  (.A(II13165), .Z(g3306) ) ;
INV     gate3213  (.A(g309), .Z(g3337) ) ;
INV     gate3214  (.A(g550), .Z(II13169) ) ;
INV     gate3215  (.A(II13169), .Z(g3338) ) ;
INV     gate3216  (.A(g499), .Z(g3365) ) ;
INV     gate3217  (.A(g629), .Z(II13173) ) ;
INV     gate3218  (.A(II13173), .Z(g3366) ) ;
INV     gate3219  (.A(g630), .Z(II13176) ) ;
INV     gate3220  (.A(II13176), .Z(g3398) ) ;
INV     gate3221  (.A(g853), .Z(II13179) ) ;
INV     gate3222  (.A(II13179), .Z(g3410) ) ;
INV     gate3223  (.A(g995), .Z(II13182) ) ;
INV     gate3224  (.A(II13182), .Z(g3460) ) ;
INV     gate3225  (.A(g992), .Z(g3461) ) ;
INV     gate3226  (.A(g1088), .Z(II13186) ) ;
INV     gate3227  (.A(II13186), .Z(g3462) ) ;
INV     gate3228  (.A(g996), .Z(g3493) ) ;
INV     gate3229  (.A(g1236), .Z(II13190) ) ;
INV     gate3230  (.A(II13190), .Z(g3494) ) ;
INV     gate3231  (.A(g1186), .Z(g3521) ) ;
INV     gate3232  (.A(g1315), .Z(II13194) ) ;
INV     gate3233  (.A(II13194), .Z(g3522) ) ;
INV     gate3234  (.A(g1316), .Z(II13197) ) ;
INV     gate3235  (.A(II13197), .Z(g3554) ) ;
INV     gate3236  (.A(g1547), .Z(II13200) ) ;
INV     gate3237  (.A(II13200), .Z(g3566) ) ;
INV     gate3238  (.A(g1689), .Z(II13203) ) ;
INV     gate3239  (.A(II13203), .Z(g3616) ) ;
INV     gate3240  (.A(g1686), .Z(g3617) ) ;
INV     gate3241  (.A(g1782), .Z(II13207) ) ;
INV     gate3242  (.A(II13207), .Z(g3618) ) ;
INV     gate3243  (.A(g1690), .Z(g3649) ) ;
INV     gate3244  (.A(g1930), .Z(II13211) ) ;
INV     gate3245  (.A(II13211), .Z(g3650) ) ;
INV     gate3246  (.A(g1880), .Z(g3677) ) ;
INV     gate3247  (.A(g2009), .Z(II13215) ) ;
INV     gate3248  (.A(II13215), .Z(g3678) ) ;
INV     gate3249  (.A(g2010), .Z(II13218) ) ;
INV     gate3250  (.A(II13218), .Z(g3710) ) ;
INV     gate3251  (.A(g2241), .Z(II13221) ) ;
INV     gate3252  (.A(II13221), .Z(g3722) ) ;
INV     gate3253  (.A(g2383), .Z(II13224) ) ;
INV     gate3254  (.A(II13224), .Z(g3772) ) ;
INV     gate3255  (.A(g2380), .Z(g3773) ) ;
INV     gate3256  (.A(g2476), .Z(II13228) ) ;
INV     gate3257  (.A(II13228), .Z(g3774) ) ;
INV     gate3258  (.A(g2384), .Z(g3805) ) ;
INV     gate3259  (.A(g2624), .Z(II13232) ) ;
INV     gate3260  (.A(II13232), .Z(g3806) ) ;
INV     gate3261  (.A(g2574), .Z(g3833) ) ;
INV     gate3262  (.A(g2703), .Z(II13236) ) ;
INV     gate3263  (.A(II13236), .Z(g3834) ) ;
INV     gate3264  (.A(g2704), .Z(II13239) ) ;
INV     gate3265  (.A(II13239), .Z(g3866) ) ;
INV     gate3266  (.A(g2879), .Z(II13242) ) ;
INV     gate3267  (.A(II13242), .Z(g3878) ) ;
INV     gate3268  (.A(g2950), .Z(g3897) ) ;
INV     gate3269  (.A(g2987), .Z(II13246) ) ;
INV     gate3270  (.A(II13246), .Z(g3900) ) ;
INV     gate3271  (.A(g3080), .Z(g3919) ) ;
INV     gate3272  (.A(g150), .Z(g3922) ) ;
INV     gate3273  (.A(g155), .Z(g3925) ) ;
INV     gate3274  (.A(g157), .Z(g3928) ) ;
INV     gate3275  (.A(g171), .Z(g3931) ) ;
INV     gate3276  (.A(g176), .Z(g3934) ) ;
INV     gate3277  (.A(g178), .Z(g3937) ) ;
INV     gate3278  (.A(g408), .Z(g3940) ) ;
INV     gate3279  (.A(g455), .Z(g3941) ) ;
INV     gate3280  (.A(g699), .Z(g3942) ) ;
INV     gate3281  (.A(g726), .Z(g3945) ) ;
INV     gate3282  (.A(g835), .Z(g3948) ) ;
INV     gate3283  (.A(g840), .Z(g3951) ) ;
INV     gate3284  (.A(g842), .Z(g3954) ) ;
INV     gate3285  (.A(g856), .Z(g3957) ) ;
INV     gate3286  (.A(g861), .Z(g3960) ) ;
INV     gate3287  (.A(g863), .Z(g3963) ) ;
INV     gate3288  (.A(g1526), .Z(g3966) ) ;
INV     gate3289  (.A(g1531), .Z(g3969) ) ;
INV     gate3290  (.A(g1533), .Z(g3972) ) ;
INV     gate3291  (.A(g1552), .Z(g3975) ) ;
INV     gate3292  (.A(g1554), .Z(g3978) ) ;
INV     gate3293  (.A(g2217), .Z(g3981) ) ;
INV     gate3294  (.A(g2222), .Z(g3984) ) ;
INV     gate3295  (.A(g2224), .Z(g3987) ) ;
INV     gate3296  (.A(g2245), .Z(g3990) ) ;
INV     gate3297  (.A(g2848), .Z(II13275) ) ;
INV     gate3298  (.A(g2848), .Z(g3994) ) ;
INV     gate3299  (.A(g3064), .Z(g3995) ) ;
INV     gate3300  (.A(g3073), .Z(g3996) ) ;
INV     gate3301  (.A(g45), .Z(g3997) ) ;
INV     gate3302  (.A(g23), .Z(g3998) ) ;
INV     gate3303  (.A(g3204), .Z(g3999) ) ;
INV     gate3304  (.A(g153), .Z(g4000) ) ;
INV     gate3305  (.A(g158), .Z(g4003) ) ;
INV     gate3306  (.A(g160), .Z(g4006) ) ;
INV     gate3307  (.A(g174), .Z(g4009) ) ;
INV     gate3308  (.A(g179), .Z(g4012) ) ;
INV     gate3309  (.A(g411), .Z(g4015) ) ;
INV     gate3310  (.A(g417), .Z(g4016) ) ;
INV     gate3311  (.A(g427), .Z(g4017) ) ;
INV     gate3312  (.A(g700), .Z(g4020) ) ;
INV     gate3313  (.A(g702), .Z(g4023) ) ;
INV     gate3314  (.A(g727), .Z(g4026) ) ;
INV     gate3315  (.A(g838), .Z(g4029) ) ;
INV     gate3316  (.A(g843), .Z(g4032) ) ;
INV     gate3317  (.A(g845), .Z(g4035) ) ;
INV     gate3318  (.A(g859), .Z(g4038) ) ;
INV     gate3319  (.A(g864), .Z(g4041) ) ;
INV     gate3320  (.A(g866), .Z(g4044) ) ;
INV     gate3321  (.A(g1095), .Z(g4047) ) ;
INV     gate3322  (.A(g1142), .Z(g4048) ) ;
INV     gate3323  (.A(g1385), .Z(g4049) ) ;
INV     gate3324  (.A(g1412), .Z(g4052) ) ;
INV     gate3325  (.A(g1529), .Z(g4055) ) ;
INV     gate3326  (.A(g1534), .Z(g4058) ) ;
INV     gate3327  (.A(g1536), .Z(g4061) ) ;
INV     gate3328  (.A(g1550), .Z(g4064) ) ;
INV     gate3329  (.A(g1555), .Z(g4067) ) ;
INV     gate3330  (.A(g1557), .Z(g4070) ) ;
INV     gate3331  (.A(g2220), .Z(g4073) ) ;
INV     gate3332  (.A(g2225), .Z(g4076) ) ;
INV     gate3333  (.A(g2227), .Z(g4079) ) ;
INV     gate3334  (.A(g2246), .Z(g4082) ) ;
INV     gate3335  (.A(g2248), .Z(g4085) ) ;
INV     gate3336  (.A(g2836), .Z(II13316) ) ;
INV     gate3337  (.A(g2836), .Z(g4089) ) ;
INV     gate3338  (.A(g2864), .Z(II13320) ) ;
INV     gate3339  (.A(g2864), .Z(g4091) ) ;
INV     gate3340  (.A(g3074), .Z(g4092) ) ;
INV     gate3341  (.A(g33), .Z(g4093) ) ;
INV     gate3342  (.A(g3207), .Z(g4094) ) ;
INV     gate3343  (.A(g130), .Z(g4095) ) ;
INV     gate3344  (.A(g156), .Z(g4098) ) ;
INV     gate3345  (.A(g161), .Z(g4101) ) ;
INV     gate3346  (.A(g163), .Z(g4104) ) ;
INV     gate3347  (.A(g177), .Z(g4107) ) ;
INV     gate3348  (.A(g414), .Z(g4110) ) ;
INV     gate3349  (.A(g420), .Z(g4111) ) ;
INV     gate3350  (.A(g428), .Z(g4112) ) ;
INV     gate3351  (.A(g698), .Z(g4115) ) ;
INV     gate3352  (.A(g703), .Z(g4118) ) ;
INV     gate3353  (.A(g705), .Z(g4121) ) ;
INV     gate3354  (.A(g725), .Z(g4124) ) ;
INV     gate3355  (.A(g841), .Z(g4127) ) ;
INV     gate3356  (.A(g846), .Z(g4130) ) ;
INV     gate3357  (.A(g848), .Z(g4133) ) ;
INV     gate3358  (.A(g862), .Z(g4136) ) ;
INV     gate3359  (.A(g867), .Z(g4139) ) ;
INV     gate3360  (.A(g1098), .Z(g4142) ) ;
INV     gate3361  (.A(g1104), .Z(g4143) ) ;
INV     gate3362  (.A(g1114), .Z(g4144) ) ;
INV     gate3363  (.A(g1386), .Z(g4147) ) ;
INV     gate3364  (.A(g1388), .Z(g4150) ) ;
INV     gate3365  (.A(g1413), .Z(g4153) ) ;
INV     gate3366  (.A(g1532), .Z(g4156) ) ;
INV     gate3367  (.A(g1537), .Z(g4159) ) ;
INV     gate3368  (.A(g1539), .Z(g4162) ) ;
INV     gate3369  (.A(g1553), .Z(g4165) ) ;
INV     gate3370  (.A(g1558), .Z(g4168) ) ;
INV     gate3371  (.A(g1560), .Z(g4171) ) ;
INV     gate3372  (.A(g1789), .Z(g4174) ) ;
INV     gate3373  (.A(g1836), .Z(g4175) ) ;
INV     gate3374  (.A(g2079), .Z(g4176) ) ;
INV     gate3375  (.A(g2106), .Z(g4179) ) ;
INV     gate3376  (.A(g2223), .Z(g4182) ) ;
INV     gate3377  (.A(g2228), .Z(g4185) ) ;
INV     gate3378  (.A(g2230), .Z(g4188) ) ;
INV     gate3379  (.A(g2244), .Z(g4191) ) ;
INV     gate3380  (.A(g2249), .Z(g4194) ) ;
INV     gate3381  (.A(g2251), .Z(g4197) ) ;
INV     gate3382  (.A(g2851), .Z(II13366) ) ;
INV     gate3383  (.A(g2851), .Z(g4201) ) ;
INV     gate3384  (.A(g42), .Z(g4202) ) ;
INV     gate3385  (.A(g20), .Z(g4203) ) ;
INV     gate3386  (.A(g3188), .Z(g4204) ) ;
INV     gate3387  (.A(g131), .Z(g4205) ) ;
INV     gate3388  (.A(g133), .Z(g4208) ) ;
INV     gate3389  (.A(g159), .Z(g4211) ) ;
INV     gate3390  (.A(g164), .Z(g4214) ) ;
INV     gate3391  (.A(g354), .Z(g4217) ) ;
INV     gate3392  (.A(g423), .Z(g4220) ) ;
INV     gate3393  (.A(g426), .Z(g4221) ) ;
INV     gate3394  (.A(g429), .Z(g4224) ) ;
INV     gate3395  (.A(g701), .Z(g4225) ) ;
INV     gate3396  (.A(g706), .Z(g4228) ) ;
INV     gate3397  (.A(g708), .Z(g4231) ) ;
INV     gate3398  (.A(g818), .Z(g4234) ) ;
INV     gate3399  (.A(g844), .Z(g4237) ) ;
INV     gate3400  (.A(g849), .Z(g4240) ) ;
INV     gate3401  (.A(g851), .Z(g4243) ) ;
INV     gate3402  (.A(g865), .Z(g4246) ) ;
INV     gate3403  (.A(g1101), .Z(g4249) ) ;
INV     gate3404  (.A(g1107), .Z(g4250) ) ;
INV     gate3405  (.A(g1115), .Z(g4251) ) ;
INV     gate3406  (.A(g1384), .Z(g4254) ) ;
INV     gate3407  (.A(g1389), .Z(g4257) ) ;
INV     gate3408  (.A(g1391), .Z(g4260) ) ;
INV     gate3409  (.A(g1411), .Z(g4263) ) ;
INV     gate3410  (.A(g1535), .Z(g4266) ) ;
INV     gate3411  (.A(g1540), .Z(g4269) ) ;
INV     gate3412  (.A(g1542), .Z(g4272) ) ;
INV     gate3413  (.A(g1556), .Z(g4275) ) ;
INV     gate3414  (.A(g1561), .Z(g4278) ) ;
INV     gate3415  (.A(g1792), .Z(g4281) ) ;
INV     gate3416  (.A(g1798), .Z(g4282) ) ;
INV     gate3417  (.A(g1808), .Z(g4283) ) ;
INV     gate3418  (.A(g2080), .Z(g4286) ) ;
INV     gate3419  (.A(g2082), .Z(g4289) ) ;
INV     gate3420  (.A(g2107), .Z(g4292) ) ;
INV     gate3421  (.A(g2226), .Z(g4295) ) ;
INV     gate3422  (.A(g2231), .Z(g4298) ) ;
INV     gate3423  (.A(g2233), .Z(g4301) ) ;
INV     gate3424  (.A(g2247), .Z(g4304) ) ;
INV     gate3425  (.A(g2252), .Z(g4307) ) ;
INV     gate3426  (.A(g2254), .Z(g4310) ) ;
INV     gate3427  (.A(g2483), .Z(g4313) ) ;
INV     gate3428  (.A(g2530), .Z(g4314) ) ;
INV     gate3429  (.A(g2773), .Z(g4315) ) ;
INV     gate3430  (.A(g2800), .Z(g4318) ) ;
INV     gate3431  (.A(g2839), .Z(II13417) ) ;
INV     gate3432  (.A(g2839), .Z(g4322) ) ;
INV     gate3433  (.A(g2867), .Z(II13421) ) ;
INV     gate3434  (.A(g2867), .Z(g4324) ) ;
INV     gate3435  (.A(g36), .Z(g4325) ) ;
INV     gate3436  (.A(g181), .Z(g4326) ) ;
INV     gate3437  (.A(g129), .Z(g4329) ) ;
INV     gate3438  (.A(g134), .Z(g4332) ) ;
INV     gate3439  (.A(g162), .Z(g4335) ) ;
INV     gate3440  (.A(g101), .Z(II13430) ) ;
INV     gate3441  (.A(II13430), .Z(g4338) ) ;
INV     gate3442  (.A(g105), .Z(II13433) ) ;
INV     gate3443  (.A(II13433), .Z(g4339) ) ;
INV     gate3444  (.A(g343), .Z(g4340) ) ;
INV     gate3445  (.A(g369), .Z(g4343) ) ;
INV     gate3446  (.A(g432), .Z(g4346) ) ;
INV     gate3447  (.A(g438), .Z(g4347) ) ;
INV     gate3448  (.A(g704), .Z(g4348) ) ;
INV     gate3449  (.A(g709), .Z(g4351) ) ;
INV     gate3450  (.A(g711), .Z(g4354) ) ;
INV     gate3451  (.A(g729), .Z(g4357) ) ;
INV     gate3452  (.A(g819), .Z(g4360) ) ;
INV     gate3453  (.A(g821), .Z(g4363) ) ;
INV     gate3454  (.A(g847), .Z(g4366) ) ;
INV     gate3455  (.A(g852), .Z(g4369) ) ;
INV     gate3456  (.A(g1041), .Z(g4372) ) ;
INV     gate3457  (.A(g1110), .Z(g4375) ) ;
INV     gate3458  (.A(g1113), .Z(g4376) ) ;
INV     gate3459  (.A(g1116), .Z(g4379) ) ;
INV     gate3460  (.A(g1387), .Z(g4380) ) ;
INV     gate3461  (.A(g1392), .Z(g4383) ) ;
INV     gate3462  (.A(g1394), .Z(g4386) ) ;
INV     gate3463  (.A(g1512), .Z(g4389) ) ;
INV     gate3464  (.A(g1538), .Z(g4392) ) ;
INV     gate3465  (.A(g1543), .Z(g4395) ) ;
INV     gate3466  (.A(g1545), .Z(g4398) ) ;
INV     gate3467  (.A(g1559), .Z(g4401) ) ;
INV     gate3468  (.A(g1795), .Z(g4404) ) ;
INV     gate3469  (.A(g1801), .Z(g4405) ) ;
INV     gate3470  (.A(g1809), .Z(g4406) ) ;
INV     gate3471  (.A(g2078), .Z(g4409) ) ;
INV     gate3472  (.A(g2083), .Z(g4412) ) ;
INV     gate3473  (.A(g2085), .Z(g4415) ) ;
INV     gate3474  (.A(g2105), .Z(g4418) ) ;
INV     gate3475  (.A(g2229), .Z(g4421) ) ;
INV     gate3476  (.A(g2234), .Z(g4424) ) ;
INV     gate3477  (.A(g2236), .Z(g4427) ) ;
INV     gate3478  (.A(g2250), .Z(g4430) ) ;
INV     gate3479  (.A(g2255), .Z(g4433) ) ;
INV     gate3480  (.A(g2486), .Z(g4436) ) ;
INV     gate3481  (.A(g2492), .Z(g4437) ) ;
INV     gate3482  (.A(g2502), .Z(g4438) ) ;
INV     gate3483  (.A(g2774), .Z(g4441) ) ;
INV     gate3484  (.A(g2776), .Z(g4444) ) ;
INV     gate3485  (.A(g2801), .Z(g4447) ) ;
INV     gate3486  (.A(g2854), .Z(II13478) ) ;
INV     gate3487  (.A(g2854), .Z(g4451) ) ;
INV     gate3488  (.A(g17), .Z(g4452) ) ;
INV     gate3489  (.A(g132), .Z(g4453) ) ;
INV     gate3490  (.A(g309), .Z(g4456) ) ;
INV     gate3491  (.A(g346), .Z(g4465) ) ;
INV     gate3492  (.A(g358), .Z(g4468) ) ;
INV     gate3493  (.A(g384), .Z(g4471) ) ;
INV     gate3494  (.A(g435), .Z(g4474) ) ;
INV     gate3495  (.A(g441), .Z(g4475) ) ;
INV     gate3496  (.A(g576), .Z(g4476) ) ;
INV     gate3497  (.A(g587), .Z(g4479) ) ;
INV     gate3498  (.A(g707), .Z(g4480) ) ;
INV     gate3499  (.A(g712), .Z(g4483) ) ;
INV     gate3500  (.A(g714), .Z(g4486) ) ;
INV     gate3501  (.A(g730), .Z(g4489) ) ;
INV     gate3502  (.A(g732), .Z(g4492) ) ;
INV     gate3503  (.A(g869), .Z(g4495) ) ;
INV     gate3504  (.A(g817), .Z(g4498) ) ;
INV     gate3505  (.A(g822), .Z(g4501) ) ;
INV     gate3506  (.A(g850), .Z(g4504) ) ;
INV     gate3507  (.A(g789), .Z(II13501) ) ;
INV     gate3508  (.A(II13501), .Z(g4507) ) ;
INV     gate3509  (.A(g793), .Z(II13504) ) ;
INV     gate3510  (.A(II13504), .Z(g4508) ) ;
INV     gate3511  (.A(g1030), .Z(g4509) ) ;
INV     gate3512  (.A(g1056), .Z(g4512) ) ;
INV     gate3513  (.A(g1119), .Z(g4515) ) ;
INV     gate3514  (.A(g1125), .Z(g4516) ) ;
INV     gate3515  (.A(g1390), .Z(g4517) ) ;
INV     gate3516  (.A(g1395), .Z(g4520) ) ;
INV     gate3517  (.A(g1397), .Z(g4523) ) ;
INV     gate3518  (.A(g1415), .Z(g4526) ) ;
INV     gate3519  (.A(g1513), .Z(g4529) ) ;
INV     gate3520  (.A(g1515), .Z(g4532) ) ;
INV     gate3521  (.A(g1541), .Z(g4535) ) ;
INV     gate3522  (.A(g1546), .Z(g4538) ) ;
INV     gate3523  (.A(g1735), .Z(g4541) ) ;
INV     gate3524  (.A(g1804), .Z(g4544) ) ;
INV     gate3525  (.A(g1807), .Z(g4545) ) ;
INV     gate3526  (.A(g1810), .Z(g4548) ) ;
INV     gate3527  (.A(g2081), .Z(g4549) ) ;
INV     gate3528  (.A(g2086), .Z(g4552) ) ;
INV     gate3529  (.A(g2088), .Z(g4555) ) ;
INV     gate3530  (.A(g2206), .Z(g4558) ) ;
INV     gate3531  (.A(g2232), .Z(g4561) ) ;
INV     gate3532  (.A(g2237), .Z(g4564) ) ;
INV     gate3533  (.A(g2239), .Z(g4567) ) ;
INV     gate3534  (.A(g2253), .Z(g4570) ) ;
INV     gate3535  (.A(g2489), .Z(g4573) ) ;
INV     gate3536  (.A(g2495), .Z(g4574) ) ;
INV     gate3537  (.A(g2503), .Z(g4575) ) ;
INV     gate3538  (.A(g2772), .Z(g4578) ) ;
INV     gate3539  (.A(g2777), .Z(g4581) ) ;
INV     gate3540  (.A(g2779), .Z(g4584) ) ;
INV     gate3541  (.A(g2799), .Z(g4587) ) ;
INV     gate3542  (.A(g2870), .Z(II13538) ) ;
INV     gate3543  (.A(g2870), .Z(g4591) ) ;
INV     gate3544  (.A(g361), .Z(g4592) ) ;
INV     gate3545  (.A(g373), .Z(g4595) ) ;
INV     gate3546  (.A(g398), .Z(g4598) ) ;
INV     gate3547  (.A(g444), .Z(g4601) ) ;
INV     gate3548  (.A(g525), .Z(g4602) ) ;
INV     gate3549  (.A(g577), .Z(g4603) ) ;
INV     gate3550  (.A(g579), .Z(g4606) ) ;
INV     gate3551  (.A(g590), .Z(g4609) ) ;
INV     gate3552  (.A(g596), .Z(g4610) ) ;
INV     gate3553  (.A(g710), .Z(g4611) ) ;
INV     gate3554  (.A(g715), .Z(g4614) ) ;
INV     gate3555  (.A(g717), .Z(g4617) ) ;
INV     gate3556  (.A(g728), .Z(g4620) ) ;
INV     gate3557  (.A(g733), .Z(g4623) ) ;
INV     gate3558  (.A(g735), .Z(g4626) ) ;
INV     gate3559  (.A(g820), .Z(g4629) ) ;
INV     gate3560  (.A(g996), .Z(g4632) ) ;
INV     gate3561  (.A(g1033), .Z(g4641) ) ;
INV     gate3562  (.A(g1045), .Z(g4644) ) ;
INV     gate3563  (.A(g1071), .Z(g4647) ) ;
INV     gate3564  (.A(g1122), .Z(g4650) ) ;
INV     gate3565  (.A(g1128), .Z(g4651) ) ;
INV     gate3566  (.A(g1262), .Z(g4652) ) ;
INV     gate3567  (.A(g1273), .Z(g4655) ) ;
INV     gate3568  (.A(g1393), .Z(g4656) ) ;
INV     gate3569  (.A(g1398), .Z(g4659) ) ;
INV     gate3570  (.A(g1400), .Z(g4662) ) ;
INV     gate3571  (.A(g1416), .Z(g4665) ) ;
INV     gate3572  (.A(g1418), .Z(g4668) ) ;
INV     gate3573  (.A(g1563), .Z(g4671) ) ;
INV     gate3574  (.A(g1511), .Z(g4674) ) ;
INV     gate3575  (.A(g1516), .Z(g4677) ) ;
INV     gate3576  (.A(g1544), .Z(g4680) ) ;
INV     gate3577  (.A(g1476), .Z(II13575) ) ;
INV     gate3578  (.A(II13575), .Z(g4683) ) ;
INV     gate3579  (.A(g1481), .Z(II13578) ) ;
INV     gate3580  (.A(II13578), .Z(g4684) ) ;
INV     gate3581  (.A(g1724), .Z(g4685) ) ;
INV     gate3582  (.A(g1750), .Z(g4688) ) ;
INV     gate3583  (.A(g1813), .Z(g4691) ) ;
INV     gate3584  (.A(g1819), .Z(g4692) ) ;
INV     gate3585  (.A(g2084), .Z(g4693) ) ;
INV     gate3586  (.A(g2089), .Z(g4696) ) ;
INV     gate3587  (.A(g2091), .Z(g4699) ) ;
INV     gate3588  (.A(g2109), .Z(g4702) ) ;
INV     gate3589  (.A(g2207), .Z(g4705) ) ;
INV     gate3590  (.A(g2209), .Z(g4708) ) ;
INV     gate3591  (.A(g2235), .Z(g4711) ) ;
INV     gate3592  (.A(g2240), .Z(g4714) ) ;
INV     gate3593  (.A(g2429), .Z(g4717) ) ;
INV     gate3594  (.A(g2498), .Z(g4720) ) ;
INV     gate3595  (.A(g2501), .Z(g4721) ) ;
INV     gate3596  (.A(g2504), .Z(g4724) ) ;
INV     gate3597  (.A(g2775), .Z(g4725) ) ;
INV     gate3598  (.A(g2780), .Z(g4728) ) ;
INV     gate3599  (.A(g2782), .Z(g4731) ) ;
INV     gate3600  (.A(g11), .Z(g4734) ) ;
INV     gate3601  (.A(g121), .Z(II13601) ) ;
INV     gate3602  (.A(II13601), .Z(g4735) ) ;
INV     gate3603  (.A(g125), .Z(II13604) ) ;
INV     gate3604  (.A(II13604), .Z(g4736) ) ;
INV     gate3605  (.A(g376), .Z(g4737) ) ;
INV     gate3606  (.A(g388), .Z(g4740) ) ;
INV     gate3607  (.A(g575), .Z(g4743) ) ;
INV     gate3608  (.A(g580), .Z(g4746) ) ;
INV     gate3609  (.A(g582), .Z(g4749) ) ;
INV     gate3610  (.A(g593), .Z(g4752) ) ;
INV     gate3611  (.A(g599), .Z(g4753) ) ;
INV     gate3612  (.A(g713), .Z(g4754) ) ;
INV     gate3613  (.A(g718), .Z(g4757) ) ;
INV     gate3614  (.A(g720), .Z(g4760) ) ;
INV     gate3615  (.A(g731), .Z(g4763) ) ;
INV     gate3616  (.A(g736), .Z(g4766) ) ;
INV     gate3617  (.A(g1048), .Z(g4769) ) ;
INV     gate3618  (.A(g1060), .Z(g4772) ) ;
INV     gate3619  (.A(g1085), .Z(g4775) ) ;
INV     gate3620  (.A(g1131), .Z(g4778) ) ;
INV     gate3621  (.A(g1211), .Z(g4779) ) ;
INV     gate3622  (.A(g1263), .Z(g4780) ) ;
INV     gate3623  (.A(g1265), .Z(g4783) ) ;
INV     gate3624  (.A(g1276), .Z(g4786) ) ;
INV     gate3625  (.A(g1282), .Z(g4787) ) ;
INV     gate3626  (.A(g1396), .Z(g4788) ) ;
INV     gate3627  (.A(g1401), .Z(g4791) ) ;
INV     gate3628  (.A(g1403), .Z(g4794) ) ;
INV     gate3629  (.A(g1414), .Z(g4797) ) ;
INV     gate3630  (.A(g1419), .Z(g4800) ) ;
INV     gate3631  (.A(g1421), .Z(g4803) ) ;
INV     gate3632  (.A(g1514), .Z(g4806) ) ;
INV     gate3633  (.A(g1690), .Z(g4809) ) ;
INV     gate3634  (.A(g1727), .Z(g4818) ) ;
INV     gate3635  (.A(g1739), .Z(g4821) ) ;
INV     gate3636  (.A(g1765), .Z(g4824) ) ;
INV     gate3637  (.A(g1816), .Z(g4827) ) ;
INV     gate3638  (.A(g1822), .Z(g4828) ) ;
INV     gate3639  (.A(g1956), .Z(g4829) ) ;
INV     gate3640  (.A(g1967), .Z(g4832) ) ;
INV     gate3641  (.A(g2087), .Z(g4833) ) ;
INV     gate3642  (.A(g2092), .Z(g4836) ) ;
INV     gate3643  (.A(g2094), .Z(g4839) ) ;
INV     gate3644  (.A(g2110), .Z(g4842) ) ;
INV     gate3645  (.A(g2112), .Z(g4845) ) ;
INV     gate3646  (.A(g2257), .Z(g4848) ) ;
INV     gate3647  (.A(g2205), .Z(g4851) ) ;
INV     gate3648  (.A(g2210), .Z(g4854) ) ;
INV     gate3649  (.A(g2238), .Z(g4857) ) ;
INV     gate3650  (.A(g2170), .Z(II13652) ) ;
INV     gate3651  (.A(II13652), .Z(g4860) ) ;
INV     gate3652  (.A(g2175), .Z(II13655) ) ;
INV     gate3653  (.A(II13655), .Z(g4861) ) ;
INV     gate3654  (.A(g2418), .Z(g4862) ) ;
INV     gate3655  (.A(g2444), .Z(g4865) ) ;
INV     gate3656  (.A(g2507), .Z(g4868) ) ;
INV     gate3657  (.A(g2513), .Z(g4869) ) ;
INV     gate3658  (.A(g2778), .Z(g4870) ) ;
INV     gate3659  (.A(g2783), .Z(g4873) ) ;
INV     gate3660  (.A(g2785), .Z(g4876) ) ;
INV     gate3661  (.A(g2803), .Z(g4879) ) ;
INV     gate3662  (.A(g391), .Z(g4882) ) ;
INV     gate3663  (.A(g448), .Z(g4885) ) ;
INV     gate3664  (.A(g578), .Z(g4888) ) ;
INV     gate3665  (.A(g583), .Z(g4891) ) ;
INV     gate3666  (.A(g585), .Z(g4894) ) ;
INV     gate3667  (.A(g602), .Z(g4897) ) ;
INV     gate3668  (.A(g605), .Z(g4898) ) ;
INV     gate3669  (.A(g716), .Z(g4899) ) ;
INV     gate3670  (.A(g721), .Z(g4902) ) ;
INV     gate3671  (.A(g723), .Z(g4905) ) ;
INV     gate3672  (.A(g734), .Z(g4908) ) ;
INV     gate3673  (.A(g809), .Z(II13677) ) ;
INV     gate3674  (.A(II13677), .Z(g4911) ) ;
INV     gate3675  (.A(g813), .Z(II13680) ) ;
INV     gate3676  (.A(II13680), .Z(g4912) ) ;
INV     gate3677  (.A(g1063), .Z(g4913) ) ;
INV     gate3678  (.A(g1075), .Z(g4916) ) ;
INV     gate3679  (.A(g1261), .Z(g4919) ) ;
INV     gate3680  (.A(g1266), .Z(g4922) ) ;
INV     gate3681  (.A(g1268), .Z(g4925) ) ;
INV     gate3682  (.A(g1279), .Z(g4928) ) ;
INV     gate3683  (.A(g1285), .Z(g4929) ) ;
INV     gate3684  (.A(g1399), .Z(g4930) ) ;
INV     gate3685  (.A(g1404), .Z(g4933) ) ;
INV     gate3686  (.A(g1406), .Z(g4936) ) ;
INV     gate3687  (.A(g1417), .Z(g4939) ) ;
INV     gate3688  (.A(g1422), .Z(g4942) ) ;
INV     gate3689  (.A(g1742), .Z(g4945) ) ;
INV     gate3690  (.A(g1754), .Z(g4948) ) ;
INV     gate3691  (.A(g1779), .Z(g4951) ) ;
INV     gate3692  (.A(g1825), .Z(g4954) ) ;
INV     gate3693  (.A(g1905), .Z(g4955) ) ;
INV     gate3694  (.A(g1957), .Z(g4956) ) ;
INV     gate3695  (.A(g1959), .Z(g4959) ) ;
INV     gate3696  (.A(g1970), .Z(g4962) ) ;
INV     gate3697  (.A(g1976), .Z(g4963) ) ;
INV     gate3698  (.A(g2090), .Z(g4964) ) ;
INV     gate3699  (.A(g2095), .Z(g4967) ) ;
INV     gate3700  (.A(g2097), .Z(g4970) ) ;
INV     gate3701  (.A(g2108), .Z(g4973) ) ;
INV     gate3702  (.A(g2113), .Z(g4976) ) ;
INV     gate3703  (.A(g2115), .Z(g4979) ) ;
INV     gate3704  (.A(g2208), .Z(g4982) ) ;
INV     gate3705  (.A(g2384), .Z(g4985) ) ;
INV     gate3706  (.A(g2421), .Z(g4994) ) ;
INV     gate3707  (.A(g2433), .Z(g4997) ) ;
INV     gate3708  (.A(g2459), .Z(g5000) ) ;
INV     gate3709  (.A(g2510), .Z(g5003) ) ;
INV     gate3710  (.A(g2516), .Z(g5004) ) ;
INV     gate3711  (.A(g2650), .Z(g5005) ) ;
INV     gate3712  (.A(g2661), .Z(g5008) ) ;
INV     gate3713  (.A(g2781), .Z(g5009) ) ;
INV     gate3714  (.A(g2786), .Z(g5012) ) ;
INV     gate3715  (.A(g2788), .Z(g5015) ) ;
INV     gate3716  (.A(g2804), .Z(g5018) ) ;
INV     gate3717  (.A(g2806), .Z(g5021) ) ;
INV     gate3718  (.A(g449), .Z(g5024) ) ;
INV     gate3719  (.A(g581), .Z(g5027) ) ;
INV     gate3720  (.A(g586), .Z(g5030) ) ;
INV     gate3721  (.A(g608), .Z(g5033) ) ;
INV     gate3722  (.A(g614), .Z(g5034) ) ;
INV     gate3723  (.A(g719), .Z(g5035) ) ;
INV     gate3724  (.A(g724), .Z(g5038) ) ;
INV     gate3725  (.A(g1078), .Z(g5041) ) ;
INV     gate3726  (.A(g1135), .Z(g5044) ) ;
INV     gate3727  (.A(g1264), .Z(g5047) ) ;
INV     gate3728  (.A(g1269), .Z(g5050) ) ;
INV     gate3729  (.A(g1271), .Z(g5053) ) ;
INV     gate3730  (.A(g1288), .Z(g5056) ) ;
INV     gate3731  (.A(g1291), .Z(g5057) ) ;
INV     gate3732  (.A(g1402), .Z(g5058) ) ;
INV     gate3733  (.A(g1407), .Z(g5061) ) ;
INV     gate3734  (.A(g1409), .Z(g5064) ) ;
INV     gate3735  (.A(g1420), .Z(g5067) ) ;
INV     gate3736  (.A(g1501), .Z(II13742) ) ;
INV     gate3737  (.A(II13742), .Z(g5070) ) ;
INV     gate3738  (.A(g1506), .Z(II13745) ) ;
INV     gate3739  (.A(II13745), .Z(g5071) ) ;
INV     gate3740  (.A(g1757), .Z(g5072) ) ;
INV     gate3741  (.A(g1769), .Z(g5075) ) ;
INV     gate3742  (.A(g1955), .Z(g5078) ) ;
INV     gate3743  (.A(g1960), .Z(g5081) ) ;
INV     gate3744  (.A(g1962), .Z(g5084) ) ;
INV     gate3745  (.A(g1973), .Z(g5087) ) ;
INV     gate3746  (.A(g1979), .Z(g5088) ) ;
INV     gate3747  (.A(g2093), .Z(g5089) ) ;
INV     gate3748  (.A(g2098), .Z(g5092) ) ;
INV     gate3749  (.A(g2100), .Z(g5095) ) ;
INV     gate3750  (.A(g2111), .Z(g5098) ) ;
INV     gate3751  (.A(g2116), .Z(g5101) ) ;
INV     gate3752  (.A(g2436), .Z(g5104) ) ;
INV     gate3753  (.A(g2448), .Z(g5107) ) ;
INV     gate3754  (.A(g2473), .Z(g5110) ) ;
INV     gate3755  (.A(g2519), .Z(g5113) ) ;
INV     gate3756  (.A(g2599), .Z(g5114) ) ;
INV     gate3757  (.A(g2651), .Z(g5115) ) ;
INV     gate3758  (.A(g2653), .Z(g5118) ) ;
INV     gate3759  (.A(g2664), .Z(g5121) ) ;
INV     gate3760  (.A(g2670), .Z(g5122) ) ;
INV     gate3761  (.A(g2784), .Z(g5123) ) ;
INV     gate3762  (.A(g2789), .Z(g5126) ) ;
INV     gate3763  (.A(g2791), .Z(g5129) ) ;
INV     gate3764  (.A(g2802), .Z(g5132) ) ;
INV     gate3765  (.A(g2807), .Z(g5135) ) ;
INV     gate3766  (.A(g2809), .Z(g5138) ) ;
INV     gate3767  (.A(g109), .Z(II13775) ) ;
INV     gate3768  (.A(II13775), .Z(g5141) ) ;
INV     gate3769  (.A(g447), .Z(g5142) ) ;
INV     gate3770  (.A(g584), .Z(g5145) ) ;
INV     gate3771  (.A(g611), .Z(g5148) ) ;
INV     gate3772  (.A(g617), .Z(g5149) ) ;
INV     gate3773  (.A(g722), .Z(g5150) ) ;
INV     gate3774  (.A(g1136), .Z(g5153) ) ;
INV     gate3775  (.A(g1267), .Z(g5156) ) ;
INV     gate3776  (.A(g1272), .Z(g5159) ) ;
INV     gate3777  (.A(g1294), .Z(g5162) ) ;
INV     gate3778  (.A(g1300), .Z(g5163) ) ;
INV     gate3779  (.A(g1405), .Z(g5164) ) ;
INV     gate3780  (.A(g1410), .Z(g5167) ) ;
INV     gate3781  (.A(g1772), .Z(g5170) ) ;
INV     gate3782  (.A(g1829), .Z(g5173) ) ;
INV     gate3783  (.A(g1958), .Z(g5176) ) ;
INV     gate3784  (.A(g1963), .Z(g5179) ) ;
INV     gate3785  (.A(g1965), .Z(g5182) ) ;
INV     gate3786  (.A(g1982), .Z(g5185) ) ;
INV     gate3787  (.A(g1985), .Z(g5186) ) ;
INV     gate3788  (.A(g2096), .Z(g5187) ) ;
INV     gate3789  (.A(g2101), .Z(g5190) ) ;
INV     gate3790  (.A(g2103), .Z(g5193) ) ;
INV     gate3791  (.A(g2114), .Z(g5196) ) ;
INV     gate3792  (.A(g2195), .Z(II13801) ) ;
INV     gate3793  (.A(II13801), .Z(g5199) ) ;
INV     gate3794  (.A(g2200), .Z(II13804) ) ;
INV     gate3795  (.A(II13804), .Z(g5200) ) ;
INV     gate3796  (.A(g2451), .Z(g5201) ) ;
INV     gate3797  (.A(g2463), .Z(g5204) ) ;
INV     gate3798  (.A(g2649), .Z(g5207) ) ;
INV     gate3799  (.A(g2654), .Z(g5210) ) ;
INV     gate3800  (.A(g2656), .Z(g5213) ) ;
INV     gate3801  (.A(g2667), .Z(g5216) ) ;
INV     gate3802  (.A(g2673), .Z(g5217) ) ;
INV     gate3803  (.A(g2787), .Z(g5218) ) ;
INV     gate3804  (.A(g2792), .Z(g5221) ) ;
INV     gate3805  (.A(g2794), .Z(g5224) ) ;
INV     gate3806  (.A(g2805), .Z(g5227) ) ;
INV     gate3807  (.A(g2810), .Z(g5230) ) ;
INV     gate3808  (.A(g620), .Z(g5233) ) ;
INV     gate3809  (.A(g797), .Z(II13820) ) ;
INV     gate3810  (.A(II13820), .Z(g5234) ) ;
INV     gate3811  (.A(g1134), .Z(g5235) ) ;
INV     gate3812  (.A(g1270), .Z(g5238) ) ;
INV     gate3813  (.A(g1297), .Z(g5241) ) ;
INV     gate3814  (.A(g1303), .Z(g5242) ) ;
INV     gate3815  (.A(g1408), .Z(g5243) ) ;
INV     gate3816  (.A(g1830), .Z(g5246) ) ;
INV     gate3817  (.A(g1961), .Z(g5249) ) ;
INV     gate3818  (.A(g1966), .Z(g5252) ) ;
INV     gate3819  (.A(g1988), .Z(g5255) ) ;
INV     gate3820  (.A(g1994), .Z(g5256) ) ;
INV     gate3821  (.A(g2099), .Z(g5257) ) ;
INV     gate3822  (.A(g2104), .Z(g5260) ) ;
INV     gate3823  (.A(g2466), .Z(g5263) ) ;
INV     gate3824  (.A(g2523), .Z(g5266) ) ;
INV     gate3825  (.A(g2652), .Z(g5269) ) ;
INV     gate3826  (.A(g2657), .Z(g5272) ) ;
INV     gate3827  (.A(g2659), .Z(g5275) ) ;
INV     gate3828  (.A(g2676), .Z(g5278) ) ;
INV     gate3829  (.A(g2679), .Z(g5279) ) ;
INV     gate3830  (.A(g2790), .Z(g5280) ) ;
INV     gate3831  (.A(g2795), .Z(g5283) ) ;
INV     gate3832  (.A(g2797), .Z(g5286) ) ;
INV     gate3833  (.A(g2808), .Z(g5289) ) ;
INV     gate3834  (.A(g2857), .Z(g5292) ) ;
INV     gate3835  (.A(g738), .Z(g5293) ) ;
INV     gate3836  (.A(g1306), .Z(g5296) ) ;
INV     gate3837  (.A(g1486), .Z(II13849) ) ;
INV     gate3838  (.A(II13849), .Z(g5297) ) ;
INV     gate3839  (.A(g1828), .Z(g5298) ) ;
INV     gate3840  (.A(g1964), .Z(g5301) ) ;
INV     gate3841  (.A(g1991), .Z(g5304) ) ;
INV     gate3842  (.A(g1997), .Z(g5305) ) ;
INV     gate3843  (.A(g2102), .Z(g5306) ) ;
INV     gate3844  (.A(g2524), .Z(g5309) ) ;
INV     gate3845  (.A(g2655), .Z(g5312) ) ;
INV     gate3846  (.A(g2660), .Z(g5315) ) ;
INV     gate3847  (.A(g2682), .Z(g5318) ) ;
INV     gate3848  (.A(g2688), .Z(g5319) ) ;
INV     gate3849  (.A(g2793), .Z(g5320) ) ;
INV     gate3850  (.A(g2798), .Z(g5323) ) ;
INV     gate3851  (.A(g2873), .Z(g5326) ) ;
INV     gate3852  (.A(g739), .Z(g5327) ) ;
INV     gate3853  (.A(g1424), .Z(g5330) ) ;
INV     gate3854  (.A(g2000), .Z(g5333) ) ;
INV     gate3855  (.A(g2180), .Z(II13868) ) ;
INV     gate3856  (.A(II13868), .Z(g5334) ) ;
INV     gate3857  (.A(g2522), .Z(g5335) ) ;
INV     gate3858  (.A(g2658), .Z(g5338) ) ;
INV     gate3859  (.A(g2685), .Z(g5341) ) ;
INV     gate3860  (.A(g2691), .Z(g5342) ) ;
INV     gate3861  (.A(g2796), .Z(g5343) ) ;
INV     gate3862  (.A(g3106), .Z(g5346) ) ;
INV     gate3863  (.A(g2877), .Z(g5349) ) ;
INV     gate3864  (.A(g737), .Z(g5352) ) ;
INV     gate3865  (.A(g1425), .Z(g5355) ) ;
INV     gate3866  (.A(g2118), .Z(g5358) ) ;
INV     gate3867  (.A(g2694), .Z(g5361) ) ;
INV     gate3868  (.A(g2817), .Z(g5362) ) ;
INV     gate3869  (.A(g3107), .Z(g5363) ) ;
INV     gate3870  (.A(g2878), .Z(g5366) ) ;
INV     gate3871  (.A(g1423), .Z(g5369) ) ;
INV     gate3872  (.A(g2119), .Z(g5372) ) ;
INV     gate3873  (.A(g2812), .Z(g5375) ) ;
INV     gate3874  (.A(g2933), .Z(g5378) ) ;
INV     gate3875  (.A(g3108), .Z(g5379) ) ;
INV     gate3876  (.A(g2117), .Z(g5382) ) ;
INV     gate3877  (.A(g2813), .Z(g5385) ) ;
INV     gate3878  (.A(g3040), .Z(II13892) ) ;
INV     gate3879  (.A(g3040), .Z(g5389) ) ;
INV     gate3880  (.A(g343), .Z(II13896) ) ;
INV     gate3881  (.A(II13896), .Z(g5390) ) ;
INV     gate3882  (.A(g2811), .Z(g5391) ) ;
INV     gate3883  (.A(g3054), .Z(g5394) ) ;
INV     gate3884  (.A(g346), .Z(II13901) ) ;
INV     gate3885  (.A(II13901), .Z(g5395) ) ;
INV     gate3886  (.A(g358), .Z(II13904) ) ;
INV     gate3887  (.A(II13904), .Z(g5396) ) ;
INV     gate3888  (.A(g1030), .Z(II13907) ) ;
INV     gate3889  (.A(II13907), .Z(g5397) ) ;
INV     gate3890  (.A(g361), .Z(II13910) ) ;
INV     gate3891  (.A(II13910), .Z(g5398) ) ;
INV     gate3892  (.A(g373), .Z(II13913) ) ;
INV     gate3893  (.A(II13913), .Z(g5399) ) ;
INV     gate3894  (.A(g1033), .Z(II13916) ) ;
INV     gate3895  (.A(II13916), .Z(g5400) ) ;
INV     gate3896  (.A(g1045), .Z(II13919) ) ;
INV     gate3897  (.A(II13919), .Z(g5401) ) ;
INV     gate3898  (.A(g1724), .Z(II13922) ) ;
INV     gate3899  (.A(II13922), .Z(g5402) ) ;
INV     gate3900  (.A(g376), .Z(II13925) ) ;
INV     gate3901  (.A(II13925), .Z(g5403) ) ;
INV     gate3902  (.A(g388), .Z(II13928) ) ;
INV     gate3903  (.A(II13928), .Z(g5404) ) ;
INV     gate3904  (.A(g1048), .Z(II13931) ) ;
INV     gate3905  (.A(II13931), .Z(g5405) ) ;
INV     gate3906  (.A(g1060), .Z(II13934) ) ;
INV     gate3907  (.A(II13934), .Z(g5406) ) ;
INV     gate3908  (.A(g1727), .Z(II13937) ) ;
INV     gate3909  (.A(II13937), .Z(g5407) ) ;
INV     gate3910  (.A(g1739), .Z(II13940) ) ;
INV     gate3911  (.A(II13940), .Z(g5408) ) ;
INV     gate3912  (.A(g2418), .Z(II13943) ) ;
INV     gate3913  (.A(II13943), .Z(g5409) ) ;
INV     gate3914  (.A(g3079), .Z(g5410) ) ;
INV     gate3915  (.A(g391), .Z(II13947) ) ;
INV     gate3916  (.A(II13947), .Z(g5411) ) ;
INV     gate3917  (.A(g1063), .Z(II13950) ) ;
INV     gate3918  (.A(II13950), .Z(g5412) ) ;
INV     gate3919  (.A(g1075), .Z(II13953) ) ;
INV     gate3920  (.A(II13953), .Z(g5413) ) ;
INV     gate3921  (.A(g1742), .Z(II13956) ) ;
INV     gate3922  (.A(II13956), .Z(g5414) ) ;
INV     gate3923  (.A(g1754), .Z(II13959) ) ;
INV     gate3924  (.A(II13959), .Z(g5415) ) ;
INV     gate3925  (.A(g2421), .Z(II13962) ) ;
INV     gate3926  (.A(II13962), .Z(g5416) ) ;
INV     gate3927  (.A(g2433), .Z(II13965) ) ;
INV     gate3928  (.A(II13965), .Z(g5417) ) ;
INV     gate3929  (.A(g1078), .Z(II13968) ) ;
INV     gate3930  (.A(II13968), .Z(g5418) ) ;
INV     gate3931  (.A(g1757), .Z(II13971) ) ;
INV     gate3932  (.A(II13971), .Z(g5419) ) ;
INV     gate3933  (.A(g1769), .Z(II13974) ) ;
INV     gate3934  (.A(II13974), .Z(g5420) ) ;
INV     gate3935  (.A(g2436), .Z(II13977) ) ;
INV     gate3936  (.A(II13977), .Z(g5421) ) ;
INV     gate3937  (.A(g2448), .Z(II13980) ) ;
INV     gate3938  (.A(II13980), .Z(g5422) ) ;
INV     gate3939  (.A(g2879), .Z(g5423) ) ;
INV     gate3940  (.A(g1772), .Z(II13984) ) ;
INV     gate3941  (.A(II13984), .Z(g5424) ) ;
INV     gate3942  (.A(g2451), .Z(II13987) ) ;
INV     gate3943  (.A(II13987), .Z(g5425) ) ;
INV     gate3944  (.A(g2463), .Z(II13990) ) ;
INV     gate3945  (.A(II13990), .Z(g5426) ) ;
INV     gate3946  (.A(g2466), .Z(II13993) ) ;
INV     gate3947  (.A(II13993), .Z(g5427) ) ;
INV     gate3948  (.A(g3210), .Z(g5428) ) ;
INV     gate3949  (.A(g3211), .Z(g5431) ) ;
INV     gate3950  (.A(g3084), .Z(g5434) ) ;
INV     gate3951  (.A(g276), .Z(II13999) ) ;
INV     gate3952  (.A(g276), .Z(II14002) ) ;
INV     gate3953  (.A(II14002), .Z(g5438) ) ;
INV     gate3954  (.A(g3085), .Z(g5469) ) ;
INV     gate3955  (.A(g963), .Z(II14006) ) ;
INV     gate3956  (.A(g963), .Z(II14009) ) ;
INV     gate3957  (.A(II14009), .Z(g5473) ) ;
INV     gate3958  (.A(g3086), .Z(g5504) ) ;
INV     gate3959  (.A(g3155), .Z(g5507) ) ;
INV     gate3960  (.A(g499), .Z(II14014) ) ;
INV     gate3961  (.A(II14014), .Z(g5508) ) ;
INV     gate3962  (.A(g1657), .Z(II14017) ) ;
INV     gate3963  (.A(g1657), .Z(II14020) ) ;
INV     gate3964  (.A(II14020), .Z(g5512) ) ;
INV     gate3965  (.A(g3087), .Z(g5543) ) ;
INV     gate3966  (.A(g3164), .Z(g5546) ) ;
INV     gate3967  (.A(g101), .Z(g5547) ) ;
INV     gate3968  (.A(g105), .Z(g5548) ) ;
INV     gate3969  (.A(g182), .Z(II14027) ) ;
INV     gate3970  (.A(g182), .Z(II14030) ) ;
INV     gate3971  (.A(II14030), .Z(g5550) ) ;
INV     gate3972  (.A(g514), .Z(g5551) ) ;
INV     gate3973  (.A(g1186), .Z(II14034) ) ;
INV     gate3974  (.A(II14034), .Z(g5552) ) ;
INV     gate3975  (.A(g2351), .Z(II14037) ) ;
INV     gate3976  (.A(g2351), .Z(II14040) ) ;
INV     gate3977  (.A(II14040), .Z(g5556) ) ;
INV     gate3978  (.A(g3091), .Z(g5587) ) ;
INV     gate3979  (.A(g3158), .Z(g5590) ) ;
INV     gate3980  (.A(g3173), .Z(g5591) ) ;
INV     gate3981  (.A(g515), .Z(g5592) ) ;
INV     gate3982  (.A(g789), .Z(g5593) ) ;
INV     gate3983  (.A(g793), .Z(g5594) ) ;
INV     gate3984  (.A(g870), .Z(II14049) ) ;
INV     gate3985  (.A(g870), .Z(II14052) ) ;
INV     gate3986  (.A(II14052), .Z(g5596) ) ;
INV     gate3987  (.A(g1200), .Z(g5597) ) ;
INV     gate3988  (.A(g1880), .Z(II14056) ) ;
INV     gate3989  (.A(II14056), .Z(g5598) ) ;
INV     gate3990  (.A(g3092), .Z(g5601) ) ;
INV     gate3991  (.A(g3167), .Z(g5604) ) ;
INV     gate3992  (.A(g3182), .Z(g5605) ) ;
INV     gate3993  (.A(g79), .Z(g5606) ) ;
INV     gate3994  (.A(g1201), .Z(g5609) ) ;
INV     gate3995  (.A(g1476), .Z(g5610) ) ;
INV     gate3996  (.A(g1481), .Z(g5611) ) ;
INV     gate3997  (.A(g1564), .Z(II14066) ) ;
INV     gate3998  (.A(g1564), .Z(II14069) ) ;
INV     gate3999  (.A(II14069), .Z(g5613) ) ;
INV     gate4000  (.A(g1894), .Z(g5614) ) ;
INV     gate4001  (.A(g2574), .Z(II14073) ) ;
INV     gate4002  (.A(II14073), .Z(g5615) ) ;
INV     gate4003  (.A(g3093), .Z(g5618) ) ;
INV     gate4004  (.A(g3161), .Z(g5621) ) ;
INV     gate4005  (.A(g3176), .Z(g5622) ) ;
INV     gate4006  (.A(g70), .Z(g5623) ) ;
INV     gate4007  (.A(g121), .Z(g5626) ) ;
INV     gate4008  (.A(g125), .Z(g5627) ) ;
INV     gate4009  (.A(g300), .Z(g5628) ) ;
INV     gate4010  (.A(g325), .Z(II14083) ) ;
INV     gate4011  (.A(g767), .Z(g5631) ) ;
INV     gate4012  (.A(g1895), .Z(g5634) ) ;
INV     gate4013  (.A(g2170), .Z(g5635) ) ;
INV     gate4014  (.A(g2175), .Z(g5636) ) ;
INV     gate4015  (.A(g2258), .Z(II14091) ) ;
INV     gate4016  (.A(g2258), .Z(II14094) ) ;
INV     gate4017  (.A(II14094), .Z(g5638) ) ;
INV     gate4018  (.A(g2588), .Z(g5639) ) ;
INV     gate4019  (.A(g3170), .Z(g5640) ) ;
INV     gate4020  (.A(g3185), .Z(g5641) ) ;
INV     gate4021  (.A(g61), .Z(g5642) ) ;
INV     gate4022  (.A(g101), .Z(g5645) ) ;
INV     gate4023  (.A(g213), .Z(g5646) ) ;
INV     gate4024  (.A(g301), .Z(g5647) ) ;
INV     gate4025  (.A(g331), .Z(II14104) ) ;
INV     gate4026  (.A(g758), .Z(g5651) ) ;
INV     gate4027  (.A(g809), .Z(g5654) ) ;
INV     gate4028  (.A(g813), .Z(g5655) ) ;
INV     gate4029  (.A(g987), .Z(g5656) ) ;
INV     gate4030  (.A(g1012), .Z(II14113) ) ;
INV     gate4031  (.A(g1453), .Z(g5659) ) ;
INV     gate4032  (.A(g2589), .Z(g5662) ) ;
INV     gate4033  (.A(g3179), .Z(g5663) ) ;
INV     gate4034  (.A(g65), .Z(g5664) ) ;
INV     gate4035  (.A(g105), .Z(g5665) ) ;
INV     gate4036  (.A(g216), .Z(g5666) ) ;
INV     gate4037  (.A(g222), .Z(g5667) ) ;
INV     gate4038  (.A(g299), .Z(g5668) ) ;
INV     gate4039  (.A(g302), .Z(g5675) ) ;
INV     gate4040  (.A(g506), .Z(g5679) ) ;
INV     gate4041  (.A(g749), .Z(g5680) ) ;
INV     gate4042  (.A(g789), .Z(g5683) ) ;
INV     gate4043  (.A(g900), .Z(g5684) ) ;
INV     gate4044  (.A(g988), .Z(g5685) ) ;
INV     gate4045  (.A(g1018), .Z(II14134) ) ;
INV     gate4046  (.A(g1444), .Z(g5689) ) ;
INV     gate4047  (.A(g1501), .Z(g5692) ) ;
INV     gate4048  (.A(g1506), .Z(g5693) ) ;
INV     gate4049  (.A(g1681), .Z(g5694) ) ;
INV     gate4050  (.A(g1706), .Z(II14143) ) ;
INV     gate4051  (.A(g2147), .Z(g5697) ) ;
INV     gate4052  (.A(g3088), .Z(g5700) ) ;
INV     gate4053  (.A(g3231), .Z(II14149) ) ;
INV     gate4054  (.A(II14149), .Z(g5701) ) ;
INV     gate4055  (.A(g56), .Z(g5702) ) ;
INV     gate4056  (.A(g109), .Z(g5703) ) ;
INV     gate4057  (.A(g219), .Z(g5704) ) ;
INV     gate4058  (.A(g225), .Z(g5705) ) ;
INV     gate4059  (.A(g231), .Z(g5706) ) ;
INV     gate4060  (.A(g109), .Z(g5707) ) ;
INV     gate4061  (.A(g303), .Z(g5708) ) ;
INV     gate4062  (.A(g305), .Z(g5712) ) ;
INV     gate4063  (.A(g113), .Z(II14163) ) ;
INV     gate4064  (.A(II14163), .Z(g5713) ) ;
INV     gate4065  (.A(g507), .Z(g5714) ) ;
INV     gate4066  (.A(g541), .Z(g5715) ) ;
INV     gate4067  (.A(g753), .Z(g5716) ) ;
INV     gate4068  (.A(g793), .Z(g5717) ) ;
INV     gate4069  (.A(g903), .Z(g5718) ) ;
INV     gate4070  (.A(g909), .Z(g5719) ) ;
INV     gate4071  (.A(g986), .Z(g5720) ) ;
INV     gate4072  (.A(g989), .Z(g5727) ) ;
INV     gate4073  (.A(g1192), .Z(g5731) ) ;
INV     gate4074  (.A(g1435), .Z(g5732) ) ;
INV     gate4075  (.A(g1476), .Z(g5735) ) ;
INV     gate4076  (.A(g1594), .Z(g5736) ) ;
INV     gate4077  (.A(g1682), .Z(g5737) ) ;
INV     gate4078  (.A(g1712), .Z(II14182) ) ;
INV     gate4079  (.A(g2138), .Z(g5741) ) ;
INV     gate4080  (.A(g2195), .Z(g5744) ) ;
INV     gate4081  (.A(g2200), .Z(g5745) ) ;
INV     gate4082  (.A(g2375), .Z(g5746) ) ;
INV     gate4083  (.A(g2400), .Z(II14191) ) ;
INV     gate4084  (.A(g3212), .Z(II14195) ) ;
INV     gate4085  (.A(II14195), .Z(g5749) ) ;
INV     gate4086  (.A(g92), .Z(g5750) ) ;
INV     gate4087  (.A(g52), .Z(g5751) ) ;
INV     gate4088  (.A(g113), .Z(g5752) ) ;
INV     gate4089  (.A(g228), .Z(g5753) ) ;
INV     gate4090  (.A(g234), .Z(g5754) ) ;
INV     gate4091  (.A(g240), .Z(g5755) ) ;
INV     gate4092  (.A(g304), .Z(g5756) ) ;
INV     gate4093  (.A(g508), .Z(g5759) ) ;
INV     gate4094  (.A(g744), .Z(g5760) ) ;
INV     gate4095  (.A(g797), .Z(g5761) ) ;
INV     gate4096  (.A(g906), .Z(g5762) ) ;
INV     gate4097  (.A(g912), .Z(g5763) ) ;
INV     gate4098  (.A(g918), .Z(g5764) ) ;
INV     gate4099  (.A(g797), .Z(g5765) ) ;
INV     gate4100  (.A(g990), .Z(g5766) ) ;
INV     gate4101  (.A(g992), .Z(g5770) ) ;
INV     gate4102  (.A(g801), .Z(II14219) ) ;
INV     gate4103  (.A(II14219), .Z(g5771) ) ;
INV     gate4104  (.A(g1193), .Z(g5772) ) ;
INV     gate4105  (.A(g1227), .Z(g5773) ) ;
INV     gate4106  (.A(g1439), .Z(g5774) ) ;
INV     gate4107  (.A(g1481), .Z(g5775) ) ;
INV     gate4108  (.A(g1597), .Z(g5776) ) ;
INV     gate4109  (.A(g1603), .Z(g5777) ) ;
INV     gate4110  (.A(g1680), .Z(g5778) ) ;
INV     gate4111  (.A(g1683), .Z(g5785) ) ;
INV     gate4112  (.A(g1886), .Z(g5789) ) ;
INV     gate4113  (.A(g2129), .Z(g5790) ) ;
INV     gate4114  (.A(g2170), .Z(g5793) ) ;
INV     gate4115  (.A(g2288), .Z(g5794) ) ;
INV     gate4116  (.A(g2376), .Z(g5795) ) ;
INV     gate4117  (.A(g2406), .Z(II14238) ) ;
INV     gate4118  (.A(g3221), .Z(II14243) ) ;
INV     gate4119  (.A(II14243), .Z(g5799) ) ;
INV     gate4120  (.A(g3227), .Z(II14246) ) ;
INV     gate4121  (.A(II14246), .Z(g5800) ) ;
INV     gate4122  (.A(g3216), .Z(II14249) ) ;
INV     gate4123  (.A(II14249), .Z(g5801) ) ;
INV     gate4124  (.A(g83), .Z(g5802) ) ;
INV     gate4125  (.A(g117), .Z(g5803) ) ;
INV     gate4126  (.A(g237), .Z(g5804) ) ;
INV     gate4127  (.A(g243), .Z(g5805) ) ;
INV     gate4128  (.A(g249), .Z(g5806) ) ;
INV     gate4129  (.A(g509), .Z(g5808) ) ;
INV     gate4130  (.A(g780), .Z(g5809) ) ;
INV     gate4131  (.A(g740), .Z(g5810) ) ;
INV     gate4132  (.A(g801), .Z(g5811) ) ;
INV     gate4133  (.A(g915), .Z(g5812) ) ;
INV     gate4134  (.A(g921), .Z(g5813) ) ;
INV     gate4135  (.A(g927), .Z(g5814) ) ;
INV     gate4136  (.A(g991), .Z(g5815) ) ;
INV     gate4137  (.A(g1194), .Z(g5818) ) ;
INV     gate4138  (.A(g1430), .Z(g5819) ) ;
INV     gate4139  (.A(g1486), .Z(g5820) ) ;
INV     gate4140  (.A(g1600), .Z(g5821) ) ;
INV     gate4141  (.A(g1606), .Z(g5822) ) ;
INV     gate4142  (.A(g1612), .Z(g5823) ) ;
INV     gate4143  (.A(g1486), .Z(g5824) ) ;
INV     gate4144  (.A(g1684), .Z(g5825) ) ;
INV     gate4145  (.A(g1686), .Z(g5829) ) ;
INV     gate4146  (.A(g1491), .Z(II14280) ) ;
INV     gate4147  (.A(II14280), .Z(g5830) ) ;
INV     gate4148  (.A(g1887), .Z(g5831) ) ;
INV     gate4149  (.A(g1921), .Z(g5832) ) ;
INV     gate4150  (.A(g2133), .Z(g5833) ) ;
INV     gate4151  (.A(g2175), .Z(g5834) ) ;
INV     gate4152  (.A(g2291), .Z(g5835) ) ;
INV     gate4153  (.A(g2297), .Z(g5836) ) ;
INV     gate4154  (.A(g2374), .Z(g5837) ) ;
INV     gate4155  (.A(g2377), .Z(g5844) ) ;
INV     gate4156  (.A(g2580), .Z(g5848) ) ;
INV     gate4157  (.A(g3228), .Z(II14295) ) ;
INV     gate4158  (.A(II14295), .Z(g5849) ) ;
INV     gate4159  (.A(g3217), .Z(II14298) ) ;
INV     gate4160  (.A(II14298), .Z(g5850) ) ;
INV     gate4161  (.A(g74), .Z(g5851) ) ;
INV     gate4162  (.A(g121), .Z(g5852) ) ;
INV     gate4163  (.A(g246), .Z(g5853) ) ;
INV     gate4164  (.A(g252), .Z(g5854) ) ;
INV     gate4165  (.A(g258), .Z(g5855) ) ;
INV     gate4166  (.A(g97), .Z(II14306) ) ;
INV     gate4167  (.A(II14306), .Z(g5856) ) ;
INV     gate4168  (.A(g538), .Z(g5857) ) ;
INV     gate4169  (.A(g771), .Z(g5858) ) ;
INV     gate4170  (.A(g805), .Z(g5859) ) ;
INV     gate4171  (.A(g924), .Z(g5860) ) ;
INV     gate4172  (.A(g930), .Z(g5861) ) ;
INV     gate4173  (.A(g936), .Z(g5862) ) ;
INV     gate4174  (.A(g1195), .Z(g5864) ) ;
INV     gate4175  (.A(g1466), .Z(g5865) ) ;
INV     gate4176  (.A(g1426), .Z(g5866) ) ;
INV     gate4177  (.A(g1491), .Z(g5867) ) ;
INV     gate4178  (.A(g1609), .Z(g5868) ) ;
INV     gate4179  (.A(g1615), .Z(g5869) ) ;
INV     gate4180  (.A(g1621), .Z(g5870) ) ;
INV     gate4181  (.A(g1685), .Z(g5871) ) ;
INV     gate4182  (.A(g1888), .Z(g5874) ) ;
INV     gate4183  (.A(g2124), .Z(g5875) ) ;
INV     gate4184  (.A(g2180), .Z(g5876) ) ;
INV     gate4185  (.A(g2294), .Z(g5877) ) ;
INV     gate4186  (.A(g2300), .Z(g5878) ) ;
INV     gate4187  (.A(g2306), .Z(g5879) ) ;
INV     gate4188  (.A(g2180), .Z(g5880) ) ;
INV     gate4189  (.A(g2378), .Z(g5881) ) ;
INV     gate4190  (.A(g2380), .Z(g5885) ) ;
INV     gate4191  (.A(g2185), .Z(II14338) ) ;
INV     gate4192  (.A(II14338), .Z(g5886) ) ;
INV     gate4193  (.A(g2581), .Z(g5887) ) ;
INV     gate4194  (.A(g2615), .Z(g5888) ) ;
INV     gate4195  (.A(g3219), .Z(II14343) ) ;
INV     gate4196  (.A(II14343), .Z(g5889) ) ;
INV     gate4197  (.A(g88), .Z(g5890) ) ;
INV     gate4198  (.A(g125), .Z(g5893) ) ;
INV     gate4199  (.A(g186), .Z(g5894) ) ;
INV     gate4200  (.A(g255), .Z(g5895) ) ;
INV     gate4201  (.A(g261), .Z(g5896) ) ;
INV     gate4202  (.A(g267), .Z(g5897) ) ;
INV     gate4203  (.A(g762), .Z(g5898) ) ;
INV     gate4204  (.A(g809), .Z(g5899) ) ;
INV     gate4205  (.A(g933), .Z(g5900) ) ;
INV     gate4206  (.A(g939), .Z(g5901) ) ;
INV     gate4207  (.A(g945), .Z(g5902) ) ;
INV     gate4208  (.A(g785), .Z(II14357) ) ;
INV     gate4209  (.A(II14357), .Z(g5903) ) ;
INV     gate4210  (.A(g1224), .Z(g5904) ) ;
INV     gate4211  (.A(g1457), .Z(g5905) ) ;
INV     gate4212  (.A(g1496), .Z(g5906) ) ;
INV     gate4213  (.A(g1618), .Z(g5907) ) ;
INV     gate4214  (.A(g1624), .Z(g5908) ) ;
INV     gate4215  (.A(g1630), .Z(g5909) ) ;
INV     gate4216  (.A(g1889), .Z(g5911) ) ;
INV     gate4217  (.A(g2160), .Z(g5912) ) ;
INV     gate4218  (.A(g2120), .Z(g5913) ) ;
INV     gate4219  (.A(g2185), .Z(g5914) ) ;
INV     gate4220  (.A(g2303), .Z(g5915) ) ;
INV     gate4221  (.A(g2309), .Z(g5916) ) ;
INV     gate4222  (.A(g2315), .Z(g5917) ) ;
INV     gate4223  (.A(g2379), .Z(g5918) ) ;
INV     gate4224  (.A(g2582), .Z(g5921) ) ;
INV     gate4225  (.A(g3234), .Z(II14378) ) ;
INV     gate4226  (.A(II14378), .Z(g5922) ) ;
INV     gate4227  (.A(g3223), .Z(II14381) ) ;
INV     gate4228  (.A(II14381), .Z(g5923) ) ;
INV     gate4229  (.A(g3218), .Z(II14384) ) ;
INV     gate4230  (.A(II14384), .Z(g5924) ) ;
INV     gate4231  (.A(g189), .Z(g5925) ) ;
INV     gate4232  (.A(g195), .Z(g5926) ) ;
INV     gate4233  (.A(g264), .Z(g5927) ) ;
INV     gate4234  (.A(g270), .Z(g5928) ) ;
INV     gate4235  (.A(g776), .Z(g5929) ) ;
INV     gate4236  (.A(g813), .Z(g5932) ) ;
INV     gate4237  (.A(g873), .Z(g5933) ) ;
INV     gate4238  (.A(g942), .Z(g5934) ) ;
INV     gate4239  (.A(g948), .Z(g5935) ) ;
INV     gate4240  (.A(g954), .Z(g5936) ) ;
INV     gate4241  (.A(g1448), .Z(g5937) ) ;
INV     gate4242  (.A(g1501), .Z(g5938) ) ;
INV     gate4243  (.A(g1627), .Z(g5939) ) ;
INV     gate4244  (.A(g1633), .Z(g5940) ) ;
INV     gate4245  (.A(g1639), .Z(g5941) ) ;
INV     gate4246  (.A(g1471), .Z(II14402) ) ;
INV     gate4247  (.A(II14402), .Z(g5942) ) ;
INV     gate4248  (.A(g1918), .Z(g5943) ) ;
INV     gate4249  (.A(g2151), .Z(g5944) ) ;
INV     gate4250  (.A(g2190), .Z(g5945) ) ;
INV     gate4251  (.A(g2312), .Z(g5946) ) ;
INV     gate4252  (.A(g2318), .Z(g5947) ) ;
INV     gate4253  (.A(g2324), .Z(g5948) ) ;
INV     gate4254  (.A(g2583), .Z(g5950) ) ;
INV     gate4255  (.A(g3233), .Z(II14413) ) ;
INV     gate4256  (.A(II14413), .Z(g5951) ) ;
INV     gate4257  (.A(g3222), .Z(II14416) ) ;
INV     gate4258  (.A(II14416), .Z(g5952) ) ;
INV     gate4259  (.A(g97), .Z(g5953) ) ;
INV     gate4260  (.A(g192), .Z(g5954) ) ;
INV     gate4261  (.A(g198), .Z(g5955) ) ;
INV     gate4262  (.A(g204), .Z(g5956) ) ;
INV     gate4263  (.A(g273), .Z(g5957) ) ;
INV     gate4264  (.A(g117), .Z(II14424) ) ;
INV     gate4265  (.A(II14424), .Z(g5958) ) ;
INV     gate4266  (.A(g876), .Z(g5959) ) ;
INV     gate4267  (.A(g882), .Z(g5960) ) ;
INV     gate4268  (.A(g951), .Z(g5961) ) ;
INV     gate4269  (.A(g957), .Z(g5962) ) ;
INV     gate4270  (.A(g1462), .Z(g5963) ) ;
INV     gate4271  (.A(g1506), .Z(g5966) ) ;
INV     gate4272  (.A(g1567), .Z(g5967) ) ;
INV     gate4273  (.A(g1636), .Z(g5968) ) ;
INV     gate4274  (.A(g1642), .Z(g5969) ) ;
INV     gate4275  (.A(g1648), .Z(g5970) ) ;
INV     gate4276  (.A(g2142), .Z(g5971) ) ;
INV     gate4277  (.A(g2195), .Z(g5972) ) ;
INV     gate4278  (.A(g2321), .Z(g5973) ) ;
INV     gate4279  (.A(g2327), .Z(g5974) ) ;
INV     gate4280  (.A(g2333), .Z(g5975) ) ;
INV     gate4281  (.A(g2165), .Z(II14442) ) ;
INV     gate4282  (.A(II14442), .Z(g5976) ) ;
INV     gate4283  (.A(g2612), .Z(g5977) ) ;
INV     gate4284  (.A(g3230), .Z(II14446) ) ;
INV     gate4285  (.A(II14446), .Z(g5978) ) ;
INV     gate4286  (.A(g3224), .Z(II14449) ) ;
INV     gate4287  (.A(II14449), .Z(g5979) ) ;
INV     gate4288  (.A(g201), .Z(g5980) ) ;
INV     gate4289  (.A(g207), .Z(g5981) ) ;
INV     gate4290  (.A(g785), .Z(g5982) ) ;
INV     gate4291  (.A(g879), .Z(g5983) ) ;
INV     gate4292  (.A(g885), .Z(g5984) ) ;
INV     gate4293  (.A(g891), .Z(g5985) ) ;
INV     gate4294  (.A(g960), .Z(g5986) ) ;
INV     gate4295  (.A(g805), .Z(II14459) ) ;
INV     gate4296  (.A(II14459), .Z(g5987) ) ;
INV     gate4297  (.A(g1570), .Z(g5988) ) ;
INV     gate4298  (.A(g1576), .Z(g5989) ) ;
INV     gate4299  (.A(g1645), .Z(g5990) ) ;
INV     gate4300  (.A(g1651), .Z(g5991) ) ;
INV     gate4301  (.A(g2156), .Z(g5992) ) ;
INV     gate4302  (.A(g2200), .Z(g5995) ) ;
INV     gate4303  (.A(g2261), .Z(g5996) ) ;
INV     gate4304  (.A(g2330), .Z(g5997) ) ;
INV     gate4305  (.A(g2336), .Z(g5998) ) ;
INV     gate4306  (.A(g2342), .Z(g5999) ) ;
INV     gate4307  (.A(g3080), .Z(II14472) ) ;
INV     gate4308  (.A(II14472), .Z(g6000) ) ;
INV     gate4309  (.A(g3225), .Z(II14475) ) ;
INV     gate4310  (.A(II14475), .Z(g6014) ) ;
INV     gate4311  (.A(g3213), .Z(II14478) ) ;
INV     gate4312  (.A(II14478), .Z(g6015) ) ;
INV     gate4313  (.A(g210), .Z(g6016) ) ;
INV     gate4314  (.A(g888), .Z(g6017) ) ;
INV     gate4315  (.A(g894), .Z(g6018) ) ;
INV     gate4316  (.A(g1471), .Z(g6019) ) ;
INV     gate4317  (.A(g1573), .Z(g6020) ) ;
INV     gate4318  (.A(g1579), .Z(g6021) ) ;
INV     gate4319  (.A(g1585), .Z(g6022) ) ;
INV     gate4320  (.A(g1654), .Z(g6023) ) ;
INV     gate4321  (.A(g1496), .Z(II14489) ) ;
INV     gate4322  (.A(II14489), .Z(g6024) ) ;
INV     gate4323  (.A(g2264), .Z(g6025) ) ;
INV     gate4324  (.A(g2270), .Z(g6026) ) ;
INV     gate4325  (.A(g2339), .Z(g6027) ) ;
INV     gate4326  (.A(g2345), .Z(g6028) ) ;
INV     gate4327  (.A(g3226), .Z(II14496) ) ;
INV     gate4328  (.A(II14496), .Z(g6029) ) ;
INV     gate4329  (.A(g3214), .Z(II14499) ) ;
INV     gate4330  (.A(II14499), .Z(g6030) ) ;
INV     gate4331  (.A(g471), .Z(II14502) ) ;
INV     gate4332  (.A(II14502), .Z(g6031) ) ;
INV     gate4333  (.A(g897), .Z(g6032) ) ;
INV     gate4334  (.A(g1582), .Z(g6033) ) ;
INV     gate4335  (.A(g1588), .Z(g6034) ) ;
INV     gate4336  (.A(g2165), .Z(g6035) ) ;
INV     gate4337  (.A(g2267), .Z(g6036) ) ;
INV     gate4338  (.A(g2273), .Z(g6037) ) ;
INV     gate4339  (.A(g2279), .Z(g6038) ) ;
INV     gate4340  (.A(g2348), .Z(g6039) ) ;
INV     gate4341  (.A(g2190), .Z(II14513) ) ;
INV     gate4342  (.A(II14513), .Z(g6040) ) ;
INV     gate4343  (.A(g3215), .Z(II14516) ) ;
INV     gate4344  (.A(II14516), .Z(g6041) ) ;
INV     gate4345  (.A(g1158), .Z(II14519) ) ;
INV     gate4346  (.A(II14519), .Z(g6042) ) ;
INV     gate4347  (.A(g1591), .Z(g6043) ) ;
INV     gate4348  (.A(g2276), .Z(g6044) ) ;
INV     gate4349  (.A(g2282), .Z(g6045) ) ;
INV     gate4350  (.A(g1852), .Z(II14525) ) ;
INV     gate4351  (.A(II14525), .Z(g6046) ) ;
INV     gate4352  (.A(g2285), .Z(g6047) ) ;
INV     gate4353  (.A(g3142), .Z(II14529) ) ;
INV     gate4354  (.A(II14529), .Z(g6048) ) ;
INV     gate4355  (.A(g354), .Z(II14532) ) ;
INV     gate4356  (.A(II14532), .Z(g6051) ) ;
INV     gate4357  (.A(g2546), .Z(II14535) ) ;
INV     gate4358  (.A(II14535), .Z(g6052) ) ;
INV     gate4359  (.A(g369), .Z(II14538) ) ;
INV     gate4360  (.A(II14538), .Z(g6053) ) ;
INV     gate4361  (.A(g455), .Z(II14541) ) ;
INV     gate4362  (.A(II14541), .Z(g6054) ) ;
INV     gate4363  (.A(g1041), .Z(II14544) ) ;
INV     gate4364  (.A(II14544), .Z(g6055) ) ;
INV     gate4365  (.A(g384), .Z(II14547) ) ;
INV     gate4366  (.A(II14547), .Z(g6056) ) ;
INV     gate4367  (.A(g458), .Z(II14550) ) ;
INV     gate4368  (.A(II14550), .Z(g6057) ) ;
INV     gate4369  (.A(g1056), .Z(II14553) ) ;
INV     gate4370  (.A(II14553), .Z(g6058) ) ;
INV     gate4371  (.A(g1142), .Z(II14556) ) ;
INV     gate4372  (.A(II14556), .Z(g6059) ) ;
INV     gate4373  (.A(g1735), .Z(II14559) ) ;
INV     gate4374  (.A(II14559), .Z(g6060) ) ;
INV     gate4375  (.A(g398), .Z(II14562) ) ;
INV     gate4376  (.A(II14562), .Z(g6061) ) ;
INV     gate4377  (.A(g461), .Z(II14565) ) ;
INV     gate4378  (.A(II14565), .Z(g6062) ) ;
INV     gate4379  (.A(g1071), .Z(II14568) ) ;
INV     gate4380  (.A(II14568), .Z(g6063) ) ;
INV     gate4381  (.A(g1145), .Z(II14571) ) ;
INV     gate4382  (.A(II14571), .Z(g6064) ) ;
INV     gate4383  (.A(g1750), .Z(II14574) ) ;
INV     gate4384  (.A(II14574), .Z(g6065) ) ;
INV     gate4385  (.A(g1836), .Z(II14577) ) ;
INV     gate4386  (.A(II14577), .Z(g6066) ) ;
INV     gate4387  (.A(g2429), .Z(II14580) ) ;
INV     gate4388  (.A(II14580), .Z(g6067) ) ;
INV     gate4389  (.A(g499), .Z(g6068) ) ;
INV     gate4390  (.A(g465), .Z(II14584) ) ;
INV     gate4391  (.A(II14584), .Z(g6079) ) ;
INV     gate4392  (.A(g1085), .Z(II14587) ) ;
INV     gate4393  (.A(II14587), .Z(g6080) ) ;
INV     gate4394  (.A(g1148), .Z(II14590) ) ;
INV     gate4395  (.A(II14590), .Z(g6081) ) ;
INV     gate4396  (.A(g1765), .Z(II14593) ) ;
INV     gate4397  (.A(II14593), .Z(g6082) ) ;
INV     gate4398  (.A(g1839), .Z(II14596) ) ;
INV     gate4399  (.A(II14596), .Z(g6083) ) ;
INV     gate4400  (.A(g2444), .Z(II14599) ) ;
INV     gate4401  (.A(II14599), .Z(g6084) ) ;
INV     gate4402  (.A(g2530), .Z(II14602) ) ;
INV     gate4403  (.A(II14602), .Z(g6085) ) ;
INV     gate4404  (.A(g468), .Z(II14605) ) ;
INV     gate4405  (.A(II14605), .Z(g6086) ) ;
INV     gate4406  (.A(g1186), .Z(g6087) ) ;
INV     gate4407  (.A(g1152), .Z(II14609) ) ;
INV     gate4408  (.A(II14609), .Z(g6098) ) ;
INV     gate4409  (.A(g1779), .Z(II14612) ) ;
INV     gate4410  (.A(II14612), .Z(g6099) ) ;
INV     gate4411  (.A(g1842), .Z(II14615) ) ;
INV     gate4412  (.A(II14615), .Z(g6100) ) ;
INV     gate4413  (.A(g2459), .Z(II14618) ) ;
INV     gate4414  (.A(II14618), .Z(g6101) ) ;
INV     gate4415  (.A(g2533), .Z(II14621) ) ;
INV     gate4416  (.A(II14621), .Z(g6102) ) ;
INV     gate4417  (.A(g1155), .Z(II14624) ) ;
INV     gate4418  (.A(II14624), .Z(g6103) ) ;
INV     gate4419  (.A(g1880), .Z(g6104) ) ;
INV     gate4420  (.A(g1846), .Z(II14628) ) ;
INV     gate4421  (.A(II14628), .Z(g6115) ) ;
INV     gate4422  (.A(g2473), .Z(II14631) ) ;
INV     gate4423  (.A(II14631), .Z(g6116) ) ;
INV     gate4424  (.A(g2536), .Z(II14634) ) ;
INV     gate4425  (.A(II14634), .Z(g6117) ) ;
INV     gate4426  (.A(g1849), .Z(II14637) ) ;
INV     gate4427  (.A(II14637), .Z(g6118) ) ;
INV     gate4428  (.A(g2574), .Z(g6119) ) ;
INV     gate4429  (.A(g2540), .Z(II14641) ) ;
INV     gate4430  (.A(II14641), .Z(g6130) ) ;
INV     gate4431  (.A(g3142), .Z(II14644) ) ;
INV     gate4432  (.A(II14644), .Z(g6131) ) ;
INV     gate4433  (.A(g2543), .Z(II14647) ) ;
INV     gate4434  (.A(II14647), .Z(g6134) ) ;
INV     gate4435  (.A(g525), .Z(II14650) ) ;
INV     gate4436  (.A(II14650), .Z(g6135) ) ;
INV     gate4437  (.A(g672), .Z(g6136) ) ;
INV     gate4438  (.A(g3220), .Z(II14654) ) ;
INV     gate4439  (.A(II14654), .Z(g6139) ) ;
INV     gate4440  (.A(g524), .Z(g6140) ) ;
INV     gate4441  (.A(g554), .Z(g6141) ) ;
INV     gate4442  (.A(g679), .Z(g6142) ) ;
INV     gate4443  (.A(g1211), .Z(II14660) ) ;
INV     gate4444  (.A(II14660), .Z(g6145) ) ;
INV     gate4445  (.A(g1358), .Z(g6146) ) ;
INV     gate4446  (.A(g3097), .Z(g6149) ) ;
INV     gate4447  (.A(g3147), .Z(II14665) ) ;
INV     gate4448  (.A(II14665), .Z(g6153) ) ;
INV     gate4449  (.A(g3232), .Z(II14668) ) ;
INV     gate4450  (.A(II14668), .Z(g6156) ) ;
INV     gate4451  (.A(g686), .Z(g6157) ) ;
INV     gate4452  (.A(g1210), .Z(g6161) ) ;
INV     gate4453  (.A(g1240), .Z(g6162) ) ;
INV     gate4454  (.A(g1365), .Z(g6163) ) ;
INV     gate4455  (.A(g1905), .Z(II14675) ) ;
INV     gate4456  (.A(II14675), .Z(g6166) ) ;
INV     gate4457  (.A(g2052), .Z(g6167) ) ;
INV     gate4458  (.A(g3098), .Z(g6170) ) ;
INV     gate4459  (.A(g557), .Z(g6173) ) ;
INV     gate4460  (.A(g633), .Z(g6177) ) ;
INV     gate4461  (.A(g692), .Z(g6180) ) ;
INV     gate4462  (.A(g291), .Z(g6183) ) ;
INV     gate4463  (.A(g1372), .Z(g6184) ) ;
INV     gate4464  (.A(g1904), .Z(g6188) ) ;
INV     gate4465  (.A(g1934), .Z(g6189) ) ;
INV     gate4466  (.A(g2059), .Z(g6190) ) ;
INV     gate4467  (.A(g2599), .Z(II14688) ) ;
INV     gate4468  (.A(II14688), .Z(g6193) ) ;
INV     gate4469  (.A(g2746), .Z(g6194) ) ;
INV     gate4470  (.A(g3099), .Z(g6197) ) ;
INV     gate4471  (.A(g542), .Z(g6200) ) ;
INV     gate4472  (.A(g646), .Z(g6201) ) ;
INV     gate4473  (.A(g289), .Z(g6204) ) ;
INV     gate4474  (.A(g1243), .Z(g6205) ) ;
INV     gate4475  (.A(g1319), .Z(g6209) ) ;
INV     gate4476  (.A(g1378), .Z(g6212) ) ;
INV     gate4477  (.A(g978), .Z(g6215) ) ;
INV     gate4478  (.A(g2066), .Z(g6216) ) ;
INV     gate4479  (.A(g2598), .Z(g6220) ) ;
INV     gate4480  (.A(g2628), .Z(g6221) ) ;
INV     gate4481  (.A(g2753), .Z(g6222) ) ;
INV     gate4482  (.A(g2818), .Z(II14704) ) ;
INV     gate4483  (.A(g2818), .Z(g6226) ) ;
INV     gate4484  (.A(g3100), .Z(g6227) ) ;
INV     gate4485  (.A(g3229), .Z(II14709) ) ;
INV     gate4486  (.A(II14709), .Z(g6230) ) ;
INV     gate4487  (.A(g138), .Z(II14712) ) ;
INV     gate4488  (.A(g138), .Z(II14715) ) ;
INV     gate4489  (.A(II14715), .Z(g6232) ) ;
INV     gate4490  (.A(g510), .Z(g6281) ) ;
INV     gate4491  (.A(g640), .Z(g6284) ) ;
INV     gate4492  (.A(g287), .Z(g6288) ) ;
INV     gate4493  (.A(g1228), .Z(g6289) ) ;
INV     gate4494  (.A(g1332), .Z(g6290) ) ;
INV     gate4495  (.A(g976), .Z(g6293) ) ;
INV     gate4496  (.A(g1937), .Z(g6294) ) ;
INV     gate4497  (.A(g2013), .Z(g6298) ) ;
INV     gate4498  (.A(g2072), .Z(g6301) ) ;
INV     gate4499  (.A(g1672), .Z(g6304) ) ;
INV     gate4500  (.A(g2760), .Z(g6305) ) ;
INV     gate4501  (.A(g14), .Z(g6309) ) ;
INV     gate4502  (.A(g3101), .Z(g6310) ) ;
INV     gate4503  (.A(g135), .Z(II14731) ) ;
INV     gate4504  (.A(g135), .Z(II14734) ) ;
INV     gate4505  (.A(II14734), .Z(g6314) ) ;
INV     gate4506  (.A(g653), .Z(g6363) ) ;
INV     gate4507  (.A(g285), .Z(g6367) ) ;
INV     gate4508  (.A(g826), .Z(II14739) ) ;
INV     gate4509  (.A(g826), .Z(II14742) ) ;
INV     gate4510  (.A(II14742), .Z(g6369) ) ;
INV     gate4511  (.A(g1196), .Z(g6418) ) ;
INV     gate4512  (.A(g1326), .Z(g6421) ) ;
INV     gate4513  (.A(g974), .Z(g6425) ) ;
INV     gate4514  (.A(g1922), .Z(g6426) ) ;
INV     gate4515  (.A(g2026), .Z(g6427) ) ;
INV     gate4516  (.A(g1670), .Z(g6430) ) ;
INV     gate4517  (.A(g2631), .Z(g6431) ) ;
INV     gate4518  (.A(g2707), .Z(g6435) ) ;
INV     gate4519  (.A(g2766), .Z(g6438) ) ;
INV     gate4520  (.A(g2366), .Z(g6441) ) ;
INV     gate4521  (.A(g2821), .Z(II14755) ) ;
INV     gate4522  (.A(g2821), .Z(g6443) ) ;
INV     gate4523  (.A(g3102), .Z(g6444) ) ;
INV     gate4524  (.A(g405), .Z(II14760) ) ;
INV     gate4525  (.A(g405), .Z(II14763) ) ;
INV     gate4526  (.A(II14763), .Z(g6448) ) ;
INV     gate4527  (.A(g545), .Z(II14766) ) ;
INV     gate4528  (.A(g545), .Z(II14769) ) ;
INV     gate4529  (.A(II14769), .Z(g6486) ) ;
INV     gate4530  (.A(g544), .Z(g6512) ) ;
INV     gate4531  (.A(g660), .Z(g6513) ) ;
INV     gate4532  (.A(g283), .Z(g6517) ) ;
INV     gate4533  (.A(g823), .Z(II14775) ) ;
INV     gate4534  (.A(g823), .Z(II14778) ) ;
INV     gate4535  (.A(II14778), .Z(g6519) ) ;
INV     gate4536  (.A(g1339), .Z(g6568) ) ;
INV     gate4537  (.A(g972), .Z(g6572) ) ;
INV     gate4538  (.A(g1520), .Z(II14783) ) ;
INV     gate4539  (.A(g1520), .Z(II14786) ) ;
INV     gate4540  (.A(II14786), .Z(g6574) ) ;
INV     gate4541  (.A(g1890), .Z(g6623) ) ;
INV     gate4542  (.A(g2020), .Z(g6626) ) ;
INV     gate4543  (.A(g1668), .Z(g6630) ) ;
INV     gate4544  (.A(g2616), .Z(g6631) ) ;
INV     gate4545  (.A(g2720), .Z(g6632) ) ;
INV     gate4546  (.A(g2364), .Z(g6635) ) ;
INV     gate4547  (.A(g1491), .Z(g6636) ) ;
INV     gate4548  (.A(g5), .Z(g6637) ) ;
INV     gate4549  (.A(g3103), .Z(g6638) ) ;
INV     gate4550  (.A(g113), .Z(g6641) ) ;
INV     gate4551  (.A(g551), .Z(II14799) ) ;
INV     gate4552  (.A(g551), .Z(II14802) ) ;
INV     gate4553  (.A(II14802), .Z(g6643) ) ;
INV     gate4554  (.A(g464), .Z(g6672) ) ;
INV     gate4555  (.A(g458), .Z(g6675) ) ;
INV     gate4556  (.A(g559), .Z(g6676) ) ;
INV     gate4557  (.A(g623), .Z(II14808) ) ;
INV     gate4558  (.A(g623), .Z(II14811) ) ;
INV     gate4559  (.A(II14811), .Z(g6678) ) ;
INV     gate4560  (.A(g666), .Z(g6707) ) ;
INV     gate4561  (.A(g281), .Z(g6711) ) ;
INV     gate4562  (.A(g1092), .Z(II14816) ) ;
INV     gate4563  (.A(g1092), .Z(II14819) ) ;
INV     gate4564  (.A(II14819), .Z(g6713) ) ;
INV     gate4565  (.A(g1231), .Z(II14822) ) ;
INV     gate4566  (.A(g1231), .Z(II14825) ) ;
INV     gate4567  (.A(II14825), .Z(g6751) ) ;
INV     gate4568  (.A(g1230), .Z(g6776) ) ;
INV     gate4569  (.A(g1346), .Z(g6777) ) ;
INV     gate4570  (.A(g970), .Z(g6781) ) ;
INV     gate4571  (.A(g1517), .Z(II14831) ) ;
INV     gate4572  (.A(g1517), .Z(II14834) ) ;
INV     gate4573  (.A(II14834), .Z(g6783) ) ;
INV     gate4574  (.A(g2033), .Z(g6832) ) ;
INV     gate4575  (.A(g1666), .Z(g6836) ) ;
INV     gate4576  (.A(g2214), .Z(II14839) ) ;
INV     gate4577  (.A(g2214), .Z(II14842) ) ;
INV     gate4578  (.A(II14842), .Z(g6838) ) ;
INV     gate4579  (.A(g2584), .Z(g6887) ) ;
INV     gate4580  (.A(g2714), .Z(g6890) ) ;
INV     gate4581  (.A(g2362), .Z(g6894) ) ;
INV     gate4582  (.A(g2824), .Z(II14848) ) ;
INV     gate4583  (.A(g2824), .Z(g6896) ) ;
INV     gate4584  (.A(g1486), .Z(g6897) ) ;
INV     gate4585  (.A(g2993), .Z(g6898) ) ;
INV     gate4586  (.A(g3006), .Z(g6901) ) ;
INV     gate4587  (.A(g3104), .Z(g6905) ) ;
INV     gate4588  (.A(g484), .Z(g6908) ) ;
INV     gate4589  (.A(g626), .Z(II14857) ) ;
INV     gate4590  (.A(g626), .Z(II14860) ) ;
INV     gate4591  (.A(II14860), .Z(g6912) ) ;
INV     gate4592  (.A(g279), .Z(g6942) ) ;
INV     gate4593  (.A(g801), .Z(g6943) ) ;
INV     gate4594  (.A(g1237), .Z(II14865) ) ;
INV     gate4595  (.A(g1237), .Z(II14868) ) ;
INV     gate4596  (.A(II14868), .Z(g6945) ) ;
INV     gate4597  (.A(g1151), .Z(g6974) ) ;
INV     gate4598  (.A(g1145), .Z(g6977) ) ;
INV     gate4599  (.A(g1245), .Z(g6978) ) ;
INV     gate4600  (.A(g1309), .Z(II14874) ) ;
INV     gate4601  (.A(g1309), .Z(II14877) ) ;
INV     gate4602  (.A(II14877), .Z(g6980) ) ;
INV     gate4603  (.A(g1352), .Z(g7009) ) ;
INV     gate4604  (.A(g968), .Z(g7013) ) ;
INV     gate4605  (.A(g1786), .Z(II14882) ) ;
INV     gate4606  (.A(g1786), .Z(II14885) ) ;
INV     gate4607  (.A(II14885), .Z(g7015) ) ;
INV     gate4608  (.A(g1925), .Z(II14888) ) ;
INV     gate4609  (.A(g1925), .Z(II14891) ) ;
INV     gate4610  (.A(II14891), .Z(g7053) ) ;
INV     gate4611  (.A(g1924), .Z(g7078) ) ;
INV     gate4612  (.A(g2040), .Z(g7079) ) ;
INV     gate4613  (.A(g1664), .Z(g7083) ) ;
INV     gate4614  (.A(g2211), .Z(II14897) ) ;
INV     gate4615  (.A(g2211), .Z(II14900) ) ;
INV     gate4616  (.A(II14900), .Z(g7085) ) ;
INV     gate4617  (.A(g2727), .Z(g7134) ) ;
INV     gate4618  (.A(g2360), .Z(g7138) ) ;
INV     gate4619  (.A(g1481), .Z(g7139) ) ;
INV     gate4620  (.A(g2170), .Z(g7140) ) ;
INV     gate4621  (.A(g2195), .Z(g7141) ) ;
INV     gate4622  (.A(g8), .Z(g7142) ) ;
INV     gate4623  (.A(g2998), .Z(g7143) ) ;
INV     gate4624  (.A(g3013), .Z(g7146) ) ;
INV     gate4625  (.A(g3105), .Z(g7149) ) ;
INV     gate4626  (.A(g3136), .Z(g7152) ) ;
INV     gate4627  (.A(g480), .Z(g7153) ) ;
INV     gate4628  (.A(g461), .Z(g7156) ) ;
INV     gate4629  (.A(g453), .Z(g7157) ) ;
INV     gate4630  (.A(g1171), .Z(g7158) ) ;
INV     gate4631  (.A(g1312), .Z(II14917) ) ;
INV     gate4632  (.A(g1312), .Z(II14920) ) ;
INV     gate4633  (.A(II14920), .Z(g7162) ) ;
INV     gate4634  (.A(g966), .Z(g7192) ) ;
INV     gate4635  (.A(g1491), .Z(g7193) ) ;
INV     gate4636  (.A(g1931), .Z(II14925) ) ;
INV     gate4637  (.A(g1931), .Z(II14928) ) ;
INV     gate4638  (.A(II14928), .Z(g7195) ) ;
INV     gate4639  (.A(g1845), .Z(g7224) ) ;
INV     gate4640  (.A(g1839), .Z(g7227) ) ;
INV     gate4641  (.A(g1939), .Z(g7228) ) ;
INV     gate4642  (.A(g2003), .Z(II14934) ) ;
INV     gate4643  (.A(g2003), .Z(II14937) ) ;
INV     gate4644  (.A(II14937), .Z(g7230) ) ;
INV     gate4645  (.A(g2046), .Z(g7259) ) ;
INV     gate4646  (.A(g1662), .Z(g7263) ) ;
INV     gate4647  (.A(g2480), .Z(II14942) ) ;
INV     gate4648  (.A(g2480), .Z(II14945) ) ;
INV     gate4649  (.A(II14945), .Z(g7265) ) ;
INV     gate4650  (.A(g2619), .Z(II14948) ) ;
INV     gate4651  (.A(g2619), .Z(II14951) ) ;
INV     gate4652  (.A(II14951), .Z(g7303) ) ;
INV     gate4653  (.A(g2618), .Z(g7328) ) ;
INV     gate4654  (.A(g2734), .Z(g7329) ) ;
INV     gate4655  (.A(g2358), .Z(g7333) ) ;
INV     gate4656  (.A(g2827), .Z(II14957) ) ;
INV     gate4657  (.A(g2827), .Z(g7335) ) ;
INV     gate4658  (.A(g1476), .Z(g7336) ) ;
INV     gate4659  (.A(g2190), .Z(g7337) ) ;
INV     gate4660  (.A(g3002), .Z(g7338) ) ;
INV     gate4661  (.A(g3024), .Z(g7342) ) ;
INV     gate4662  (.A(g3139), .Z(g7345) ) ;
INV     gate4663  (.A(g97), .Z(g7346) ) ;
INV     gate4664  (.A(g490), .Z(g7347) ) ;
INV     gate4665  (.A(g451), .Z(g7348) ) ;
INV     gate4666  (.A(g1167), .Z(g7349) ) ;
INV     gate4667  (.A(g1148), .Z(g7352) ) ;
INV     gate4668  (.A(g1140), .Z(g7353) ) ;
INV     gate4669  (.A(g1865), .Z(g7354) ) ;
INV     gate4670  (.A(g2006), .Z(II14973) ) ;
INV     gate4671  (.A(g2006), .Z(II14976) ) ;
INV     gate4672  (.A(II14976), .Z(g7358) ) ;
INV     gate4673  (.A(g1660), .Z(g7388) ) ;
INV     gate4674  (.A(g2185), .Z(g7389) ) ;
INV     gate4675  (.A(g2625), .Z(II14981) ) ;
INV     gate4676  (.A(g2625), .Z(II14984) ) ;
INV     gate4677  (.A(II14984), .Z(g7391) ) ;
INV     gate4678  (.A(g2539), .Z(g7420) ) ;
INV     gate4679  (.A(g2533), .Z(g7423) ) ;
INV     gate4680  (.A(g2633), .Z(g7424) ) ;
INV     gate4681  (.A(g2697), .Z(II14990) ) ;
INV     gate4682  (.A(g2697), .Z(II14993) ) ;
INV     gate4683  (.A(II14993), .Z(g7426) ) ;
INV     gate4684  (.A(g2740), .Z(g7455) ) ;
INV     gate4685  (.A(g2356), .Z(g7459) ) ;
INV     gate4686  (.A(g1471), .Z(g7460) ) ;
INV     gate4687  (.A(g2175), .Z(g7461) ) ;
INV     gate4688  (.A(g2912), .Z(g7462) ) ;
INV     gate4689  (.A(g2), .Z(g7465) ) ;
INV     gate4690  (.A(g3010), .Z(g7466) ) ;
INV     gate4691  (.A(g3036), .Z(g7471) ) ;
INV     gate4692  (.A(g493), .Z(g7475) ) ;
INV     gate4693  (.A(g785), .Z(g7476) ) ;
INV     gate4694  (.A(g1177), .Z(g7477) ) ;
INV     gate4695  (.A(g1138), .Z(g7478) ) ;
INV     gate4696  (.A(g1861), .Z(g7479) ) ;
INV     gate4697  (.A(g1842), .Z(g7482) ) ;
INV     gate4698  (.A(g1834), .Z(g7483) ) ;
INV     gate4699  (.A(g2559), .Z(g7484) ) ;
INV     gate4700  (.A(g2700), .Z(II15012) ) ;
INV     gate4701  (.A(g2700), .Z(II15015) ) ;
INV     gate4702  (.A(II15015), .Z(g7488) ) ;
INV     gate4703  (.A(g2354), .Z(g7518) ) ;
INV     gate4704  (.A(g2830), .Z(II15019) ) ;
INV     gate4705  (.A(g2830), .Z(g7520) ) ;
INV     gate4706  (.A(g2200), .Z(g7521) ) ;
INV     gate4707  (.A(g2917), .Z(g7522) ) ;
INV     gate4708  (.A(g3018), .Z(g7527) ) ;
INV     gate4709  (.A(g465), .Z(g7529) ) ;
INV     gate4710  (.A(g496), .Z(g7530) ) ;
INV     gate4711  (.A(g1180), .Z(g7531) ) ;
INV     gate4712  (.A(g1471), .Z(g7532) ) ;
INV     gate4713  (.A(g1871), .Z(g7533) ) ;
INV     gate4714  (.A(g1832), .Z(g7534) ) ;
INV     gate4715  (.A(g2555), .Z(g7535) ) ;
INV     gate4716  (.A(g2536), .Z(g7538) ) ;
INV     gate4717  (.A(g2528), .Z(g7539) ) ;
INV     gate4718  (.A(g1506), .Z(g7540) ) ;
INV     gate4719  (.A(g2180), .Z(g7541) ) ;
INV     gate4720  (.A(g2883), .Z(g7542) ) ;
INV     gate4721  (.A(g2920), .Z(g7545) ) ;
INV     gate4722  (.A(g2990), .Z(g7548) ) ;
INV     gate4723  (.A(g3028), .Z(g7549) ) ;
INV     gate4724  (.A(g3114), .Z(g7553) ) ;
INV     gate4725  (.A(g117), .Z(g7554) ) ;
INV     gate4726  (.A(g1152), .Z(g7555) ) ;
INV     gate4727  (.A(g1183), .Z(g7556) ) ;
INV     gate4728  (.A(g1874), .Z(g7557) ) ;
INV     gate4729  (.A(g2165), .Z(g7558) ) ;
INV     gate4730  (.A(g2565), .Z(g7559) ) ;
INV     gate4731  (.A(g2526), .Z(g7560) ) ;
INV     gate4732  (.A(g1501), .Z(g7561) ) ;
INV     gate4733  (.A(g2888), .Z(g7562) ) ;
INV     gate4734  (.A(g2896), .Z(g7566) ) ;
INV     gate4735  (.A(g3032), .Z(g7570) ) ;
INV     gate4736  (.A(g3120), .Z(g7573) ) ;
INV     gate4737  (.A(g3128), .Z(g7574) ) ;
INV     gate4738  (.A(g468), .Z(g7576) ) ;
INV     gate4739  (.A(g805), .Z(g7577) ) ;
INV     gate4740  (.A(g1846), .Z(g7578) ) ;
INV     gate4741  (.A(g1877), .Z(g7579) ) ;
INV     gate4742  (.A(g2568), .Z(g7580) ) ;
INV     gate4743  (.A(g1496), .Z(g7581) ) ;
INV     gate4744  (.A(g2185), .Z(g7582) ) ;
INV     gate4745  (.A(g2892), .Z(g7583) ) ;
INV     gate4746  (.A(g2903), .Z(g7587) ) ;
INV     gate4747  (.A(g1155), .Z(g7590) ) ;
INV     gate4748  (.A(g1496), .Z(g7591) ) ;
INV     gate4749  (.A(g2540), .Z(g7592) ) ;
INV     gate4750  (.A(g2571), .Z(g7593) ) ;
INV     gate4751  (.A(g2165), .Z(g7594) ) ;
INV     gate4752  (.A(g2900), .Z(g7595) ) ;
INV     gate4753  (.A(g2908), .Z(g7600) ) ;
INV     gate4754  (.A(g3133), .Z(g7603) ) ;
INV     gate4755  (.A(g471), .Z(g7604) ) ;
INV     gate4756  (.A(g1849), .Z(g7605) ) ;
INV     gate4757  (.A(g2190), .Z(g7606) ) ;
INV     gate4758  (.A(g2924), .Z(g7607) ) ;
INV     gate4759  (.A(g312), .Z(g7610) ) ;
INV     gate4760  (.A(g1158), .Z(g7613) ) ;
INV     gate4761  (.A(g2543), .Z(g7614) ) ;
INV     gate4762  (.A(g3123), .Z(g7615) ) ;
INV     gate4763  (.A(g313), .Z(g7616) ) ;
INV     gate4764  (.A(g999), .Z(g7619) ) ;
INV     gate4765  (.A(g1852), .Z(g7622) ) ;
INV     gate4766  (.A(g314), .Z(g7623) ) ;
INV     gate4767  (.A(g315), .Z(g7626) ) ;
INV     gate4768  (.A(g403), .Z(g7629) ) ;
INV     gate4769  (.A(g1000), .Z(g7632) ) ;
INV     gate4770  (.A(g1693), .Z(g7635) ) ;
INV     gate4771  (.A(g2546), .Z(g7638) ) ;
INV     gate4772  (.A(g3094), .Z(g7639) ) ;
INV     gate4773  (.A(g3125), .Z(g7642) ) ;
INV     gate4774  (.A(g316), .Z(g7643) ) ;
INV     gate4775  (.A(g318), .Z(g7646) ) ;
INV     gate4776  (.A(g404), .Z(g7649) ) ;
INV     gate4777  (.A(g1001), .Z(g7652) ) ;
INV     gate4778  (.A(g1002), .Z(g7655) ) ;
INV     gate4779  (.A(g1090), .Z(g7658) ) ;
INV     gate4780  (.A(g1694), .Z(g7661) ) ;
INV     gate4781  (.A(g2387), .Z(g7664) ) ;
INV     gate4782  (.A(g3095), .Z(g7667) ) ;
INV     gate4783  (.A(g317), .Z(g7670) ) ;
INV     gate4784  (.A(g319), .Z(g7673) ) ;
INV     gate4785  (.A(g402), .Z(g7676) ) ;
INV     gate4786  (.A(g1003), .Z(g7679) ) ;
INV     gate4787  (.A(g1005), .Z(g7682) ) ;
INV     gate4788  (.A(g1091), .Z(g7685) ) ;
INV     gate4789  (.A(g1695), .Z(g7688) ) ;
INV     gate4790  (.A(g1696), .Z(g7691) ) ;
INV     gate4791  (.A(g1784), .Z(g7694) ) ;
INV     gate4792  (.A(g2388), .Z(g7697) ) ;
INV     gate4793  (.A(g3096), .Z(g7700) ) ;
INV     gate4794  (.A(g320), .Z(g7703) ) ;
INV     gate4795  (.A(g1004), .Z(g7706) ) ;
INV     gate4796  (.A(g1006), .Z(g7709) ) ;
INV     gate4797  (.A(g1089), .Z(g7712) ) ;
INV     gate4798  (.A(g1697), .Z(g7715) ) ;
INV     gate4799  (.A(g1699), .Z(g7718) ) ;
INV     gate4800  (.A(g1785), .Z(g7721) ) ;
INV     gate4801  (.A(g2389), .Z(g7724) ) ;
INV     gate4802  (.A(g2390), .Z(g7727) ) ;
INV     gate4803  (.A(g2478), .Z(g7730) ) ;
INV     gate4804  (.A(g1007), .Z(g7733) ) ;
INV     gate4805  (.A(g1698), .Z(g7736) ) ;
INV     gate4806  (.A(g1700), .Z(g7739) ) ;
INV     gate4807  (.A(g1783), .Z(g7742) ) ;
INV     gate4808  (.A(g2391), .Z(g7745) ) ;
INV     gate4809  (.A(g2393), .Z(g7748) ) ;
INV     gate4810  (.A(g2479), .Z(g7751) ) ;
INV     gate4811  (.A(g322), .Z(g7754) ) ;
INV     gate4812  (.A(g1701), .Z(g7757) ) ;
INV     gate4813  (.A(g2392), .Z(g7760) ) ;
INV     gate4814  (.A(g2394), .Z(g7763) ) ;
INV     gate4815  (.A(g2477), .Z(g7766) ) ;
INV     gate4816  (.A(g323), .Z(g7769) ) ;
INV     gate4817  (.A(g659), .Z(g7772) ) ;
INV     gate4818  (.A(g1009), .Z(g7776) ) ;
INV     gate4819  (.A(g2395), .Z(g7779) ) ;
INV     gate4820  (.A(g321), .Z(g7782) ) ;
INV     gate4821  (.A(g1010), .Z(g7785) ) ;
INV     gate4822  (.A(g1345), .Z(g7788) ) ;
INV     gate4823  (.A(g1703), .Z(g7792) ) ;
INV     gate4824  (.A(g1008), .Z(g7796) ) ;
INV     gate4825  (.A(g1704), .Z(g7799) ) ;
INV     gate4826  (.A(g2039), .Z(g7802) ) ;
INV     gate4827  (.A(g2397), .Z(g7806) ) ;
INV     gate4828  (.A(g1702), .Z(g7809) ) ;
INV     gate4829  (.A(g2398), .Z(g7812) ) ;
INV     gate4830  (.A(g2733), .Z(g7815) ) ;
INV     gate4831  (.A(g479), .Z(g7819) ) ;
INV     gate4832  (.A(g510), .Z(g7822) ) ;
INV     gate4833  (.A(g2396), .Z(g7823) ) ;
INV     gate4834  (.A(g2987), .Z(g7826) ) ;
INV     gate4835  (.A(g478), .Z(g7827) ) ;
INV     gate4836  (.A(g1166), .Z(g7830) ) ;
INV     gate4837  (.A(g1196), .Z(g7833) ) ;
INV     gate4838  (.A(g2953), .Z(g7834) ) ;
INV     gate4839  (.A(g3044), .Z(g7837) ) ;
INV     gate4840  (.A(g477), .Z(g7838) ) ;
INV     gate4841  (.A(g630), .Z(g7841) ) ;
INV     gate4842  (.A(g1165), .Z(g7842) ) ;
INV     gate4843  (.A(g1860), .Z(g7845) ) ;
INV     gate4844  (.A(g1890), .Z(g7848) ) ;
INV     gate4845  (.A(g2956), .Z(g7849) ) ;
INV     gate4846  (.A(g2981), .Z(g7852) ) ;
INV     gate4847  (.A(g3045), .Z(g7856) ) ;
INV     gate4848  (.A(g3055), .Z(g7857) ) ;
INV     gate4849  (.A(g1164), .Z(g7858) ) ;
INV     gate4850  (.A(g1316), .Z(g7861) ) ;
INV     gate4851  (.A(g1859), .Z(g7862) ) ;
INV     gate4852  (.A(g2554), .Z(g7865) ) ;
INV     gate4853  (.A(g2584), .Z(g7868) ) ;
INV     gate4854  (.A(g2959), .Z(g7869) ) ;
INV     gate4855  (.A(g2874), .Z(g7872) ) ;
INV     gate4856  (.A(g3046), .Z(g7877) ) ;
INV     gate4857  (.A(g3056), .Z(g7878) ) ;
INV     gate4858  (.A(g3065), .Z(g7879) ) ;
INV     gate4859  (.A(g3201), .Z(g7880) ) ;
INV     gate4860  (.A(g1858), .Z(g7888) ) ;
INV     gate4861  (.A(g2010), .Z(g7891) ) ;
INV     gate4862  (.A(g2553), .Z(g7892) ) ;
INV     gate4863  (.A(g3047), .Z(g7897) ) ;
INV     gate4864  (.A(g3057), .Z(g7898) ) ;
INV     gate4865  (.A(g3066), .Z(g7899) ) ;
INV     gate4866  (.A(g3075), .Z(g7900) ) ;
INV     gate4867  (.A(g3151), .Z(II15222) ) ;
INV     gate4868  (.A(II15222), .Z(g7901) ) ;
INV     gate4869  (.A(g488), .Z(g7906) ) ;
INV     gate4870  (.A(g474), .Z(II15226) ) ;
INV     gate4871  (.A(g474), .Z(g7910) ) ;
INV     gate4872  (.A(g499), .Z(II15230) ) ;
INV     gate4873  (.A(II15230), .Z(g7911) ) ;
INV     gate4874  (.A(g2552), .Z(g7912) ) ;
INV     gate4875  (.A(g2704), .Z(g7915) ) ;
INV     gate4876  (.A(g2935), .Z(g7916) ) ;
INV     gate4877  (.A(g2963), .Z(g7919) ) ;
INV     gate4878  (.A(g3048), .Z(g7924) ) ;
INV     gate4879  (.A(g3058), .Z(g7925) ) ;
INV     gate4880  (.A(g3067), .Z(g7926) ) ;
INV     gate4881  (.A(g3076), .Z(g7927) ) ;
INV     gate4882  (.A(g3204), .Z(g7928) ) ;
INV     gate4883  (.A(g2950), .Z(II15256) ) ;
INV     gate4884  (.A(II15256), .Z(g7936) ) ;
INV     gate4885  (.A(g165), .Z(g7949) ) ;
INV     gate4886  (.A(g142), .Z(g7950) ) ;
INV     gate4887  (.A(g487), .Z(g7953) ) ;
INV     gate4888  (.A(g481), .Z(II15262) ) ;
INV     gate4889  (.A(g481), .Z(g7957) ) ;
INV     gate4890  (.A(g1175), .Z(g7958) ) ;
INV     gate4891  (.A(g1161), .Z(II15267) ) ;
INV     gate4892  (.A(g1161), .Z(g7962) ) ;
INV     gate4893  (.A(g1186), .Z(II15271) ) ;
INV     gate4894  (.A(II15271), .Z(g7963) ) ;
INV     gate4895  (.A(g2938), .Z(g7964) ) ;
INV     gate4896  (.A(g2966), .Z(g7967) ) ;
INV     gate4897  (.A(g3049), .Z(g7971) ) ;
INV     gate4898  (.A(g3059), .Z(g7972) ) ;
INV     gate4899  (.A(g3068), .Z(g7973) ) ;
INV     gate4900  (.A(g3077), .Z(g7974) ) ;
INV     gate4901  (.A(g39), .Z(g7975) ) ;
INV     gate4902  (.A(g3109), .Z(II15288) ) ;
INV     gate4903  (.A(II15288), .Z(g7976) ) ;
INV     gate4904  (.A(g3191), .Z(g7989) ) ;
INV     gate4905  (.A(g143), .Z(g7990) ) ;
INV     gate4906  (.A(g145), .Z(g7993) ) ;
INV     gate4907  (.A(g486), .Z(g7996) ) ;
INV     gate4908  (.A(g485), .Z(g7999) ) ;
INV     gate4909  (.A(g853), .Z(g8000) ) ;
INV     gate4910  (.A(g830), .Z(g8001) ) ;
INV     gate4911  (.A(g1174), .Z(g8004) ) ;
INV     gate4912  (.A(g1168), .Z(II15299) ) ;
INV     gate4913  (.A(g1168), .Z(g8008) ) ;
INV     gate4914  (.A(g1869), .Z(g8009) ) ;
INV     gate4915  (.A(g1855), .Z(II15304) ) ;
INV     gate4916  (.A(g1855), .Z(g8013) ) ;
INV     gate4917  (.A(g1880), .Z(II15308) ) ;
INV     gate4918  (.A(II15308), .Z(g8014) ) ;
INV     gate4919  (.A(g2941), .Z(g8015) ) ;
INV     gate4920  (.A(g2969), .Z(g8018) ) ;
INV     gate4921  (.A(g2930), .Z(II15313) ) ;
INV     gate4922  (.A(g2930), .Z(g8022) ) ;
INV     gate4923  (.A(g2842), .Z(II15317) ) ;
INV     gate4924  (.A(g2842), .Z(g8024) ) ;
INV     gate4925  (.A(g3050), .Z(g8025) ) ;
INV     gate4926  (.A(g3060), .Z(g8026) ) ;
INV     gate4927  (.A(g3069), .Z(g8027) ) ;
INV     gate4928  (.A(g3078), .Z(g8028) ) ;
INV     gate4929  (.A(g3083), .Z(g8029) ) ;
INV     gate4930  (.A(g3117), .Z(II15326) ) ;
INV     gate4931  (.A(g3117), .Z(II15329) ) ;
INV     gate4932  (.A(II15329), .Z(g8031) ) ;
INV     gate4933  (.A(g3194), .Z(g8044) ) ;
INV     gate4934  (.A(g3207), .Z(g8045) ) ;
INV     gate4935  (.A(g141), .Z(g8053) ) ;
INV     gate4936  (.A(g146), .Z(g8056) ) ;
INV     gate4937  (.A(g148), .Z(g8059) ) ;
INV     gate4938  (.A(g169), .Z(g8062) ) ;
INV     gate4939  (.A(g831), .Z(g8065) ) ;
INV     gate4940  (.A(g833), .Z(g8068) ) ;
INV     gate4941  (.A(g1173), .Z(g8071) ) ;
INV     gate4942  (.A(g1172), .Z(g8074) ) ;
INV     gate4943  (.A(g1547), .Z(g8075) ) ;
INV     gate4944  (.A(g1524), .Z(g8076) ) ;
INV     gate4945  (.A(g1868), .Z(g8079) ) ;
INV     gate4946  (.A(g1862), .Z(II15345) ) ;
INV     gate4947  (.A(g1862), .Z(g8083) ) ;
INV     gate4948  (.A(g2563), .Z(g8084) ) ;
INV     gate4949  (.A(g2549), .Z(II15350) ) ;
INV     gate4950  (.A(g2549), .Z(g8088) ) ;
INV     gate4951  (.A(g2574), .Z(II15354) ) ;
INV     gate4952  (.A(II15354), .Z(g8089) ) ;
INV     gate4953  (.A(g2944), .Z(g8090) ) ;
INV     gate4954  (.A(g2972), .Z(g8093) ) ;
INV     gate4955  (.A(g2858), .Z(II15359) ) ;
INV     gate4956  (.A(g2858), .Z(g8097) ) ;
INV     gate4957  (.A(g3051), .Z(g8098) ) ;
INV     gate4958  (.A(g3061), .Z(g8099) ) ;
INV     gate4959  (.A(g3070), .Z(g8100) ) ;
INV     gate4960  (.A(g2997), .Z(g8101) ) ;
INV     gate4961  (.A(g27), .Z(g8102) ) ;
INV     gate4962  (.A(g185), .Z(g8103) ) ;
INV     gate4963  (.A(g3129), .Z(II15369) ) ;
INV     gate4964  (.A(g3129), .Z(II15372) ) ;
INV     gate4965  (.A(II15372), .Z(g8107) ) ;
INV     gate4966  (.A(g3197), .Z(g8120) ) ;
INV     gate4967  (.A(g144), .Z(g8123) ) ;
INV     gate4968  (.A(g149), .Z(g8126) ) ;
INV     gate4969  (.A(g151), .Z(g8129) ) ;
INV     gate4970  (.A(g170), .Z(g8132) ) ;
INV     gate4971  (.A(g172), .Z(g8135) ) ;
INV     gate4972  (.A(g829), .Z(g8138) ) ;
INV     gate4973  (.A(g834), .Z(g8141) ) ;
INV     gate4974  (.A(g836), .Z(g8144) ) ;
INV     gate4975  (.A(g857), .Z(g8147) ) ;
INV     gate4976  (.A(g1525), .Z(g8150) ) ;
INV     gate4977  (.A(g1527), .Z(g8153) ) ;
INV     gate4978  (.A(g1867), .Z(g8156) ) ;
INV     gate4979  (.A(g1866), .Z(g8159) ) ;
INV     gate4980  (.A(g2241), .Z(g8160) ) ;
INV     gate4981  (.A(g2218), .Z(g8161) ) ;
INV     gate4982  (.A(g2562), .Z(g8164) ) ;
INV     gate4983  (.A(g2556), .Z(II15392) ) ;
INV     gate4984  (.A(g2556), .Z(g8168) ) ;
INV     gate4985  (.A(g2947), .Z(g8169) ) ;
INV     gate4986  (.A(g2975), .Z(g8172) ) ;
INV     gate4987  (.A(g2845), .Z(II15398) ) ;
INV     gate4988  (.A(g2845), .Z(g8176) ) ;
INV     gate4989  (.A(g3043), .Z(g8177) ) ;
INV     gate4990  (.A(g3052), .Z(g8178) ) ;
INV     gate4991  (.A(g3062), .Z(g8179) ) ;
INV     gate4992  (.A(g3071), .Z(g8180) ) ;
INV     gate4993  (.A(g48), .Z(g8181) ) ;
INV     gate4994  (.A(g3198), .Z(g8182) ) ;
INV     gate4995  (.A(g3188), .Z(g8183) ) ;
INV     gate4996  (.A(g147), .Z(g8191) ) ;
INV     gate4997  (.A(g152), .Z(g8194) ) ;
INV     gate4998  (.A(g154), .Z(g8197) ) ;
INV     gate4999  (.A(g168), .Z(g8200) ) ;
INV     gate5000  (.A(g173), .Z(g8203) ) ;
INV     gate5001  (.A(g175), .Z(g8206) ) ;
INV     gate5002  (.A(g832), .Z(g8209) ) ;
INV     gate5003  (.A(g837), .Z(g8212) ) ;
INV     gate5004  (.A(g839), .Z(g8215) ) ;
INV     gate5005  (.A(g858), .Z(g8218) ) ;
INV     gate5006  (.A(g860), .Z(g8221) ) ;
INV     gate5007  (.A(g1523), .Z(g8224) ) ;
INV     gate5008  (.A(g1528), .Z(g8227) ) ;
INV     gate5009  (.A(g1530), .Z(g8230) ) ;
INV     gate5010  (.A(g1551), .Z(g8233) ) ;
INV     gate5011  (.A(g2219), .Z(g8236) ) ;
INV     gate5012  (.A(g2221), .Z(g8239) ) ;
INV     gate5013  (.A(g2561), .Z(g8242) ) ;
INV     gate5014  (.A(g2560), .Z(g8245) ) ;
INV     gate5015  (.A(g2978), .Z(g8246) ) ;
INV     gate5016  (.A(g2833), .Z(II15429) ) ;
INV     gate5017  (.A(g2833), .Z(g8250) ) ;
INV     gate5018  (.A(g2861), .Z(II15433) ) ;
INV     gate5019  (.A(g2861), .Z(g8252) ) ;
INV     gate5020  (.A(g3053), .Z(g8253) ) ;
INV     gate5021  (.A(g3063), .Z(g8254) ) ;
INV     gate5022  (.A(g3072), .Z(g8255) ) ;
INV     gate5023  (.A(g30), .Z(g8256) ) ;
INV     gate5024  (.A(g3201), .Z(g8257) ) ;
INV     gate5025  (.A(g3235), .Z(II15442) ) ;
INV     gate5026  (.A(g3236), .Z(II15445) ) ;
INV     gate5027  (.A(g3237), .Z(II15448) ) ;
INV     gate5028  (.A(g3238), .Z(II15451) ) ;
INV     gate5029  (.A(g3239), .Z(II15454) ) ;
INV     gate5030  (.A(g3240), .Z(II15457) ) ;
INV     gate5031  (.A(g3241), .Z(II15460) ) ;
INV     gate5032  (.A(g3242), .Z(II15463) ) ;
INV     gate5033  (.A(g3243), .Z(II15466) ) ;
INV     gate5034  (.A(g3244), .Z(II15469) ) ;
INV     gate5035  (.A(g3245), .Z(II15472) ) ;
INV     gate5036  (.A(g3246), .Z(II15475) ) ;
INV     gate5037  (.A(g3247), .Z(II15478) ) ;
INV     gate5038  (.A(g3248), .Z(II15481) ) ;
INV     gate5039  (.A(g3249), .Z(II15484) ) ;
INV     gate5040  (.A(g3250), .Z(II15487) ) ;
INV     gate5041  (.A(g3251), .Z(II15490) ) ;
INV     gate5042  (.A(g3252), .Z(II15493) ) ;
INV     gate5043  (.A(g3253), .Z(g8276) ) ;
INV     gate5044  (.A(g3305), .Z(g8277) ) ;
INV     gate5045  (.A(g3337), .Z(g8278) ) ;
INV     gate5046  (.A(g7911), .Z(II15499) ) ;
INV     gate5047  (.A(g3365), .Z(g8285) ) ;
INV     gate5048  (.A(g3461), .Z(g8286) ) ;
INV     gate5049  (.A(g3493), .Z(g8287) ) ;
INV     gate5050  (.A(g7963), .Z(II15505) ) ;
INV     gate5051  (.A(g3521), .Z(g8294) ) ;
INV     gate5052  (.A(g3617), .Z(g8295) ) ;
INV     gate5053  (.A(g3649), .Z(g8296) ) ;
INV     gate5054  (.A(g8014), .Z(II15511) ) ;
INV     gate5055  (.A(g3677), .Z(g8303) ) ;
INV     gate5056  (.A(g3773), .Z(g8304) ) ;
INV     gate5057  (.A(g3805), .Z(g8305) ) ;
INV     gate5058  (.A(g8089), .Z(II15517) ) ;
INV     gate5059  (.A(g3833), .Z(g8312) ) ;
INV     gate5060  (.A(g3897), .Z(g8313) ) ;
INV     gate5061  (.A(g3919), .Z(g8317) ) ;
INV     gate5062  (.A(g3254), .Z(II15523) ) ;
INV     gate5063  (.A(II15523), .Z(g8321) ) ;
INV     gate5064  (.A(g6314), .Z(II15526) ) ;
INV     gate5065  (.A(II15526), .Z(g8324) ) ;
INV     gate5066  (.A(g3410), .Z(II15532) ) ;
INV     gate5067  (.A(II15532), .Z(g8330) ) ;
INV     gate5068  (.A(g6519), .Z(II15535) ) ;
INV     gate5069  (.A(II15535), .Z(g8333) ) ;
INV     gate5070  (.A(g6369), .Z(II15538) ) ;
INV     gate5071  (.A(II15538), .Z(g8336) ) ;
INV     gate5072  (.A(g3410), .Z(II15543) ) ;
INV     gate5073  (.A(II15543), .Z(g8341) ) ;
INV     gate5074  (.A(g6783), .Z(II15546) ) ;
INV     gate5075  (.A(II15546), .Z(g8344) ) ;
INV     gate5076  (.A(g6574), .Z(II15549) ) ;
INV     gate5077  (.A(II15549), .Z(g8347) ) ;
INV     gate5078  (.A(g3566), .Z(II15553) ) ;
INV     gate5079  (.A(II15553), .Z(g8351) ) ;
INV     gate5080  (.A(g6783), .Z(II15556) ) ;
INV     gate5081  (.A(II15556), .Z(g8354) ) ;
INV     gate5082  (.A(g7015), .Z(II15559) ) ;
INV     gate5083  (.A(II15559), .Z(g8357) ) ;
INV     gate5084  (.A(g5778), .Z(II15562) ) ;
INV     gate5085  (.A(II15562), .Z(g8360) ) ;
INV     gate5086  (.A(g6838), .Z(II15565) ) ;
INV     gate5087  (.A(II15565), .Z(g8363) ) ;
INV     gate5088  (.A(g3722), .Z(II15568) ) ;
INV     gate5089  (.A(II15568), .Z(g8366) ) ;
INV     gate5090  (.A(g7085), .Z(II15571) ) ;
INV     gate5091  (.A(II15571), .Z(g8369) ) ;
INV     gate5092  (.A(g6838), .Z(II15574) ) ;
INV     gate5093  (.A(II15574), .Z(g8372) ) ;
INV     gate5094  (.A(g7265), .Z(II15577) ) ;
INV     gate5095  (.A(II15577), .Z(g8375) ) ;
INV     gate5096  (.A(g5837), .Z(II15580) ) ;
INV     gate5097  (.A(II15580), .Z(g8378) ) ;
INV     gate5098  (.A(g3254), .Z(II15584) ) ;
INV     gate5099  (.A(II15584), .Z(g8382) ) ;
INV     gate5100  (.A(g3410), .Z(II15590) ) ;
INV     gate5101  (.A(II15590), .Z(g8388) ) ;
INV     gate5102  (.A(g6519), .Z(II15593) ) ;
INV     gate5103  (.A(II15593), .Z(g8391) ) ;
INV     gate5104  (.A(g3566), .Z(II15599) ) ;
INV     gate5105  (.A(II15599), .Z(g8397) ) ;
INV     gate5106  (.A(g6783), .Z(II15602) ) ;
INV     gate5107  (.A(II15602), .Z(g8400) ) ;
INV     gate5108  (.A(g6574), .Z(II15605) ) ;
INV     gate5109  (.A(II15605), .Z(g8403) ) ;
INV     gate5110  (.A(g3566), .Z(II15610) ) ;
INV     gate5111  (.A(II15610), .Z(g8408) ) ;
INV     gate5112  (.A(g7085), .Z(II15613) ) ;
INV     gate5113  (.A(II15613), .Z(g8411) ) ;
INV     gate5114  (.A(g6838), .Z(II15616) ) ;
INV     gate5115  (.A(II15616), .Z(g8414) ) ;
INV     gate5116  (.A(g3722), .Z(II15620) ) ;
INV     gate5117  (.A(II15620), .Z(g8418) ) ;
INV     gate5118  (.A(g7085), .Z(II15623) ) ;
INV     gate5119  (.A(II15623), .Z(g8421) ) ;
INV     gate5120  (.A(g7265), .Z(II15626) ) ;
INV     gate5121  (.A(II15626), .Z(g8424) ) ;
INV     gate5122  (.A(g5837), .Z(II15629) ) ;
INV     gate5123  (.A(II15629), .Z(g8427) ) ;
INV     gate5124  (.A(g3410), .Z(II15636) ) ;
INV     gate5125  (.A(II15636), .Z(g8434) ) ;
INV     gate5126  (.A(g3566), .Z(II15642) ) ;
INV     gate5127  (.A(II15642), .Z(g8440) ) ;
INV     gate5128  (.A(g6783), .Z(II15645) ) ;
INV     gate5129  (.A(II15645), .Z(g8443) ) ;
INV     gate5130  (.A(g3722), .Z(II15651) ) ;
INV     gate5131  (.A(II15651), .Z(g8449) ) ;
INV     gate5132  (.A(g7085), .Z(II15654) ) ;
INV     gate5133  (.A(II15654), .Z(g8452) ) ;
INV     gate5134  (.A(g6838), .Z(II15657) ) ;
INV     gate5135  (.A(II15657), .Z(g8455) ) ;
INV     gate5136  (.A(g3722), .Z(II15662) ) ;
INV     gate5137  (.A(II15662), .Z(g8460) ) ;
INV     gate5138  (.A(g3566), .Z(II15671) ) ;
INV     gate5139  (.A(II15671), .Z(g8469) ) ;
INV     gate5140  (.A(g3722), .Z(II15677) ) ;
INV     gate5141  (.A(II15677), .Z(g8475) ) ;
INV     gate5142  (.A(g7085), .Z(II15680) ) ;
INV     gate5143  (.A(II15680), .Z(g8478) ) ;
INV     gate5144  (.A(g3722), .Z(II15696) ) ;
INV     gate5145  (.A(II15696), .Z(g8494) ) ;
INV     gate5146  (.A(g6139), .Z(g8514) ) ;
INV     gate5147  (.A(g6156), .Z(g8530) ) ;
INV     gate5148  (.A(g6230), .Z(g8568) ) ;
INV     gate5149  (.A(g6000), .Z(II15771) ) ;
INV     gate5150  (.A(II15771), .Z(g8569) ) ;
INV     gate5151  (.A(g6000), .Z(II15779) ) ;
INV     gate5152  (.A(II15779), .Z(g8575) ) ;
INV     gate5153  (.A(g6000), .Z(II15784) ) ;
INV     gate5154  (.A(II15784), .Z(g8578) ) ;
INV     gate5155  (.A(g6000), .Z(II15787) ) ;
INV     gate5156  (.A(II15787), .Z(g8579) ) ;
INV     gate5157  (.A(g6281), .Z(g8580) ) ;
INV     gate5158  (.A(g6418), .Z(g8587) ) ;
INV     gate5159  (.A(g6623), .Z(g8594) ) ;
INV     gate5160  (.A(g3338), .Z(II15794) ) ;
INV     gate5161  (.A(II15794), .Z(g8602) ) ;
INV     gate5162  (.A(g6887), .Z(g8605) ) ;
INV     gate5163  (.A(g3494), .Z(II15800) ) ;
INV     gate5164  (.A(II15800), .Z(g8614) ) ;
INV     gate5165  (.A(g8107), .Z(II15803) ) ;
INV     gate5166  (.A(II15803), .Z(g8617) ) ;
INV     gate5167  (.A(g5550), .Z(II15806) ) ;
INV     gate5168  (.A(II15806), .Z(g8620) ) ;
INV     gate5169  (.A(g3338), .Z(II15810) ) ;
INV     gate5170  (.A(II15810), .Z(g8622) ) ;
INV     gate5171  (.A(g3650), .Z(II15815) ) ;
INV     gate5172  (.A(II15815), .Z(g8627) ) ;
INV     gate5173  (.A(g5596), .Z(II15818) ) ;
INV     gate5174  (.A(II15818), .Z(g8630) ) ;
INV     gate5175  (.A(g3494), .Z(II15822) ) ;
INV     gate5176  (.A(II15822), .Z(g8632) ) ;
INV     gate5177  (.A(g3806), .Z(II15827) ) ;
INV     gate5178  (.A(II15827), .Z(g8637) ) ;
INV     gate5179  (.A(g8031), .Z(II15830) ) ;
INV     gate5180  (.A(II15830), .Z(g8640) ) ;
INV     gate5181  (.A(g3338), .Z(II15833) ) ;
INV     gate5182  (.A(II15833), .Z(g8643) ) ;
INV     gate5183  (.A(g3366), .Z(II15836) ) ;
INV     gate5184  (.A(II15836), .Z(g8646) ) ;
INV     gate5185  (.A(g5613), .Z(II15839) ) ;
INV     gate5186  (.A(II15839), .Z(g8649) ) ;
INV     gate5187  (.A(g3650), .Z(II15843) ) ;
INV     gate5188  (.A(II15843), .Z(g8651) ) ;
INV     gate5189  (.A(g3878), .Z(II15847) ) ;
INV     gate5190  (.A(II15847), .Z(g8655) ) ;
INV     gate5191  (.A(g5627), .Z(II15850) ) ;
INV     gate5192  (.A(II15850), .Z(g8658) ) ;
INV     gate5193  (.A(g3494), .Z(II15853) ) ;
INV     gate5194  (.A(II15853), .Z(g8659) ) ;
INV     gate5195  (.A(g3522), .Z(II15856) ) ;
INV     gate5196  (.A(II15856), .Z(g8662) ) ;
INV     gate5197  (.A(g5638), .Z(II15859) ) ;
INV     gate5198  (.A(II15859), .Z(g8665) ) ;
INV     gate5199  (.A(g3806), .Z(II15863) ) ;
INV     gate5200  (.A(II15863), .Z(g8667) ) ;
INV     gate5201  (.A(g3878), .Z(II15866) ) ;
INV     gate5202  (.A(II15866), .Z(g8670) ) ;
INV     gate5203  (.A(g7976), .Z(II15869) ) ;
INV     gate5204  (.A(II15869), .Z(g8673) ) ;
INV     gate5205  (.A(g5655), .Z(II15873) ) ;
INV     gate5206  (.A(II15873), .Z(g8677) ) ;
INV     gate5207  (.A(g3650), .Z(II15876) ) ;
INV     gate5208  (.A(II15876), .Z(g8678) ) ;
INV     gate5209  (.A(g3678), .Z(II15879) ) ;
INV     gate5210  (.A(II15879), .Z(g8681) ) ;
INV     gate5211  (.A(g3878), .Z(II15882) ) ;
INV     gate5212  (.A(II15882), .Z(g8684) ) ;
INV     gate5213  (.A(g5693), .Z(II15887) ) ;
INV     gate5214  (.A(II15887), .Z(g8689) ) ;
INV     gate5215  (.A(g3806), .Z(II15890) ) ;
INV     gate5216  (.A(II15890), .Z(g8690) ) ;
INV     gate5217  (.A(g3834), .Z(II15893) ) ;
INV     gate5218  (.A(II15893), .Z(g8693) ) ;
INV     gate5219  (.A(g3878), .Z(II15896) ) ;
INV     gate5220  (.A(II15896), .Z(g8696) ) ;
INV     gate5221  (.A(g5626), .Z(II15899) ) ;
INV     gate5222  (.A(II15899), .Z(g8699) ) ;
INV     gate5223  (.A(g6486), .Z(II15902) ) ;
INV     gate5224  (.A(II15902), .Z(g8700) ) ;
INV     gate5225  (.A(g5745), .Z(II15909) ) ;
INV     gate5226  (.A(II15909), .Z(g8707) ) ;
INV     gate5227  (.A(g3878), .Z(II15912) ) ;
INV     gate5228  (.A(II15912), .Z(g8708) ) ;
INV     gate5229  (.A(g3878), .Z(II15915) ) ;
INV     gate5230  (.A(II15915), .Z(g8711) ) ;
INV     gate5231  (.A(g6643), .Z(II15918) ) ;
INV     gate5232  (.A(II15918), .Z(g8714) ) ;
INV     gate5233  (.A(g5654), .Z(II15922) ) ;
INV     gate5234  (.A(II15922), .Z(g8718) ) ;
INV     gate5235  (.A(g6751), .Z(II15925) ) ;
INV     gate5236  (.A(II15925), .Z(g8719) ) ;
INV     gate5237  (.A(g5423), .Z(II15932) ) ;
INV     gate5238  (.A(II15932), .Z(g8726) ) ;
INV     gate5239  (.A(g3878), .Z(II15935) ) ;
INV     gate5240  (.A(II15935), .Z(g8745) ) ;
INV     gate5241  (.A(g3338), .Z(II15938) ) ;
INV     gate5242  (.A(II15938), .Z(g8748) ) ;
INV     gate5243  (.A(g6945), .Z(II15942) ) ;
INV     gate5244  (.A(II15942), .Z(g8752) ) ;
INV     gate5245  (.A(g5692), .Z(II15946) ) ;
INV     gate5246  (.A(II15946), .Z(g8756) ) ;
INV     gate5247  (.A(g7053), .Z(II15949) ) ;
INV     gate5248  (.A(II15949), .Z(g8757) ) ;
INV     gate5249  (.A(g3878), .Z(II15955) ) ;
INV     gate5250  (.A(II15955), .Z(g8763) ) ;
INV     gate5251  (.A(g3878), .Z(II15958) ) ;
INV     gate5252  (.A(II15958), .Z(g8766) ) ;
INV     gate5253  (.A(g6051), .Z(II15961) ) ;
INV     gate5254  (.A(II15961), .Z(g8769) ) ;
INV     gate5255  (.A(g7554), .Z(II15964) ) ;
INV     gate5256  (.A(II15964), .Z(g8770) ) ;
INV     gate5257  (.A(g3494), .Z(II15967) ) ;
INV     gate5258  (.A(II15967), .Z(g8771) ) ;
INV     gate5259  (.A(g7195), .Z(II15971) ) ;
INV     gate5260  (.A(II15971), .Z(g8775) ) ;
INV     gate5261  (.A(g5744), .Z(II15975) ) ;
INV     gate5262  (.A(II15975), .Z(g8779) ) ;
INV     gate5263  (.A(g7303), .Z(II15978) ) ;
INV     gate5264  (.A(II15978), .Z(g8780) ) ;
INV     gate5265  (.A(g3878), .Z(II15983) ) ;
INV     gate5266  (.A(II15983), .Z(g8785) ) ;
INV     gate5267  (.A(g3878), .Z(II15986) ) ;
INV     gate5268  (.A(II15986), .Z(g8788) ) ;
INV     gate5269  (.A(g6053), .Z(II15989) ) ;
INV     gate5270  (.A(II15989), .Z(g8791) ) ;
INV     gate5271  (.A(g6055), .Z(II15992) ) ;
INV     gate5272  (.A(II15992), .Z(g8792) ) ;
INV     gate5273  (.A(g7577), .Z(II15995) ) ;
INV     gate5274  (.A(II15995), .Z(g8793) ) ;
INV     gate5275  (.A(g3650), .Z(II15998) ) ;
INV     gate5276  (.A(II15998), .Z(g8794) ) ;
INV     gate5277  (.A(g7391), .Z(II16002) ) ;
INV     gate5278  (.A(II16002), .Z(g8798) ) ;
INV     gate5279  (.A(g3878), .Z(II16006) ) ;
INV     gate5280  (.A(II16006), .Z(g8802) ) ;
INV     gate5281  (.A(g3878), .Z(II16009) ) ;
INV     gate5282  (.A(II16009), .Z(g8805) ) ;
INV     gate5283  (.A(g5390), .Z(II16012) ) ;
INV     gate5284  (.A(II16012), .Z(g8808) ) ;
INV     gate5285  (.A(g6056), .Z(II16015) ) ;
INV     gate5286  (.A(II16015), .Z(g8809) ) ;
INV     gate5287  (.A(g6058), .Z(II16018) ) ;
INV     gate5288  (.A(II16018), .Z(g8810) ) ;
INV     gate5289  (.A(g6060), .Z(II16021) ) ;
INV     gate5290  (.A(II16021), .Z(g8811) ) ;
INV     gate5291  (.A(g7591), .Z(II16024) ) ;
INV     gate5292  (.A(II16024), .Z(g8812) ) ;
INV     gate5293  (.A(g3806), .Z(II16027) ) ;
INV     gate5294  (.A(II16027), .Z(g8813) ) ;
INV     gate5295  (.A(g3878), .Z(II16031) ) ;
INV     gate5296  (.A(II16031), .Z(g8817) ) ;
INV     gate5297  (.A(g5396), .Z(II16034) ) ;
INV     gate5298  (.A(II16034), .Z(g8820) ) ;
INV     gate5299  (.A(g6061), .Z(II16037) ) ;
INV     gate5300  (.A(II16037), .Z(g8821) ) ;
INV     gate5301  (.A(g4602), .Z(g8822) ) ;
INV     gate5302  (.A(g6486), .Z(II16041) ) ;
INV     gate5303  (.A(II16041), .Z(g8823) ) ;
INV     gate5304  (.A(g5397), .Z(II16044) ) ;
INV     gate5305  (.A(II16044), .Z(g8824) ) ;
INV     gate5306  (.A(g6063), .Z(II16047) ) ;
INV     gate5307  (.A(II16047), .Z(g8825) ) ;
INV     gate5308  (.A(g6065), .Z(II16050) ) ;
INV     gate5309  (.A(II16050), .Z(g8826) ) ;
INV     gate5310  (.A(g6067), .Z(II16053) ) ;
INV     gate5311  (.A(II16053), .Z(g8827) ) ;
INV     gate5312  (.A(g7606), .Z(II16056) ) ;
INV     gate5313  (.A(II16056), .Z(g8828) ) ;
INV     gate5314  (.A(g3878), .Z(II16059) ) ;
INV     gate5315  (.A(II16059), .Z(g8829) ) ;
INV     gate5316  (.A(g3900), .Z(II16062) ) ;
INV     gate5317  (.A(II16062), .Z(g8832) ) ;
INV     gate5318  (.A(g7936), .Z(II16065) ) ;
INV     gate5319  (.A(II16065), .Z(g8835) ) ;
INV     gate5320  (.A(g5438), .Z(II16068) ) ;
INV     gate5321  (.A(II16068), .Z(g8836) ) ;
INV     gate5322  (.A(g5395), .Z(II16071) ) ;
INV     gate5323  (.A(II16071), .Z(g8839) ) ;
INV     gate5324  (.A(g5399), .Z(II16074) ) ;
INV     gate5325  (.A(II16074), .Z(g8840) ) ;
INV     gate5326  (.A(g6086), .Z(II16079) ) ;
INV     gate5327  (.A(II16079), .Z(g8843) ) ;
INV     gate5328  (.A(g5401), .Z(II16082) ) ;
INV     gate5329  (.A(II16082), .Z(g8844) ) ;
INV     gate5330  (.A(g6080), .Z(II16085) ) ;
INV     gate5331  (.A(II16085), .Z(g8845) ) ;
INV     gate5332  (.A(g4779), .Z(g8846) ) ;
INV     gate5333  (.A(g6751), .Z(II16089) ) ;
INV     gate5334  (.A(II16089), .Z(g8847) ) ;
INV     gate5335  (.A(g5402), .Z(II16092) ) ;
INV     gate5336  (.A(II16092), .Z(g8850) ) ;
INV     gate5337  (.A(g6082), .Z(II16095) ) ;
INV     gate5338  (.A(II16095), .Z(g8851) ) ;
INV     gate5339  (.A(g6084), .Z(II16098) ) ;
INV     gate5340  (.A(II16098), .Z(g8852) ) ;
INV     gate5341  (.A(g3878), .Z(II16101) ) ;
INV     gate5342  (.A(II16101), .Z(g8853) ) ;
INV     gate5343  (.A(g6448), .Z(II16104) ) ;
INV     gate5344  (.A(II16104), .Z(g8856) ) ;
INV     gate5345  (.A(g5398), .Z(II16107) ) ;
INV     gate5346  (.A(II16107), .Z(g8859) ) ;
INV     gate5347  (.A(g5404), .Z(II16110) ) ;
INV     gate5348  (.A(II16110), .Z(g8860) ) ;
INV     gate5349  (.A(g7936), .Z(II16114) ) ;
INV     gate5350  (.A(II16114), .Z(g8862) ) ;
INV     gate5351  (.A(g5473), .Z(II16117) ) ;
INV     gate5352  (.A(II16117), .Z(g8863) ) ;
INV     gate5353  (.A(g5400), .Z(II16120) ) ;
INV     gate5354  (.A(II16120), .Z(g8866) ) ;
INV     gate5355  (.A(g5406), .Z(II16123) ) ;
INV     gate5356  (.A(II16123), .Z(g8867) ) ;
INV     gate5357  (.A(g6103), .Z(II16128) ) ;
INV     gate5358  (.A(II16128), .Z(g8870) ) ;
INV     gate5359  (.A(g5408), .Z(II16131) ) ;
INV     gate5360  (.A(II16131), .Z(g8871) ) ;
INV     gate5361  (.A(g6099), .Z(II16134) ) ;
INV     gate5362  (.A(II16134), .Z(g8872) ) ;
INV     gate5363  (.A(g4955), .Z(g8873) ) ;
INV     gate5364  (.A(g7053), .Z(II16138) ) ;
INV     gate5365  (.A(II16138), .Z(g8874) ) ;
INV     gate5366  (.A(g5409), .Z(II16141) ) ;
INV     gate5367  (.A(II16141), .Z(g8877) ) ;
INV     gate5368  (.A(g6101), .Z(II16144) ) ;
INV     gate5369  (.A(II16144), .Z(g8878) ) ;
INV     gate5370  (.A(g3878), .Z(II16147) ) ;
INV     gate5371  (.A(II16147), .Z(g8879) ) ;
INV     gate5372  (.A(g3900), .Z(II16150) ) ;
INV     gate5373  (.A(II16150), .Z(g8882) ) ;
INV     gate5374  (.A(g3306), .Z(II16153) ) ;
INV     gate5375  (.A(II16153), .Z(g8885) ) ;
INV     gate5376  (.A(g5438), .Z(II16156) ) ;
INV     gate5377  (.A(II16156), .Z(g8888) ) ;
INV     gate5378  (.A(g5403), .Z(II16159) ) ;
INV     gate5379  (.A(II16159), .Z(g8891) ) ;
INV     gate5380  (.A(g6031), .Z(II16163) ) ;
INV     gate5381  (.A(II16163), .Z(g8893) ) ;
INV     gate5382  (.A(g6713), .Z(II16166) ) ;
INV     gate5383  (.A(II16166), .Z(g8894) ) ;
INV     gate5384  (.A(g5405), .Z(II16169) ) ;
INV     gate5385  (.A(II16169), .Z(g8897) ) ;
INV     gate5386  (.A(g5413), .Z(II16172) ) ;
INV     gate5387  (.A(II16172), .Z(g8898) ) ;
INV     gate5388  (.A(g7936), .Z(II16176) ) ;
INV     gate5389  (.A(II16176), .Z(g8900) ) ;
INV     gate5390  (.A(g5512), .Z(II16179) ) ;
INV     gate5391  (.A(II16179), .Z(g8901) ) ;
INV     gate5392  (.A(g5407), .Z(II16182) ) ;
INV     gate5393  (.A(II16182), .Z(g8904) ) ;
INV     gate5394  (.A(g5415), .Z(II16185) ) ;
INV     gate5395  (.A(II16185), .Z(g8905) ) ;
INV     gate5396  (.A(g6118), .Z(II16190) ) ;
INV     gate5397  (.A(II16190), .Z(g8908) ) ;
INV     gate5398  (.A(g5417), .Z(II16193) ) ;
INV     gate5399  (.A(II16193), .Z(g8909) ) ;
INV     gate5400  (.A(g6116), .Z(II16196) ) ;
INV     gate5401  (.A(II16196), .Z(g8910) ) ;
INV     gate5402  (.A(g5114), .Z(g8911) ) ;
INV     gate5403  (.A(g7303), .Z(II16200) ) ;
INV     gate5404  (.A(II16200), .Z(g8912) ) ;
INV     gate5405  (.A(g3878), .Z(II16203) ) ;
INV     gate5406  (.A(II16203), .Z(g8915) ) ;
INV     gate5407  (.A(g6448), .Z(II16206) ) ;
INV     gate5408  (.A(II16206), .Z(g8918) ) ;
INV     gate5409  (.A(g5438), .Z(II16209) ) ;
INV     gate5410  (.A(II16209), .Z(g8921) ) ;
INV     gate5411  (.A(g5411), .Z(II16212) ) ;
INV     gate5412  (.A(II16212), .Z(g8924) ) ;
INV     gate5413  (.A(g3462), .Z(II16215) ) ;
INV     gate5414  (.A(II16215), .Z(g8925) ) ;
INV     gate5415  (.A(g5473), .Z(II16218) ) ;
INV     gate5416  (.A(II16218), .Z(g8928) ) ;
INV     gate5417  (.A(g5412), .Z(II16221) ) ;
INV     gate5418  (.A(II16221), .Z(g8931) ) ;
INV     gate5419  (.A(g6042), .Z(II16225) ) ;
INV     gate5420  (.A(II16225), .Z(g8933) ) ;
INV     gate5421  (.A(g7015), .Z(II16228) ) ;
INV     gate5422  (.A(II16228), .Z(g8934) ) ;
INV     gate5423  (.A(g5414), .Z(II16231) ) ;
INV     gate5424  (.A(II16231), .Z(g8937) ) ;
INV     gate5425  (.A(g5420), .Z(II16234) ) ;
INV     gate5426  (.A(II16234), .Z(g8938) ) ;
INV     gate5427  (.A(g7936), .Z(II16238) ) ;
INV     gate5428  (.A(II16238), .Z(g8940) ) ;
INV     gate5429  (.A(g5556), .Z(II16241) ) ;
INV     gate5430  (.A(II16241), .Z(g8941) ) ;
INV     gate5431  (.A(g5416), .Z(II16244) ) ;
INV     gate5432  (.A(II16244), .Z(g8944) ) ;
INV     gate5433  (.A(g5422), .Z(II16247) ) ;
INV     gate5434  (.A(II16247), .Z(g8945) ) ;
INV     gate5435  (.A(g6134), .Z(II16252) ) ;
INV     gate5436  (.A(II16252), .Z(g8948) ) ;
INV     gate5437  (.A(g3900), .Z(II16255) ) ;
INV     gate5438  (.A(II16255), .Z(g8949) ) ;
INV     gate5439  (.A(g3306), .Z(II16258) ) ;
INV     gate5440  (.A(II16258), .Z(g8952) ) ;
INV     gate5441  (.A(g6448), .Z(II16261) ) ;
INV     gate5442  (.A(II16261), .Z(g8955) ) ;
INV     gate5443  (.A(g6713), .Z(II16264) ) ;
INV     gate5444  (.A(II16264), .Z(g8958) ) ;
INV     gate5445  (.A(g5473), .Z(II16267) ) ;
INV     gate5446  (.A(II16267), .Z(g8961) ) ;
INV     gate5447  (.A(g5418), .Z(II16270) ) ;
INV     gate5448  (.A(II16270), .Z(g8964) ) ;
INV     gate5449  (.A(g3618), .Z(II16273) ) ;
INV     gate5450  (.A(II16273), .Z(g8965) ) ;
INV     gate5451  (.A(g5512), .Z(II16276) ) ;
INV     gate5452  (.A(II16276), .Z(g8968) ) ;
INV     gate5453  (.A(g5419), .Z(II16279) ) ;
INV     gate5454  (.A(II16279), .Z(g8971) ) ;
INV     gate5455  (.A(g6046), .Z(II16283) ) ;
INV     gate5456  (.A(II16283), .Z(g8973) ) ;
INV     gate5457  (.A(g7265), .Z(II16286) ) ;
INV     gate5458  (.A(II16286), .Z(g8974) ) ;
INV     gate5459  (.A(g5421), .Z(II16289) ) ;
INV     gate5460  (.A(II16289), .Z(g8977) ) ;
INV     gate5461  (.A(g5426), .Z(II16292) ) ;
INV     gate5462  (.A(II16292), .Z(g8978) ) ;
INV     gate5463  (.A(g3306), .Z(II16296) ) ;
INV     gate5464  (.A(II16296), .Z(g8980) ) ;
INV     gate5465  (.A(g6486), .Z(g8983) ) ;
INV     gate5466  (.A(g3462), .Z(II16300) ) ;
INV     gate5467  (.A(II16300), .Z(g8984) ) ;
INV     gate5468  (.A(g6713), .Z(II16303) ) ;
INV     gate5469  (.A(II16303), .Z(g8987) ) ;
INV     gate5470  (.A(g7015), .Z(II16306) ) ;
INV     gate5471  (.A(II16306), .Z(g8990) ) ;
INV     gate5472  (.A(g5512), .Z(II16309) ) ;
INV     gate5473  (.A(II16309), .Z(g8993) ) ;
INV     gate5474  (.A(g5424), .Z(II16312) ) ;
INV     gate5475  (.A(II16312), .Z(g8996) ) ;
INV     gate5476  (.A(g3774), .Z(II16315) ) ;
INV     gate5477  (.A(II16315), .Z(g8997) ) ;
INV     gate5478  (.A(g5556), .Z(II16318) ) ;
INV     gate5479  (.A(II16318), .Z(g9000) ) ;
INV     gate5480  (.A(g5425), .Z(II16321) ) ;
INV     gate5481  (.A(II16321), .Z(g9003) ) ;
INV     gate5482  (.A(g6052), .Z(II16325) ) ;
INV     gate5483  (.A(II16325), .Z(g9005) ) ;
INV     gate5484  (.A(g3900), .Z(II16328) ) ;
INV     gate5485  (.A(II16328), .Z(g9006) ) ;
INV     gate5486  (.A(g3462), .Z(II16332) ) ;
INV     gate5487  (.A(II16332), .Z(g9010) ) ;
INV     gate5488  (.A(g3618), .Z(II16335) ) ;
INV     gate5489  (.A(II16335), .Z(g9013) ) ;
INV     gate5490  (.A(g7015), .Z(II16338) ) ;
INV     gate5491  (.A(II16338), .Z(g9016) ) ;
INV     gate5492  (.A(g7265), .Z(II16341) ) ;
INV     gate5493  (.A(II16341), .Z(g9019) ) ;
INV     gate5494  (.A(g5556), .Z(II16344) ) ;
INV     gate5495  (.A(II16344), .Z(g9022) ) ;
INV     gate5496  (.A(g5427), .Z(II16347) ) ;
INV     gate5497  (.A(II16347), .Z(g9025) ) ;
INV     gate5498  (.A(g5679), .Z(g9027) ) ;
INV     gate5499  (.A(g3618), .Z(II16354) ) ;
INV     gate5500  (.A(II16354), .Z(g9035) ) ;
INV     gate5501  (.A(g3774), .Z(II16357) ) ;
INV     gate5502  (.A(II16357), .Z(g9038) ) ;
INV     gate5503  (.A(g7265), .Z(II16360) ) ;
INV     gate5504  (.A(II16360), .Z(g9041) ) ;
INV     gate5505  (.A(g3900), .Z(II16363) ) ;
INV     gate5506  (.A(II16363), .Z(g9044) ) ;
INV     gate5507  (.A(g5731), .Z(g9050) ) ;
INV     gate5508  (.A(g3774), .Z(II16372) ) ;
INV     gate5509  (.A(II16372), .Z(g9058) ) ;
INV     gate5510  (.A(g5789), .Z(g9067) ) ;
INV     gate5511  (.A(g5848), .Z(g9084) ) ;
INV     gate5512  (.A(g3366), .Z(II16432) ) ;
INV     gate5513  (.A(II16432), .Z(g9128) ) ;
INV     gate5514  (.A(g3522), .Z(II16438) ) ;
INV     gate5515  (.A(II16438), .Z(g9134) ) ;
INV     gate5516  (.A(g3678), .Z(II16444) ) ;
INV     gate5517  (.A(II16444), .Z(g9140) ) ;
INV     gate5518  (.A(g3834), .Z(II16450) ) ;
INV     gate5519  (.A(II16450), .Z(g9146) ) ;
INV     gate5520  (.A(g7936), .Z(II16453) ) ;
INV     gate5521  (.A(II16453), .Z(g9149) ) ;
INV     gate5522  (.A(g5893), .Z(g9150) ) ;
INV     gate5523  (.A(g7936), .Z(II16457) ) ;
INV     gate5524  (.A(II16457), .Z(g9159) ) ;
INV     gate5525  (.A(g6170), .Z(g9160) ) ;
INV     gate5526  (.A(g5852), .Z(g9161) ) ;
INV     gate5527  (.A(g5438), .Z(II16462) ) ;
INV     gate5528  (.A(II16462), .Z(g9170) ) ;
INV     gate5529  (.A(g6000), .Z(II16465) ) ;
INV     gate5530  (.A(II16465), .Z(g9173) ) ;
INV     gate5531  (.A(g5932), .Z(g9174) ) ;
INV     gate5532  (.A(g7936), .Z(II16469) ) ;
INV     gate5533  (.A(II16469), .Z(g9183) ) ;
INV     gate5534  (.A(g7901), .Z(II16472) ) ;
INV     gate5535  (.A(II16472), .Z(g9184) ) ;
INV     gate5536  (.A(g5803), .Z(g9187) ) ;
INV     gate5537  (.A(g6448), .Z(II16476) ) ;
INV     gate5538  (.A(II16476), .Z(g9196) ) ;
INV     gate5539  (.A(g5438), .Z(II16479) ) ;
INV     gate5540  (.A(II16479), .Z(g9199) ) ;
INV     gate5541  (.A(g6000), .Z(II16482) ) ;
INV     gate5542  (.A(II16482), .Z(g9202) ) ;
INV     gate5543  (.A(g5899), .Z(g9203) ) ;
INV     gate5544  (.A(g5473), .Z(II16486) ) ;
INV     gate5545  (.A(II16486), .Z(g9212) ) ;
INV     gate5546  (.A(g6000), .Z(II16489) ) ;
INV     gate5547  (.A(II16489), .Z(g9215) ) ;
INV     gate5548  (.A(g5966), .Z(g9216) ) ;
INV     gate5549  (.A(g7936), .Z(II16493) ) ;
INV     gate5550  (.A(II16493), .Z(g9225) ) ;
INV     gate5551  (.A(g5434), .Z(g9226) ) ;
INV     gate5552  (.A(g5587), .Z(g9227) ) ;
INV     gate5553  (.A(g7667), .Z(g9228) ) ;
INV     gate5554  (.A(g7901), .Z(II16499) ) ;
INV     gate5555  (.A(II16499), .Z(g9229) ) ;
INV     gate5556  (.A(g5752), .Z(g9232) ) ;
INV     gate5557  (.A(g3306), .Z(II16504) ) ;
INV     gate5558  (.A(II16504), .Z(g9242) ) ;
INV     gate5559  (.A(g6448), .Z(II16507) ) ;
INV     gate5560  (.A(II16507), .Z(g9245) ) ;
INV     gate5561  (.A(g5859), .Z(g9248) ) ;
INV     gate5562  (.A(g6713), .Z(II16511) ) ;
INV     gate5563  (.A(II16511), .Z(g9257) ) ;
INV     gate5564  (.A(g5473), .Z(II16514) ) ;
INV     gate5565  (.A(II16514), .Z(g9260) ) ;
INV     gate5566  (.A(g6000), .Z(II16517) ) ;
INV     gate5567  (.A(II16517), .Z(g9263) ) ;
INV     gate5568  (.A(g5938), .Z(g9264) ) ;
INV     gate5569  (.A(g5512), .Z(II16521) ) ;
INV     gate5570  (.A(II16521), .Z(g9273) ) ;
INV     gate5571  (.A(g6000), .Z(II16524) ) ;
INV     gate5572  (.A(II16524), .Z(g9276) ) ;
INV     gate5573  (.A(g5995), .Z(g9277) ) ;
INV     gate5574  (.A(g6197), .Z(g9286) ) ;
INV     gate5575  (.A(g6638), .Z(g9287) ) ;
INV     gate5576  (.A(g5363), .Z(g9288) ) ;
INV     gate5577  (.A(g5379), .Z(g9289) ) ;
INV     gate5578  (.A(g7901), .Z(II16532) ) ;
INV     gate5579  (.A(II16532), .Z(g9290) ) ;
INV     gate5580  (.A(g5703), .Z(g9293) ) ;
INV     gate5581  (.A(g3306), .Z(II16538) ) ;
INV     gate5582  (.A(II16538), .Z(g9303) ) ;
INV     gate5583  (.A(g5438), .Z(II16541) ) ;
INV     gate5584  (.A(II16541), .Z(g9306) ) ;
INV     gate5585  (.A(g6054), .Z(II16544) ) ;
INV     gate5586  (.A(II16544), .Z(g9309) ) ;
INV     gate5587  (.A(g5811), .Z(g9310) ) ;
INV     gate5588  (.A(g3462), .Z(II16549) ) ;
INV     gate5589  (.A(II16549), .Z(g9320) ) ;
INV     gate5590  (.A(g6713), .Z(II16552) ) ;
INV     gate5591  (.A(II16552), .Z(g9323) ) ;
INV     gate5592  (.A(g5906), .Z(g9326) ) ;
INV     gate5593  (.A(g7015), .Z(II16556) ) ;
INV     gate5594  (.A(II16556), .Z(g9335) ) ;
INV     gate5595  (.A(g5512), .Z(II16559) ) ;
INV     gate5596  (.A(II16559), .Z(g9338) ) ;
INV     gate5597  (.A(g6000), .Z(II16562) ) ;
INV     gate5598  (.A(II16562), .Z(g9341) ) ;
INV     gate5599  (.A(g5972), .Z(g9342) ) ;
INV     gate5600  (.A(g5556), .Z(II16566) ) ;
INV     gate5601  (.A(II16566), .Z(g9351) ) ;
INV     gate5602  (.A(g6000), .Z(II16569) ) ;
INV     gate5603  (.A(II16569), .Z(g9354) ) ;
INV     gate5604  (.A(g7639), .Z(g9355) ) ;
INV     gate5605  (.A(g5665), .Z(g9356) ) ;
INV     gate5606  (.A(g6448), .Z(II16578) ) ;
INV     gate5607  (.A(II16578), .Z(g9368) ) ;
INV     gate5608  (.A(g5438), .Z(II16581) ) ;
INV     gate5609  (.A(II16581), .Z(g9371) ) ;
INV     gate5610  (.A(g5761), .Z(g9374) ) ;
INV     gate5611  (.A(g3462), .Z(II16587) ) ;
INV     gate5612  (.A(II16587), .Z(g9384) ) ;
INV     gate5613  (.A(g5473), .Z(II16590) ) ;
INV     gate5614  (.A(II16590), .Z(g9387) ) ;
INV     gate5615  (.A(g6059), .Z(II16593) ) ;
INV     gate5616  (.A(II16593), .Z(g9390) ) ;
INV     gate5617  (.A(g5867), .Z(g9391) ) ;
INV     gate5618  (.A(g3618), .Z(II16598) ) ;
INV     gate5619  (.A(II16598), .Z(g9401) ) ;
INV     gate5620  (.A(g7015), .Z(II16601) ) ;
INV     gate5621  (.A(II16601), .Z(g9404) ) ;
INV     gate5622  (.A(g5945), .Z(g9407) ) ;
INV     gate5623  (.A(g7265), .Z(II16605) ) ;
INV     gate5624  (.A(II16605), .Z(g9416) ) ;
INV     gate5625  (.A(g5556), .Z(II16608) ) ;
INV     gate5626  (.A(II16608), .Z(g9419) ) ;
INV     gate5627  (.A(g6000), .Z(II16611) ) ;
INV     gate5628  (.A(II16611), .Z(g9422) ) ;
INV     gate5629  (.A(g5428), .Z(g9423) ) ;
INV     gate5630  (.A(g5469), .Z(g9424) ) ;
INV     gate5631  (.A(g5346), .Z(g9425) ) ;
INV     gate5632  (.A(g5543), .Z(g9426) ) ;
INV     gate5633  (.A(g5645), .Z(g9427) ) ;
INV     gate5634  (.A(g3306), .Z(II16624) ) ;
INV     gate5635  (.A(II16624), .Z(g9443) ) ;
INV     gate5636  (.A(g6448), .Z(II16627) ) ;
INV     gate5637  (.A(II16627), .Z(g9446) ) ;
INV     gate5638  (.A(g6057), .Z(II16630) ) ;
INV     gate5639  (.A(II16630), .Z(g9449) ) ;
INV     gate5640  (.A(g6486), .Z(II16633) ) ;
INV     gate5641  (.A(II16633), .Z(g9450) ) ;
INV     gate5642  (.A(g5717), .Z(g9453) ) ;
INV     gate5643  (.A(g6713), .Z(II16641) ) ;
INV     gate5644  (.A(II16641), .Z(g9465) ) ;
INV     gate5645  (.A(g5473), .Z(II16644) ) ;
INV     gate5646  (.A(II16644), .Z(g9468) ) ;
INV     gate5647  (.A(g5820), .Z(g9471) ) ;
INV     gate5648  (.A(g3618), .Z(II16650) ) ;
INV     gate5649  (.A(II16650), .Z(g9481) ) ;
INV     gate5650  (.A(g5512), .Z(II16653) ) ;
INV     gate5651  (.A(II16653), .Z(g9484) ) ;
INV     gate5652  (.A(g6066), .Z(II16656) ) ;
INV     gate5653  (.A(II16656), .Z(g9487) ) ;
INV     gate5654  (.A(g5914), .Z(g9488) ) ;
INV     gate5655  (.A(g3774), .Z(II16661) ) ;
INV     gate5656  (.A(II16661), .Z(g9498) ) ;
INV     gate5657  (.A(g7265), .Z(II16664) ) ;
INV     gate5658  (.A(II16664), .Z(g9501) ) ;
INV     gate5659  (.A(g6149), .Z(g9504) ) ;
INV     gate5660  (.A(g6227), .Z(g9505) ) ;
INV     gate5661  (.A(g6444), .Z(g9506) ) ;
INV     gate5662  (.A(g5953), .Z(g9507) ) ;
INV     gate5663  (.A(g3306), .Z(II16677) ) ;
INV     gate5664  (.A(II16677), .Z(g9524) ) ;
INV     gate5665  (.A(g5508), .Z(g9527) ) ;
INV     gate5666  (.A(g6643), .Z(II16681) ) ;
INV     gate5667  (.A(II16681), .Z(g9528) ) ;
INV     gate5668  (.A(g6486), .Z(II16684) ) ;
INV     gate5669  (.A(II16684), .Z(g9531) ) ;
INV     gate5670  (.A(g5683), .Z(g9569) ) ;
INV     gate5671  (.A(g3462), .Z(II16694) ) ;
INV     gate5672  (.A(II16694), .Z(g9585) ) ;
INV     gate5673  (.A(g6713), .Z(II16697) ) ;
INV     gate5674  (.A(II16697), .Z(g9588) ) ;
INV     gate5675  (.A(g6064), .Z(II16700) ) ;
INV     gate5676  (.A(II16700), .Z(g9591) ) ;
INV     gate5677  (.A(g6751), .Z(II16703) ) ;
INV     gate5678  (.A(II16703), .Z(g9592) ) ;
INV     gate5679  (.A(g5775), .Z(g9595) ) ;
INV     gate5680  (.A(g7015), .Z(II16711) ) ;
INV     gate5681  (.A(II16711), .Z(g9607) ) ;
INV     gate5682  (.A(g5512), .Z(II16714) ) ;
INV     gate5683  (.A(II16714), .Z(g9610) ) ;
INV     gate5684  (.A(g5876), .Z(g9613) ) ;
INV     gate5685  (.A(g3774), .Z(II16720) ) ;
INV     gate5686  (.A(II16720), .Z(g9623) ) ;
INV     gate5687  (.A(g5556), .Z(II16723) ) ;
INV     gate5688  (.A(II16723), .Z(g9626) ) ;
INV     gate5689  (.A(g6085), .Z(II16726) ) ;
INV     gate5690  (.A(II16726), .Z(g9629) ) ;
INV     gate5691  (.A(g6062), .Z(II16741) ) ;
INV     gate5692  (.A(II16741), .Z(g9640) ) ;
INV     gate5693  (.A(g3338), .Z(II16744) ) ;
INV     gate5694  (.A(II16744), .Z(g9641) ) ;
INV     gate5695  (.A(g6643), .Z(II16747) ) ;
INV     gate5696  (.A(II16747), .Z(g9644) ) ;
INV     gate5697  (.A(g5982), .Z(g9649) ) ;
INV     gate5698  (.A(g3462), .Z(II16759) ) ;
INV     gate5699  (.A(II16759), .Z(g9666) ) ;
INV     gate5700  (.A(g5552), .Z(g9669) ) ;
INV     gate5701  (.A(g6945), .Z(II16763) ) ;
INV     gate5702  (.A(II16763), .Z(g9670) ) ;
INV     gate5703  (.A(g6751), .Z(II16766) ) ;
INV     gate5704  (.A(II16766), .Z(g9673) ) ;
INV     gate5705  (.A(g5735), .Z(g9711) ) ;
INV     gate5706  (.A(g3618), .Z(II16776) ) ;
INV     gate5707  (.A(II16776), .Z(g9727) ) ;
INV     gate5708  (.A(g7015), .Z(II16779) ) ;
INV     gate5709  (.A(II16779), .Z(g9730) ) ;
INV     gate5710  (.A(g6083), .Z(II16782) ) ;
INV     gate5711  (.A(II16782), .Z(g9733) ) ;
INV     gate5712  (.A(g7053), .Z(II16785) ) ;
INV     gate5713  (.A(II16785), .Z(g9734) ) ;
INV     gate5714  (.A(g5834), .Z(g9737) ) ;
INV     gate5715  (.A(g7265), .Z(II16793) ) ;
INV     gate5716  (.A(II16793), .Z(g9749) ) ;
INV     gate5717  (.A(g5556), .Z(II16796) ) ;
INV     gate5718  (.A(II16796), .Z(g9752) ) ;
INV     gate5719  (.A(g5431), .Z(g9755) ) ;
INV     gate5720  (.A(g5504), .Z(g9756) ) ;
INV     gate5721  (.A(g5601), .Z(g9757) ) ;
INV     gate5722  (.A(g5618), .Z(g9758) ) ;
INV     gate5723  (.A(g3338), .Z(II16811) ) ;
INV     gate5724  (.A(II16811), .Z(g9767) ) ;
INV     gate5725  (.A(g6486), .Z(II16814) ) ;
INV     gate5726  (.A(II16814), .Z(g9770) ) ;
INV     gate5727  (.A(g6081), .Z(II16832) ) ;
INV     gate5728  (.A(II16832), .Z(g9786) ) ;
INV     gate5729  (.A(g3494), .Z(II16835) ) ;
INV     gate5730  (.A(II16835), .Z(g9787) ) ;
INV     gate5731  (.A(g6945), .Z(II16838) ) ;
INV     gate5732  (.A(II16838), .Z(g9790) ) ;
INV     gate5733  (.A(g6019), .Z(g9795) ) ;
INV     gate5734  (.A(g3618), .Z(II16850) ) ;
INV     gate5735  (.A(II16850), .Z(g9812) ) ;
INV     gate5736  (.A(g5598), .Z(g9815) ) ;
INV     gate5737  (.A(g7195), .Z(II16854) ) ;
INV     gate5738  (.A(II16854), .Z(g9816) ) ;
INV     gate5739  (.A(g7053), .Z(II16857) ) ;
INV     gate5740  (.A(II16857), .Z(g9819) ) ;
INV     gate5741  (.A(g5793), .Z(g9857) ) ;
INV     gate5742  (.A(g3774), .Z(II16867) ) ;
INV     gate5743  (.A(II16867), .Z(g9873) ) ;
INV     gate5744  (.A(g7265), .Z(II16870) ) ;
INV     gate5745  (.A(II16870), .Z(g9876) ) ;
INV     gate5746  (.A(g6102), .Z(II16873) ) ;
INV     gate5747  (.A(II16873), .Z(g9879) ) ;
INV     gate5748  (.A(g7303), .Z(II16876) ) ;
INV     gate5749  (.A(II16876), .Z(g9880) ) ;
INV     gate5750  (.A(g6310), .Z(g9884) ) ;
INV     gate5751  (.A(g6905), .Z(g9885) ) ;
INV     gate5752  (.A(g7149), .Z(g9886) ) ;
INV     gate5753  (.A(g6643), .Z(II16897) ) ;
INV     gate5754  (.A(II16897), .Z(g9895) ) ;
INV     gate5755  (.A(g6486), .Z(II16900) ) ;
INV     gate5756  (.A(II16900), .Z(g9898) ) ;
INV     gate5757  (.A(g3494), .Z(II16915) ) ;
INV     gate5758  (.A(II16915), .Z(g9913) ) ;
INV     gate5759  (.A(g6751), .Z(II16918) ) ;
INV     gate5760  (.A(II16918), .Z(g9916) ) ;
INV     gate5761  (.A(g6100), .Z(II16936) ) ;
INV     gate5762  (.A(II16936), .Z(g9932) ) ;
INV     gate5763  (.A(g3650), .Z(II16939) ) ;
INV     gate5764  (.A(II16939), .Z(g9933) ) ;
INV     gate5765  (.A(g7195), .Z(II16942) ) ;
INV     gate5766  (.A(II16942), .Z(g9936) ) ;
INV     gate5767  (.A(g6035), .Z(g9941) ) ;
INV     gate5768  (.A(g3774), .Z(II16954) ) ;
INV     gate5769  (.A(II16954), .Z(g9958) ) ;
INV     gate5770  (.A(g5615), .Z(g9961) ) ;
INV     gate5771  (.A(g7391), .Z(II16958) ) ;
INV     gate5772  (.A(II16958), .Z(g9962) ) ;
INV     gate5773  (.A(g7303), .Z(II16961) ) ;
INV     gate5774  (.A(II16961), .Z(g9965) ) ;
INV     gate5775  (.A(g3900), .Z(II16972) ) ;
INV     gate5776  (.A(II16972), .Z(g10004) ) ;
INV     gate5777  (.A(g5292), .Z(g10015) ) ;
INV     gate5778  (.A(g7936), .Z(II16984) ) ;
INV     gate5779  (.A(II16984), .Z(g10016) ) ;
INV     gate5780  (.A(g6079), .Z(II16987) ) ;
INV     gate5781  (.A(II16987), .Z(g10017) ) ;
INV     gate5782  (.A(g3338), .Z(II16990) ) ;
INV     gate5783  (.A(II16990), .Z(g10018) ) ;
INV     gate5784  (.A(g6643), .Z(II16993) ) ;
INV     gate5785  (.A(II16993), .Z(g10021) ) ;
INV     gate5786  (.A(g6945), .Z(II17009) ) ;
INV     gate5787  (.A(II17009), .Z(g10049) ) ;
INV     gate5788  (.A(g6751), .Z(II17012) ) ;
INV     gate5789  (.A(II17012), .Z(g10052) ) ;
INV     gate5790  (.A(g3650), .Z(II17027) ) ;
INV     gate5791  (.A(II17027), .Z(g10067) ) ;
INV     gate5792  (.A(g7053), .Z(II17030) ) ;
INV     gate5793  (.A(II17030), .Z(g10070) ) ;
INV     gate5794  (.A(g6117), .Z(II17048) ) ;
INV     gate5795  (.A(II17048), .Z(g10086) ) ;
INV     gate5796  (.A(g3806), .Z(II17051) ) ;
INV     gate5797  (.A(II17051), .Z(g10087) ) ;
INV     gate5798  (.A(g7391), .Z(II17054) ) ;
INV     gate5799  (.A(II17054), .Z(g10090) ) ;
INV     gate5800  (.A(g3900), .Z(II17066) ) ;
INV     gate5801  (.A(II17066), .Z(g10096) ) ;
INV     gate5802  (.A(g7700), .Z(g10099) ) ;
NOR3    gate5803  (.A(g3151), .B(g3142), .C(g3147), .Z(g7528) ) ;
INV     gate5804  (.A(g7528), .Z(II17070) ) ;
INV     gate5805  (.A(II17070), .Z(g10100) ) ;
INV     gate5806  (.A(g3338), .Z(II17081) ) ;
INV     gate5807  (.A(II17081), .Z(g10109) ) ;
INV     gate5808  (.A(g5326), .Z(g10124) ) ;
INV     gate5809  (.A(g7936), .Z(II17097) ) ;
INV     gate5810  (.A(II17097), .Z(g10125) ) ;
INV     gate5811  (.A(g6098), .Z(II17100) ) ;
INV     gate5812  (.A(II17100), .Z(g10126) ) ;
INV     gate5813  (.A(g3494), .Z(II17103) ) ;
INV     gate5814  (.A(II17103), .Z(g10127) ) ;
INV     gate5815  (.A(g6945), .Z(II17106) ) ;
INV     gate5816  (.A(II17106), .Z(g10130) ) ;
INV     gate5817  (.A(g7195), .Z(II17122) ) ;
INV     gate5818  (.A(II17122), .Z(g10158) ) ;
INV     gate5819  (.A(g7053), .Z(II17125) ) ;
INV     gate5820  (.A(II17125), .Z(g10161) ) ;
INV     gate5821  (.A(g3806), .Z(II17140) ) ;
INV     gate5822  (.A(II17140), .Z(g10176) ) ;
INV     gate5823  (.A(g7303), .Z(II17143) ) ;
INV     gate5824  (.A(II17143), .Z(g10179) ) ;
INV     gate5825  (.A(g3900), .Z(II17159) ) ;
INV     gate5826  (.A(II17159), .Z(g10189) ) ;
INV     gate5827  (.A(g3494), .Z(II17184) ) ;
INV     gate5828  (.A(II17184), .Z(g10214) ) ;
INV     gate5829  (.A(g5349), .Z(g10229) ) ;
INV     gate5830  (.A(g7936), .Z(II17200) ) ;
INV     gate5831  (.A(II17200), .Z(g10230) ) ;
INV     gate5832  (.A(g6115), .Z(II17203) ) ;
INV     gate5833  (.A(II17203), .Z(g10231) ) ;
INV     gate5834  (.A(g3650), .Z(II17206) ) ;
INV     gate5835  (.A(II17206), .Z(g10232) ) ;
INV     gate5836  (.A(g7195), .Z(II17209) ) ;
INV     gate5837  (.A(II17209), .Z(g10235) ) ;
INV     gate5838  (.A(g7391), .Z(II17225) ) ;
INV     gate5839  (.A(II17225), .Z(g10263) ) ;
INV     gate5840  (.A(g7303), .Z(II17228) ) ;
INV     gate5841  (.A(II17228), .Z(g10266) ) ;
INV     gate5842  (.A(g3900), .Z(II17235) ) ;
INV     gate5843  (.A(II17235), .Z(g10273) ) ;
INV     gate5844  (.A(g3900), .Z(II17238) ) ;
INV     gate5845  (.A(II17238), .Z(g10276) ) ;
INV     gate5846  (.A(g3650), .Z(II17278) ) ;
INV     gate5847  (.A(II17278), .Z(g10316) ) ;
INV     gate5848  (.A(g5366), .Z(g10331) ) ;
INV     gate5849  (.A(g7936), .Z(II17294) ) ;
INV     gate5850  (.A(II17294), .Z(g10332) ) ;
INV     gate5851  (.A(g6130), .Z(II17297) ) ;
INV     gate5852  (.A(II17297), .Z(g10333) ) ;
INV     gate5853  (.A(g3806), .Z(II17300) ) ;
INV     gate5854  (.A(II17300), .Z(g10334) ) ;
INV     gate5855  (.A(g7391), .Z(II17303) ) ;
INV     gate5856  (.A(II17303), .Z(g10337) ) ;
INV     gate5857  (.A(g3900), .Z(II17311) ) ;
INV     gate5858  (.A(II17311), .Z(g10357) ) ;
INV     gate5859  (.A(g3806), .Z(II17363) ) ;
INV     gate5860  (.A(II17363), .Z(g10409) ) ;
INV     gate5861  (.A(g3900), .Z(II17370) ) ;
INV     gate5862  (.A(II17370), .Z(g10416) ) ;
INV     gate5863  (.A(g3900), .Z(II17373) ) ;
INV     gate5864  (.A(II17373), .Z(g10419) ) ;
INV     gate5865  (.A(g7910), .Z(g10424) ) ;
INV     gate5866  (.A(g7826), .Z(g10481) ) ;
INV     gate5867  (.A(g3900), .Z(II17433) ) ;
INV     gate5868  (.A(II17433), .Z(g10482) ) ;
INV     gate5869  (.A(g7957), .Z(g10486) ) ;
INV     gate5870  (.A(g7962), .Z(g10500) ) ;
INV     gate5871  (.A(g3900), .Z(II17483) ) ;
INV     gate5872  (.A(II17483), .Z(g10542) ) ;
INV     gate5873  (.A(g3900), .Z(II17486) ) ;
INV     gate5874  (.A(II17486), .Z(g10545) ) ;
INV     gate5875  (.A(g7999), .Z(g10549) ) ;
INV     gate5876  (.A(g8008), .Z(g10560) ) ;
INV     gate5877  (.A(g8013), .Z(g10574) ) ;
INV     gate5878  (.A(g3900), .Z(II17527) ) ;
INV     gate5879  (.A(II17527), .Z(g10601) ) ;
INV     gate5880  (.A(g8074), .Z(g10606) ) ;
INV     gate5881  (.A(g8083), .Z(g10617) ) ;
INV     gate5882  (.A(g8088), .Z(g10631) ) ;
INV     gate5883  (.A(g3900), .Z(II17557) ) ;
INV     gate5884  (.A(II17557), .Z(g10646) ) ;
INV     gate5885  (.A(g8159), .Z(g10653) ) ;
INV     gate5886  (.A(g8168), .Z(g10664) ) ;
INV     gate5887  (.A(g8245), .Z(g10683) ) ;
INV     gate5888  (.A(g4326), .Z(g10694) ) ;
INV     gate5889  (.A(g4495), .Z(g10714) ) ;
INV     gate5890  (.A(g6173), .Z(g10730) ) ;
INV     gate5891  (.A(g4671), .Z(g10735) ) ;
INV     gate5892  (.A(g6205), .Z(g10749) ) ;
INV     gate5893  (.A(g4848), .Z(g10754) ) ;
INV     gate5894  (.A(g6048), .Z(g10765) ) ;
INV     gate5895  (.A(g6676), .Z(g10766) ) ;
INV     gate5896  (.A(g6294), .Z(g10767) ) ;
INV     gate5897  (.A(g6978), .Z(g10772) ) ;
INV     gate5898  (.A(g6431), .Z(g10773) ) ;
NOR2    gate5899  (.A(g2984), .B(g2985), .Z(g7575) ) ;
INV     gate5900  (.A(g7575), .Z(II17627) ) ;
INV     gate5901  (.A(II17627), .Z(g10779) ) ;
INV     gate5902  (.A(g7228), .Z(g10783) ) ;
INV     gate5903  (.A(g6183), .Z(II17632) ) ;
INV     gate5904  (.A(II17632), .Z(g10787) ) ;
INV     gate5905  (.A(g7424), .Z(g10788) ) ;
INV     gate5906  (.A(g6204), .Z(II17637) ) ;
INV     gate5907  (.A(II17637), .Z(g10792) ) ;
INV     gate5908  (.A(g6215), .Z(II17641) ) ;
INV     gate5909  (.A(II17641), .Z(g10796) ) ;
INV     gate5910  (.A(g6288), .Z(II17645) ) ;
INV     gate5911  (.A(II17645), .Z(g10800) ) ;
INV     gate5912  (.A(g6293), .Z(II17649) ) ;
INV     gate5913  (.A(II17649), .Z(g10804) ) ;
INV     gate5914  (.A(g6304), .Z(II17653) ) ;
INV     gate5915  (.A(II17653), .Z(g10808) ) ;
INV     gate5916  (.A(g5701), .Z(g10809) ) ;
INV     gate5917  (.A(g6367), .Z(II17658) ) ;
INV     gate5918  (.A(II17658), .Z(g10813) ) ;
INV     gate5919  (.A(g6425), .Z(II17662) ) ;
INV     gate5920  (.A(II17662), .Z(g10817) ) ;
INV     gate5921  (.A(g6430), .Z(II17666) ) ;
INV     gate5922  (.A(II17666), .Z(g10821) ) ;
INV     gate5923  (.A(g6441), .Z(II17670) ) ;
INV     gate5924  (.A(II17670), .Z(g10825) ) ;
INV     gate5925  (.A(g8107), .Z(II17673) ) ;
INV     gate5926  (.A(II17673), .Z(g10826) ) ;
INV     gate5927  (.A(g5749), .Z(g10829) ) ;
INV     gate5928  (.A(g6517), .Z(II17677) ) ;
INV     gate5929  (.A(II17677), .Z(g10830) ) ;
INV     gate5930  (.A(g6572), .Z(II17681) ) ;
INV     gate5931  (.A(II17681), .Z(g10834) ) ;
INV     gate5932  (.A(g6630), .Z(II17685) ) ;
INV     gate5933  (.A(II17685), .Z(g10838) ) ;
INV     gate5934  (.A(g6635), .Z(II17689) ) ;
INV     gate5935  (.A(II17689), .Z(g10842) ) ;
INV     gate5936  (.A(g8107), .Z(II17692) ) ;
INV     gate5937  (.A(II17692), .Z(g10843) ) ;
INV     gate5938  (.A(g5799), .Z(g10846) ) ;
INV     gate5939  (.A(g5800), .Z(g10847) ) ;
INV     gate5940  (.A(g5801), .Z(g10848) ) ;
INV     gate5941  (.A(g6711), .Z(II17698) ) ;
INV     gate5942  (.A(II17698), .Z(g10849) ) ;
INV     gate5943  (.A(g6781), .Z(II17701) ) ;
INV     gate5944  (.A(II17701), .Z(g10850) ) ;
INV     gate5945  (.A(g6836), .Z(II17705) ) ;
INV     gate5946  (.A(II17705), .Z(g10854) ) ;
INV     gate5947  (.A(g6894), .Z(II17709) ) ;
INV     gate5948  (.A(II17709), .Z(g10858) ) ;
INV     gate5949  (.A(g8031), .Z(II17712) ) ;
INV     gate5950  (.A(II17712), .Z(g10859) ) ;
INV     gate5951  (.A(g8107), .Z(II17715) ) ;
INV     gate5952  (.A(II17715), .Z(g10862) ) ;
INV     gate5953  (.A(g6131), .Z(g10865) ) ;
INV     gate5954  (.A(g5849), .Z(g10866) ) ;
INV     gate5955  (.A(g5850), .Z(g10867) ) ;
INV     gate5956  (.A(g6641), .Z(II17721) ) ;
INV     gate5957  (.A(II17721), .Z(g10868) ) ;
INV     gate5958  (.A(g6942), .Z(II17724) ) ;
INV     gate5959  (.A(II17724), .Z(g10869) ) ;
INV     gate5960  (.A(g7013), .Z(II17727) ) ;
INV     gate5961  (.A(II17727), .Z(g10870) ) ;
INV     gate5962  (.A(g7083), .Z(II17730) ) ;
INV     gate5963  (.A(II17730), .Z(g10871) ) ;
INV     gate5964  (.A(g7138), .Z(II17734) ) ;
INV     gate5965  (.A(II17734), .Z(g10875) ) ;
INV     gate5966  (.A(g6000), .Z(II17737) ) ;
INV     gate5967  (.A(II17737), .Z(g10876) ) ;
INV     gate5968  (.A(g8031), .Z(II17740) ) ;
INV     gate5969  (.A(II17740), .Z(g10877) ) ;
INV     gate5970  (.A(g8107), .Z(II17743) ) ;
INV     gate5971  (.A(II17743), .Z(g10880) ) ;
INV     gate5972  (.A(g8107), .Z(II17746) ) ;
INV     gate5973  (.A(II17746), .Z(g10883) ) ;
INV     gate5974  (.A(g5889), .Z(g10886) ) ;
INV     gate5975  (.A(g7157), .Z(II17750) ) ;
INV     gate5976  (.A(II17750), .Z(g10887) ) ;
INV     gate5977  (.A(g6943), .Z(II17753) ) ;
INV     gate5978  (.A(II17753), .Z(g10888) ) ;
INV     gate5979  (.A(g7192), .Z(II17756) ) ;
INV     gate5980  (.A(II17756), .Z(g10889) ) ;
INV     gate5981  (.A(g7263), .Z(II17759) ) ;
INV     gate5982  (.A(II17759), .Z(g10890) ) ;
INV     gate5983  (.A(g7333), .Z(II17762) ) ;
INV     gate5984  (.A(II17762), .Z(g10891) ) ;
INV     gate5985  (.A(g7976), .Z(II17765) ) ;
INV     gate5986  (.A(II17765), .Z(g10892) ) ;
INV     gate5987  (.A(g8031), .Z(II17768) ) ;
INV     gate5988  (.A(II17768), .Z(g10895) ) ;
INV     gate5989  (.A(g8107), .Z(II17771) ) ;
INV     gate5990  (.A(II17771), .Z(g10898) ) ;
INV     gate5991  (.A(g8107), .Z(II17774) ) ;
INV     gate5992  (.A(II17774), .Z(g10901) ) ;
INV     gate5993  (.A(g5922), .Z(g10904) ) ;
INV     gate5994  (.A(g5923), .Z(g10905) ) ;
INV     gate5995  (.A(g5924), .Z(g10906) ) ;
INV     gate5996  (.A(g7348), .Z(II17780) ) ;
INV     gate5997  (.A(II17780), .Z(g10907) ) ;
INV     gate5998  (.A(g7353), .Z(II17783) ) ;
INV     gate5999  (.A(II17783), .Z(g10908) ) ;
INV     gate6000  (.A(g7193), .Z(II17786) ) ;
INV     gate6001  (.A(II17786), .Z(g10909) ) ;
INV     gate6002  (.A(g7388), .Z(II17789) ) ;
INV     gate6003  (.A(II17789), .Z(g10910) ) ;
INV     gate6004  (.A(g7459), .Z(II17792) ) ;
INV     gate6005  (.A(II17792), .Z(g10911) ) ;
INV     gate6006  (.A(g7976), .Z(II17795) ) ;
INV     gate6007  (.A(II17795), .Z(g10912) ) ;
INV     gate6008  (.A(g8031), .Z(II17798) ) ;
INV     gate6009  (.A(II17798), .Z(g10915) ) ;
INV     gate6010  (.A(g8107), .Z(II17801) ) ;
INV     gate6011  (.A(II17801), .Z(g10918) ) ;
INV     gate6012  (.A(g8031), .Z(II17804) ) ;
INV     gate6013  (.A(II17804), .Z(g10921) ) ;
INV     gate6014  (.A(g8107), .Z(II17807) ) ;
INV     gate6015  (.A(II17807), .Z(g10924) ) ;
INV     gate6016  (.A(g6153), .Z(g10927) ) ;
INV     gate6017  (.A(g5951), .Z(g10928) ) ;
INV     gate6018  (.A(g5952), .Z(g10929) ) ;
INV     gate6019  (.A(g5707), .Z(II17813) ) ;
INV     gate6020  (.A(II17813), .Z(g10930) ) ;
INV     gate6021  (.A(g7346), .Z(II17816) ) ;
INV     gate6022  (.A(II17816), .Z(g10931) ) ;
INV     gate6023  (.A(g6448), .Z(II17819) ) ;
INV     gate6024  (.A(II17819), .Z(g10932) ) ;
INV     gate6025  (.A(g7478), .Z(II17822) ) ;
INV     gate6026  (.A(II17822), .Z(g10933) ) ;
INV     gate6027  (.A(g7483), .Z(II17825) ) ;
INV     gate6028  (.A(II17825), .Z(g10934) ) ;
INV     gate6029  (.A(g7389), .Z(II17828) ) ;
INV     gate6030  (.A(II17828), .Z(g10935) ) ;
INV     gate6031  (.A(g7518), .Z(II17831) ) ;
INV     gate6032  (.A(II17831), .Z(g10936) ) ;
INV     gate6033  (.A(g7976), .Z(II17834) ) ;
INV     gate6034  (.A(II17834), .Z(g10937) ) ;
INV     gate6035  (.A(g8031), .Z(II17837) ) ;
INV     gate6036  (.A(II17837), .Z(g10940) ) ;
INV     gate6037  (.A(g8107), .Z(II17840) ) ;
INV     gate6038  (.A(II17840), .Z(g10943) ) ;
INV     gate6039  (.A(g8031), .Z(II17843) ) ;
INV     gate6040  (.A(II17843), .Z(g10946) ) ;
INV     gate6041  (.A(g8107), .Z(II17846) ) ;
INV     gate6042  (.A(II17846), .Z(g10949) ) ;
INV     gate6043  (.A(g8103), .Z(II17849) ) ;
INV     gate6044  (.A(II17849), .Z(g10952) ) ;
INV     gate6045  (.A(g5978), .Z(g10961) ) ;
INV     gate6046  (.A(g5979), .Z(g10962) ) ;
INV     gate6047  (.A(g6232), .Z(II17854) ) ;
INV     gate6048  (.A(II17854), .Z(g10963) ) ;
INV     gate6049  (.A(g6448), .Z(II17857) ) ;
INV     gate6050  (.A(II17857), .Z(g10966) ) ;
INV     gate6051  (.A(g5765), .Z(II17860) ) ;
INV     gate6052  (.A(II17860), .Z(g10967) ) ;
INV     gate6053  (.A(g7476), .Z(II17863) ) ;
INV     gate6054  (.A(II17863), .Z(g10968) ) ;
INV     gate6055  (.A(g6713), .Z(II17866) ) ;
INV     gate6056  (.A(II17866), .Z(g10969) ) ;
INV     gate6057  (.A(g7534), .Z(II17869) ) ;
INV     gate6058  (.A(II17869), .Z(g10972) ) ;
INV     gate6059  (.A(g7539), .Z(II17872) ) ;
INV     gate6060  (.A(II17872), .Z(g10973) ) ;
INV     gate6061  (.A(g7976), .Z(II17875) ) ;
INV     gate6062  (.A(II17875), .Z(g10974) ) ;
INV     gate6063  (.A(g8031), .Z(II17878) ) ;
INV     gate6064  (.A(II17878), .Z(g10977) ) ;
INV     gate6065  (.A(g7976), .Z(II17881) ) ;
INV     gate6066  (.A(II17881), .Z(g10980) ) ;
INV     gate6067  (.A(g8031), .Z(II17884) ) ;
INV     gate6068  (.A(II17884), .Z(g10983) ) ;
INV     gate6069  (.A(g6014), .Z(g10986) ) ;
INV     gate6070  (.A(g6015), .Z(g10987) ) ;
INV     gate6071  (.A(g6314), .Z(II17889) ) ;
INV     gate6072  (.A(II17889), .Z(g10988) ) ;
INV     gate6073  (.A(g6232), .Z(II17892) ) ;
INV     gate6074  (.A(II17892), .Z(g10991) ) ;
INV     gate6075  (.A(g6448), .Z(II17895) ) ;
INV     gate6076  (.A(II17895), .Z(g10994) ) ;
INV     gate6077  (.A(g6643), .Z(II17898) ) ;
INV     gate6078  (.A(II17898), .Z(g10995) ) ;
INV     gate6079  (.A(g6369), .Z(II17901) ) ;
INV     gate6080  (.A(II17901), .Z(g10996) ) ;
INV     gate6081  (.A(g6713), .Z(II17904) ) ;
INV     gate6082  (.A(II17904), .Z(g10999) ) ;
INV     gate6083  (.A(g5824), .Z(II17907) ) ;
INV     gate6084  (.A(II17907), .Z(g11002) ) ;
INV     gate6085  (.A(g7532), .Z(II17910) ) ;
INV     gate6086  (.A(II17910), .Z(g11003) ) ;
INV     gate6087  (.A(g7015), .Z(II17913) ) ;
INV     gate6088  (.A(II17913), .Z(g11004) ) ;
INV     gate6089  (.A(g7560), .Z(II17916) ) ;
INV     gate6090  (.A(II17916), .Z(g11007) ) ;
INV     gate6091  (.A(g7976), .Z(II17919) ) ;
INV     gate6092  (.A(II17919), .Z(g11008) ) ;
INV     gate6093  (.A(g8031), .Z(II17922) ) ;
INV     gate6094  (.A(II17922), .Z(g11011) ) ;
INV     gate6095  (.A(g7976), .Z(II17925) ) ;
INV     gate6096  (.A(II17925), .Z(g11014) ) ;
INV     gate6097  (.A(g8031), .Z(II17928) ) ;
INV     gate6098  (.A(II17928), .Z(g11017) ) ;
INV     gate6099  (.A(g6029), .Z(g11020) ) ;
INV     gate6100  (.A(g6030), .Z(g11021) ) ;
INV     gate6101  (.A(g3254), .Z(II17933) ) ;
INV     gate6102  (.A(II17933), .Z(g11022) ) ;
INV     gate6103  (.A(g6314), .Z(II17936) ) ;
INV     gate6104  (.A(II17936), .Z(g11025) ) ;
INV     gate6105  (.A(g6232), .Z(II17939) ) ;
INV     gate6106  (.A(II17939), .Z(g11028) ) ;
INV     gate6107  (.A(g5548), .Z(II17942) ) ;
INV     gate6108  (.A(II17942), .Z(g11031) ) ;
INV     gate6109  (.A(g5668), .Z(II17945) ) ;
INV     gate6110  (.A(II17945), .Z(g11032) ) ;
INV     gate6111  (.A(g6643), .Z(II17948) ) ;
INV     gate6112  (.A(II17948), .Z(g11035) ) ;
INV     gate6113  (.A(g6519), .Z(II17951) ) ;
INV     gate6114  (.A(II17951), .Z(g11036) ) ;
INV     gate6115  (.A(g6369), .Z(II17954) ) ;
INV     gate6116  (.A(II17954), .Z(g11039) ) ;
INV     gate6117  (.A(g6713), .Z(II17957) ) ;
INV     gate6118  (.A(II17957), .Z(g11042) ) ;
INV     gate6119  (.A(g6945), .Z(II17960) ) ;
INV     gate6120  (.A(II17960), .Z(g11045) ) ;
INV     gate6121  (.A(g6574), .Z(II17963) ) ;
INV     gate6122  (.A(II17963), .Z(g11048) ) ;
INV     gate6123  (.A(g7015), .Z(II17966) ) ;
INV     gate6124  (.A(II17966), .Z(g11051) ) ;
INV     gate6125  (.A(g5880), .Z(II17969) ) ;
INV     gate6126  (.A(II17969), .Z(g11054) ) ;
INV     gate6127  (.A(g7558), .Z(II17972) ) ;
INV     gate6128  (.A(II17972), .Z(g11055) ) ;
INV     gate6129  (.A(g7265), .Z(II17975) ) ;
INV     gate6130  (.A(II17975), .Z(g11056) ) ;
NOR2    gate6131  (.A(g2992), .B(g2991), .Z(g7795) ) ;
INV     gate6132  (.A(g7795), .Z(II17978) ) ;
INV     gate6133  (.A(II17978), .Z(g11059) ) ;
INV     gate6134  (.A(g7976), .Z(II17981) ) ;
INV     gate6135  (.A(II17981), .Z(g11063) ) ;
INV     gate6136  (.A(g7976), .Z(II17984) ) ;
INV     gate6137  (.A(II17984), .Z(g11066) ) ;
INV     gate6138  (.A(g8257), .Z(g11069) ) ;
INV     gate6139  (.A(g6041), .Z(g11078) ) ;
INV     gate6140  (.A(g3254), .Z(II17989) ) ;
INV     gate6141  (.A(II17989), .Z(g11079) ) ;
INV     gate6142  (.A(g6314), .Z(II17992) ) ;
INV     gate6143  (.A(II17992), .Z(g11082) ) ;
INV     gate6144  (.A(g6232), .Z(II17995) ) ;
INV     gate6145  (.A(II17995), .Z(g11085) ) ;
INV     gate6146  (.A(g5668), .Z(II17998) ) ;
INV     gate6147  (.A(II17998), .Z(g11088) ) ;
INV     gate6148  (.A(g6643), .Z(II18001) ) ;
INV     gate6149  (.A(II18001), .Z(g11091) ) ;
INV     gate6150  (.A(g3410), .Z(II18004) ) ;
INV     gate6151  (.A(II18004), .Z(g11092) ) ;
INV     gate6152  (.A(g6519), .Z(II18007) ) ;
INV     gate6153  (.A(II18007), .Z(g11095) ) ;
INV     gate6154  (.A(g6369), .Z(II18010) ) ;
INV     gate6155  (.A(II18010), .Z(g11098) ) ;
INV     gate6156  (.A(g5594), .Z(II18013) ) ;
INV     gate6157  (.A(II18013), .Z(g11101) ) ;
INV     gate6158  (.A(g5720), .Z(II18016) ) ;
INV     gate6159  (.A(II18016), .Z(g11102) ) ;
INV     gate6160  (.A(g6945), .Z(II18019) ) ;
INV     gate6161  (.A(II18019), .Z(g11105) ) ;
INV     gate6162  (.A(g6783), .Z(II18022) ) ;
INV     gate6163  (.A(II18022), .Z(g11108) ) ;
INV     gate6164  (.A(g6574), .Z(II18025) ) ;
INV     gate6165  (.A(II18025), .Z(g11111) ) ;
INV     gate6166  (.A(g7015), .Z(II18028) ) ;
INV     gate6167  (.A(II18028), .Z(g11114) ) ;
INV     gate6168  (.A(g7195), .Z(II18031) ) ;
INV     gate6169  (.A(II18031), .Z(g11117) ) ;
INV     gate6170  (.A(g6838), .Z(II18034) ) ;
INV     gate6171  (.A(II18034), .Z(g11120) ) ;
INV     gate6172  (.A(g7265), .Z(II18037) ) ;
INV     gate6173  (.A(II18037), .Z(g11123) ) ;
INV     gate6174  (.A(g7976), .Z(II18040) ) ;
INV     gate6175  (.A(II18040), .Z(g11126) ) ;
INV     gate6176  (.A(g7976), .Z(II18043) ) ;
INV     gate6177  (.A(II18043), .Z(g11129) ) ;
INV     gate6178  (.A(g3254), .Z(II18046) ) ;
INV     gate6179  (.A(II18046), .Z(g11132) ) ;
INV     gate6180  (.A(g6314), .Z(II18049) ) ;
INV     gate6181  (.A(II18049), .Z(g11135) ) ;
INV     gate6182  (.A(g6232), .Z(II18052) ) ;
INV     gate6183  (.A(II18052), .Z(g11138) ) ;
INV     gate6184  (.A(g5668), .Z(II18055) ) ;
INV     gate6185  (.A(II18055), .Z(g11141) ) ;
INV     gate6186  (.A(g6643), .Z(II18058) ) ;
INV     gate6187  (.A(II18058), .Z(g11144) ) ;
INV     gate6188  (.A(g3410), .Z(II18061) ) ;
INV     gate6189  (.A(II18061), .Z(g11145) ) ;
INV     gate6190  (.A(g6519), .Z(II18064) ) ;
INV     gate6191  (.A(II18064), .Z(g11148) ) ;
INV     gate6192  (.A(g6369), .Z(II18067) ) ;
INV     gate6193  (.A(II18067), .Z(g11151) ) ;
INV     gate6194  (.A(g5720), .Z(II18070) ) ;
INV     gate6195  (.A(II18070), .Z(g11154) ) ;
INV     gate6196  (.A(g6945), .Z(II18073) ) ;
INV     gate6197  (.A(II18073), .Z(g11157) ) ;
INV     gate6198  (.A(g3566), .Z(II18076) ) ;
INV     gate6199  (.A(II18076), .Z(g11160) ) ;
INV     gate6200  (.A(g6783), .Z(II18079) ) ;
INV     gate6201  (.A(II18079), .Z(g11163) ) ;
INV     gate6202  (.A(g6574), .Z(II18082) ) ;
INV     gate6203  (.A(II18082), .Z(g11166) ) ;
INV     gate6204  (.A(g5611), .Z(II18085) ) ;
INV     gate6205  (.A(II18085), .Z(g11169) ) ;
INV     gate6206  (.A(g5778), .Z(II18088) ) ;
INV     gate6207  (.A(II18088), .Z(g11170) ) ;
INV     gate6208  (.A(g7195), .Z(II18091) ) ;
INV     gate6209  (.A(II18091), .Z(g11173) ) ;
INV     gate6210  (.A(g7085), .Z(II18094) ) ;
INV     gate6211  (.A(II18094), .Z(g11176) ) ;
INV     gate6212  (.A(g6838), .Z(II18097) ) ;
INV     gate6213  (.A(II18097), .Z(g11179) ) ;
INV     gate6214  (.A(g7265), .Z(II18100) ) ;
INV     gate6215  (.A(II18100), .Z(g11182) ) ;
INV     gate6216  (.A(g7391), .Z(II18103) ) ;
INV     gate6217  (.A(II18103), .Z(g11185) ) ;
INV     gate6218  (.A(g3999), .Z(g11190) ) ;
INV     gate6219  (.A(g3254), .Z(II18121) ) ;
INV     gate6220  (.A(II18121), .Z(g11199) ) ;
INV     gate6221  (.A(g6314), .Z(II18124) ) ;
INV     gate6222  (.A(II18124), .Z(g11202) ) ;
INV     gate6223  (.A(g6232), .Z(II18127) ) ;
INV     gate6224  (.A(II18127), .Z(g11205) ) ;
INV     gate6225  (.A(g5547), .Z(II18130) ) ;
INV     gate6226  (.A(II18130), .Z(g11208) ) ;
INV     gate6227  (.A(g6448), .Z(II18133) ) ;
INV     gate6228  (.A(II18133), .Z(g11209) ) ;
INV     gate6229  (.A(g5668), .Z(II18136) ) ;
INV     gate6230  (.A(II18136), .Z(g11210) ) ;
INV     gate6231  (.A(g6643), .Z(II18139) ) ;
INV     gate6232  (.A(II18139), .Z(g11213) ) ;
INV     gate6233  (.A(g3410), .Z(II18142) ) ;
INV     gate6234  (.A(II18142), .Z(g11216) ) ;
INV     gate6235  (.A(g6519), .Z(II18145) ) ;
INV     gate6236  (.A(II18145), .Z(g11219) ) ;
INV     gate6237  (.A(g6369), .Z(II18148) ) ;
INV     gate6238  (.A(II18148), .Z(g11222) ) ;
INV     gate6239  (.A(g5720), .Z(II18151) ) ;
INV     gate6240  (.A(II18151), .Z(g11225) ) ;
INV     gate6241  (.A(g6945), .Z(II18154) ) ;
INV     gate6242  (.A(II18154), .Z(g11228) ) ;
INV     gate6243  (.A(g3566), .Z(II18157) ) ;
INV     gate6244  (.A(II18157), .Z(g11231) ) ;
INV     gate6245  (.A(g6783), .Z(II18160) ) ;
INV     gate6246  (.A(II18160), .Z(g11234) ) ;
INV     gate6247  (.A(g6574), .Z(II18163) ) ;
INV     gate6248  (.A(II18163), .Z(g11237) ) ;
INV     gate6249  (.A(g5778), .Z(II18166) ) ;
INV     gate6250  (.A(II18166), .Z(g11240) ) ;
INV     gate6251  (.A(g7195), .Z(II18169) ) ;
INV     gate6252  (.A(II18169), .Z(g11243) ) ;
INV     gate6253  (.A(g3722), .Z(II18172) ) ;
INV     gate6254  (.A(II18172), .Z(g11246) ) ;
INV     gate6255  (.A(g7085), .Z(II18175) ) ;
INV     gate6256  (.A(II18175), .Z(g11249) ) ;
INV     gate6257  (.A(g6838), .Z(II18178) ) ;
INV     gate6258  (.A(II18178), .Z(g11252) ) ;
INV     gate6259  (.A(g5636), .Z(II18181) ) ;
INV     gate6260  (.A(II18181), .Z(g11255) ) ;
INV     gate6261  (.A(g5837), .Z(II18184) ) ;
INV     gate6262  (.A(II18184), .Z(g11256) ) ;
INV     gate6263  (.A(g7391), .Z(II18187) ) ;
INV     gate6264  (.A(II18187), .Z(g11259) ) ;
INV     gate6265  (.A(g6232), .Z(II18211) ) ;
INV     gate6266  (.A(II18211), .Z(g11265) ) ;
INV     gate6267  (.A(g3254), .Z(II18214) ) ;
INV     gate6268  (.A(II18214), .Z(g11268) ) ;
INV     gate6269  (.A(g6314), .Z(II18217) ) ;
INV     gate6270  (.A(II18217), .Z(g11271) ) ;
INV     gate6271  (.A(g6232), .Z(II18220) ) ;
INV     gate6272  (.A(II18220), .Z(g11274) ) ;
INV     gate6273  (.A(g6448), .Z(II18223) ) ;
INV     gate6274  (.A(II18223), .Z(g11277) ) ;
INV     gate6275  (.A(g5668), .Z(II18226) ) ;
INV     gate6276  (.A(II18226), .Z(g11278) ) ;
INV     gate6277  (.A(g3410), .Z(II18229) ) ;
INV     gate6278  (.A(II18229), .Z(g11281) ) ;
INV     gate6279  (.A(g6519), .Z(II18232) ) ;
INV     gate6280  (.A(II18232), .Z(g11284) ) ;
INV     gate6281  (.A(g6369), .Z(II18235) ) ;
INV     gate6282  (.A(II18235), .Z(g11287) ) ;
INV     gate6283  (.A(g5593), .Z(II18238) ) ;
INV     gate6284  (.A(II18238), .Z(g11290) ) ;
INV     gate6285  (.A(g6713), .Z(II18241) ) ;
INV     gate6286  (.A(II18241), .Z(g11291) ) ;
INV     gate6287  (.A(g5720), .Z(II18244) ) ;
INV     gate6288  (.A(II18244), .Z(g11294) ) ;
INV     gate6289  (.A(g6945), .Z(II18247) ) ;
INV     gate6290  (.A(II18247), .Z(g11297) ) ;
INV     gate6291  (.A(g3566), .Z(II18250) ) ;
INV     gate6292  (.A(II18250), .Z(g11300) ) ;
INV     gate6293  (.A(g6783), .Z(II18253) ) ;
INV     gate6294  (.A(II18253), .Z(g11303) ) ;
INV     gate6295  (.A(g6574), .Z(II18256) ) ;
INV     gate6296  (.A(II18256), .Z(g11306) ) ;
INV     gate6297  (.A(g5778), .Z(II18259) ) ;
INV     gate6298  (.A(II18259), .Z(g11309) ) ;
INV     gate6299  (.A(g7195), .Z(II18262) ) ;
INV     gate6300  (.A(II18262), .Z(g11312) ) ;
INV     gate6301  (.A(g3722), .Z(II18265) ) ;
INV     gate6302  (.A(II18265), .Z(g11315) ) ;
INV     gate6303  (.A(g7085), .Z(II18268) ) ;
INV     gate6304  (.A(II18268), .Z(g11318) ) ;
INV     gate6305  (.A(g6838), .Z(II18271) ) ;
INV     gate6306  (.A(II18271), .Z(g11321) ) ;
INV     gate6307  (.A(g5837), .Z(II18274) ) ;
INV     gate6308  (.A(II18274), .Z(g11324) ) ;
INV     gate6309  (.A(g7391), .Z(II18277) ) ;
INV     gate6310  (.A(II18277), .Z(g11327) ) ;
INV     gate6311  (.A(g4094), .Z(g11332) ) ;
INV     gate6312  (.A(g6314), .Z(II18295) ) ;
INV     gate6313  (.A(II18295), .Z(g11341) ) ;
INV     gate6314  (.A(g6232), .Z(II18298) ) ;
INV     gate6315  (.A(II18298), .Z(g11344) ) ;
INV     gate6316  (.A(g3254), .Z(II18302) ) ;
INV     gate6317  (.A(II18302), .Z(g11348) ) ;
INV     gate6318  (.A(g6314), .Z(II18305) ) ;
INV     gate6319  (.A(II18305), .Z(g11351) ) ;
INV     gate6320  (.A(g6448), .Z(II18308) ) ;
INV     gate6321  (.A(II18308), .Z(g11354) ) ;
INV     gate6322  (.A(g5668), .Z(II18311) ) ;
INV     gate6323  (.A(II18311), .Z(g11355) ) ;
INV     gate6324  (.A(g6369), .Z(II18314) ) ;
INV     gate6325  (.A(II18314), .Z(g11358) ) ;
INV     gate6326  (.A(g3410), .Z(II18317) ) ;
INV     gate6327  (.A(II18317), .Z(g11361) ) ;
INV     gate6328  (.A(g6519), .Z(II18320) ) ;
INV     gate6329  (.A(II18320), .Z(g11364) ) ;
INV     gate6330  (.A(g6369), .Z(II18323) ) ;
INV     gate6331  (.A(II18323), .Z(g11367) ) ;
INV     gate6332  (.A(g6713), .Z(II18326) ) ;
INV     gate6333  (.A(II18326), .Z(g11370) ) ;
INV     gate6334  (.A(g5720), .Z(II18329) ) ;
INV     gate6335  (.A(II18329), .Z(g11373) ) ;
INV     gate6336  (.A(g3566), .Z(II18332) ) ;
INV     gate6337  (.A(II18332), .Z(g11376) ) ;
INV     gate6338  (.A(g6783), .Z(II18335) ) ;
INV     gate6339  (.A(II18335), .Z(g11379) ) ;
INV     gate6340  (.A(g6574), .Z(II18338) ) ;
INV     gate6341  (.A(II18338), .Z(g11382) ) ;
INV     gate6342  (.A(g5610), .Z(II18341) ) ;
INV     gate6343  (.A(II18341), .Z(g11385) ) ;
INV     gate6344  (.A(g7015), .Z(II18344) ) ;
INV     gate6345  (.A(II18344), .Z(g11386) ) ;
INV     gate6346  (.A(g5778), .Z(II18347) ) ;
INV     gate6347  (.A(II18347), .Z(g11389) ) ;
INV     gate6348  (.A(g7195), .Z(II18350) ) ;
INV     gate6349  (.A(II18350), .Z(g11392) ) ;
INV     gate6350  (.A(g3722), .Z(II18353) ) ;
INV     gate6351  (.A(II18353), .Z(g11395) ) ;
INV     gate6352  (.A(g7085), .Z(II18356) ) ;
INV     gate6353  (.A(II18356), .Z(g11398) ) ;
INV     gate6354  (.A(g6838), .Z(II18359) ) ;
INV     gate6355  (.A(II18359), .Z(g11401) ) ;
INV     gate6356  (.A(g5837), .Z(II18362) ) ;
INV     gate6357  (.A(II18362), .Z(g11404) ) ;
INV     gate6358  (.A(g7391), .Z(II18365) ) ;
INV     gate6359  (.A(II18365), .Z(g11407) ) ;
INV     gate6360  (.A(g3254), .Z(II18375) ) ;
INV     gate6361  (.A(II18375), .Z(g11411) ) ;
INV     gate6362  (.A(g6314), .Z(II18378) ) ;
INV     gate6363  (.A(II18378), .Z(g11414) ) ;
INV     gate6364  (.A(g6232), .Z(II18381) ) ;
INV     gate6365  (.A(II18381), .Z(g11417) ) ;
INV     gate6366  (.A(g3254), .Z(II18386) ) ;
INV     gate6367  (.A(II18386), .Z(g11422) ) ;
INV     gate6368  (.A(g6519), .Z(II18389) ) ;
INV     gate6369  (.A(II18389), .Z(g11425) ) ;
INV     gate6370  (.A(g6369), .Z(II18392) ) ;
INV     gate6371  (.A(II18392), .Z(g11428) ) ;
INV     gate6372  (.A(g3410), .Z(II18396) ) ;
INV     gate6373  (.A(II18396), .Z(g11432) ) ;
INV     gate6374  (.A(g6519), .Z(II18399) ) ;
INV     gate6375  (.A(II18399), .Z(g11435) ) ;
INV     gate6376  (.A(g6713), .Z(II18402) ) ;
INV     gate6377  (.A(II18402), .Z(g11438) ) ;
INV     gate6378  (.A(g5720), .Z(II18405) ) ;
INV     gate6379  (.A(II18405), .Z(g11441) ) ;
INV     gate6380  (.A(g6574), .Z(II18408) ) ;
INV     gate6381  (.A(II18408), .Z(g11444) ) ;
INV     gate6382  (.A(g3566), .Z(II18411) ) ;
INV     gate6383  (.A(II18411), .Z(g11447) ) ;
INV     gate6384  (.A(g6783), .Z(II18414) ) ;
INV     gate6385  (.A(II18414), .Z(g11450) ) ;
INV     gate6386  (.A(g6574), .Z(II18417) ) ;
INV     gate6387  (.A(II18417), .Z(g11453) ) ;
INV     gate6388  (.A(g7015), .Z(II18420) ) ;
INV     gate6389  (.A(II18420), .Z(g11456) ) ;
INV     gate6390  (.A(g5778), .Z(II18423) ) ;
INV     gate6391  (.A(II18423), .Z(g11459) ) ;
INV     gate6392  (.A(g3722), .Z(II18426) ) ;
INV     gate6393  (.A(II18426), .Z(g11462) ) ;
INV     gate6394  (.A(g7085), .Z(II18429) ) ;
INV     gate6395  (.A(II18429), .Z(g11465) ) ;
INV     gate6396  (.A(g6838), .Z(II18432) ) ;
INV     gate6397  (.A(II18432), .Z(g11468) ) ;
INV     gate6398  (.A(g5635), .Z(II18435) ) ;
INV     gate6399  (.A(II18435), .Z(g11471) ) ;
INV     gate6400  (.A(g7265), .Z(II18438) ) ;
INV     gate6401  (.A(II18438), .Z(g11472) ) ;
INV     gate6402  (.A(g5837), .Z(II18441) ) ;
INV     gate6403  (.A(II18441), .Z(g11475) ) ;
INV     gate6404  (.A(g7391), .Z(II18444) ) ;
INV     gate6405  (.A(II18444), .Z(g11478) ) ;
INV     gate6406  (.A(g4204), .Z(g11481) ) ;
INV     gate6407  (.A(g8276), .Z(g11490) ) ;
INV     gate6408  (.A(g10868), .Z(II18449) ) ;
INV     gate6409  (.A(g10930), .Z(II18452) ) ;
INV     gate6410  (.A(g11031), .Z(II18455) ) ;
INV     gate6411  (.A(g11208), .Z(II18458) ) ;
INV     gate6412  (.A(g10931), .Z(II18461) ) ;
INV     gate6413  (.A(g8620), .Z(II18464) ) ;
INV     gate6414  (.A(g8769), .Z(II18467) ) ;
INV     gate6415  (.A(g8808), .Z(II18470) ) ;
INV     gate6416  (.A(g8839), .Z(II18473) ) ;
INV     gate6417  (.A(g8791), .Z(II18476) ) ;
INV     gate6418  (.A(g8820), .Z(II18479) ) ;
INV     gate6419  (.A(g8859), .Z(II18482) ) ;
INV     gate6420  (.A(g8809), .Z(II18485) ) ;
INV     gate6421  (.A(g8840), .Z(II18488) ) ;
INV     gate6422  (.A(g8891), .Z(II18491) ) ;
INV     gate6423  (.A(g8821), .Z(II18494) ) ;
INV     gate6424  (.A(g8860), .Z(II18497) ) ;
INV     gate6425  (.A(g8924), .Z(II18500) ) ;
INV     gate6426  (.A(g8658), .Z(II18503) ) ;
INV     gate6427  (.A(g8699), .Z(II18506) ) ;
INV     gate6428  (.A(g8770), .Z(II18509) ) ;
INV     gate6429  (.A(g9309), .Z(II18512) ) ;
INV     gate6430  (.A(g8843), .Z(II18515) ) ;
INV     gate6431  (.A(g8893), .Z(II18518) ) ;
INV     gate6432  (.A(g9449), .Z(II18521) ) ;
INV     gate6433  (.A(g9640), .Z(II18524) ) ;
INV     gate6434  (.A(g10017), .Z(II18527) ) ;
INV     gate6435  (.A(g10888), .Z(II18530) ) ;
INV     gate6436  (.A(g10967), .Z(II18533) ) ;
INV     gate6437  (.A(g11101), .Z(II18536) ) ;
INV     gate6438  (.A(g11290), .Z(II18539) ) ;
INV     gate6439  (.A(g10968), .Z(II18542) ) ;
INV     gate6440  (.A(g8630), .Z(II18545) ) ;
INV     gate6441  (.A(g8792), .Z(II18548) ) ;
INV     gate6442  (.A(g8824), .Z(II18551) ) ;
INV     gate6443  (.A(g8866), .Z(II18554) ) ;
INV     gate6444  (.A(g8810), .Z(II18557) ) ;
INV     gate6445  (.A(g8844), .Z(II18560) ) ;
INV     gate6446  (.A(g8897), .Z(II18563) ) ;
INV     gate6447  (.A(g8825), .Z(II18566) ) ;
INV     gate6448  (.A(g8867), .Z(II18569) ) ;
INV     gate6449  (.A(g8931), .Z(II18572) ) ;
INV     gate6450  (.A(g8845), .Z(II18575) ) ;
INV     gate6451  (.A(g8898), .Z(II18578) ) ;
INV     gate6452  (.A(g8964), .Z(II18581) ) ;
INV     gate6453  (.A(g8677), .Z(II18584) ) ;
INV     gate6454  (.A(g8718), .Z(II18587) ) ;
INV     gate6455  (.A(g8793), .Z(II18590) ) ;
INV     gate6456  (.A(g9390), .Z(II18593) ) ;
INV     gate6457  (.A(g8870), .Z(II18596) ) ;
INV     gate6458  (.A(g8933), .Z(II18599) ) ;
INV     gate6459  (.A(g9591), .Z(II18602) ) ;
INV     gate6460  (.A(g9786), .Z(II18605) ) ;
INV     gate6461  (.A(g10126), .Z(II18608) ) ;
INV     gate6462  (.A(g10909), .Z(II18611) ) ;
INV     gate6463  (.A(g11002), .Z(II18614) ) ;
INV     gate6464  (.A(g11169), .Z(II18617) ) ;
INV     gate6465  (.A(g11385), .Z(II18620) ) ;
INV     gate6466  (.A(g11003), .Z(II18623) ) ;
INV     gate6467  (.A(g8649), .Z(II18626) ) ;
INV     gate6468  (.A(g8811), .Z(II18629) ) ;
INV     gate6469  (.A(g8850), .Z(II18632) ) ;
INV     gate6470  (.A(g8904), .Z(II18635) ) ;
INV     gate6471  (.A(g8826), .Z(II18638) ) ;
INV     gate6472  (.A(g8871), .Z(II18641) ) ;
INV     gate6473  (.A(g8937), .Z(II18644) ) ;
INV     gate6474  (.A(g8851), .Z(II18647) ) ;
INV     gate6475  (.A(g8905), .Z(II18650) ) ;
INV     gate6476  (.A(g8971), .Z(II18653) ) ;
INV     gate6477  (.A(g8872), .Z(II18656) ) ;
INV     gate6478  (.A(g8938), .Z(II18659) ) ;
INV     gate6479  (.A(g8996), .Z(II18662) ) ;
INV     gate6480  (.A(g8689), .Z(II18665) ) ;
INV     gate6481  (.A(g8756), .Z(II18668) ) ;
INV     gate6482  (.A(g8812), .Z(II18671) ) ;
INV     gate6483  (.A(g9487), .Z(II18674) ) ;
INV     gate6484  (.A(g8908), .Z(II18677) ) ;
INV     gate6485  (.A(g8973), .Z(II18680) ) ;
INV     gate6486  (.A(g9733), .Z(II18683) ) ;
INV     gate6487  (.A(g9932), .Z(II18686) ) ;
INV     gate6488  (.A(g10231), .Z(II18689) ) ;
INV     gate6489  (.A(g10935), .Z(II18692) ) ;
INV     gate6490  (.A(g11054), .Z(II18695) ) ;
INV     gate6491  (.A(g11255), .Z(II18698) ) ;
INV     gate6492  (.A(g11471), .Z(II18701) ) ;
INV     gate6493  (.A(g11055), .Z(II18704) ) ;
INV     gate6494  (.A(g8665), .Z(II18707) ) ;
INV     gate6495  (.A(g8827), .Z(II18710) ) ;
INV     gate6496  (.A(g8877), .Z(II18713) ) ;
INV     gate6497  (.A(g8944), .Z(II18716) ) ;
INV     gate6498  (.A(g8852), .Z(II18719) ) ;
INV     gate6499  (.A(g8909), .Z(II18722) ) ;
INV     gate6500  (.A(g8977), .Z(II18725) ) ;
INV     gate6501  (.A(g8878), .Z(II18728) ) ;
INV     gate6502  (.A(g8945), .Z(II18731) ) ;
INV     gate6503  (.A(g9003), .Z(II18734) ) ;
INV     gate6504  (.A(g8910), .Z(II18737) ) ;
INV     gate6505  (.A(g8978), .Z(II18740) ) ;
INV     gate6506  (.A(g9025), .Z(II18743) ) ;
INV     gate6507  (.A(g8707), .Z(II18746) ) ;
INV     gate6508  (.A(g8779), .Z(II18749) ) ;
INV     gate6509  (.A(g8828), .Z(II18752) ) ;
INV     gate6510  (.A(g9629), .Z(II18755) ) ;
INV     gate6511  (.A(g8948), .Z(II18758) ) ;
INV     gate6512  (.A(g9005), .Z(II18761) ) ;
INV     gate6513  (.A(g9879), .Z(II18764) ) ;
INV     gate6514  (.A(g10086), .Z(II18767) ) ;
INV     gate6515  (.A(g10333), .Z(II18770) ) ;
INV     gate6516  (.A(g10830), .Z(II18773) ) ;
INV     gate6517  (.A(II18773), .Z(g11599) ) ;
INV     gate6518  (.A(g9050), .Z(II18777) ) ;
INV     gate6519  (.A(II18777), .Z(g11603) ) ;
INV     gate6520  (.A(g10870), .Z(II18780) ) ;
INV     gate6521  (.A(II18780), .Z(g11606) ) ;
INV     gate6522  (.A(g9067), .Z(II18784) ) ;
INV     gate6523  (.A(II18784), .Z(g11608) ) ;
INV     gate6524  (.A(g10910), .Z(II18787) ) ;
INV     gate6525  (.A(II18787), .Z(g11611) ) ;
INV     gate6526  (.A(g9084), .Z(II18791) ) ;
INV     gate6527  (.A(II18791), .Z(g11613) ) ;
INV     gate6528  (.A(g10973), .Z(II18794) ) ;
INV     gate6529  (.A(II18794), .Z(g11616) ) ;
INV     gate6530  (.A(g10601), .Z(g11620) ) ;
INV     gate6531  (.A(g10961), .Z(g11623) ) ;
INV     gate6532  (.A(g10813), .Z(II18810) ) ;
INV     gate6533  (.A(II18810), .Z(g11628) ) ;
INV     gate6534  (.A(g10850), .Z(II18813) ) ;
INV     gate6535  (.A(II18813), .Z(g11629) ) ;
INV     gate6536  (.A(g9067), .Z(II18817) ) ;
INV     gate6537  (.A(II18817), .Z(g11633) ) ;
INV     gate6538  (.A(g10890), .Z(II18820) ) ;
INV     gate6539  (.A(II18820), .Z(g11636) ) ;
INV     gate6540  (.A(g9084), .Z(II18824) ) ;
INV     gate6541  (.A(II18824), .Z(g11638) ) ;
INV     gate6542  (.A(g10936), .Z(II18827) ) ;
INV     gate6543  (.A(II18827), .Z(g11641) ) ;
INV     gate6544  (.A(g10646), .Z(g11642) ) ;
INV     gate6545  (.A(g10834), .Z(II18835) ) ;
INV     gate6546  (.A(II18835), .Z(g11651) ) ;
INV     gate6547  (.A(g10871), .Z(II18838) ) ;
INV     gate6548  (.A(II18838), .Z(g11652) ) ;
INV     gate6549  (.A(g9084), .Z(II18842) ) ;
INV     gate6550  (.A(II18842), .Z(g11656) ) ;
INV     gate6551  (.A(g10911), .Z(II18845) ) ;
INV     gate6552  (.A(II18845), .Z(g11659) ) ;
INV     gate6553  (.A(g10854), .Z(II18854) ) ;
INV     gate6554  (.A(II18854), .Z(g11670) ) ;
INV     gate6555  (.A(g10891), .Z(II18857) ) ;
INV     gate6556  (.A(II18857), .Z(g11671) ) ;
INV     gate6557  (.A(g10875), .Z(II18866) ) ;
INV     gate6558  (.A(II18866), .Z(g11682) ) ;
INV     gate6559  (.A(g10928), .Z(g11706) ) ;
INV     gate6560  (.A(g10826), .Z(g11732) ) ;
INV     gate6561  (.A(g10843), .Z(g11734) ) ;
INV     gate6562  (.A(g10859), .Z(g11735) ) ;
INV     gate6563  (.A(g10862), .Z(g11736) ) ;
INV     gate6564  (.A(g10809), .Z(g11737) ) ;
INV     gate6565  (.A(g10877), .Z(g11740) ) ;
INV     gate6566  (.A(g10880), .Z(g11741) ) ;
INV     gate6567  (.A(g10883), .Z(g11742) ) ;
INV     gate6568  (.A(g8530), .Z(g11743) ) ;
INV     gate6569  (.A(g10892), .Z(g11745) ) ;
INV     gate6570  (.A(g10895), .Z(g11746) ) ;
INV     gate6571  (.A(g10898), .Z(g11747) ) ;
INV     gate6572  (.A(g10901), .Z(g11748) ) ;
AND3    gate6573  (.A(g7595), .B(g7600), .C(II17599), .Z(g10711) ) ;
INV     gate6574  (.A(g10711), .Z(II18929) ) ;
INV     gate6575  (.A(II18929), .Z(g11749) ) ;
INV     gate6576  (.A(g8514), .Z(g11758) ) ;
INV     gate6577  (.A(g10912), .Z(g11761) ) ;
INV     gate6578  (.A(g10915), .Z(g11762) ) ;
INV     gate6579  (.A(g10918), .Z(g11763) ) ;
INV     gate6580  (.A(g10921), .Z(g11764) ) ;
INV     gate6581  (.A(g10924), .Z(g11765) ) ;
INV     gate6582  (.A(g10886), .Z(g11766) ) ;
INV     gate6583  (.A(g9149), .Z(II18943) ) ;
INV     gate6584  (.A(II18943), .Z(g11769) ) ;
INV     gate6585  (.A(g10932), .Z(g11770) ) ;
INV     gate6586  (.A(g10937), .Z(g11774) ) ;
INV     gate6587  (.A(g10940), .Z(g11775) ) ;
INV     gate6588  (.A(g10943), .Z(g11776) ) ;
INV     gate6589  (.A(g10946), .Z(g11777) ) ;
INV     gate6590  (.A(g10949), .Z(g11778) ) ;
INV     gate6591  (.A(g10906), .Z(g11779) ) ;
INV     gate6592  (.A(g10963), .Z(g11782) ) ;
INV     gate6593  (.A(g10966), .Z(g11783) ) ;
INV     gate6594  (.A(g9159), .Z(II18962) ) ;
INV     gate6595  (.A(II18962), .Z(g11786) ) ;
INV     gate6596  (.A(g10969), .Z(g11787) ) ;
INV     gate6597  (.A(g8726), .Z(II18969) ) ;
INV     gate6598  (.A(II18969), .Z(g11791) ) ;
INV     gate6599  (.A(g10974), .Z(g11794) ) ;
INV     gate6600  (.A(g10977), .Z(g11795) ) ;
INV     gate6601  (.A(g10980), .Z(g11796) ) ;
INV     gate6602  (.A(g10983), .Z(g11797) ) ;
INV     gate6603  (.A(g10867), .Z(g11798) ) ;
INV     gate6604  (.A(g10988), .Z(g11801) ) ;
INV     gate6605  (.A(g10991), .Z(g11802) ) ;
INV     gate6606  (.A(g10994), .Z(g11803) ) ;
INV     gate6607  (.A(g10995), .Z(g11804) ) ;
INV     gate6608  (.A(g10996), .Z(g11808) ) ;
INV     gate6609  (.A(g10999), .Z(g11809) ) ;
INV     gate6610  (.A(g9183), .Z(II18990) ) ;
INV     gate6611  (.A(II18990), .Z(g11812) ) ;
INV     gate6612  (.A(g11004), .Z(g11813) ) ;
INV     gate6613  (.A(g11008), .Z(g11817) ) ;
INV     gate6614  (.A(g11011), .Z(g11818) ) ;
INV     gate6615  (.A(g11014), .Z(g11819) ) ;
INV     gate6616  (.A(g11017), .Z(g11820) ) ;
INV     gate6617  (.A(g10848), .Z(g11821) ) ;
INV     gate6618  (.A(g11022), .Z(g11824) ) ;
INV     gate6619  (.A(g11025), .Z(g11825) ) ;
INV     gate6620  (.A(g11028), .Z(g11826) ) ;
INV     gate6621  (.A(g11032), .Z(g11827) ) ;
INV     gate6622  (.A(g11035), .Z(g11829) ) ;
INV     gate6623  (.A(g11036), .Z(g11834) ) ;
INV     gate6624  (.A(g11039), .Z(g11835) ) ;
INV     gate6625  (.A(g11042), .Z(g11836) ) ;
INV     gate6626  (.A(g11045), .Z(g11837) ) ;
INV     gate6627  (.A(g11048), .Z(g11841) ) ;
INV     gate6628  (.A(g11051), .Z(g11842) ) ;
INV     gate6629  (.A(g9225), .Z(II19025) ) ;
INV     gate6630  (.A(II19025), .Z(g11845) ) ;
INV     gate6631  (.A(g11056), .Z(g11846) ) ;
INV     gate6632  (.A(g8726), .Z(II19030) ) ;
INV     gate6633  (.A(II19030), .Z(g11848) ) ;
INV     gate6634  (.A(g11063), .Z(g11852) ) ;
INV     gate6635  (.A(g11066), .Z(g11853) ) ;
INV     gate6636  (.A(g11078), .Z(g11854) ) ;
INV     gate6637  (.A(g11079), .Z(g11856) ) ;
INV     gate6638  (.A(g11082), .Z(g11857) ) ;
INV     gate6639  (.A(g11085), .Z(g11858) ) ;
INV     gate6640  (.A(g11088), .Z(g11859) ) ;
INV     gate6641  (.A(g11091), .Z(g11862) ) ;
INV     gate6642  (.A(g11092), .Z(g11866) ) ;
INV     gate6643  (.A(g11095), .Z(g11867) ) ;
INV     gate6644  (.A(g11098), .Z(g11868) ) ;
INV     gate6645  (.A(g11102), .Z(g11869) ) ;
INV     gate6646  (.A(g11105), .Z(g11871) ) ;
INV     gate6647  (.A(g11108), .Z(g11876) ) ;
INV     gate6648  (.A(g11111), .Z(g11877) ) ;
INV     gate6649  (.A(g11114), .Z(g11878) ) ;
INV     gate6650  (.A(g11117), .Z(g11879) ) ;
INV     gate6651  (.A(g11120), .Z(g11883) ) ;
INV     gate6652  (.A(g11123), .Z(g11884) ) ;
INV     gate6653  (.A(g11126), .Z(g11886) ) ;
INV     gate6654  (.A(g11129), .Z(g11887) ) ;
INV     gate6655  (.A(g11021), .Z(g11888) ) ;
INV     gate6656  (.A(g11132), .Z(g11891) ) ;
INV     gate6657  (.A(g11135), .Z(g11892) ) ;
INV     gate6658  (.A(g11138), .Z(g11893) ) ;
INV     gate6659  (.A(g11141), .Z(g11894) ) ;
INV     gate6660  (.A(g11144), .Z(g11895) ) ;
INV     gate6661  (.A(g11145), .Z(g11898) ) ;
INV     gate6662  (.A(g11148), .Z(g11899) ) ;
INV     gate6663  (.A(g11151), .Z(g11900) ) ;
INV     gate6664  (.A(g11154), .Z(g11901) ) ;
INV     gate6665  (.A(g11157), .Z(g11904) ) ;
INV     gate6666  (.A(g11160), .Z(g11908) ) ;
INV     gate6667  (.A(g11163), .Z(g11909) ) ;
INV     gate6668  (.A(g11166), .Z(g11910) ) ;
INV     gate6669  (.A(g11170), .Z(g11911) ) ;
INV     gate6670  (.A(g11173), .Z(g11913) ) ;
INV     gate6671  (.A(g11176), .Z(g11918) ) ;
INV     gate6672  (.A(g11179), .Z(g11919) ) ;
INV     gate6673  (.A(g11182), .Z(g11920) ) ;
INV     gate6674  (.A(g11185), .Z(g11921) ) ;
INV     gate6675  (.A(g8726), .Z(II19105) ) ;
INV     gate6676  (.A(II19105), .Z(g11923) ) ;
INV     gate6677  (.A(g10987), .Z(g11927) ) ;
INV     gate6678  (.A(g11199), .Z(g11929) ) ;
INV     gate6679  (.A(g11202), .Z(g11930) ) ;
INV     gate6680  (.A(g11205), .Z(g11931) ) ;
INV     gate6681  (.A(g11209), .Z(g11932) ) ;
INV     gate6682  (.A(g11210), .Z(g11933) ) ;
INV     gate6683  (.A(g11213), .Z(g11936) ) ;
INV     gate6684  (.A(g9202), .Z(II19119) ) ;
INV     gate6685  (.A(II19119), .Z(g11937) ) ;
INV     gate6686  (.A(g11216), .Z(g11941) ) ;
INV     gate6687  (.A(g11219), .Z(g11942) ) ;
INV     gate6688  (.A(g11222), .Z(g11943) ) ;
INV     gate6689  (.A(g11225), .Z(g11944) ) ;
INV     gate6690  (.A(g11228), .Z(g11945) ) ;
INV     gate6691  (.A(g11231), .Z(g11948) ) ;
INV     gate6692  (.A(g11234), .Z(g11949) ) ;
INV     gate6693  (.A(g11237), .Z(g11950) ) ;
INV     gate6694  (.A(g11240), .Z(g11951) ) ;
INV     gate6695  (.A(g11243), .Z(g11954) ) ;
INV     gate6696  (.A(g11246), .Z(g11958) ) ;
INV     gate6697  (.A(g11249), .Z(g11959) ) ;
INV     gate6698  (.A(g11252), .Z(g11960) ) ;
INV     gate6699  (.A(g11256), .Z(g11961) ) ;
INV     gate6700  (.A(g11259), .Z(g11963) ) ;
INV     gate6701  (.A(g11265), .Z(g11968) ) ;
INV     gate6702  (.A(g11268), .Z(g11969) ) ;
INV     gate6703  (.A(g11271), .Z(g11970) ) ;
INV     gate6704  (.A(g11274), .Z(g11971) ) ;
INV     gate6705  (.A(g11277), .Z(g11972) ) ;
INV     gate6706  (.A(g11278), .Z(g11973) ) ;
INV     gate6707  (.A(g10549), .Z(II19160) ) ;
INV     gate6708  (.A(II19160), .Z(g11976) ) ;
INV     gate6709  (.A(g11281), .Z(g11982) ) ;
INV     gate6710  (.A(g11284), .Z(g11983) ) ;
INV     gate6711  (.A(g11287), .Z(g11984) ) ;
INV     gate6712  (.A(g11291), .Z(g11985) ) ;
INV     gate6713  (.A(g11294), .Z(g11986) ) ;
INV     gate6714  (.A(g11297), .Z(g11989) ) ;
INV     gate6715  (.A(g9263), .Z(II19174) ) ;
INV     gate6716  (.A(II19174), .Z(g11990) ) ;
INV     gate6717  (.A(g11300), .Z(g11994) ) ;
INV     gate6718  (.A(g11303), .Z(g11995) ) ;
INV     gate6719  (.A(g11306), .Z(g11996) ) ;
INV     gate6720  (.A(g11309), .Z(g11997) ) ;
INV     gate6721  (.A(g11312), .Z(g11998) ) ;
INV     gate6722  (.A(g11315), .Z(g12001) ) ;
INV     gate6723  (.A(g11318), .Z(g12002) ) ;
INV     gate6724  (.A(g11321), .Z(g12003) ) ;
INV     gate6725  (.A(g11324), .Z(g12004) ) ;
INV     gate6726  (.A(g11327), .Z(g12007) ) ;
INV     gate6727  (.A(g8726), .Z(II19195) ) ;
INV     gate6728  (.A(II19195), .Z(g12009) ) ;
INV     gate6729  (.A(g10772), .Z(g12013) ) ;
INV     gate6730  (.A(g10100), .Z(g12017) ) ;
INV     gate6731  (.A(g11341), .Z(g12020) ) ;
INV     gate6732  (.A(g11344), .Z(g12021) ) ;
INV     gate6733  (.A(g11348), .Z(g12022) ) ;
INV     gate6734  (.A(g11351), .Z(g12023) ) ;
INV     gate6735  (.A(g11354), .Z(g12024) ) ;
INV     gate6736  (.A(g11355), .Z(g12025) ) ;
INV     gate6737  (.A(g10424), .Z(II19208) ) ;
INV     gate6738  (.A(II19208), .Z(g12027) ) ;
INV     gate6739  (.A(g10486), .Z(II19211) ) ;
INV     gate6740  (.A(II19211), .Z(g12030) ) ;
INV     gate6741  (.A(g11358), .Z(g12037) ) ;
INV     gate6742  (.A(g11361), .Z(g12038) ) ;
INV     gate6743  (.A(g11364), .Z(g12039) ) ;
INV     gate6744  (.A(g11367), .Z(g12040) ) ;
INV     gate6745  (.A(g11370), .Z(g12041) ) ;
INV     gate6746  (.A(g11373), .Z(g12042) ) ;
INV     gate6747  (.A(g10606), .Z(II19226) ) ;
INV     gate6748  (.A(II19226), .Z(g12045) ) ;
INV     gate6749  (.A(g11376), .Z(g12051) ) ;
INV     gate6750  (.A(g11379), .Z(g12052) ) ;
INV     gate6751  (.A(g11382), .Z(g12053) ) ;
INV     gate6752  (.A(g11386), .Z(g12054) ) ;
INV     gate6753  (.A(g11389), .Z(g12055) ) ;
INV     gate6754  (.A(g11392), .Z(g12058) ) ;
INV     gate6755  (.A(g9341), .Z(II19240) ) ;
INV     gate6756  (.A(II19240), .Z(g12059) ) ;
INV     gate6757  (.A(g11395), .Z(g12063) ) ;
INV     gate6758  (.A(g11398), .Z(g12064) ) ;
INV     gate6759  (.A(g11401), .Z(g12065) ) ;
INV     gate6760  (.A(g11404), .Z(g12066) ) ;
INV     gate6761  (.A(g11407), .Z(g12067) ) ;
INV     gate6762  (.A(g10783), .Z(g12071) ) ;
INV     gate6763  (.A(g11411), .Z(g12075) ) ;
INV     gate6764  (.A(g11414), .Z(g12076) ) ;
INV     gate6765  (.A(g11417), .Z(g12077) ) ;
INV     gate6766  (.A(g11422), .Z(g12078) ) ;
INV     gate6767  (.A(g11425), .Z(g12084) ) ;
INV     gate6768  (.A(g11428), .Z(g12085) ) ;
INV     gate6769  (.A(g11432), .Z(g12086) ) ;
INV     gate6770  (.A(g11435), .Z(g12087) ) ;
INV     gate6771  (.A(g11438), .Z(g12088) ) ;
INV     gate6772  (.A(g11441), .Z(g12089) ) ;
INV     gate6773  (.A(g10500), .Z(II19271) ) ;
INV     gate6774  (.A(II19271), .Z(g12091) ) ;
INV     gate6775  (.A(g10560), .Z(II19274) ) ;
INV     gate6776  (.A(II19274), .Z(g12094) ) ;
INV     gate6777  (.A(g11444), .Z(g12101) ) ;
INV     gate6778  (.A(g11447), .Z(g12102) ) ;
INV     gate6779  (.A(g11450), .Z(g12103) ) ;
INV     gate6780  (.A(g11453), .Z(g12104) ) ;
INV     gate6781  (.A(g11456), .Z(g12105) ) ;
INV     gate6782  (.A(g11459), .Z(g12106) ) ;
INV     gate6783  (.A(g10653), .Z(II19289) ) ;
INV     gate6784  (.A(II19289), .Z(g12109) ) ;
INV     gate6785  (.A(g11462), .Z(g12115) ) ;
INV     gate6786  (.A(g11465), .Z(g12116) ) ;
INV     gate6787  (.A(g11468), .Z(g12117) ) ;
INV     gate6788  (.A(g11472), .Z(g12118) ) ;
INV     gate6789  (.A(g11475), .Z(g12119) ) ;
INV     gate6790  (.A(g11478), .Z(g12122) ) ;
INV     gate6791  (.A(g9422), .Z(II19303) ) ;
INV     gate6792  (.A(II19303), .Z(g12123) ) ;
INV     gate6793  (.A(g8726), .Z(II19307) ) ;
INV     gate6794  (.A(II19307), .Z(g12125) ) ;
INV     gate6795  (.A(g10788), .Z(g12130) ) ;
INV     gate6796  (.A(g8321), .Z(g12134) ) ;
INV     gate6797  (.A(g8324), .Z(g12135) ) ;
INV     gate6798  (.A(g10424), .Z(II19315) ) ;
INV     gate6799  (.A(II19315), .Z(g12136) ) ;
INV     gate6800  (.A(g10486), .Z(II19318) ) ;
INV     gate6801  (.A(II19318), .Z(g12139) ) ;
INV     gate6802  (.A(g10549), .Z(II19321) ) ;
INV     gate6803  (.A(II19321), .Z(g12142) ) ;
INV     gate6804  (.A(g8330), .Z(g12147) ) ;
INV     gate6805  (.A(g8333), .Z(g12148) ) ;
INV     gate6806  (.A(g8336), .Z(g12149) ) ;
INV     gate6807  (.A(g8341), .Z(g12150) ) ;
INV     gate6808  (.A(g8344), .Z(g12156) ) ;
INV     gate6809  (.A(g8347), .Z(g12157) ) ;
INV     gate6810  (.A(g8351), .Z(g12158) ) ;
INV     gate6811  (.A(g8354), .Z(g12159) ) ;
INV     gate6812  (.A(g8357), .Z(g12160) ) ;
INV     gate6813  (.A(g8360), .Z(g12161) ) ;
INV     gate6814  (.A(g10574), .Z(II19342) ) ;
INV     gate6815  (.A(II19342), .Z(g12163) ) ;
INV     gate6816  (.A(g10617), .Z(II19345) ) ;
INV     gate6817  (.A(II19345), .Z(g12166) ) ;
INV     gate6818  (.A(g8363), .Z(g12173) ) ;
INV     gate6819  (.A(g8366), .Z(g12174) ) ;
INV     gate6820  (.A(g8369), .Z(g12175) ) ;
INV     gate6821  (.A(g8372), .Z(g12176) ) ;
INV     gate6822  (.A(g8375), .Z(g12177) ) ;
INV     gate6823  (.A(g8378), .Z(g12178) ) ;
INV     gate6824  (.A(g10683), .Z(II19360) ) ;
INV     gate6825  (.A(II19360), .Z(g12181) ) ;
INV     gate6826  (.A(g8285), .Z(g12187) ) ;
INV     gate6827  (.A(g8382), .Z(g12191) ) ;
INV     gate6828  (.A(g8388), .Z(g12196) ) ;
INV     gate6829  (.A(g8391), .Z(g12197) ) ;
INV     gate6830  (.A(g10500), .Z(II19374) ) ;
INV     gate6831  (.A(II19374), .Z(g12198) ) ;
INV     gate6832  (.A(g10560), .Z(II19377) ) ;
INV     gate6833  (.A(II19377), .Z(g12201) ) ;
INV     gate6834  (.A(g10606), .Z(II19380) ) ;
INV     gate6835  (.A(II19380), .Z(g12204) ) ;
INV     gate6836  (.A(g8397), .Z(g12209) ) ;
INV     gate6837  (.A(g8400), .Z(g12210) ) ;
INV     gate6838  (.A(g8403), .Z(g12211) ) ;
INV     gate6839  (.A(g8408), .Z(g12212) ) ;
INV     gate6840  (.A(g8411), .Z(g12218) ) ;
INV     gate6841  (.A(g8414), .Z(g12219) ) ;
INV     gate6842  (.A(g8418), .Z(g12220) ) ;
INV     gate6843  (.A(g8421), .Z(g12221) ) ;
INV     gate6844  (.A(g8424), .Z(g12222) ) ;
INV     gate6845  (.A(g8427), .Z(g12223) ) ;
INV     gate6846  (.A(g10631), .Z(II19401) ) ;
INV     gate6847  (.A(II19401), .Z(g12225) ) ;
INV     gate6848  (.A(g10664), .Z(II19404) ) ;
INV     gate6849  (.A(II19404), .Z(g12228) ) ;
INV     gate6850  (.A(g8294), .Z(g12235) ) ;
INV     gate6851  (.A(g10486), .Z(II19412) ) ;
INV     gate6852  (.A(II19412), .Z(g12239) ) ;
INV     gate6853  (.A(g10549), .Z(II19415) ) ;
INV     gate6854  (.A(II19415), .Z(g12242) ) ;
INV     gate6855  (.A(g8434), .Z(g12246) ) ;
INV     gate6856  (.A(g8440), .Z(g12251) ) ;
INV     gate6857  (.A(g8443), .Z(g12252) ) ;
INV     gate6858  (.A(g10574), .Z(II19426) ) ;
INV     gate6859  (.A(II19426), .Z(g12253) ) ;
INV     gate6860  (.A(g10617), .Z(II19429) ) ;
INV     gate6861  (.A(II19429), .Z(g12256) ) ;
INV     gate6862  (.A(g10653), .Z(II19432) ) ;
INV     gate6863  (.A(II19432), .Z(g12259) ) ;
INV     gate6864  (.A(g8449), .Z(g12264) ) ;
INV     gate6865  (.A(g8452), .Z(g12265) ) ;
INV     gate6866  (.A(g8455), .Z(g12266) ) ;
INV     gate6867  (.A(g8460), .Z(g12267) ) ;
INV     gate6868  (.A(g8303), .Z(g12275) ) ;
INV     gate6869  (.A(g10424), .Z(II19449) ) ;
INV     gate6870  (.A(II19449), .Z(g12279) ) ;
INV     gate6871  (.A(g10560), .Z(II19452) ) ;
INV     gate6872  (.A(II19452), .Z(g12282) ) ;
INV     gate6873  (.A(g10606), .Z(II19455) ) ;
INV     gate6874  (.A(II19455), .Z(g12285) ) ;
INV     gate6875  (.A(g8469), .Z(g12289) ) ;
INV     gate6876  (.A(g8475), .Z(g12294) ) ;
INV     gate6877  (.A(g8478), .Z(g12295) ) ;
INV     gate6878  (.A(g10631), .Z(II19466) ) ;
INV     gate6879  (.A(II19466), .Z(g12296) ) ;
INV     gate6880  (.A(g10664), .Z(II19469) ) ;
INV     gate6881  (.A(II19469), .Z(g12299) ) ;
INV     gate6882  (.A(g10683), .Z(II19472) ) ;
INV     gate6883  (.A(II19472), .Z(g12302) ) ;
INV     gate6884  (.A(g8312), .Z(g12308) ) ;
INV     gate6885  (.A(g10549), .Z(II19479) ) ;
INV     gate6886  (.A(II19479), .Z(g12312) ) ;
INV     gate6887  (.A(g10500), .Z(II19482) ) ;
INV     gate6888  (.A(II19482), .Z(g12315) ) ;
INV     gate6889  (.A(g10617), .Z(II19485) ) ;
INV     gate6890  (.A(II19485), .Z(g12318) ) ;
INV     gate6891  (.A(g10653), .Z(II19488) ) ;
INV     gate6892  (.A(II19488), .Z(g12321) ) ;
INV     gate6893  (.A(g8494), .Z(g12325) ) ;
INV     gate6894  (.A(g10829), .Z(g12332) ) ;
INV     gate6895  (.A(g10424), .Z(II19500) ) ;
INV     gate6896  (.A(II19500), .Z(g12333) ) ;
INV     gate6897  (.A(g10486), .Z(II19503) ) ;
INV     gate6898  (.A(II19503), .Z(g12336) ) ;
INV     gate6899  (.A(g10606), .Z(II19507) ) ;
INV     gate6900  (.A(II19507), .Z(g12340) ) ;
INV     gate6901  (.A(g10574), .Z(II19510) ) ;
INV     gate6902  (.A(II19510), .Z(g12343) ) ;
INV     gate6903  (.A(g10664), .Z(II19513) ) ;
INV     gate6904  (.A(II19513), .Z(g12346) ) ;
INV     gate6905  (.A(g10683), .Z(II19516) ) ;
INV     gate6906  (.A(II19516), .Z(g12349) ) ;
NAND4   gate6907  (.A(g8182), .B(g8120), .C(g8044), .D(g7989), .Z(g8381) ) ;
INV     gate6908  (.A(g8381), .Z(g12354) ) ;
INV     gate6909  (.A(g10866), .Z(g12362) ) ;
INV     gate6910  (.A(g10500), .Z(II19523) ) ;
INV     gate6911  (.A(II19523), .Z(g12363) ) ;
INV     gate6912  (.A(g10560), .Z(II19526) ) ;
INV     gate6913  (.A(II19526), .Z(g12366) ) ;
INV     gate6914  (.A(g10653), .Z(II19530) ) ;
INV     gate6915  (.A(II19530), .Z(g12370) ) ;
INV     gate6916  (.A(g10631), .Z(II19533) ) ;
INV     gate6917  (.A(II19533), .Z(g12373) ) ;
INV     gate6918  (.A(g10847), .Z(g12378) ) ;
INV     gate6919  (.A(g10549), .Z(II19539) ) ;
INV     gate6920  (.A(II19539), .Z(g12379) ) ;
INV     gate6921  (.A(g10574), .Z(II19542) ) ;
INV     gate6922  (.A(II19542), .Z(g12382) ) ;
INV     gate6923  (.A(g10617), .Z(II19545) ) ;
INV     gate6924  (.A(II19545), .Z(g12385) ) ;
INV     gate6925  (.A(g10683), .Z(II19549) ) ;
INV     gate6926  (.A(II19549), .Z(g12389) ) ;
NOR4    gate6927  (.A(g3198), .B(g8120), .C(g3194), .D(g3191), .Z(g8430) ) ;
INV     gate6928  (.A(g8430), .Z(II19552) ) ;
INV     gate6929  (.A(II19552), .Z(g12392) ) ;
INV     gate6930  (.A(g11020), .Z(g12408) ) ;
INV     gate6931  (.A(g10606), .Z(II19557) ) ;
INV     gate6932  (.A(II19557), .Z(g12409) ) ;
INV     gate6933  (.A(g10631), .Z(II19560) ) ;
INV     gate6934  (.A(II19560), .Z(g12412) ) ;
INV     gate6935  (.A(g10664), .Z(II19563) ) ;
INV     gate6936  (.A(II19563), .Z(g12415) ) ;
INV     gate6937  (.A(g10986), .Z(g12420) ) ;
INV     gate6938  (.A(g10653), .Z(II19569) ) ;
INV     gate6939  (.A(II19569), .Z(g12421) ) ;
INV     gate6940  (.A(g10962), .Z(g12424) ) ;
INV     gate6941  (.A(g8835), .Z(II19573) ) ;
INV     gate6942  (.A(II19573), .Z(g12425) ) ;
INV     gate6943  (.A(g10683), .Z(II19576) ) ;
INV     gate6944  (.A(II19576), .Z(g12426) ) ;
INV     gate6945  (.A(g10905), .Z(g12430) ) ;
INV     gate6946  (.A(g8862), .Z(II19582) ) ;
INV     gate6947  (.A(II19582), .Z(g12432) ) ;
INV     gate6948  (.A(g10929), .Z(g12434) ) ;
INV     gate6949  (.A(g9173), .Z(II19587) ) ;
INV     gate6950  (.A(II19587), .Z(g12435) ) ;
INV     gate6951  (.A(g8900), .Z(II19591) ) ;
INV     gate6952  (.A(II19591), .Z(g12437) ) ;
INV     gate6953  (.A(g10846), .Z(g12438) ) ;
NOR3    gate6954  (.A(g5711), .B(g5758), .C(g5807), .Z(g10810) ) ;
INV     gate6955  (.A(g10810), .Z(II19595) ) ;
INV     gate6956  (.A(II19595), .Z(g12439) ) ;
INV     gate6957  (.A(g9215), .Z(II19598) ) ;
INV     gate6958  (.A(II19598), .Z(g12440) ) ;
INV     gate6959  (.A(g8940), .Z(II19602) ) ;
INV     gate6960  (.A(II19602), .Z(g12442) ) ;
NOR3    gate6961  (.A(g5678), .B(g5710), .C(g5757), .Z(g10797) ) ;
INV     gate6962  (.A(g10797), .Z(II19605) ) ;
INV     gate6963  (.A(II19605), .Z(g12443) ) ;
NOR3    gate6964  (.A(g5769), .B(g5817), .C(g5863), .Z(g10831) ) ;
INV     gate6965  (.A(g10831), .Z(II19608) ) ;
INV     gate6966  (.A(II19608), .Z(g12444) ) ;
INV     gate6967  (.A(g9276), .Z(II19611) ) ;
INV     gate6968  (.A(II19611), .Z(g12445) ) ;
NOR3    gate6969  (.A(g5650), .B(g5677), .C(g5709), .Z(g10789) ) ;
INV     gate6970  (.A(g10789), .Z(II19615) ) ;
INV     gate6971  (.A(II19615), .Z(g12447) ) ;
NOR3    gate6972  (.A(g5730), .B(g5768), .C(g5816), .Z(g10814) ) ;
INV     gate6973  (.A(g10814), .Z(II19618) ) ;
INV     gate6974  (.A(II19618), .Z(g12448) ) ;
NOR3    gate6975  (.A(g5828), .B(g5873), .C(g5910), .Z(g10851) ) ;
INV     gate6976  (.A(g10851), .Z(II19621) ) ;
INV     gate6977  (.A(II19621), .Z(g12449) ) ;
INV     gate6978  (.A(g9354), .Z(II19624) ) ;
INV     gate6979  (.A(II19624), .Z(g12450) ) ;
NOR3    gate6980  (.A(g5630), .B(g5649), .C(g5676), .Z(g10784) ) ;
INV     gate6981  (.A(g10784), .Z(II19628) ) ;
INV     gate6982  (.A(II19628), .Z(g12452) ) ;
NOR3    gate6983  (.A(g5688), .B(g5729), .C(g5767), .Z(g10801) ) ;
INV     gate6984  (.A(g10801), .Z(II19631) ) ;
INV     gate6985  (.A(II19631), .Z(g12453) ) ;
NOR3    gate6986  (.A(g5788), .B(g5827), .C(g5872), .Z(g10835) ) ;
INV     gate6987  (.A(g10835), .Z(II19634) ) ;
INV     gate6988  (.A(II19634), .Z(g12454) ) ;
NOR3    gate6989  (.A(g5884), .B(g5920), .C(g5949), .Z(g10872) ) ;
INV     gate6990  (.A(g10872), .Z(II19637) ) ;
INV     gate6991  (.A(II19637), .Z(g12455) ) ;
INV     gate6992  (.A(g8602), .Z(g12456) ) ;
NOR3    gate6993  (.A(g5658), .B(g5687), .C(g5728), .Z(g10793) ) ;
INV     gate6994  (.A(g10793), .Z(II19642) ) ;
INV     gate6995  (.A(II19642), .Z(g12460) ) ;
NOR3    gate6996  (.A(g5740), .B(g5787), .C(g5826), .Z(g10818) ) ;
INV     gate6997  (.A(g10818), .Z(II19645) ) ;
INV     gate6998  (.A(II19645), .Z(g12461) ) ;
NOR3    gate6999  (.A(g5847), .B(g5883), .C(g5919), .Z(g10855) ) ;
INV     gate7000  (.A(g10855), .Z(II19648) ) ;
INV     gate7001  (.A(II19648), .Z(g12462) ) ;
INV     gate7002  (.A(g10730), .Z(g12463) ) ;
INV     gate7003  (.A(g8614), .Z(g12466) ) ;
NOR3    gate7004  (.A(g5696), .B(g5739), .C(g5786), .Z(g10805) ) ;
INV     gate7005  (.A(g10805), .Z(II19654) ) ;
INV     gate7006  (.A(II19654), .Z(g12470) ) ;
NOR3    gate7007  (.A(g5798), .B(g5846), .C(g5882), .Z(g10839) ) ;
INV     gate7008  (.A(g10839), .Z(II19657) ) ;
INV     gate7009  (.A(II19657), .Z(g12471) ) ;
INV     gate7010  (.A(g8617), .Z(g12472) ) ;
INV     gate7011  (.A(g8580), .Z(g12473) ) ;
INV     gate7012  (.A(g8622), .Z(g12476) ) ;
INV     gate7013  (.A(g10749), .Z(g12478) ) ;
INV     gate7014  (.A(g8627), .Z(g12481) ) ;
NOR3    gate7015  (.A(g5748), .B(g5797), .C(g5845), .Z(g10822) ) ;
INV     gate7016  (.A(g10822), .Z(II19667) ) ;
INV     gate7017  (.A(II19667), .Z(g12485) ) ;
INV     gate7018  (.A(g8587), .Z(g12490) ) ;
INV     gate7019  (.A(g8632), .Z(g12493) ) ;
INV     gate7020  (.A(g10767), .Z(g12495) ) ;
INV     gate7021  (.A(g8637), .Z(g12498) ) ;
INV     gate7022  (.A(g8640), .Z(g12502) ) ;
INV     gate7023  (.A(g8643), .Z(g12504) ) ;
INV     gate7024  (.A(g8646), .Z(g12505) ) ;
INV     gate7025  (.A(g8594), .Z(g12510) ) ;
INV     gate7026  (.A(g8651), .Z(g12513) ) ;
INV     gate7027  (.A(g10773), .Z(g12515) ) ;
INV     gate7028  (.A(g8655), .Z(g12518) ) ;
INV     gate7029  (.A(g10016), .Z(II19689) ) ;
INV     gate7030  (.A(II19689), .Z(g12519) ) ;
INV     gate7031  (.A(g8659), .Z(g12521) ) ;
INV     gate7032  (.A(g8662), .Z(g12522) ) ;
INV     gate7033  (.A(g8605), .Z(g12527) ) ;
INV     gate7034  (.A(g8667), .Z(g12530) ) ;
INV     gate7035  (.A(g8670), .Z(g12532) ) ;
INV     gate7036  (.A(g8673), .Z(g12533) ) ;
INV     gate7037  (.A(g10125), .Z(II19702) ) ;
INV     gate7038  (.A(II19702), .Z(g12534) ) ;
INV     gate7039  (.A(g8678), .Z(g12536) ) ;
INV     gate7040  (.A(g8681), .Z(g12537) ) ;
INV     gate7041  (.A(g8684), .Z(g12542) ) ;
INV     gate7042  (.A(g10230), .Z(II19711) ) ;
INV     gate7043  (.A(II19711), .Z(g12543) ) ;
INV     gate7044  (.A(g8690), .Z(g12545) ) ;
INV     gate7045  (.A(g8693), .Z(g12546) ) ;
INV     gate7046  (.A(g8696), .Z(g12547) ) ;
INV     gate7047  (.A(g8726), .Z(II19718) ) ;
INV     gate7048  (.A(II19718), .Z(g12548) ) ;
INV     gate7049  (.A(g8700), .Z(g12551) ) ;
INV     gate7050  (.A(g10332), .Z(II19722) ) ;
INV     gate7051  (.A(II19722), .Z(g12552) ) ;
INV     gate7052  (.A(g8708), .Z(g12553) ) ;
INV     gate7053  (.A(g8711), .Z(g12554) ) ;
INV     gate7054  (.A(g8726), .Z(II19727) ) ;
INV     gate7055  (.A(II19727), .Z(g12555) ) ;
INV     gate7056  (.A(g8714), .Z(g12558) ) ;
INV     gate7057  (.A(g8719), .Z(g12559) ) ;
INV     gate7058  (.A(g8745), .Z(g12560) ) ;
INV     gate7059  (.A(g8726), .Z(II19733) ) ;
INV     gate7060  (.A(II19733), .Z(g12561) ) ;
INV     gate7061  (.A(g9184), .Z(II19736) ) ;
INV     gate7062  (.A(II19736), .Z(g12564) ) ;
INV     gate7063  (.A(g10694), .Z(II19739) ) ;
INV     gate7064  (.A(II19739), .Z(g12565) ) ;
INV     gate7065  (.A(g8748), .Z(g12596) ) ;
INV     gate7066  (.A(g8752), .Z(g12597) ) ;
INV     gate7067  (.A(g8757), .Z(g12598) ) ;
INV     gate7068  (.A(g8763), .Z(g12599) ) ;
INV     gate7069  (.A(g8766), .Z(g12600) ) ;
INV     gate7070  (.A(g8726), .Z(II19747) ) ;
INV     gate7071  (.A(II19747), .Z(g12601) ) ;
INV     gate7072  (.A(g8726), .Z(II19750) ) ;
INV     gate7073  (.A(II19750), .Z(g12604) ) ;
INV     gate7074  (.A(g9229), .Z(II19753) ) ;
INV     gate7075  (.A(II19753), .Z(g12607) ) ;
INV     gate7076  (.A(g10424), .Z(II19756) ) ;
INV     gate7077  (.A(II19756), .Z(g12608) ) ;
INV     gate7078  (.A(g10714), .Z(II19759) ) ;
INV     gate7079  (.A(II19759), .Z(g12611) ) ;
INV     gate7080  (.A(g8771), .Z(g12642) ) ;
INV     gate7081  (.A(g8775), .Z(g12643) ) ;
INV     gate7082  (.A(g8780), .Z(g12644) ) ;
INV     gate7083  (.A(g8785), .Z(g12645) ) ;
INV     gate7084  (.A(g8788), .Z(g12646) ) ;
INV     gate7085  (.A(g8726), .Z(II19767) ) ;
INV     gate7086  (.A(II19767), .Z(g12647) ) ;
NAND2   gate7087  (.A(g7772), .B(g3366), .Z(g10038) ) ;
INV     gate7088  (.A(g10038), .Z(II19771) ) ;
INV     gate7089  (.A(II19771), .Z(g12651) ) ;
INV     gate7090  (.A(g10500), .Z(II19774) ) ;
INV     gate7091  (.A(II19774), .Z(g12654) ) ;
INV     gate7092  (.A(g10735), .Z(II19777) ) ;
INV     gate7093  (.A(II19777), .Z(g12657) ) ;
INV     gate7094  (.A(g8794), .Z(g12688) ) ;
INV     gate7095  (.A(g8798), .Z(g12689) ) ;
INV     gate7096  (.A(g8802), .Z(g12690) ) ;
INV     gate7097  (.A(g8805), .Z(g12691) ) ;
INV     gate7098  (.A(g8726), .Z(II19784) ) ;
INV     gate7099  (.A(II19784), .Z(g12692) ) ;
INV     gate7100  (.A(g8726), .Z(II19787) ) ;
INV     gate7101  (.A(II19787), .Z(g12695) ) ;
INV     gate7102  (.A(g10486), .Z(II19791) ) ;
INV     gate7103  (.A(II19791), .Z(g12699) ) ;
NAND2   gate7104  (.A(g3398), .B(g6678), .Z(g10676) ) ;
INV     gate7105  (.A(g10676), .Z(II19794) ) ;
INV     gate7106  (.A(II19794), .Z(g12702) ) ;
NAND2   gate7107  (.A(g7788), .B(g3522), .Z(g10147) ) ;
INV     gate7108  (.A(g10147), .Z(II19797) ) ;
INV     gate7109  (.A(II19797), .Z(g12705) ) ;
INV     gate7110  (.A(g10574), .Z(II19800) ) ;
INV     gate7111  (.A(II19800), .Z(g12708) ) ;
INV     gate7112  (.A(g10754), .Z(II19803) ) ;
INV     gate7113  (.A(II19803), .Z(g12711) ) ;
INV     gate7114  (.A(g8813), .Z(g12742) ) ;
INV     gate7115  (.A(g8817), .Z(g12743) ) ;
INV     gate7116  (.A(g8726), .Z(II19808) ) ;
INV     gate7117  (.A(II19808), .Z(g12744) ) ;
INV     gate7118  (.A(g8823), .Z(g12748) ) ;
NAND2   gate7119  (.A(g3398), .B(g6912), .Z(g10649) ) ;
INV     gate7120  (.A(g10649), .Z(II19813) ) ;
INV     gate7121  (.A(II19813), .Z(g12749) ) ;
NAND2   gate7122  (.A(g3398), .B(g6678), .Z(g10703) ) ;
INV     gate7123  (.A(g10703), .Z(II19816) ) ;
INV     gate7124  (.A(II19816), .Z(g12752) ) ;
INV     gate7125  (.A(g10560), .Z(II19820) ) ;
INV     gate7126  (.A(II19820), .Z(g12756) ) ;
NAND2   gate7127  (.A(g3554), .B(g6980), .Z(g10705) ) ;
INV     gate7128  (.A(g10705), .Z(II19823) ) ;
INV     gate7129  (.A(II19823), .Z(g12759) ) ;
NAND2   gate7130  (.A(g7802), .B(g3678), .Z(g10252) ) ;
INV     gate7131  (.A(g10252), .Z(II19826) ) ;
INV     gate7132  (.A(II19826), .Z(g12762) ) ;
INV     gate7133  (.A(g10631), .Z(II19829) ) ;
INV     gate7134  (.A(II19829), .Z(g12765) ) ;
INV     gate7135  (.A(g8829), .Z(g12768) ) ;
INV     gate7136  (.A(g8726), .Z(II19833) ) ;
INV     gate7137  (.A(II19833), .Z(g12769) ) ;
INV     gate7138  (.A(g8726), .Z(II19836) ) ;
INV     gate7139  (.A(II19836), .Z(g12772) ) ;
INV     gate7140  (.A(g8832), .Z(g12775) ) ;
INV     gate7141  (.A(g10766), .Z(g12776) ) ;
INV     gate7142  (.A(g8836), .Z(g12782) ) ;
NAND2   gate7143  (.A(g3398), .B(g3366), .Z(g8533) ) ;
INV     gate7144  (.A(g8533), .Z(II19844) ) ;
INV     gate7145  (.A(II19844), .Z(g12783) ) ;
NAND2   gate7146  (.A(g3398), .B(g6912), .Z(g10677) ) ;
INV     gate7147  (.A(g10677), .Z(II19847) ) ;
INV     gate7148  (.A(II19847), .Z(g12786) ) ;
INV     gate7149  (.A(g8847), .Z(g12790) ) ;
NAND2   gate7150  (.A(g3554), .B(g7162), .Z(g10679) ) ;
INV     gate7151  (.A(g10679), .Z(II19852) ) ;
INV     gate7152  (.A(II19852), .Z(g12791) ) ;
NAND2   gate7153  (.A(g3554), .B(g6980), .Z(g10723) ) ;
INV     gate7154  (.A(g10723), .Z(II19855) ) ;
INV     gate7155  (.A(II19855), .Z(g12794) ) ;
INV     gate7156  (.A(g10617), .Z(II19859) ) ;
INV     gate7157  (.A(II19859), .Z(g12798) ) ;
NAND2   gate7158  (.A(g3710), .B(g7230), .Z(g10725) ) ;
INV     gate7159  (.A(g10725), .Z(II19862) ) ;
INV     gate7160  (.A(II19862), .Z(g12801) ) ;
NAND2   gate7161  (.A(g7815), .B(g3834), .Z(g10354) ) ;
INV     gate7162  (.A(g10354), .Z(II19865) ) ;
INV     gate7163  (.A(II19865), .Z(g12804) ) ;
INV     gate7164  (.A(g8853), .Z(g12807) ) ;
INV     gate7165  (.A(g8726), .Z(II19869) ) ;
INV     gate7166  (.A(II19869), .Z(g12808) ) ;
INV     gate7167  (.A(g8317), .Z(II19872) ) ;
INV     gate7168  (.A(II19872), .Z(g12811) ) ;
INV     gate7169  (.A(g8856), .Z(g12815) ) ;
NAND2   gate7170  (.A(g3398), .B(g3366), .Z(g8547) ) ;
INV     gate7171  (.A(g8547), .Z(II19877) ) ;
INV     gate7172  (.A(II19877), .Z(g12816) ) ;
INV     gate7173  (.A(g8863), .Z(g12821) ) ;
NAND2   gate7174  (.A(g3554), .B(g3522), .Z(g8550) ) ;
INV     gate7175  (.A(g8550), .Z(II19883) ) ;
INV     gate7176  (.A(II19883), .Z(g12822) ) ;
NAND2   gate7177  (.A(g3554), .B(g7162), .Z(g10706) ) ;
INV     gate7178  (.A(g10706), .Z(II19886) ) ;
INV     gate7179  (.A(II19886), .Z(g12825) ) ;
INV     gate7180  (.A(g8874), .Z(g12829) ) ;
NAND2   gate7181  (.A(g3710), .B(g7358), .Z(g10708) ) ;
INV     gate7182  (.A(g10708), .Z(II19891) ) ;
INV     gate7183  (.A(II19891), .Z(g12830) ) ;
NAND2   gate7184  (.A(g3710), .B(g7230), .Z(g10744) ) ;
INV     gate7185  (.A(g10744), .Z(II19894) ) ;
INV     gate7186  (.A(II19894), .Z(g12833) ) ;
INV     gate7187  (.A(g10664), .Z(II19898) ) ;
INV     gate7188  (.A(II19898), .Z(g12837) ) ;
NAND2   gate7189  (.A(g3866), .B(g7426), .Z(g10746) ) ;
INV     gate7190  (.A(g10746), .Z(II19901) ) ;
INV     gate7191  (.A(II19901), .Z(g12840) ) ;
INV     gate7192  (.A(g8879), .Z(g12843) ) ;
INV     gate7193  (.A(g8726), .Z(II19905) ) ;
INV     gate7194  (.A(II19905), .Z(g12844) ) ;
INV     gate7195  (.A(g8882), .Z(g12847) ) ;
INV     gate7196  (.A(g11059), .Z(g12848) ) ;
INV     gate7197  (.A(g8885), .Z(g12850) ) ;
INV     gate7198  (.A(g8888), .Z(g12851) ) ;
INV     gate7199  (.A(g8894), .Z(g12853) ) ;
NAND2   gate7200  (.A(g3554), .B(g3522), .Z(g8560) ) ;
INV     gate7201  (.A(g8560), .Z(II19915) ) ;
INV     gate7202  (.A(II19915), .Z(g12854) ) ;
INV     gate7203  (.A(g8901), .Z(g12859) ) ;
NAND2   gate7204  (.A(g3710), .B(g3678), .Z(g8563) ) ;
INV     gate7205  (.A(g8563), .Z(II19921) ) ;
INV     gate7206  (.A(II19921), .Z(g12860) ) ;
NAND2   gate7207  (.A(g3710), .B(g7358), .Z(g10726) ) ;
INV     gate7208  (.A(g10726), .Z(II19924) ) ;
INV     gate7209  (.A(II19924), .Z(g12863) ) ;
INV     gate7210  (.A(g8912), .Z(g12867) ) ;
NAND2   gate7211  (.A(g3866), .B(g7488), .Z(g10728) ) ;
INV     gate7212  (.A(g10728), .Z(II19929) ) ;
INV     gate7213  (.A(II19929), .Z(g12868) ) ;
NAND2   gate7214  (.A(g3866), .B(g7426), .Z(g10763) ) ;
INV     gate7215  (.A(g10763), .Z(II19932) ) ;
INV     gate7216  (.A(II19932), .Z(g12871) ) ;
INV     gate7217  (.A(g8915), .Z(g12874) ) ;
INV     gate7218  (.A(g10779), .Z(g12875) ) ;
INV     gate7219  (.A(g8918), .Z(g12881) ) ;
INV     gate7220  (.A(g8921), .Z(g12882) ) ;
INV     gate7221  (.A(g8925), .Z(g12891) ) ;
INV     gate7222  (.A(g8928), .Z(g12892) ) ;
INV     gate7223  (.A(g8934), .Z(g12894) ) ;
NAND2   gate7224  (.A(g3710), .B(g3678), .Z(g8571) ) ;
INV     gate7225  (.A(g8571), .Z(II19952) ) ;
INV     gate7226  (.A(II19952), .Z(g12895) ) ;
INV     gate7227  (.A(g8941), .Z(g12900) ) ;
NAND2   gate7228  (.A(g3866), .B(g3834), .Z(g8574) ) ;
INV     gate7229  (.A(g8574), .Z(II19958) ) ;
INV     gate7230  (.A(II19958), .Z(g12901) ) ;
NAND2   gate7231  (.A(g3866), .B(g7488), .Z(g10747) ) ;
INV     gate7232  (.A(g10747), .Z(II19961) ) ;
INV     gate7233  (.A(II19961), .Z(g12904) ) ;
INV     gate7234  (.A(g8949), .Z(g12907) ) ;
INV     gate7235  (.A(g10904), .Z(g12909) ) ;
INV     gate7236  (.A(g8952), .Z(g12914) ) ;
INV     gate7237  (.A(g8955), .Z(g12915) ) ;
INV     gate7238  (.A(g8958), .Z(g12921) ) ;
INV     gate7239  (.A(g8961), .Z(g12922) ) ;
INV     gate7240  (.A(g8965), .Z(g12931) ) ;
INV     gate7241  (.A(g8968), .Z(g12932) ) ;
INV     gate7242  (.A(g8974), .Z(g12934) ) ;
NAND2   gate7243  (.A(g3866), .B(g3834), .Z(g8577) ) ;
INV     gate7244  (.A(g8577), .Z(II19986) ) ;
INV     gate7245  (.A(II19986), .Z(g12935) ) ;
INV     gate7246  (.A(g8980), .Z(g12940) ) ;
INV     gate7247  (.A(g8984), .Z(g12943) ) ;
INV     gate7248  (.A(g8987), .Z(g12944) ) ;
INV     gate7249  (.A(g8990), .Z(g12950) ) ;
INV     gate7250  (.A(g8993), .Z(g12951) ) ;
INV     gate7251  (.A(g8997), .Z(g12960) ) ;
INV     gate7252  (.A(g9000), .Z(g12961) ) ;
INV     gate7253  (.A(g8313), .Z(II20009) ) ;
INV     gate7254  (.A(II20009), .Z(g12962) ) ;
INV     gate7255  (.A(g9006), .Z(g12965) ) ;
INV     gate7256  (.A(g9010), .Z(g12969) ) ;
INV     gate7257  (.A(g9013), .Z(g12972) ) ;
INV     gate7258  (.A(g9016), .Z(g12973) ) ;
INV     gate7259  (.A(g9019), .Z(g12979) ) ;
INV     gate7260  (.A(g9022), .Z(g12980) ) ;
INV     gate7261  (.A(g9035), .Z(g12993) ) ;
INV     gate7262  (.A(g9038), .Z(g12996) ) ;
INV     gate7263  (.A(g9041), .Z(g12997) ) ;
INV     gate7264  (.A(g9044), .Z(g12998) ) ;
INV     gate7265  (.A(g9058), .Z(g13003) ) ;
AND3    gate7266  (.A(g7466), .B(g7342), .C(II17429), .Z(g10480) ) ;
INV     gate7267  (.A(g10480), .Z(II20062) ) ;
INV     gate7268  (.A(II20062), .Z(g13011) ) ;
INV     gate7269  (.A(g10810), .Z(g13025) ) ;
INV     gate7270  (.A(g10797), .Z(g13033) ) ;
INV     gate7271  (.A(g10831), .Z(g13036) ) ;
INV     gate7272  (.A(g10789), .Z(g13043) ) ;
INV     gate7273  (.A(g10814), .Z(g13046) ) ;
INV     gate7274  (.A(g10851), .Z(g13049) ) ;
INV     gate7275  (.A(g10784), .Z(g13057) ) ;
INV     gate7276  (.A(g10801), .Z(g13060) ) ;
INV     gate7277  (.A(g10835), .Z(g13063) ) ;
INV     gate7278  (.A(g10872), .Z(g13066) ) ;
INV     gate7279  (.A(g10876), .Z(II20117) ) ;
INV     gate7280  (.A(II20117), .Z(g13070) ) ;
INV     gate7281  (.A(g10793), .Z(g13073) ) ;
INV     gate7282  (.A(g10818), .Z(g13076) ) ;
INV     gate7283  (.A(g10855), .Z(g13079) ) ;
INV     gate7284  (.A(g10805), .Z(g13092) ) ;
INV     gate7285  (.A(g10839), .Z(g13095) ) ;
INV     gate7286  (.A(g9128), .Z(g13101) ) ;
INV     gate7287  (.A(g10822), .Z(g13107) ) ;
INV     gate7288  (.A(g9134), .Z(g13117) ) ;
INV     gate7289  (.A(g9140), .Z(g13130) ) ;
INV     gate7290  (.A(g9146), .Z(g13141) ) ;
INV     gate7291  (.A(g9170), .Z(g13148) ) ;
INV     gate7292  (.A(g9184), .Z(g13151) ) ;
INV     gate7293  (.A(g9196), .Z(g13152) ) ;
INV     gate7294  (.A(g9199), .Z(g13153) ) ;
INV     gate7295  (.A(g9212), .Z(g13154) ) ;
INV     gate7296  (.A(g9229), .Z(g13157) ) ;
INV     gate7297  (.A(g9242), .Z(g13158) ) ;
INV     gate7298  (.A(g9245), .Z(g13159) ) ;
INV     gate7299  (.A(g9257), .Z(g13161) ) ;
INV     gate7300  (.A(g9260), .Z(g13162) ) ;
INV     gate7301  (.A(g9273), .Z(g13163) ) ;
INV     gate7302  (.A(g9290), .Z(g13166) ) ;
INV     gate7303  (.A(g9303), .Z(g13167) ) ;
INV     gate7304  (.A(g9306), .Z(g13168) ) ;
INV     gate7305  (.A(g9320), .Z(g13169) ) ;
INV     gate7306  (.A(g9323), .Z(g13170) ) ;
INV     gate7307  (.A(g9335), .Z(g13172) ) ;
INV     gate7308  (.A(g9338), .Z(g13173) ) ;
INV     gate7309  (.A(g9351), .Z(g13174) ) ;
INV     gate7310  (.A(g9368), .Z(g13176) ) ;
INV     gate7311  (.A(g9371), .Z(g13177) ) ;
INV     gate7312  (.A(g9384), .Z(g13178) ) ;
INV     gate7313  (.A(g9387), .Z(g13179) ) ;
INV     gate7314  (.A(g9401), .Z(g13180) ) ;
INV     gate7315  (.A(g9404), .Z(g13181) ) ;
INV     gate7316  (.A(g9416), .Z(g13183) ) ;
INV     gate7317  (.A(g9419), .Z(g13184) ) ;
INV     gate7318  (.A(g9443), .Z(g13185) ) ;
INV     gate7319  (.A(g9446), .Z(g13186) ) ;
INV     gate7320  (.A(g9450), .Z(g13187) ) ;
INV     gate7321  (.A(g9465), .Z(g13188) ) ;
INV     gate7322  (.A(g9468), .Z(g13189) ) ;
INV     gate7323  (.A(g9481), .Z(g13190) ) ;
INV     gate7324  (.A(g9484), .Z(g13191) ) ;
INV     gate7325  (.A(g9498), .Z(g13192) ) ;
INV     gate7326  (.A(g9501), .Z(g13193) ) ;
INV     gate7327  (.A(g9524), .Z(g13195) ) ;
INV     gate7328  (.A(g9528), .Z(g13196) ) ;
INV     gate7329  (.A(g9531), .Z(g13197) ) ;
INV     gate7330  (.A(g9585), .Z(g13198) ) ;
INV     gate7331  (.A(g9588), .Z(g13199) ) ;
INV     gate7332  (.A(g9592), .Z(g13200) ) ;
INV     gate7333  (.A(g9607), .Z(g13201) ) ;
INV     gate7334  (.A(g9610), .Z(g13202) ) ;
INV     gate7335  (.A(g9623), .Z(g13203) ) ;
INV     gate7336  (.A(g9626), .Z(g13204) ) ;
INV     gate7337  (.A(g9641), .Z(g13205) ) ;
INV     gate7338  (.A(g9644), .Z(g13206) ) ;
INV     gate7339  (.A(g9666), .Z(g13207) ) ;
INV     gate7340  (.A(g9670), .Z(g13208) ) ;
INV     gate7341  (.A(g9673), .Z(g13209) ) ;
INV     gate7342  (.A(g9727), .Z(g13210) ) ;
INV     gate7343  (.A(g9730), .Z(g13211) ) ;
INV     gate7344  (.A(g9734), .Z(g13212) ) ;
INV     gate7345  (.A(g9749), .Z(g13213) ) ;
INV     gate7346  (.A(g9752), .Z(g13214) ) ;
INV     gate7347  (.A(g9027), .Z(II20264) ) ;
INV     gate7348  (.A(II20264), .Z(g13215) ) ;
INV     gate7349  (.A(g9767), .Z(g13218) ) ;
INV     gate7350  (.A(g9770), .Z(g13219) ) ;
INV     gate7351  (.A(g9787), .Z(g13220) ) ;
INV     gate7352  (.A(g9790), .Z(g13221) ) ;
INV     gate7353  (.A(g9812), .Z(g13222) ) ;
INV     gate7354  (.A(g9816), .Z(g13223) ) ;
INV     gate7355  (.A(g9819), .Z(g13224) ) ;
INV     gate7356  (.A(g9873), .Z(g13225) ) ;
INV     gate7357  (.A(g9876), .Z(g13226) ) ;
INV     gate7358  (.A(g9880), .Z(g13227) ) ;
INV     gate7359  (.A(g9027), .Z(II20278) ) ;
INV     gate7360  (.A(II20278), .Z(g13229) ) ;
INV     gate7361  (.A(g9895), .Z(g13232) ) ;
INV     gate7362  (.A(g9898), .Z(g13233) ) ;
INV     gate7363  (.A(g9050), .Z(II20283) ) ;
INV     gate7364  (.A(II20283), .Z(g13234) ) ;
INV     gate7365  (.A(g9913), .Z(g13237) ) ;
INV     gate7366  (.A(g9916), .Z(g13238) ) ;
INV     gate7367  (.A(g9933), .Z(g13239) ) ;
INV     gate7368  (.A(g9936), .Z(g13240) ) ;
INV     gate7369  (.A(g9958), .Z(g13241) ) ;
INV     gate7370  (.A(g9962), .Z(g13242) ) ;
INV     gate7371  (.A(g9965), .Z(g13243) ) ;
INV     gate7372  (.A(g10004), .Z(g13244) ) ;
INV     gate7373  (.A(g10015), .Z(II20295) ) ;
INV     gate7374  (.A(II20295), .Z(g13246) ) ;
INV     gate7375  (.A(g10800), .Z(II20299) ) ;
INV     gate7376  (.A(II20299), .Z(g13248) ) ;
INV     gate7377  (.A(g10018), .Z(g13249) ) ;
INV     gate7378  (.A(g10021), .Z(g13250) ) ;
INV     gate7379  (.A(g9050), .Z(II20305) ) ;
INV     gate7380  (.A(II20305), .Z(g13252) ) ;
INV     gate7381  (.A(g10049), .Z(g13255) ) ;
INV     gate7382  (.A(g10052), .Z(g13256) ) ;
INV     gate7383  (.A(g9067), .Z(II20310) ) ;
INV     gate7384  (.A(II20310), .Z(g13257) ) ;
INV     gate7385  (.A(g10067), .Z(g13260) ) ;
INV     gate7386  (.A(g10070), .Z(g13261) ) ;
INV     gate7387  (.A(g10087), .Z(g13262) ) ;
INV     gate7388  (.A(g10090), .Z(g13263) ) ;
INV     gate7389  (.A(g10096), .Z(g13264) ) ;
INV     gate7390  (.A(g8568), .Z(g13265) ) ;
INV     gate7391  (.A(g10792), .Z(II20320) ) ;
INV     gate7392  (.A(II20320), .Z(g13267) ) ;
INV     gate7393  (.A(g10109), .Z(g13268) ) ;
INV     gate7394  (.A(g10124), .Z(II20324) ) ;
INV     gate7395  (.A(II20324), .Z(g13269) ) ;
INV     gate7396  (.A(g10817), .Z(II20328) ) ;
INV     gate7397  (.A(II20328), .Z(g13271) ) ;
INV     gate7398  (.A(g10127), .Z(g13272) ) ;
INV     gate7399  (.A(g10130), .Z(g13273) ) ;
INV     gate7400  (.A(g9067), .Z(II20334) ) ;
INV     gate7401  (.A(II20334), .Z(g13275) ) ;
INV     gate7402  (.A(g10158), .Z(g13278) ) ;
INV     gate7403  (.A(g10161), .Z(g13279) ) ;
INV     gate7404  (.A(g9084), .Z(II20339) ) ;
INV     gate7405  (.A(II20339), .Z(g13280) ) ;
INV     gate7406  (.A(g10176), .Z(g13283) ) ;
INV     gate7407  (.A(g10179), .Z(g13284) ) ;
INV     gate7408  (.A(g10189), .Z(g13285) ) ;
INV     gate7409  (.A(g10787), .Z(II20347) ) ;
INV     gate7410  (.A(II20347), .Z(g13290) ) ;
INV     gate7411  (.A(g10804), .Z(II20351) ) ;
INV     gate7412  (.A(II20351), .Z(g13292) ) ;
INV     gate7413  (.A(g10214), .Z(g13293) ) ;
INV     gate7414  (.A(g10229), .Z(II20355) ) ;
INV     gate7415  (.A(II20355), .Z(g13294) ) ;
INV     gate7416  (.A(g10838), .Z(II20359) ) ;
INV     gate7417  (.A(II20359), .Z(g13296) ) ;
INV     gate7418  (.A(g10232), .Z(g13297) ) ;
INV     gate7419  (.A(g10235), .Z(g13298) ) ;
INV     gate7420  (.A(g9084), .Z(II20365) ) ;
INV     gate7421  (.A(II20365), .Z(g13300) ) ;
INV     gate7422  (.A(g10263), .Z(g13303) ) ;
INV     gate7423  (.A(g10266), .Z(g13304) ) ;
INV     gate7424  (.A(g10273), .Z(g13308) ) ;
INV     gate7425  (.A(g10276), .Z(g13309) ) ;
INV     gate7426  (.A(g8569), .Z(II20376) ) ;
INV     gate7427  (.A(II20376), .Z(g13317) ) ;
INV     gate7428  (.A(g11213), .Z(II20379) ) ;
INV     gate7429  (.A(II20379), .Z(g13318) ) ;
INV     gate7430  (.A(g10907), .Z(II20382) ) ;
INV     gate7431  (.A(II20382), .Z(g13319) ) ;
INV     gate7432  (.A(g10796), .Z(II20386) ) ;
INV     gate7433  (.A(II20386), .Z(g13321) ) ;
INV     gate7434  (.A(g10821), .Z(II20390) ) ;
INV     gate7435  (.A(II20390), .Z(g13323) ) ;
INV     gate7436  (.A(g10316), .Z(g13324) ) ;
INV     gate7437  (.A(g10331), .Z(II20394) ) ;
INV     gate7438  (.A(II20394), .Z(g13325) ) ;
INV     gate7439  (.A(g10858), .Z(II20398) ) ;
INV     gate7440  (.A(II20398), .Z(g13327) ) ;
INV     gate7441  (.A(g10334), .Z(g13328) ) ;
INV     gate7442  (.A(g10337), .Z(g13329) ) ;
INV     gate7443  (.A(g10357), .Z(g13330) ) ;
INV     gate7444  (.A(g9027), .Z(II20407) ) ;
INV     gate7445  (.A(II20407), .Z(g13336) ) ;
INV     gate7446  (.A(g10887), .Z(II20410) ) ;
INV     gate7447  (.A(II20410), .Z(g13339) ) ;
INV     gate7448  (.A(g8575), .Z(II20414) ) ;
INV     gate7449  (.A(II20414), .Z(g13341) ) ;
INV     gate7450  (.A(g10933), .Z(II20417) ) ;
INV     gate7451  (.A(II20417), .Z(g13342) ) ;
INV     gate7452  (.A(g10808), .Z(II20421) ) ;
INV     gate7453  (.A(II20421), .Z(g13344) ) ;
INV     gate7454  (.A(g10842), .Z(II20425) ) ;
INV     gate7455  (.A(II20425), .Z(g13346) ) ;
INV     gate7456  (.A(g10409), .Z(g13347) ) ;
INV     gate7457  (.A(g10416), .Z(g13351) ) ;
INV     gate7458  (.A(g10419), .Z(g13352) ) ;
INV     gate7459  (.A(g9027), .Z(II20441) ) ;
INV     gate7460  (.A(II20441), .Z(g13356) ) ;
INV     gate7461  (.A(g10869), .Z(II20444) ) ;
INV     gate7462  (.A(II20444), .Z(g13359) ) ;
INV     gate7463  (.A(g9050), .Z(II20448) ) ;
INV     gate7464  (.A(II20448), .Z(g13361) ) ;
INV     gate7465  (.A(g10908), .Z(II20451) ) ;
INV     gate7466  (.A(II20451), .Z(g13364) ) ;
INV     gate7467  (.A(g8578), .Z(II20455) ) ;
INV     gate7468  (.A(II20455), .Z(g13366) ) ;
INV     gate7469  (.A(g10972), .Z(II20458) ) ;
INV     gate7470  (.A(II20458), .Z(g13367) ) ;
INV     gate7471  (.A(g10825), .Z(II20462) ) ;
INV     gate7472  (.A(II20462), .Z(g13369) ) ;
INV     gate7473  (.A(g10482), .Z(g13373) ) ;
INV     gate7474  (.A(g9027), .Z(II20476) ) ;
INV     gate7475  (.A(II20476), .Z(g13381) ) ;
INV     gate7476  (.A(g10849), .Z(II20479) ) ;
INV     gate7477  (.A(II20479), .Z(g13384) ) ;
INV     gate7478  (.A(g9050), .Z(II20483) ) ;
INV     gate7479  (.A(II20483), .Z(g13386) ) ;
INV     gate7480  (.A(g10889), .Z(II20486) ) ;
INV     gate7481  (.A(II20486), .Z(g13389) ) ;
INV     gate7482  (.A(g9067), .Z(II20490) ) ;
INV     gate7483  (.A(II20490), .Z(g13391) ) ;
INV     gate7484  (.A(g10934), .Z(II20493) ) ;
INV     gate7485  (.A(II20493), .Z(g13394) ) ;
INV     gate7486  (.A(g8579), .Z(II20497) ) ;
INV     gate7487  (.A(II20497), .Z(g13396) ) ;
INV     gate7488  (.A(g11007), .Z(II20500) ) ;
INV     gate7489  (.A(II20500), .Z(g13397) ) ;
INV     gate7490  (.A(g10542), .Z(g13398) ) ;
INV     gate7491  (.A(g10545), .Z(g13400) ) ;
INV     gate7492  (.A(g11769), .Z(II20514) ) ;
INV     gate7493  (.A(g12425), .Z(II20517) ) ;
INV     gate7494  (.A(g13246), .Z(II20520) ) ;
INV     gate7495  (.A(g13317), .Z(II20523) ) ;
INV     gate7496  (.A(g12519), .Z(II20526) ) ;
INV     gate7497  (.A(g13319), .Z(II20529) ) ;
INV     gate7498  (.A(g13339), .Z(II20532) ) ;
INV     gate7499  (.A(g13359), .Z(II20535) ) ;
INV     gate7500  (.A(g13384), .Z(II20538) ) ;
INV     gate7501  (.A(g11599), .Z(II20541) ) ;
INV     gate7502  (.A(g11628), .Z(II20544) ) ;
INV     gate7503  (.A(g13248), .Z(II20547) ) ;
INV     gate7504  (.A(g13267), .Z(II20550) ) ;
INV     gate7505  (.A(g13290), .Z(II20553) ) ;
INV     gate7506  (.A(g12435), .Z(II20556) ) ;
INV     gate7507  (.A(g11937), .Z(II20559) ) ;
INV     gate7508  (.A(g11786), .Z(II20562) ) ;
INV     gate7509  (.A(g12432), .Z(II20565) ) ;
INV     gate7510  (.A(g13269), .Z(II20568) ) ;
INV     gate7511  (.A(g13341), .Z(II20571) ) ;
INV     gate7512  (.A(g12534), .Z(II20574) ) ;
INV     gate7513  (.A(g13342), .Z(II20577) ) ;
INV     gate7514  (.A(g13364), .Z(II20580) ) ;
INV     gate7515  (.A(g13389), .Z(II20583) ) ;
INV     gate7516  (.A(g11606), .Z(II20586) ) ;
INV     gate7517  (.A(g11629), .Z(II20589) ) ;
INV     gate7518  (.A(g11651), .Z(II20592) ) ;
INV     gate7519  (.A(g13271), .Z(II20595) ) ;
INV     gate7520  (.A(g13292), .Z(II20598) ) ;
INV     gate7521  (.A(g13321), .Z(II20601) ) ;
INV     gate7522  (.A(g12440), .Z(II20604) ) ;
INV     gate7523  (.A(g11990), .Z(II20607) ) ;
INV     gate7524  (.A(g11812), .Z(II20610) ) ;
INV     gate7525  (.A(g12437), .Z(II20613) ) ;
INV     gate7526  (.A(g13294), .Z(II20616) ) ;
INV     gate7527  (.A(g13366), .Z(II20619) ) ;
INV     gate7528  (.A(g12543), .Z(II20622) ) ;
INV     gate7529  (.A(g13367), .Z(II20625) ) ;
INV     gate7530  (.A(g13394), .Z(II20628) ) ;
INV     gate7531  (.A(g11611), .Z(II20631) ) ;
INV     gate7532  (.A(g11636), .Z(II20634) ) ;
INV     gate7533  (.A(g11652), .Z(II20637) ) ;
INV     gate7534  (.A(g11670), .Z(II20640) ) ;
INV     gate7535  (.A(g13296), .Z(II20643) ) ;
INV     gate7536  (.A(g13323), .Z(II20646) ) ;
INV     gate7537  (.A(g13344), .Z(II20649) ) ;
INV     gate7538  (.A(g12445), .Z(II20652) ) ;
INV     gate7539  (.A(g12059), .Z(II20655) ) ;
INV     gate7540  (.A(g11845), .Z(II20658) ) ;
INV     gate7541  (.A(g12442), .Z(II20661) ) ;
INV     gate7542  (.A(g13325), .Z(II20664) ) ;
INV     gate7543  (.A(g13396), .Z(II20667) ) ;
INV     gate7544  (.A(g12552), .Z(II20670) ) ;
INV     gate7545  (.A(g13397), .Z(II20673) ) ;
INV     gate7546  (.A(g11616), .Z(II20676) ) ;
INV     gate7547  (.A(g11641), .Z(II20679) ) ;
INV     gate7548  (.A(g11659), .Z(II20682) ) ;
INV     gate7549  (.A(g11671), .Z(II20685) ) ;
INV     gate7550  (.A(g11682), .Z(II20688) ) ;
INV     gate7551  (.A(g13327), .Z(II20691) ) ;
INV     gate7552  (.A(g13346), .Z(II20694) ) ;
INV     gate7553  (.A(g13369), .Z(II20697) ) ;
INV     gate7554  (.A(g12450), .Z(II20700) ) ;
INV     gate7555  (.A(g12123), .Z(II20703) ) ;
INV     gate7556  (.A(g11490), .Z(II20706) ) ;
INV     gate7557  (.A(II20706), .Z(g13469) ) ;
INV     gate7558  (.A(g13070), .Z(II20709) ) ;
NOR3    gate7559  (.A(g8841), .B(g8861), .C(g8892), .Z(g13228) ) ;
INV     gate7560  (.A(g13228), .Z(g13519) ) ;
NOR3    gate7561  (.A(g8868), .B(g8899), .C(g8932), .Z(g13251) ) ;
INV     gate7562  (.A(g13251), .Z(g13530) ) ;
NOR3    gate7563  (.A(g8906), .B(g8939), .C(g8972), .Z(g13274) ) ;
INV     gate7564  (.A(g13274), .Z(g13541) ) ;
NOR3    gate7565  (.A(g8946), .B(g8979), .C(g9004), .Z(g13299) ) ;
INV     gate7566  (.A(g13299), .Z(g13552) ) ;
NOR3    gate7567  (.A(g10423), .B(g10485), .C(g10548), .Z(g12192) ) ;
INV     gate7568  (.A(g12192), .Z(g13565) ) ;
NOR3    gate7569  (.A(g9063), .B(g9077), .C(g9093), .Z(g11627) ) ;
INV     gate7570  (.A(g11627), .Z(g13568) ) ;
NOR3    gate7571  (.A(g8676), .B(g8687), .C(g8703), .Z(g13149) ) ;
INV     gate7572  (.A(g13149), .Z(II20791) ) ;
INV     gate7573  (.A(II20791), .Z(g13571) ) ;
NOR3    gate7574  (.A(g8601), .B(g8612), .C(g8621), .Z(g13111) ) ;
INV     gate7575  (.A(g13111), .Z(II20794) ) ;
INV     gate7576  (.A(II20794), .Z(g13572) ) ;
NOR3    gate7577  (.A(g10499), .B(g10559), .C(g10605), .Z(g12247) ) ;
INV     gate7578  (.A(g12247), .Z(g13573) ) ;
NOR3    gate7579  (.A(g9080), .B(g9096), .C(g9105), .Z(g11650) ) ;
INV     gate7580  (.A(g11650), .Z(g13576) ) ;
NOR3    gate7581  (.A(g8688), .B(g8705), .C(g8722), .Z(g13155) ) ;
INV     gate7582  (.A(g13155), .Z(II20799) ) ;
INV     gate7583  (.A(II20799), .Z(g13579) ) ;
NOR3    gate7584  (.A(g8704), .B(g8717), .C(g8751), .Z(g13160) ) ;
INV     gate7585  (.A(g13160), .Z(II20802) ) ;
INV     gate7586  (.A(II20802), .Z(g13580) ) ;
NOR3    gate7587  (.A(g8613), .B(g8625), .C(g8631), .Z(g13124) ) ;
INV     gate7588  (.A(g13124), .Z(II20805) ) ;
INV     gate7589  (.A(II20805), .Z(g13581) ) ;
NOR3    gate7590  (.A(g10573), .B(g10616), .C(g10652), .Z(g12290) ) ;
INV     gate7591  (.A(g12290), .Z(g13582) ) ;
NOR3    gate7592  (.A(g9099), .B(g9108), .C(g9115), .Z(g11669) ) ;
INV     gate7593  (.A(g11669), .Z(g13585) ) ;
NOR3    gate7594  (.A(g8706), .B(g8724), .C(g8760), .Z(g13164) ) ;
INV     gate7595  (.A(g13164), .Z(II20810) ) ;
INV     gate7596  (.A(II20810), .Z(g13588) ) ;
INV     gate7597  (.A(g13265), .Z(II20813) ) ;
INV     gate7598  (.A(II20813), .Z(g13589) ) ;
NOR3    gate7599  (.A(g10108), .B(g10198), .C(g10283), .Z(g12487) ) ;
INV     gate7600  (.A(g12487), .Z(II20816) ) ;
INV     gate7601  (.A(II20816), .Z(g13598) ) ;
NOR3    gate7602  (.A(g8723), .B(g8755), .C(g8774), .Z(g13171) ) ;
INV     gate7603  (.A(g13171), .Z(II20820) ) ;
INV     gate7604  (.A(II20820), .Z(g13600) ) ;
NOR3    gate7605  (.A(g8626), .B(g8635), .C(g8650), .Z(g13135) ) ;
INV     gate7606  (.A(g13135), .Z(II20823) ) ;
INV     gate7607  (.A(II20823), .Z(g13601) ) ;
NOR3    gate7608  (.A(g10630), .B(g10663), .C(g10682), .Z(g12326) ) ;
INV     gate7609  (.A(g12326), .Z(g13602) ) ;
NOR3    gate7610  (.A(g9111), .B(g9118), .C(g9123), .Z(g11681) ) ;
INV     gate7611  (.A(g11681), .Z(g13605) ) ;
NOR3    gate7612  (.A(g8725), .B(g8762), .C(g8783), .Z(g13175) ) ;
INV     gate7613  (.A(g13175), .Z(II20828) ) ;
INV     gate7614  (.A(II20828), .Z(g13608) ) ;
NOR3    gate7615  (.A(g10213), .B(g10300), .C(g10376), .Z(g12507) ) ;
INV     gate7616  (.A(g12507), .Z(II20832) ) ;
INV     gate7617  (.A(II20832), .Z(g13610) ) ;
NOR3    gate7618  (.A(g8761), .B(g8778), .C(g8797), .Z(g13182) ) ;
INV     gate7619  (.A(g13182), .Z(II20836) ) ;
INV     gate7620  (.A(II20836), .Z(g13612) ) ;
NOR3    gate7621  (.A(g8636), .B(g8654), .C(g8666), .Z(g13143) ) ;
INV     gate7622  (.A(g13143), .Z(II20839) ) ;
INV     gate7623  (.A(II20839), .Z(g13613) ) ;
NOR3    gate7624  (.A(g9119), .B(g9124), .C(g9127), .Z(g11690) ) ;
INV     gate7625  (.A(g11690), .Z(g13614) ) ;
NOR3    gate7626  (.A(g10315), .B(g10393), .C(g10455), .Z(g12524) ) ;
INV     gate7627  (.A(g12524), .Z(II20844) ) ;
INV     gate7628  (.A(II20844), .Z(g13620) ) ;
NOR3    gate7629  (.A(g8784), .B(g8801), .C(g8816), .Z(g13194) ) ;
INV     gate7630  (.A(g13194), .Z(II20848) ) ;
INV     gate7631  (.A(II20848), .Z(g13622) ) ;
NOR3    gate7632  (.A(g9009), .B(g9033), .C(g9048), .Z(g12457) ) ;
INV     gate7633  (.A(g12457), .Z(II20852) ) ;
INV     gate7634  (.A(II20852), .Z(g13624) ) ;
NOR3    gate7635  (.A(g9125), .B(g9131), .C(g9133), .Z(g11697) ) ;
INV     gate7636  (.A(g11697), .Z(g13626) ) ;
NOR3    gate7637  (.A(g10408), .B(g10472), .C(g10531), .Z(g12539) ) ;
INV     gate7638  (.A(g12539), .Z(II20858) ) ;
INV     gate7639  (.A(II20858), .Z(g13632) ) ;
NOR3    gate7640  (.A(g9034), .B(g9056), .C(g9065), .Z(g12467) ) ;
INV     gate7641  (.A(g12467), .Z(II20863) ) ;
INV     gate7642  (.A(II20863), .Z(g13635) ) ;
NOR3    gate7643  (.A(g9132), .B(g9137), .C(g9139), .Z(g11703) ) ;
INV     gate7644  (.A(g11703), .Z(g13637) ) ;
INV     gate7645  (.A(g13215), .Z(g13644) ) ;
NOR3    gate7646  (.A(g9057), .B(g9073), .C(g9082), .Z(g12482) ) ;
INV     gate7647  (.A(g12482), .Z(II20873) ) ;
INV     gate7648  (.A(II20873), .Z(g13647) ) ;
NOR3    gate7649  (.A(g9138), .B(g9143), .C(g9145), .Z(g11711) ) ;
INV     gate7650  (.A(g11711), .Z(g13649) ) ;
INV     gate7651  (.A(g12452), .Z(g13657) ) ;
INV     gate7652  (.A(g13229), .Z(g13669) ) ;
INV     gate7653  (.A(g13234), .Z(g13670) ) ;
NOR3    gate7654  (.A(g9074), .B(g9090), .C(g9101), .Z(g12499) ) ;
INV     gate7655  (.A(g12499), .Z(II20886) ) ;
INV     gate7656  (.A(II20886), .Z(g13673) ) ;
INV     gate7657  (.A(g12447), .Z(g13677) ) ;
INV     gate7658  (.A(g12460), .Z(g13687) ) ;
INV     gate7659  (.A(g13252), .Z(g13699) ) ;
INV     gate7660  (.A(g13257), .Z(g13700) ) ;
INV     gate7661  (.A(g12443), .Z(g13706) ) ;
INV     gate7662  (.A(g12453), .Z(g13714) ) ;
INV     gate7663  (.A(g12470), .Z(g13724) ) ;
INV     gate7664  (.A(g13275), .Z(g13736) ) ;
INV     gate7665  (.A(g13280), .Z(g13737) ) ;
AND3    gate7666  (.A(g7471), .B(g7570), .C(II20100), .Z(g13055) ) ;
INV     gate7667  (.A(g13055), .Z(II20909) ) ;
INV     gate7668  (.A(II20909), .Z(g13741) ) ;
INV     gate7669  (.A(g12439), .Z(g13750) ) ;
INV     gate7670  (.A(g12448), .Z(g13756) ) ;
INV     gate7671  (.A(g12461), .Z(g13764) ) ;
INV     gate7672  (.A(g12485), .Z(g13774) ) ;
INV     gate7673  (.A(g13300), .Z(g13786) ) ;
INV     gate7674  (.A(g12444), .Z(g13791) ) ;
INV     gate7675  (.A(g12454), .Z(g13797) ) ;
INV     gate7676  (.A(g12471), .Z(g13805) ) ;
INV     gate7677  (.A(g13336), .Z(g13817) ) ;
INV     gate7678  (.A(g12449), .Z(g13819) ) ;
INV     gate7679  (.A(g12462), .Z(g13825) ) ;
INV     gate7680  (.A(g13356), .Z(g13836) ) ;
INV     gate7681  (.A(g13361), .Z(g13838) ) ;
INV     gate7682  (.A(g12455), .Z(g13840) ) ;
NOR3    gate7683  (.A(g9241), .B(g9301), .C(g9364), .Z(g11744) ) ;
INV     gate7684  (.A(g11744), .Z(g13848) ) ;
INV     gate7685  (.A(g13381), .Z(g13849) ) ;
INV     gate7686  (.A(g13386), .Z(g13850) ) ;
INV     gate7687  (.A(g13391), .Z(g13852) ) ;
NOR3    gate7688  (.A(g9302), .B(g9365), .C(g9438), .Z(g11759) ) ;
INV     gate7689  (.A(g11759), .Z(g13856) ) ;
NOR3    gate7690  (.A(g9319), .B(g9382), .C(g9461), .Z(g11760) ) ;
INV     gate7691  (.A(g11760), .Z(g13857) ) ;
INV     gate7692  (.A(g11603), .Z(g13858) ) ;
INV     gate7693  (.A(g11608), .Z(g13859) ) ;
INV     gate7694  (.A(g11613), .Z(g13861) ) ;
NAND2   gate7695  (.A(g10481), .B(g9144), .Z(g11713) ) ;
INV     gate7696  (.A(g11713), .Z(II20959) ) ;
INV     gate7697  (.A(II20959), .Z(g13863) ) ;
NOR3    gate7698  (.A(g9366), .B(g9439), .C(g9518), .Z(g11767) ) ;
INV     gate7699  (.A(g11767), .Z(g13864) ) ;
NOR3    gate7700  (.A(g9383), .B(g9462), .C(g9580), .Z(g11772) ) ;
INV     gate7701  (.A(g11772), .Z(g13866) ) ;
NOR3    gate7702  (.A(g9400), .B(g9479), .C(g9603), .Z(g11773) ) ;
INV     gate7703  (.A(g11773), .Z(g13867) ) ;
INV     gate7704  (.A(g11633), .Z(g13868) ) ;
INV     gate7705  (.A(g11638), .Z(g13869) ) ;
NOR3    gate7706  (.A(g9440), .B(g9519), .C(g9630), .Z(g11780) ) ;
INV     gate7707  (.A(g11780), .Z(g13872) ) ;
NOR3    gate7708  (.A(g11347), .B(g11420), .C(g8327), .Z(g12698) ) ;
INV     gate7709  (.A(g12698), .Z(g13873) ) ;
NOR3    gate7710  (.A(g9463), .B(g9581), .C(g9660), .Z(g11784) ) ;
INV     gate7711  (.A(g11784), .Z(g13879) ) ;
NOR3    gate7712  (.A(g9480), .B(g9604), .C(g9722), .Z(g11789) ) ;
INV     gate7713  (.A(g11789), .Z(g13881) ) ;
NOR3    gate7714  (.A(g9497), .B(g9621), .C(g9745), .Z(g11790) ) ;
INV     gate7715  (.A(g11790), .Z(g13882) ) ;
INV     gate7716  (.A(g11656), .Z(g13883) ) ;
NOR3    gate7717  (.A(g9520), .B(g9631), .C(g9759), .Z(g11799) ) ;
INV     gate7718  (.A(g11799), .Z(g13885) ) ;
NOR3    gate7719  (.A(g11421), .B(g8328), .C(g8385), .Z(g12747) ) ;
INV     gate7720  (.A(g12747), .Z(g13886) ) ;
NOR3    gate7721  (.A(g9582), .B(g9661), .C(g9776), .Z(g11806) ) ;
INV     gate7722  (.A(g11806), .Z(g13894) ) ;
NOR3    gate7723  (.A(g11431), .B(g8339), .C(g8394), .Z(g12755) ) ;
INV     gate7724  (.A(g12755), .Z(g13895) ) ;
NOR3    gate7725  (.A(g9605), .B(g9723), .C(g9806), .Z(g11810) ) ;
INV     gate7726  (.A(g11810), .Z(g13901) ) ;
NOR3    gate7727  (.A(g9622), .B(g9746), .C(g9868), .Z(g11815) ) ;
INV     gate7728  (.A(g11815), .Z(g13903) ) ;
NOR3    gate7729  (.A(g9632), .B(g9760), .C(g9888), .Z(g11822) ) ;
INV     gate7730  (.A(g11822), .Z(g13906) ) ;
NOR3    gate7731  (.A(g8329), .B(g8386), .C(g8431), .Z(g12781) ) ;
INV     gate7732  (.A(g12781), .Z(g13907) ) ;
NOR3    gate7733  (.A(g9647), .B(g9773), .C(g9901), .Z(g11830) ) ;
INV     gate7734  (.A(g11830), .Z(g13918) ) ;
NOR3    gate7735  (.A(g9648), .B(g9775), .C(g9904), .Z(g11831) ) ;
INV     gate7736  (.A(g11831), .Z(g13922) ) ;
NOR3    gate7737  (.A(g9662), .B(g9777), .C(g9905), .Z(g11832) ) ;
INV     gate7738  (.A(g11832), .Z(g13926) ) ;
NOR3    gate7739  (.A(g8340), .B(g8395), .C(g8437), .Z(g12789) ) ;
INV     gate7740  (.A(g12789), .Z(g13927) ) ;
NOR3    gate7741  (.A(g9724), .B(g9807), .C(g9922), .Z(g11839) ) ;
INV     gate7742  (.A(g11839), .Z(g13935) ) ;
NOR3    gate7743  (.A(g8350), .B(g8406), .C(g8446), .Z(g12797) ) ;
INV     gate7744  (.A(g12797), .Z(g13936) ) ;
NOR3    gate7745  (.A(g9747), .B(g9869), .C(g9952), .Z(g11843) ) ;
INV     gate7746  (.A(g11843), .Z(g13942) ) ;
NOR3    gate7747  (.A(g9761), .B(g9889), .C(g10009), .Z(g11855) ) ;
INV     gate7748  (.A(g11855), .Z(g13945) ) ;
NOR3    gate7749  (.A(g8387), .B(g8432), .C(g8463), .Z(g12814) ) ;
INV     gate7750  (.A(g12814), .Z(g13946) ) ;
NAND2   gate7751  (.A(g8278), .B(g5438), .Z(g12503) ) ;
INV     gate7752  (.A(g12503), .Z(II21012) ) ;
INV     gate7753  (.A(II21012), .Z(g13954) ) ;
NOR3    gate7754  (.A(g9774), .B(g9902), .C(g10035), .Z(g11863) ) ;
INV     gate7755  (.A(g11863), .Z(g13958) ) ;
NOR3    gate7756  (.A(g9778), .B(g9906), .C(g10042), .Z(g11864) ) ;
INV     gate7757  (.A(g11864), .Z(g13962) ) ;
NOR3    gate7758  (.A(g8396), .B(g8438), .C(g8466), .Z(g12820) ) ;
INV     gate7759  (.A(g12820), .Z(g13963) ) ;
NOR3    gate7760  (.A(g9793), .B(g9919), .C(g10055), .Z(g11872) ) ;
INV     gate7761  (.A(g11872), .Z(g13974) ) ;
NOR3    gate7762  (.A(g9794), .B(g9921), .C(g10058), .Z(g11873) ) ;
INV     gate7763  (.A(g11873), .Z(g13978) ) ;
NOR3    gate7764  (.A(g9808), .B(g9923), .C(g10059), .Z(g11874) ) ;
INV     gate7765  (.A(g11874), .Z(g13982) ) ;
NOR3    gate7766  (.A(g8407), .B(g8447), .C(g8472), .Z(g12828) ) ;
INV     gate7767  (.A(g12828), .Z(g13983) ) ;
NOR3    gate7768  (.A(g9870), .B(g9953), .C(g10076), .Z(g11881) ) ;
INV     gate7769  (.A(g11881), .Z(g13991) ) ;
NOR3    gate7770  (.A(g8417), .B(g8458), .C(g8481), .Z(g12836) ) ;
INV     gate7771  (.A(g12836), .Z(g13992) ) ;
NOR3    gate7772  (.A(g9887), .B(g10007), .C(g10101), .Z(g11889) ) ;
INV     gate7773  (.A(g11889), .Z(g13999) ) ;
NOR3    gate7774  (.A(g9890), .B(g10010), .C(g10103), .Z(g11890) ) ;
INV     gate7775  (.A(g11890), .Z(g14000) ) ;
NOR3    gate7776  (.A(g8433), .B(g8464), .C(g8485), .Z(g12849) ) ;
INV     gate7777  (.A(g12849), .Z(g14001) ) ;
NAND2   gate7778  (.A(g8278), .B(g6448), .Z(g12486) ) ;
INV     gate7779  (.A(g12486), .Z(II21037) ) ;
INV     gate7780  (.A(II21037), .Z(g14008) ) ;
NOR3    gate7781  (.A(g9903), .B(g10036), .C(g10112), .Z(g11896) ) ;
INV     gate7782  (.A(g11896), .Z(g14011) ) ;
NOR3    gate7783  (.A(g9907), .B(g10043), .C(g10118), .Z(g11897) ) ;
INV     gate7784  (.A(g11897), .Z(g14015) ) ;
NOR3    gate7785  (.A(g8439), .B(g8467), .C(g8488), .Z(g12852) ) ;
INV     gate7786  (.A(g12852), .Z(g14016) ) ;
NAND2   gate7787  (.A(g8287), .B(g5473), .Z(g12520) ) ;
INV     gate7788  (.A(g12520), .Z(II21045) ) ;
INV     gate7789  (.A(II21045), .Z(g14024) ) ;
NOR3    gate7790  (.A(g9920), .B(g10056), .C(g10144), .Z(g11905) ) ;
INV     gate7791  (.A(g11905), .Z(g14028) ) ;
NOR3    gate7792  (.A(g9924), .B(g10060), .C(g10151), .Z(g11906) ) ;
INV     gate7793  (.A(g11906), .Z(g14032) ) ;
NOR3    gate7794  (.A(g8448), .B(g8473), .C(g8491), .Z(g12858) ) ;
INV     gate7795  (.A(g12858), .Z(g14033) ) ;
NOR3    gate7796  (.A(g9939), .B(g10073), .C(g10164), .Z(g11914) ) ;
INV     gate7797  (.A(g11914), .Z(g14044) ) ;
NOR3    gate7798  (.A(g9940), .B(g10075), .C(g10167), .Z(g11915) ) ;
INV     gate7799  (.A(g11915), .Z(g14048) ) ;
NOR3    gate7800  (.A(g9954), .B(g10077), .C(g10168), .Z(g11916) ) ;
INV     gate7801  (.A(g11916), .Z(g14052) ) ;
NOR3    gate7802  (.A(g8459), .B(g8482), .C(g8497), .Z(g12866) ) ;
INV     gate7803  (.A(g12866), .Z(g14053) ) ;
NOR3    gate7804  (.A(g10008), .B(g10102), .C(g10192), .Z(g11928) ) ;
INV     gate7805  (.A(g11928), .Z(g14061) ) ;
NOR3    gate7806  (.A(g8465), .B(g8486), .C(g8502), .Z(g12880) ) ;
INV     gate7807  (.A(g12880), .Z(g14062) ) ;
NAND2   gate7808  (.A(g8278), .B(g3306), .Z(g13147) ) ;
INV     gate7809  (.A(g13147), .Z(II21064) ) ;
INV     gate7810  (.A(II21064), .Z(g14068) ) ;
NOR3    gate7811  (.A(g10011), .B(g10104), .C(g10193), .Z(g11934) ) ;
INV     gate7812  (.A(g11934), .Z(g14071) ) ;
NOR3    gate7813  (.A(g10014), .B(g10106), .C(g10196), .Z(g11935) ) ;
INV     gate7814  (.A(g11935), .Z(g14079) ) ;
NOR3    gate7815  (.A(g10037), .B(g10113), .C(g10201), .Z(g11938) ) ;
INV     gate7816  (.A(g11938), .Z(g14086) ) ;
NOR3    gate7817  (.A(g10041), .B(g10116), .C(g10206), .Z(g11939) ) ;
INV     gate7818  (.A(g11939), .Z(g14090) ) ;
NOR3    gate7819  (.A(g10044), .B(g10119), .C(g10208), .Z(g11940) ) ;
INV     gate7820  (.A(g11940), .Z(g14091) ) ;
NOR3    gate7821  (.A(g8468), .B(g8489), .C(g8505), .Z(g12890) ) ;
INV     gate7822  (.A(g12890), .Z(g14092) ) ;
NAND2   gate7823  (.A(g8287), .B(g6713), .Z(g12506) ) ;
INV     gate7824  (.A(g12506), .Z(II21075) ) ;
INV     gate7825  (.A(II21075), .Z(g14099) ) ;
NOR3    gate7826  (.A(g10057), .B(g10145), .C(g10217), .Z(g11946) ) ;
INV     gate7827  (.A(g11946), .Z(g14102) ) ;
NOR3    gate7828  (.A(g10061), .B(g10152), .C(g10223), .Z(g11947) ) ;
INV     gate7829  (.A(g11947), .Z(g14106) ) ;
NOR3    gate7830  (.A(g8474), .B(g8492), .C(g8508), .Z(g12893) ) ;
INV     gate7831  (.A(g12893), .Z(g14107) ) ;
NAND2   gate7832  (.A(g8296), .B(g5512), .Z(g12535) ) ;
INV     gate7833  (.A(g12535), .Z(II21083) ) ;
INV     gate7834  (.A(II21083), .Z(g14115) ) ;
NOR3    gate7835  (.A(g10074), .B(g10165), .C(g10249), .Z(g11955) ) ;
INV     gate7836  (.A(g11955), .Z(g14119) ) ;
NOR3    gate7837  (.A(g10078), .B(g10169), .C(g10256), .Z(g11956) ) ;
INV     gate7838  (.A(g11956), .Z(g14123) ) ;
NOR3    gate7839  (.A(g8483), .B(g8498), .C(g8511), .Z(g12899) ) ;
INV     gate7840  (.A(g12899), .Z(g14124) ) ;
NOR3    gate7841  (.A(g10093), .B(g10182), .C(g10269), .Z(g11964) ) ;
INV     gate7842  (.A(g11964), .Z(g14135) ) ;
NOR3    gate7843  (.A(g10094), .B(g10184), .C(g10272), .Z(g11965) ) ;
INV     gate7844  (.A(g11965), .Z(g14139) ) ;
INV     gate7845  (.A(g11749), .Z(II21096) ) ;
INV     gate7846  (.A(II21096), .Z(g14144) ) ;
NOR3    gate7847  (.A(g8484), .B(g8500), .C(g8515), .Z(g12912) ) ;
INV     gate7848  (.A(g12912), .Z(g14148) ) ;
NOR3    gate7849  (.A(g8487), .B(g8503), .C(g8518), .Z(g12913) ) ;
INV     gate7850  (.A(g12913), .Z(g14153) ) ;
NOR3    gate7851  (.A(g10105), .B(g10194), .C(g10279), .Z(g11974) ) ;
INV     gate7852  (.A(g11974), .Z(g14158) ) ;
NOR3    gate7853  (.A(g10107), .B(g10197), .C(g10282), .Z(g11975) ) ;
INV     gate7854  (.A(g11975), .Z(g14165) ) ;
NOR3    gate7855  (.A(g10114), .B(g10202), .C(g10288), .Z(g11979) ) ;
INV     gate7856  (.A(g11979), .Z(g14171) ) ;
NOR3    gate7857  (.A(g10115), .B(g10204), .C(g10291), .Z(g11980) ) ;
INV     gate7858  (.A(g11980), .Z(g14175) ) ;
NOR3    gate7859  (.A(g10117), .B(g10207), .C(g10294), .Z(g11981) ) ;
INV     gate7860  (.A(g11981), .Z(g14176) ) ;
NOR3    gate7861  (.A(g8490), .B(g8506), .C(g8521), .Z(g12920) ) ;
INV     gate7862  (.A(g12920), .Z(g14177) ) ;
NAND2   gate7863  (.A(g8287), .B(g3462), .Z(g13150) ) ;
INV     gate7864  (.A(g13150), .Z(II21108) ) ;
INV     gate7865  (.A(II21108), .Z(g14183) ) ;
NOR3    gate7866  (.A(g10120), .B(g10209), .C(g10295), .Z(g11987) ) ;
INV     gate7867  (.A(g11987), .Z(g14186) ) ;
NOR3    gate7868  (.A(g10123), .B(g10211), .C(g10298), .Z(g11988) ) ;
INV     gate7869  (.A(g11988), .Z(g14194) ) ;
NOR3    gate7870  (.A(g10146), .B(g10218), .C(g10303), .Z(g11991) ) ;
INV     gate7871  (.A(g11991), .Z(g14201) ) ;
NOR3    gate7872  (.A(g10150), .B(g10221), .C(g10308), .Z(g11992) ) ;
INV     gate7873  (.A(g11992), .Z(g14205) ) ;
NOR3    gate7874  (.A(g10153), .B(g10224), .C(g10310), .Z(g11993) ) ;
INV     gate7875  (.A(g11993), .Z(g14206) ) ;
NOR3    gate7876  (.A(g8493), .B(g8509), .C(g8524), .Z(g12930) ) ;
INV     gate7877  (.A(g12930), .Z(g14207) ) ;
NAND2   gate7878  (.A(g8296), .B(g7015), .Z(g12523) ) ;
INV     gate7879  (.A(g12523), .Z(II21119) ) ;
INV     gate7880  (.A(II21119), .Z(g14214) ) ;
NOR3    gate7881  (.A(g10166), .B(g10250), .C(g10319), .Z(g11999) ) ;
INV     gate7882  (.A(g11999), .Z(g14217) ) ;
NOR3    gate7883  (.A(g10170), .B(g10257), .C(g10325), .Z(g12000) ) ;
INV     gate7884  (.A(g12000), .Z(g14221) ) ;
NOR3    gate7885  (.A(g8499), .B(g8512), .C(g8527), .Z(g12933) ) ;
INV     gate7886  (.A(g12933), .Z(g14222) ) ;
NAND2   gate7887  (.A(g8305), .B(g5556), .Z(g12544) ) ;
INV     gate7888  (.A(g12544), .Z(II21127) ) ;
INV     gate7889  (.A(II21127), .Z(g14230) ) ;
NOR3    gate7890  (.A(g10183), .B(g10270), .C(g10351), .Z(g12008) ) ;
INV     gate7891  (.A(g12008), .Z(g14234) ) ;
NOR3    gate7892  (.A(g8501), .B(g8516), .C(g8531), .Z(g12939) ) ;
INV     gate7893  (.A(g12939), .Z(g14238) ) ;
NOR3    gate7894  (.A(g10195), .B(g10280), .C(g10360), .Z(g12026) ) ;
INV     gate7895  (.A(g12026), .Z(g14244) ) ;
NOR3    gate7896  (.A(g10200), .B(g10286), .C(g10365), .Z(g12034) ) ;
INV     gate7897  (.A(g12034), .Z(g14249) ) ;
NOR3    gate7898  (.A(g10203), .B(g10289), .C(g10367), .Z(g12035) ) ;
INV     gate7899  (.A(g12035), .Z(g14252) ) ;
NOR3    gate7900  (.A(g10205), .B(g10292), .C(g10370), .Z(g12036) ) ;
INV     gate7901  (.A(g12036), .Z(g14256) ) ;
INV     gate7902  (.A(g11749), .Z(II21137) ) ;
INV     gate7903  (.A(II21137), .Z(g14259) ) ;
NOR3    gate7904  (.A(g8504), .B(g8519), .C(g8534), .Z(g12941) ) ;
INV     gate7905  (.A(g12941), .Z(g14263) ) ;
NOR3    gate7906  (.A(g8507), .B(g8522), .C(g8537), .Z(g12942) ) ;
INV     gate7907  (.A(g12942), .Z(g14268) ) ;
NOR3    gate7908  (.A(g10210), .B(g10296), .C(g10372), .Z(g12043) ) ;
INV     gate7909  (.A(g12043), .Z(g14273) ) ;
NOR3    gate7910  (.A(g10212), .B(g10299), .C(g10375), .Z(g12044) ) ;
INV     gate7911  (.A(g12044), .Z(g14280) ) ;
NOR3    gate7912  (.A(g10219), .B(g10304), .C(g10381), .Z(g12048) ) ;
INV     gate7913  (.A(g12048), .Z(g14286) ) ;
NOR3    gate7914  (.A(g10220), .B(g10306), .C(g10384), .Z(g12049) ) ;
INV     gate7915  (.A(g12049), .Z(g14290) ) ;
NOR3    gate7916  (.A(g10222), .B(g10309), .C(g10387), .Z(g12050) ) ;
INV     gate7917  (.A(g12050), .Z(g14291) ) ;
NOR3    gate7918  (.A(g8510), .B(g8525), .C(g8540), .Z(g12949) ) ;
INV     gate7919  (.A(g12949), .Z(g14292) ) ;
NAND2   gate7920  (.A(g8296), .B(g3618), .Z(g13156) ) ;
INV     gate7921  (.A(g13156), .Z(II21149) ) ;
INV     gate7922  (.A(II21149), .Z(g14298) ) ;
NOR3    gate7923  (.A(g10225), .B(g10311), .C(g10388), .Z(g12056) ) ;
INV     gate7924  (.A(g12056), .Z(g14301) ) ;
NOR3    gate7925  (.A(g10228), .B(g10313), .C(g10391), .Z(g12057) ) ;
INV     gate7926  (.A(g12057), .Z(g14309) ) ;
NOR3    gate7927  (.A(g10251), .B(g10320), .C(g10396), .Z(g12060) ) ;
INV     gate7928  (.A(g12060), .Z(g14316) ) ;
NOR3    gate7929  (.A(g10255), .B(g10323), .C(g10401), .Z(g12061) ) ;
INV     gate7930  (.A(g12061), .Z(g14320) ) ;
NOR3    gate7931  (.A(g10258), .B(g10326), .C(g10403), .Z(g12062) ) ;
INV     gate7932  (.A(g12062), .Z(g14321) ) ;
NOR3    gate7933  (.A(g8513), .B(g8528), .C(g8543), .Z(g12959) ) ;
INV     gate7934  (.A(g12959), .Z(g14322) ) ;
NAND2   gate7935  (.A(g8305), .B(g7265), .Z(g12538) ) ;
INV     gate7936  (.A(g12538), .Z(II21160) ) ;
INV     gate7937  (.A(II21160), .Z(g14329) ) ;
NOR3    gate7938  (.A(g10271), .B(g10352), .C(g10412), .Z(g12068) ) ;
INV     gate7939  (.A(g12068), .Z(g14332) ) ;
AND4    gate7940  (.A(g10693), .B(g2883), .C(g7562), .D(g10711), .Z(g13110) ) ;
INV     gate7941  (.A(g13110), .Z(II21165) ) ;
INV     gate7942  (.A(II21165), .Z(g14337) ) ;
NOR3    gate7943  (.A(g8517), .B(g8532), .C(g8546), .Z(g12967) ) ;
INV     gate7944  (.A(g12967), .Z(g14342) ) ;
NOR3    gate7945  (.A(g10281), .B(g10361), .C(g10422), .Z(g12079) ) ;
INV     gate7946  (.A(g12079), .Z(g14347) ) ;
NOR3    gate7947  (.A(g10287), .B(g10366), .C(g10433), .Z(g12081) ) ;
INV     gate7948  (.A(g12081), .Z(g14352) ) ;
NOR3    gate7949  (.A(g10290), .B(g10368), .C(g10435), .Z(g12082) ) ;
INV     gate7950  (.A(g12082), .Z(g14355) ) ;
NOR3    gate7951  (.A(g10293), .B(g10371), .C(g10438), .Z(g12083) ) ;
INV     gate7952  (.A(g12083), .Z(g14359) ) ;
NOR3    gate7953  (.A(g8520), .B(g8535), .C(g8548), .Z(g12968) ) ;
INV     gate7954  (.A(g12968), .Z(g14360) ) ;
NOR3    gate7955  (.A(g10297), .B(g10373), .C(g10439), .Z(g12090) ) ;
INV     gate7956  (.A(g12090), .Z(g14366) ) ;
NOR3    gate7957  (.A(g10302), .B(g10379), .C(g10444), .Z(g12098) ) ;
INV     gate7958  (.A(g12098), .Z(g14371) ) ;
NOR3    gate7959  (.A(g10305), .B(g10382), .C(g10446), .Z(g12099) ) ;
INV     gate7960  (.A(g12099), .Z(g14374) ) ;
NOR3    gate7961  (.A(g10307), .B(g10385), .C(g10449), .Z(g12100) ) ;
INV     gate7962  (.A(g12100), .Z(g14378) ) ;
INV     gate7963  (.A(g11749), .Z(II21178) ) ;
INV     gate7964  (.A(II21178), .Z(g14381) ) ;
NOR3    gate7965  (.A(g8523), .B(g8538), .C(g8551), .Z(g12970) ) ;
INV     gate7966  (.A(g12970), .Z(g14385) ) ;
NOR3    gate7967  (.A(g8526), .B(g8541), .C(g8554), .Z(g12971) ) ;
INV     gate7968  (.A(g12971), .Z(g14390) ) ;
NOR3    gate7969  (.A(g10312), .B(g10389), .C(g10451), .Z(g12107) ) ;
INV     gate7970  (.A(g12107), .Z(g14395) ) ;
NOR3    gate7971  (.A(g10314), .B(g10392), .C(g10454), .Z(g12108) ) ;
INV     gate7972  (.A(g12108), .Z(g14402) ) ;
NOR3    gate7973  (.A(g10321), .B(g10397), .C(g10460), .Z(g12112) ) ;
INV     gate7974  (.A(g12112), .Z(g14408) ) ;
NOR3    gate7975  (.A(g10322), .B(g10399), .C(g10463), .Z(g12113) ) ;
INV     gate7976  (.A(g12113), .Z(g14412) ) ;
NOR3    gate7977  (.A(g10324), .B(g10402), .C(g10466), .Z(g12114) ) ;
INV     gate7978  (.A(g12114), .Z(g14413) ) ;
NOR3    gate7979  (.A(g8529), .B(g8544), .C(g8557), .Z(g12978) ) ;
INV     gate7980  (.A(g12978), .Z(g14414) ) ;
NAND2   gate7981  (.A(g8305), .B(g3774), .Z(g13165) ) ;
INV     gate7982  (.A(g13165), .Z(II21190) ) ;
INV     gate7983  (.A(II21190), .Z(g14420) ) ;
NOR3    gate7984  (.A(g10327), .B(g10404), .C(g10467), .Z(g12120) ) ;
INV     gate7985  (.A(g12120), .Z(g14423) ) ;
NOR3    gate7986  (.A(g10330), .B(g10406), .C(g10470), .Z(g12121) ) ;
INV     gate7987  (.A(g12121), .Z(g14431) ) ;
NOR3    gate7988  (.A(g10353), .B(g10413), .C(g10475), .Z(g12124) ) ;
INV     gate7989  (.A(g12124), .Z(g14438) ) ;
NOR3    gate7990  (.A(g9367), .B(g9441), .C(g9521), .Z(g11768) ) ;
INV     gate7991  (.A(g11768), .Z(g14442) ) ;
NOR3    gate7992  (.A(g10369), .B(g10436), .C(g10496), .Z(g12146) ) ;
INV     gate7993  (.A(g12146), .Z(g14450) ) ;
NOR3    gate7994  (.A(g8536), .B(g8549), .C(g8559), .Z(g12991) ) ;
INV     gate7995  (.A(g12991), .Z(g14454) ) ;
NOR3    gate7996  (.A(g10374), .B(g10440), .C(g10498), .Z(g12151) ) ;
INV     gate7997  (.A(g12151), .Z(g14459) ) ;
NOR3    gate7998  (.A(g10380), .B(g10445), .C(g10509), .Z(g12153) ) ;
INV     gate7999  (.A(g12153), .Z(g14464) ) ;
NOR3    gate8000  (.A(g10383), .B(g10447), .C(g10511), .Z(g12154) ) ;
INV     gate8001  (.A(g12154), .Z(g14467) ) ;
NOR3    gate8002  (.A(g10386), .B(g10450), .C(g10514), .Z(g12155) ) ;
INV     gate8003  (.A(g12155), .Z(g14471) ) ;
NOR3    gate8004  (.A(g8539), .B(g8552), .C(g8561), .Z(g12992) ) ;
INV     gate8005  (.A(g12992), .Z(g14472) ) ;
NOR3    gate8006  (.A(g10390), .B(g10452), .C(g10515), .Z(g12162) ) ;
INV     gate8007  (.A(g12162), .Z(g14478) ) ;
NOR3    gate8008  (.A(g10395), .B(g10458), .C(g10520), .Z(g12170) ) ;
INV     gate8009  (.A(g12170), .Z(g14483) ) ;
NOR3    gate8010  (.A(g10398), .B(g10461), .C(g10522), .Z(g12171) ) ;
INV     gate8011  (.A(g12171), .Z(g14486) ) ;
NOR3    gate8012  (.A(g10400), .B(g10464), .C(g10525), .Z(g12172) ) ;
INV     gate8013  (.A(g12172), .Z(g14490) ) ;
INV     gate8014  (.A(g11749), .Z(II21208) ) ;
INV     gate8015  (.A(II21208), .Z(g14493) ) ;
NOR3    gate8016  (.A(g8542), .B(g8555), .C(g8564), .Z(g12994) ) ;
INV     gate8017  (.A(g12994), .Z(g14497) ) ;
NOR3    gate8018  (.A(g8545), .B(g8558), .C(g8567), .Z(g12995) ) ;
INV     gate8019  (.A(g12995), .Z(g14502) ) ;
NOR3    gate8020  (.A(g10405), .B(g10468), .C(g10527), .Z(g12179) ) ;
INV     gate8021  (.A(g12179), .Z(g14507) ) ;
NOR3    gate8022  (.A(g10407), .B(g10471), .C(g10530), .Z(g12180) ) ;
INV     gate8023  (.A(g12180), .Z(g14514) ) ;
NOR3    gate8024  (.A(g10414), .B(g10476), .C(g10536), .Z(g12184) ) ;
INV     gate8025  (.A(g12184), .Z(g14520) ) ;
NOR3    gate8026  (.A(g10415), .B(g10478), .C(g10539), .Z(g12185) ) ;
INV     gate8027  (.A(g12185), .Z(g14524) ) ;
NOR3    gate8028  (.A(g10437), .B(g10497), .C(g10558), .Z(g12195) ) ;
INV     gate8029  (.A(g12195), .Z(g14525) ) ;
NOR3    gate8030  (.A(g9464), .B(g9583), .C(g9663), .Z(g11785) ) ;
INV     gate8031  (.A(g11785), .Z(g14529) ) ;
NOR3    gate8032  (.A(g10448), .B(g10512), .C(g10570), .Z(g12208) ) ;
INV     gate8033  (.A(g12208), .Z(g14537) ) ;
NOR3    gate8034  (.A(g8553), .B(g8562), .C(g8570), .Z(g13001) ) ;
INV     gate8035  (.A(g13001), .Z(g14541) ) ;
NOR3    gate8036  (.A(g10453), .B(g10516), .C(g10572), .Z(g12213) ) ;
INV     gate8037  (.A(g12213), .Z(g14546) ) ;
NOR3    gate8038  (.A(g10459), .B(g10521), .C(g10583), .Z(g12215) ) ;
INV     gate8039  (.A(g12215), .Z(g14551) ) ;
NOR3    gate8040  (.A(g10462), .B(g10523), .C(g10585), .Z(g12216) ) ;
INV     gate8041  (.A(g12216), .Z(g14554) ) ;
NOR3    gate8042  (.A(g10465), .B(g10526), .C(g10588), .Z(g12217) ) ;
INV     gate8043  (.A(g12217), .Z(g14558) ) ;
NOR3    gate8044  (.A(g8556), .B(g8565), .C(g8572), .Z(g13002) ) ;
INV     gate8045  (.A(g13002), .Z(g14559) ) ;
NOR3    gate8046  (.A(g10469), .B(g10528), .C(g10589), .Z(g12224) ) ;
INV     gate8047  (.A(g12224), .Z(g14565) ) ;
NOR3    gate8048  (.A(g10474), .B(g10534), .C(g10594), .Z(g12232) ) ;
INV     gate8049  (.A(g12232), .Z(g14570) ) ;
NOR3    gate8050  (.A(g10477), .B(g10537), .C(g10596), .Z(g12233) ) ;
INV     gate8051  (.A(g12233), .Z(g14573) ) ;
NOR3    gate8052  (.A(g10479), .B(g10540), .C(g10599), .Z(g12234) ) ;
INV     gate8053  (.A(g12234), .Z(g14577) ) ;
NOR3    gate8054  (.A(g10513), .B(g10571), .C(g10615), .Z(g12250) ) ;
INV     gate8055  (.A(g12250), .Z(g14580) ) ;
NOR3    gate8056  (.A(g9606), .B(g9725), .C(g9809), .Z(g11811) ) ;
INV     gate8057  (.A(g11811), .Z(g14584) ) ;
NOR3    gate8058  (.A(g10524), .B(g10586), .C(g10627), .Z(g12263) ) ;
INV     gate8059  (.A(g12263), .Z(g14592) ) ;
NOR3    gate8060  (.A(g8566), .B(g8573), .C(g8576), .Z(g13022) ) ;
INV     gate8061  (.A(g13022), .Z(g14596) ) ;
NOR3    gate8062  (.A(g10529), .B(g10590), .C(g10629), .Z(g12268) ) ;
INV     gate8063  (.A(g12268), .Z(g14601) ) ;
NOR3    gate8064  (.A(g10535), .B(g10595), .C(g10640), .Z(g12270) ) ;
INV     gate8065  (.A(g12270), .Z(g14606) ) ;
NOR3    gate8066  (.A(g10538), .B(g10597), .C(g10642), .Z(g12271) ) ;
INV     gate8067  (.A(g12271), .Z(g14609) ) ;
NOR3    gate8068  (.A(g10541), .B(g10600), .C(g10645), .Z(g12272) ) ;
INV     gate8069  (.A(g12272), .Z(g14613) ) ;
NOR3    gate8070  (.A(g10587), .B(g10628), .C(g10662), .Z(g12293) ) ;
INV     gate8071  (.A(g12293), .Z(g14614) ) ;
NOR3    gate8072  (.A(g9748), .B(g9871), .C(g9955), .Z(g11844) ) ;
INV     gate8073  (.A(g11844), .Z(g14618) ) ;
NOR3    gate8074  (.A(g10598), .B(g10643), .C(g10674), .Z(g12306) ) ;
INV     gate8075  (.A(g12306), .Z(g14626) ) ;
NOR3    gate8076  (.A(g9026), .B(g9047), .C(g9061), .Z(g13378) ) ;
INV     gate8077  (.A(g13378), .Z(II21241) ) ;
INV     gate8078  (.A(II21241), .Z(g14630) ) ;
NOR3    gate8079  (.A(g10644), .B(g10675), .C(g10692), .Z(g12329) ) ;
INV     gate8080  (.A(g12329), .Z(g14637) ) ;
NOR3    gate8081  (.A(g9635), .B(g9763), .C(g9891), .Z(g11823) ) ;
INV     gate8082  (.A(g11823), .Z(g14641) ) ;
NOR3    gate8083  (.A(g9062), .B(g9075), .C(g9091), .Z(g11624) ) ;
INV     gate8084  (.A(g11624), .Z(II21246) ) ;
INV     gate8085  (.A(II21246), .Z(g14642) ) ;
NOR3    gate8086  (.A(g9049), .B(g9064), .C(g9078), .Z(g11600) ) ;
INV     gate8087  (.A(g11600), .Z(II21249) ) ;
INV     gate8088  (.A(II21249), .Z(g14650) ) ;
NOR3    gate8089  (.A(g9076), .B(g9092), .C(g9102), .Z(g11644) ) ;
INV     gate8090  (.A(g11644), .Z(II21252) ) ;
INV     gate8091  (.A(II21252), .Z(g14657) ) ;
NOR3    gate8092  (.A(g9781), .B(g9909), .C(g10045), .Z(g11865) ) ;
INV     gate8093  (.A(g11865), .Z(g14668) ) ;
NOR3    gate8094  (.A(g9079), .B(g9094), .C(g9103), .Z(g11647) ) ;
INV     gate8095  (.A(g11647), .Z(II21256) ) ;
INV     gate8096  (.A(II21256), .Z(g14669) ) ;
NOR3    gate8097  (.A(g9066), .B(g9081), .C(g9097), .Z(g11630) ) ;
INV     gate8098  (.A(g11630), .Z(II21259) ) ;
INV     gate8099  (.A(II21259), .Z(g14677) ) ;
INV     gate8100  (.A(g11713), .Z(II21262) ) ;
INV     gate8101  (.A(II21262), .Z(g14684) ) ;
NOR3    gate8102  (.A(g10495), .B(g10557), .C(g10604), .Z(g12245) ) ;
INV     gate8103  (.A(g12245), .Z(g14685) ) ;
NOR3    gate8104  (.A(g9095), .B(g9104), .C(g9112), .Z(g11663) ) ;
INV     gate8105  (.A(g11663), .Z(II21267) ) ;
INV     gate8106  (.A(II21267), .Z(g14691) ) ;
NOR3    gate8107  (.A(g9927), .B(g10063), .C(g10154), .Z(g11907) ) ;
INV     gate8108  (.A(g11907), .Z(g14702) ) ;
NOR3    gate8109  (.A(g9098), .B(g9106), .C(g9113), .Z(g11666) ) ;
INV     gate8110  (.A(g11666), .Z(II21271) ) ;
INV     gate8111  (.A(II21271), .Z(g14703) ) ;
NOR3    gate8112  (.A(g9083), .B(g9100), .C(g9109), .Z(g11653) ) ;
INV     gate8113  (.A(g11653), .Z(II21274) ) ;
INV     gate8114  (.A(II21274), .Z(g14711) ) ;
INV     gate8115  (.A(g12430), .Z(II21277) ) ;
INV     gate8116  (.A(II21277), .Z(g14718) ) ;
NOR3    gate8117  (.A(g10569), .B(g10614), .C(g10651), .Z(g12288) ) ;
INV     gate8118  (.A(g12288), .Z(g14719) ) ;
NOR3    gate8119  (.A(g9107), .B(g9114), .C(g9120), .Z(g11675) ) ;
INV     gate8120  (.A(g11675), .Z(II21282) ) ;
INV     gate8121  (.A(II21282), .Z(g14725) ) ;
NOR3    gate8122  (.A(g10081), .B(g10172), .C(g10259), .Z(g11957) ) ;
INV     gate8123  (.A(g11957), .Z(g14736) ) ;
NOR3    gate8124  (.A(g9110), .B(g9116), .C(g9121), .Z(g11678) ) ;
INV     gate8125  (.A(g11678), .Z(II21286) ) ;
INV     gate8126  (.A(II21286), .Z(g14737) ) ;
INV     gate8127  (.A(g12434), .Z(II21289) ) ;
INV     gate8128  (.A(II21289), .Z(g14745) ) ;
INV     gate8129  (.A(g11888), .Z(II21292) ) ;
INV     gate8130  (.A(II21292), .Z(g14746) ) ;
NOR3    gate8131  (.A(g10626), .B(g10661), .C(g10681), .Z(g12324) ) ;
INV     gate8132  (.A(g12324), .Z(g14747) ) ;
NOR3    gate8133  (.A(g9117), .B(g9122), .C(g9126), .Z(g11687) ) ;
INV     gate8134  (.A(g11687), .Z(II21297) ) ;
INV     gate8135  (.A(II21297), .Z(g14753) ) ;
INV     gate8136  (.A(g11791), .Z(g14764) ) ;
INV     gate8137  (.A(g12438), .Z(II21301) ) ;
INV     gate8138  (.A(II21301), .Z(g14765) ) ;
INV     gate8139  (.A(g11927), .Z(II21304) ) ;
INV     gate8140  (.A(II21304), .Z(g14766) ) ;
NOR3    gate8141  (.A(g10673), .B(g10691), .C(g10710), .Z(g12352) ) ;
INV     gate8142  (.A(g12352), .Z(g14768) ) ;
INV     gate8143  (.A(g12332), .Z(II21310) ) ;
INV     gate8144  (.A(II21310), .Z(g14774) ) ;
INV     gate8145  (.A(g11743), .Z(II21313) ) ;
INV     gate8146  (.A(II21313), .Z(g14775) ) ;
NOR3    gate8147  (.A(g10199), .B(g10284), .C(g10362), .Z(g12033) ) ;
INV     gate8148  (.A(g12033), .Z(g14776) ) ;
INV     gate8149  (.A(g11848), .Z(g14794) ) ;
INV     gate8150  (.A(g12362), .Z(II21318) ) ;
INV     gate8151  (.A(II21318), .Z(g14795) ) ;
INV     gate8152  (.A(g11758), .Z(II21321) ) ;
INV     gate8153  (.A(II21321), .Z(g14796) ) ;
NOR3    gate8154  (.A(g10285), .B(g10363), .C(g10430), .Z(g12080) ) ;
INV     gate8155  (.A(g12080), .Z(g14797) ) ;
NOR3    gate8156  (.A(g10301), .B(g10377), .C(g10441), .Z(g12097) ) ;
INV     gate8157  (.A(g12097), .Z(g14811) ) ;
INV     gate8158  (.A(g12378), .Z(II21326) ) ;
INV     gate8159  (.A(II21326), .Z(g14829) ) ;
INV     gate8160  (.A(g11766), .Z(II21329) ) ;
INV     gate8161  (.A(II21329), .Z(g14830) ) ;
NOR3    gate8162  (.A(g9639), .B(g9764), .C(g9892), .Z(g11828) ) ;
INV     gate8163  (.A(g11828), .Z(g14831) ) ;
NOR3    gate8164  (.A(g10364), .B(g10431), .C(g10492), .Z(g12145) ) ;
INV     gate8165  (.A(g12145), .Z(g14837) ) ;
NOR3    gate8166  (.A(g10378), .B(g10442), .C(g10506), .Z(g12152) ) ;
INV     gate8167  (.A(g12152), .Z(g14849) ) ;
NOR3    gate8168  (.A(g10394), .B(g10456), .C(g10517), .Z(g12169) ) ;
INV     gate8169  (.A(g12169), .Z(g14863) ) ;
INV     gate8170  (.A(g11923), .Z(g14881) ) ;
INV     gate8171  (.A(g12408), .Z(II21337) ) ;
INV     gate8172  (.A(II21337), .Z(g14882) ) ;
INV     gate8173  (.A(g11779), .Z(II21340) ) ;
INV     gate8174  (.A(II21340), .Z(g14883) ) ;
NOR3    gate8175  (.A(g9765), .B(g9893), .C(g10012), .Z(g11860) ) ;
INV     gate8176  (.A(g11860), .Z(g14885) ) ;
NOR3    gate8177  (.A(g10432), .B(g10493), .C(g10555), .Z(g12193) ) ;
INV     gate8178  (.A(g12193), .Z(g14895) ) ;
NOR3    gate8179  (.A(g9785), .B(g9910), .C(g10046), .Z(g11870) ) ;
INV     gate8180  (.A(g11870), .Z(g14904) ) ;
NOR3    gate8181  (.A(g10443), .B(g10507), .C(g10566), .Z(g12207) ) ;
INV     gate8182  (.A(g12207), .Z(g14910) ) ;
NOR3    gate8183  (.A(g10457), .B(g10518), .C(g10580), .Z(g12214) ) ;
INV     gate8184  (.A(g12214), .Z(g14922) ) ;
NOR3    gate8185  (.A(g10473), .B(g10532), .C(g10591), .Z(g12231) ) ;
INV     gate8186  (.A(g12231), .Z(g14936) ) ;
INV     gate8187  (.A(g12420), .Z(II21351) ) ;
INV     gate8188  (.A(II21351), .Z(g14954) ) ;
INV     gate8189  (.A(g11798), .Z(II21354) ) ;
INV     gate8190  (.A(II21354), .Z(g14955) ) ;
INV     gate8191  (.A(g11976), .Z(g14959) ) ;
NAND2   gate8192  (.A(g9534), .B(g6678), .Z(g13026) ) ;
INV     gate8193  (.A(g13026), .Z(II21361) ) ;
INV     gate8194  (.A(II21361), .Z(g14960) ) ;
NAND2   gate8195  (.A(g9534), .B(g6678), .Z(g13028) ) ;
INV     gate8196  (.A(g13028), .Z(II21364) ) ;
INV     gate8197  (.A(II21364), .Z(g14963) ) ;
NOR3    gate8198  (.A(g9911), .B(g10047), .C(g10121), .Z(g11902) ) ;
INV     gate8199  (.A(g11902), .Z(g14966) ) ;
NOR3    gate8200  (.A(g10508), .B(g10567), .C(g10612), .Z(g12248) ) ;
INV     gate8201  (.A(g12248), .Z(g14976) ) ;
NOR3    gate8202  (.A(g9931), .B(g10064), .C(g10155), .Z(g11912) ) ;
INV     gate8203  (.A(g11912), .Z(g14985) ) ;
NOR3    gate8204  (.A(g10519), .B(g10581), .C(g10623), .Z(g12262) ) ;
INV     gate8205  (.A(g12262), .Z(g14991) ) ;
NOR3    gate8206  (.A(g10533), .B(g10592), .C(g10637), .Z(g12269) ) ;
INV     gate8207  (.A(g12269), .Z(g15003) ) ;
INV     gate8208  (.A(g12009), .Z(g15017) ) ;
INV     gate8209  (.A(g12424), .Z(II21374) ) ;
INV     gate8210  (.A(II21374), .Z(g15018) ) ;
INV     gate8211  (.A(g11821), .Z(II21377) ) ;
INV     gate8212  (.A(II21377), .Z(g15019) ) ;
INV     gate8213  (.A(g13157), .Z(II21381) ) ;
INV     gate8214  (.A(II21381), .Z(g15021) ) ;
NOR3    gate8215  (.A(g9442), .B(g9522), .C(g9633), .Z(g11781) ) ;
INV     gate8216  (.A(g11781), .Z(g15022) ) ;
INV     gate8217  (.A(g12027), .Z(g15032) ) ;
INV     gate8218  (.A(g12030), .Z(g15033) ) ;
NOR2    gate8219  (.A(g10038), .B(g6284), .Z(g12883) ) ;
INV     gate8220  (.A(g12883), .Z(II21389) ) ;
INV     gate8221  (.A(II21389), .Z(g15034) ) ;
NAND2   gate8222  (.A(g9534), .B(g6912), .Z(g13020) ) ;
INV     gate8223  (.A(g13020), .Z(II21392) ) ;
INV     gate8224  (.A(II21392), .Z(g15037) ) ;
NAND2   gate8225  (.A(g9534), .B(g6678), .Z(g13034) ) ;
INV     gate8226  (.A(g13034), .Z(II21395) ) ;
INV     gate8227  (.A(II21395), .Z(g15040) ) ;
NAND2   gate8228  (.A(g9534), .B(g6912), .Z(g13021) ) ;
INV     gate8229  (.A(g13021), .Z(II21398) ) ;
INV     gate8230  (.A(II21398), .Z(g15043) ) ;
INV     gate8231  (.A(g12045), .Z(g15048) ) ;
NAND2   gate8232  (.A(g9676), .B(g6980), .Z(g13037) ) ;
INV     gate8233  (.A(g13037), .Z(II21404) ) ;
INV     gate8234  (.A(II21404), .Z(g15049) ) ;
NAND2   gate8235  (.A(g9676), .B(g6980), .Z(g13039) ) ;
INV     gate8236  (.A(g13039), .Z(II21407) ) ;
INV     gate8237  (.A(II21407), .Z(g15052) ) ;
NOR3    gate8238  (.A(g10065), .B(g10156), .C(g10226), .Z(g11952) ) ;
INV     gate8239  (.A(g11952), .Z(g15055) ) ;
NOR3    gate8240  (.A(g10582), .B(g10624), .C(g10659), .Z(g12291) ) ;
INV     gate8241  (.A(g12291), .Z(g15065) ) ;
NOR3    gate8242  (.A(g10085), .B(g10173), .C(g10260), .Z(g11962) ) ;
INV     gate8243  (.A(g11962), .Z(g15074) ) ;
NOR3    gate8244  (.A(g10593), .B(g10638), .C(g10670), .Z(g12305) ) ;
INV     gate8245  (.A(g12305), .Z(g15080) ) ;
INV     gate8246  (.A(g11854), .Z(II21415) ) ;
INV     gate8247  (.A(II21415), .Z(g15092) ) ;
INV     gate8248  (.A(g13166), .Z(II21420) ) ;
INV     gate8249  (.A(II21420), .Z(g15095) ) ;
NOR3    gate8250  (.A(g9523), .B(g9634), .C(g9762), .Z(g11800) ) ;
INV     gate8251  (.A(g11800), .Z(g15096) ) ;
NAND2   gate8252  (.A(g9534), .B(g3366), .Z(g11661) ) ;
INV     gate8253  (.A(g11661), .Z(II21426) ) ;
INV     gate8254  (.A(II21426), .Z(g15106) ) ;
NAND2   gate8255  (.A(g9534), .B(g6912), .Z(g13027) ) ;
INV     gate8256  (.A(g13027), .Z(II21429) ) ;
INV     gate8257  (.A(II21429), .Z(g15109) ) ;
NAND2   gate8258  (.A(g9534), .B(g6678), .Z(g13044) ) ;
INV     gate8259  (.A(g13044), .Z(II21432) ) ;
INV     gate8260  (.A(II21432), .Z(g15112) ) ;
NAND2   gate8261  (.A(g9534), .B(g3366), .Z(g11662) ) ;
INV     gate8262  (.A(g11662), .Z(II21435) ) ;
INV     gate8263  (.A(II21435), .Z(g15115) ) ;
NOR3    gate8264  (.A(g9584), .B(g9664), .C(g9779), .Z(g11807) ) ;
INV     gate8265  (.A(g11807), .Z(g15118) ) ;
INV     gate8266  (.A(g12091), .Z(g15128) ) ;
INV     gate8267  (.A(g12094), .Z(g15129) ) ;
NOR2    gate8268  (.A(g10147), .B(g6421), .Z(g12923) ) ;
INV     gate8269  (.A(g12923), .Z(II21443) ) ;
INV     gate8270  (.A(II21443), .Z(g15130) ) ;
NAND2   gate8271  (.A(g9676), .B(g7162), .Z(g13029) ) ;
INV     gate8272  (.A(g13029), .Z(II21446) ) ;
INV     gate8273  (.A(II21446), .Z(g15133) ) ;
NAND2   gate8274  (.A(g9676), .B(g6980), .Z(g13047) ) ;
INV     gate8275  (.A(g13047), .Z(II21449) ) ;
INV     gate8276  (.A(II21449), .Z(g15136) ) ;
NAND2   gate8277  (.A(g9676), .B(g7162), .Z(g13030) ) ;
INV     gate8278  (.A(g13030), .Z(II21452) ) ;
INV     gate8279  (.A(II21452), .Z(g15139) ) ;
INV     gate8280  (.A(g12109), .Z(g15144) ) ;
NAND2   gate8281  (.A(g9822), .B(g7230), .Z(g13050) ) ;
INV     gate8282  (.A(g13050), .Z(II21458) ) ;
INV     gate8283  (.A(II21458), .Z(g15145) ) ;
NAND2   gate8284  (.A(g9822), .B(g7230), .Z(g13052) ) ;
INV     gate8285  (.A(g13052), .Z(II21461) ) ;
INV     gate8286  (.A(II21461), .Z(g15148) ) ;
NOR3    gate8287  (.A(g10174), .B(g10261), .C(g10328), .Z(g12005) ) ;
INV     gate8288  (.A(g12005), .Z(g15151) ) ;
NOR3    gate8289  (.A(g10639), .B(g10671), .C(g10689), .Z(g12327) ) ;
INV     gate8290  (.A(g12327), .Z(g15161) ) ;
INV     gate8291  (.A(g12125), .Z(g15170) ) ;
INV     gate8292  (.A(g12136), .Z(g15174) ) ;
INV     gate8293  (.A(g12139), .Z(g15175) ) ;
INV     gate8294  (.A(g12142), .Z(g15176) ) ;
NOR3    gate8295  (.A(g10650), .B(g10678), .C(g10704), .Z(g12339) ) ;
INV     gate8296  (.A(g12339), .Z(g15177) ) ;
NAND2   gate8297  (.A(g9534), .B(g3366), .Z(g11672) ) ;
INV     gate8298  (.A(g11672), .Z(II21476) ) ;
INV     gate8299  (.A(II21476), .Z(g15179) ) ;
NAND2   gate8300  (.A(g9534), .B(g6912), .Z(g13035) ) ;
INV     gate8301  (.A(g13035), .Z(II21479) ) ;
INV     gate8302  (.A(II21479), .Z(g15182) ) ;
NAND2   gate8303  (.A(g9534), .B(g6678), .Z(g13058) ) ;
INV     gate8304  (.A(g13058), .Z(II21482) ) ;
INV     gate8305  (.A(II21482), .Z(g15185) ) ;
NOR3    gate8306  (.A(g9665), .B(g9780), .C(g9908), .Z(g11833) ) ;
INV     gate8307  (.A(g11833), .Z(g15188) ) ;
NAND2   gate8308  (.A(g9676), .B(g3522), .Z(g11673) ) ;
INV     gate8309  (.A(g11673), .Z(II21488) ) ;
INV     gate8310  (.A(II21488), .Z(g15198) ) ;
NAND2   gate8311  (.A(g9676), .B(g7162), .Z(g13038) ) ;
INV     gate8312  (.A(g13038), .Z(II21491) ) ;
INV     gate8313  (.A(II21491), .Z(g15201) ) ;
NAND2   gate8314  (.A(g9676), .B(g6980), .Z(g13061) ) ;
INV     gate8315  (.A(g13061), .Z(II21494) ) ;
INV     gate8316  (.A(II21494), .Z(g15204) ) ;
NAND2   gate8317  (.A(g9676), .B(g3522), .Z(g11674) ) ;
INV     gate8318  (.A(g11674), .Z(II21497) ) ;
INV     gate8319  (.A(II21497), .Z(g15207) ) ;
NOR3    gate8320  (.A(g9726), .B(g9810), .C(g9925), .Z(g11840) ) ;
INV     gate8321  (.A(g11840), .Z(g15210) ) ;
INV     gate8322  (.A(g12163), .Z(g15220) ) ;
INV     gate8323  (.A(g12166), .Z(g15221) ) ;
NOR2    gate8324  (.A(g10252), .B(g6626), .Z(g12952) ) ;
INV     gate8325  (.A(g12952), .Z(II21505) ) ;
INV     gate8326  (.A(II21505), .Z(g15222) ) ;
NAND2   gate8327  (.A(g9822), .B(g7358), .Z(g13040) ) ;
INV     gate8328  (.A(g13040), .Z(II21508) ) ;
INV     gate8329  (.A(II21508), .Z(g15225) ) ;
NAND2   gate8330  (.A(g9822), .B(g7230), .Z(g13064) ) ;
INV     gate8331  (.A(g13064), .Z(II21511) ) ;
INV     gate8332  (.A(II21511), .Z(g15228) ) ;
NAND2   gate8333  (.A(g9822), .B(g7358), .Z(g13041) ) ;
INV     gate8334  (.A(g13041), .Z(II21514) ) ;
INV     gate8335  (.A(II21514), .Z(g15231) ) ;
INV     gate8336  (.A(g12181), .Z(g15236) ) ;
NAND2   gate8337  (.A(g9968), .B(g7426), .Z(g13067) ) ;
INV     gate8338  (.A(g13067), .Z(II21520) ) ;
INV     gate8339  (.A(II21520), .Z(g15237) ) ;
NAND2   gate8340  (.A(g9968), .B(g7426), .Z(g13069) ) ;
INV     gate8341  (.A(g13069), .Z(II21523) ) ;
INV     gate8342  (.A(II21523), .Z(g15240) ) ;
NAND2   gate8343  (.A(g9534), .B(g3366), .Z(g11683) ) ;
INV     gate8344  (.A(g11683), .Z(II21531) ) ;
INV     gate8345  (.A(II21531), .Z(g15248) ) ;
NAND2   gate8346  (.A(g9534), .B(g6912), .Z(g13045) ) ;
INV     gate8347  (.A(g13045), .Z(II21534) ) ;
INV     gate8348  (.A(II21534), .Z(g15251) ) ;
NAND2   gate8349  (.A(g9534), .B(g6678), .Z(g13071) ) ;
INV     gate8350  (.A(g13071), .Z(II21537) ) ;
INV     gate8351  (.A(II21537), .Z(g15254) ) ;
INV     gate8352  (.A(g12198), .Z(g15260) ) ;
INV     gate8353  (.A(g12201), .Z(g15261) ) ;
INV     gate8354  (.A(g12204), .Z(g15262) ) ;
NOR3    gate8355  (.A(g10680), .B(g10707), .C(g10724), .Z(g12369) ) ;
INV     gate8356  (.A(g12369), .Z(g15263) ) ;
NAND2   gate8357  (.A(g9676), .B(g3522), .Z(g11684) ) ;
INV     gate8358  (.A(g11684), .Z(II21548) ) ;
INV     gate8359  (.A(II21548), .Z(g15265) ) ;
NAND2   gate8360  (.A(g9676), .B(g7162), .Z(g13048) ) ;
INV     gate8361  (.A(g13048), .Z(II21551) ) ;
INV     gate8362  (.A(II21551), .Z(g15268) ) ;
NAND2   gate8363  (.A(g9676), .B(g6980), .Z(g13074) ) ;
INV     gate8364  (.A(g13074), .Z(II21554) ) ;
INV     gate8365  (.A(II21554), .Z(g15271) ) ;
NOR3    gate8366  (.A(g9811), .B(g9926), .C(g10062), .Z(g11875) ) ;
INV     gate8367  (.A(g11875), .Z(g15274) ) ;
NAND2   gate8368  (.A(g9822), .B(g3678), .Z(g11685) ) ;
INV     gate8369  (.A(g11685), .Z(II21560) ) ;
INV     gate8370  (.A(II21560), .Z(g15284) ) ;
NAND2   gate8371  (.A(g9822), .B(g7358), .Z(g13051) ) ;
INV     gate8372  (.A(g13051), .Z(II21563) ) ;
INV     gate8373  (.A(II21563), .Z(g15287) ) ;
NAND2   gate8374  (.A(g9822), .B(g7230), .Z(g13077) ) ;
INV     gate8375  (.A(g13077), .Z(II21566) ) ;
INV     gate8376  (.A(II21566), .Z(g15290) ) ;
NAND2   gate8377  (.A(g9822), .B(g3678), .Z(g11686) ) ;
INV     gate8378  (.A(g11686), .Z(II21569) ) ;
INV     gate8379  (.A(II21569), .Z(g15293) ) ;
NOR3    gate8380  (.A(g9872), .B(g9956), .C(g10079), .Z(g11882) ) ;
INV     gate8381  (.A(g11882), .Z(g15296) ) ;
INV     gate8382  (.A(g12225), .Z(g15306) ) ;
INV     gate8383  (.A(g12228), .Z(g15307) ) ;
NOR2    gate8384  (.A(g10354), .B(g6890), .Z(g12981) ) ;
INV     gate8385  (.A(g12981), .Z(II21577) ) ;
INV     gate8386  (.A(II21577), .Z(g15308) ) ;
NAND2   gate8387  (.A(g9968), .B(g7488), .Z(g13053) ) ;
INV     gate8388  (.A(g13053), .Z(II21580) ) ;
INV     gate8389  (.A(II21580), .Z(g15311) ) ;
NAND2   gate8390  (.A(g9968), .B(g7426), .Z(g13080) ) ;
INV     gate8391  (.A(g13080), .Z(II21583) ) ;
INV     gate8392  (.A(II21583), .Z(g15314) ) ;
NAND2   gate8393  (.A(g9968), .B(g7488), .Z(g13054) ) ;
INV     gate8394  (.A(g13054), .Z(II21586) ) ;
INV     gate8395  (.A(II21586), .Z(g15317) ) ;
INV     gate8396  (.A(g12239), .Z(g15322) ) ;
INV     gate8397  (.A(g12242), .Z(g15323) ) ;
NAND2   gate8398  (.A(g9534), .B(g3366), .Z(g11691) ) ;
INV     gate8399  (.A(g11691), .Z(II21595) ) ;
INV     gate8400  (.A(II21595), .Z(g15326) ) ;
NAND2   gate8401  (.A(g9534), .B(g6912), .Z(g13059) ) ;
INV     gate8402  (.A(g13059), .Z(II21598) ) ;
INV     gate8403  (.A(II21598), .Z(g15329) ) ;
NAND2   gate8404  (.A(g9534), .B(g6678), .Z(g13087) ) ;
INV     gate8405  (.A(g13087), .Z(II21601) ) ;
INV     gate8406  (.A(II21601), .Z(g15332) ) ;
NAND2   gate8407  (.A(g9676), .B(g3522), .Z(g11692) ) ;
INV     gate8408  (.A(g11692), .Z(II21609) ) ;
INV     gate8409  (.A(II21609), .Z(g15340) ) ;
NAND2   gate8410  (.A(g9676), .B(g7162), .Z(g13062) ) ;
INV     gate8411  (.A(g13062), .Z(II21612) ) ;
INV     gate8412  (.A(II21612), .Z(g15343) ) ;
NAND2   gate8413  (.A(g9676), .B(g6980), .Z(g13090) ) ;
INV     gate8414  (.A(g13090), .Z(II21615) ) ;
INV     gate8415  (.A(II21615), .Z(g15346) ) ;
INV     gate8416  (.A(g12253), .Z(g15352) ) ;
INV     gate8417  (.A(g12256), .Z(g15353) ) ;
INV     gate8418  (.A(g12259), .Z(g15354) ) ;
NOR3    gate8419  (.A(g10709), .B(g10727), .C(g10745), .Z(g12388) ) ;
INV     gate8420  (.A(g12388), .Z(g15355) ) ;
NAND2   gate8421  (.A(g9822), .B(g3678), .Z(g11693) ) ;
INV     gate8422  (.A(g11693), .Z(II21626) ) ;
INV     gate8423  (.A(II21626), .Z(g15357) ) ;
NAND2   gate8424  (.A(g9822), .B(g7358), .Z(g13065) ) ;
INV     gate8425  (.A(g13065), .Z(II21629) ) ;
INV     gate8426  (.A(II21629), .Z(g15360) ) ;
NAND2   gate8427  (.A(g9822), .B(g7230), .Z(g13093) ) ;
INV     gate8428  (.A(g13093), .Z(II21632) ) ;
INV     gate8429  (.A(II21632), .Z(g15363) ) ;
NOR3    gate8430  (.A(g9957), .B(g10080), .C(g10171), .Z(g11917) ) ;
INV     gate8431  (.A(g11917), .Z(g15366) ) ;
NAND2   gate8432  (.A(g9968), .B(g3834), .Z(g11694) ) ;
INV     gate8433  (.A(g11694), .Z(II21638) ) ;
INV     gate8434  (.A(II21638), .Z(g15376) ) ;
NAND2   gate8435  (.A(g9968), .B(g7488), .Z(g13068) ) ;
INV     gate8436  (.A(g13068), .Z(II21641) ) ;
INV     gate8437  (.A(II21641), .Z(g15379) ) ;
NAND2   gate8438  (.A(g9968), .B(g7426), .Z(g13096) ) ;
INV     gate8439  (.A(g13096), .Z(II21644) ) ;
INV     gate8440  (.A(II21644), .Z(g15382) ) ;
NAND2   gate8441  (.A(g9968), .B(g3834), .Z(g11695) ) ;
INV     gate8442  (.A(g11695), .Z(II21647) ) ;
INV     gate8443  (.A(II21647), .Z(g15385) ) ;
INV     gate8444  (.A(g12279), .Z(g15390) ) ;
NAND2   gate8445  (.A(g9534), .B(g3366), .Z(g11696) ) ;
INV     gate8446  (.A(g11696), .Z(II21655) ) ;
INV     gate8447  (.A(II21655), .Z(g15393) ) ;
NAND2   gate8448  (.A(g9534), .B(g6912), .Z(g13072) ) ;
INV     gate8449  (.A(g13072), .Z(II21658) ) ;
INV     gate8450  (.A(II21658), .Z(g15396) ) ;
NAND2   gate8451  (.A(g9534), .B(g6678), .Z(g13098) ) ;
INV     gate8452  (.A(g13098), .Z(II21661) ) ;
INV     gate8453  (.A(II21661), .Z(g15399) ) ;
NAND2   gate8454  (.A(g9534), .B(g6678), .Z(g13100) ) ;
INV     gate8455  (.A(g13100), .Z(II21666) ) ;
INV     gate8456  (.A(II21666), .Z(g15404) ) ;
INV     gate8457  (.A(g12282), .Z(g15408) ) ;
INV     gate8458  (.A(g12285), .Z(g15409) ) ;
NAND2   gate8459  (.A(g9676), .B(g3522), .Z(g11698) ) ;
INV     gate8460  (.A(g11698), .Z(II21674) ) ;
INV     gate8461  (.A(II21674), .Z(g15412) ) ;
NAND2   gate8462  (.A(g9676), .B(g7162), .Z(g13075) ) ;
INV     gate8463  (.A(g13075), .Z(II21677) ) ;
INV     gate8464  (.A(II21677), .Z(g15415) ) ;
NAND2   gate8465  (.A(g9676), .B(g6980), .Z(g13102) ) ;
INV     gate8466  (.A(g13102), .Z(II21680) ) ;
INV     gate8467  (.A(II21680), .Z(g15418) ) ;
NAND2   gate8468  (.A(g9822), .B(g3678), .Z(g11699) ) ;
INV     gate8469  (.A(g11699), .Z(II21688) ) ;
INV     gate8470  (.A(II21688), .Z(g15426) ) ;
NAND2   gate8471  (.A(g9822), .B(g7358), .Z(g13078) ) ;
INV     gate8472  (.A(g13078), .Z(II21691) ) ;
INV     gate8473  (.A(II21691), .Z(g15429) ) ;
NAND2   gate8474  (.A(g9822), .B(g7230), .Z(g13105) ) ;
INV     gate8475  (.A(g13105), .Z(II21694) ) ;
INV     gate8476  (.A(II21694), .Z(g15432) ) ;
INV     gate8477  (.A(g12296), .Z(g15438) ) ;
INV     gate8478  (.A(g12299), .Z(g15439) ) ;
INV     gate8479  (.A(g12302), .Z(g15440) ) ;
NOR3    gate8480  (.A(g10729), .B(g10748), .C(g10764), .Z(g12418) ) ;
INV     gate8481  (.A(g12418), .Z(g15441) ) ;
NAND2   gate8482  (.A(g9968), .B(g3834), .Z(g11700) ) ;
INV     gate8483  (.A(g11700), .Z(II21705) ) ;
INV     gate8484  (.A(II21705), .Z(g15443) ) ;
NAND2   gate8485  (.A(g9968), .B(g7488), .Z(g13081) ) ;
INV     gate8486  (.A(g13081), .Z(II21708) ) ;
INV     gate8487  (.A(II21708), .Z(g15446) ) ;
NAND2   gate8488  (.A(g9968), .B(g7426), .Z(g13108) ) ;
INV     gate8489  (.A(g13108), .Z(II21711) ) ;
INV     gate8490  (.A(II21711), .Z(g15449) ) ;
INV     gate8491  (.A(g12312), .Z(g15458) ) ;
NAND2   gate8492  (.A(g9534), .B(g3366), .Z(g11701) ) ;
INV     gate8493  (.A(g11701), .Z(II21720) ) ;
INV     gate8494  (.A(II21720), .Z(g15461) ) ;
NAND2   gate8495  (.A(g9534), .B(g6912), .Z(g13088) ) ;
INV     gate8496  (.A(g13088), .Z(II21723) ) ;
INV     gate8497  (.A(II21723), .Z(g15464) ) ;
NAND2   gate8498  (.A(g9534), .B(g6678), .Z(g13112) ) ;
INV     gate8499  (.A(g13112), .Z(II21726) ) ;
INV     gate8500  (.A(II21726), .Z(g15467) ) ;
NAND2   gate8501  (.A(g9534), .B(g6912), .Z(g13089) ) ;
INV     gate8502  (.A(g13089), .Z(II21730) ) ;
INV     gate8503  (.A(II21730), .Z(g15471) ) ;
INV     gate8504  (.A(g12315), .Z(g15474) ) ;
NAND2   gate8505  (.A(g9676), .B(g3522), .Z(g11702) ) ;
INV     gate8506  (.A(g11702), .Z(II21736) ) ;
INV     gate8507  (.A(II21736), .Z(g15477) ) ;
NAND2   gate8508  (.A(g9676), .B(g7162), .Z(g13091) ) ;
INV     gate8509  (.A(g13091), .Z(II21739) ) ;
INV     gate8510  (.A(II21739), .Z(g15480) ) ;
NAND2   gate8511  (.A(g9676), .B(g6980), .Z(g13114) ) ;
INV     gate8512  (.A(g13114), .Z(II21742) ) ;
INV     gate8513  (.A(II21742), .Z(g15483) ) ;
NAND2   gate8514  (.A(g9676), .B(g6980), .Z(g13116) ) ;
INV     gate8515  (.A(g13116), .Z(II21747) ) ;
INV     gate8516  (.A(II21747), .Z(g15488) ) ;
INV     gate8517  (.A(g12318), .Z(g15492) ) ;
INV     gate8518  (.A(g12321), .Z(g15493) ) ;
NAND2   gate8519  (.A(g9822), .B(g3678), .Z(g11704) ) ;
INV     gate8520  (.A(g11704), .Z(II21755) ) ;
INV     gate8521  (.A(II21755), .Z(g15496) ) ;
NAND2   gate8522  (.A(g9822), .B(g7358), .Z(g13094) ) ;
INV     gate8523  (.A(g13094), .Z(II21758) ) ;
INV     gate8524  (.A(II21758), .Z(g15499) ) ;
NAND2   gate8525  (.A(g9822), .B(g7230), .Z(g13118) ) ;
INV     gate8526  (.A(g13118), .Z(II21761) ) ;
INV     gate8527  (.A(II21761), .Z(g15502) ) ;
NAND2   gate8528  (.A(g9968), .B(g3834), .Z(g11705) ) ;
INV     gate8529  (.A(g11705), .Z(II21769) ) ;
INV     gate8530  (.A(II21769), .Z(g15510) ) ;
NAND2   gate8531  (.A(g9968), .B(g7488), .Z(g13097) ) ;
INV     gate8532  (.A(g13097), .Z(II21772) ) ;
INV     gate8533  (.A(II21772), .Z(g15513) ) ;
NAND2   gate8534  (.A(g9968), .B(g7426), .Z(g13121) ) ;
INV     gate8535  (.A(g13121), .Z(II21775) ) ;
INV     gate8536  (.A(II21775), .Z(g15516) ) ;
NAND2   gate8537  (.A(g8317), .B(g2993), .Z(g13305) ) ;
INV     gate8538  (.A(g13305), .Z(II21780) ) ;
INV     gate8539  (.A(II21780), .Z(g15521) ) ;
INV     gate8540  (.A(g12333), .Z(g15524) ) ;
INV     gate8541  (.A(g12336), .Z(g15525) ) ;
NAND2   gate8542  (.A(g9534), .B(g3366), .Z(g11707) ) ;
INV     gate8543  (.A(g11707), .Z(II21787) ) ;
INV     gate8544  (.A(II21787), .Z(g15528) ) ;
NAND2   gate8545  (.A(g9534), .B(g6912), .Z(g13099) ) ;
INV     gate8546  (.A(g13099), .Z(II21790) ) ;
INV     gate8547  (.A(II21790), .Z(g15531) ) ;
NAND2   gate8548  (.A(g9534), .B(g6678), .Z(g13123) ) ;
INV     gate8549  (.A(g13123), .Z(II21793) ) ;
INV     gate8550  (.A(II21793), .Z(g15534) ) ;
NAND2   gate8551  (.A(g9534), .B(g3366), .Z(g11708) ) ;
INV     gate8552  (.A(g11708), .Z(II21796) ) ;
INV     gate8553  (.A(II21796), .Z(g15537) ) ;
INV     gate8554  (.A(g12340), .Z(g15544) ) ;
NAND2   gate8555  (.A(g9676), .B(g3522), .Z(g11709) ) ;
INV     gate8556  (.A(g11709), .Z(II21803) ) ;
INV     gate8557  (.A(II21803), .Z(g15547) ) ;
NAND2   gate8558  (.A(g9676), .B(g7162), .Z(g13103) ) ;
INV     gate8559  (.A(g13103), .Z(II21806) ) ;
INV     gate8560  (.A(II21806), .Z(g15550) ) ;
NAND2   gate8561  (.A(g9676), .B(g6980), .Z(g13125) ) ;
INV     gate8562  (.A(g13125), .Z(II21809) ) ;
INV     gate8563  (.A(II21809), .Z(g15553) ) ;
NAND2   gate8564  (.A(g9676), .B(g7162), .Z(g13104) ) ;
INV     gate8565  (.A(g13104), .Z(II21813) ) ;
INV     gate8566  (.A(II21813), .Z(g15557) ) ;
INV     gate8567  (.A(g12343), .Z(g15560) ) ;
NAND2   gate8568  (.A(g9822), .B(g3678), .Z(g11710) ) ;
INV     gate8569  (.A(g11710), .Z(II21819) ) ;
INV     gate8570  (.A(II21819), .Z(g15563) ) ;
NAND2   gate8571  (.A(g9822), .B(g7358), .Z(g13106) ) ;
INV     gate8572  (.A(g13106), .Z(II21822) ) ;
INV     gate8573  (.A(II21822), .Z(g15566) ) ;
NAND2   gate8574  (.A(g9822), .B(g7230), .Z(g13127) ) ;
INV     gate8575  (.A(g13127), .Z(II21825) ) ;
INV     gate8576  (.A(II21825), .Z(g15569) ) ;
NAND2   gate8577  (.A(g9822), .B(g7230), .Z(g13129) ) ;
INV     gate8578  (.A(g13129), .Z(II21830) ) ;
INV     gate8579  (.A(II21830), .Z(g15574) ) ;
INV     gate8580  (.A(g12346), .Z(g15578) ) ;
INV     gate8581  (.A(g12349), .Z(g15579) ) ;
NAND2   gate8582  (.A(g9968), .B(g3834), .Z(g11712) ) ;
INV     gate8583  (.A(g11712), .Z(II21838) ) ;
INV     gate8584  (.A(II21838), .Z(g15582) ) ;
NAND2   gate8585  (.A(g9968), .B(g7488), .Z(g13109) ) ;
INV     gate8586  (.A(g13109), .Z(II21841) ) ;
INV     gate8587  (.A(II21841), .Z(g15585) ) ;
NAND2   gate8588  (.A(g9968), .B(g7426), .Z(g13131) ) ;
INV     gate8589  (.A(g13131), .Z(II21844) ) ;
INV     gate8590  (.A(II21844), .Z(g15588) ) ;
NAND2   gate8591  (.A(g9534), .B(g3366), .Z(g11716) ) ;
INV     gate8592  (.A(g11716), .Z(II21852) ) ;
INV     gate8593  (.A(II21852), .Z(g15596) ) ;
NAND2   gate8594  (.A(g9534), .B(g6912), .Z(g13113) ) ;
INV     gate8595  (.A(g13113), .Z(II21855) ) ;
INV     gate8596  (.A(II21855), .Z(g15599) ) ;
INV     gate8597  (.A(g12363), .Z(g15602) ) ;
INV     gate8598  (.A(g12366), .Z(g15603) ) ;
NAND2   gate8599  (.A(g9676), .B(g3522), .Z(g11717) ) ;
INV     gate8600  (.A(g11717), .Z(II21862) ) ;
INV     gate8601  (.A(II21862), .Z(g15606) ) ;
NAND2   gate8602  (.A(g9676), .B(g7162), .Z(g13115) ) ;
INV     gate8603  (.A(g13115), .Z(II21865) ) ;
INV     gate8604  (.A(II21865), .Z(g15609) ) ;
NAND2   gate8605  (.A(g9676), .B(g6980), .Z(g13134) ) ;
INV     gate8606  (.A(g13134), .Z(II21868) ) ;
INV     gate8607  (.A(II21868), .Z(g15612) ) ;
NAND2   gate8608  (.A(g9676), .B(g3522), .Z(g11718) ) ;
INV     gate8609  (.A(g11718), .Z(II21871) ) ;
INV     gate8610  (.A(II21871), .Z(g15615) ) ;
INV     gate8611  (.A(g12370), .Z(g15622) ) ;
NAND2   gate8612  (.A(g9822), .B(g3678), .Z(g11719) ) ;
INV     gate8613  (.A(g11719), .Z(II21878) ) ;
INV     gate8614  (.A(II21878), .Z(g15625) ) ;
NAND2   gate8615  (.A(g9822), .B(g7358), .Z(g13119) ) ;
INV     gate8616  (.A(g13119), .Z(II21881) ) ;
INV     gate8617  (.A(II21881), .Z(g15628) ) ;
NAND2   gate8618  (.A(g9822), .B(g7230), .Z(g13136) ) ;
INV     gate8619  (.A(g13136), .Z(II21884) ) ;
INV     gate8620  (.A(II21884), .Z(g15631) ) ;
NAND2   gate8621  (.A(g9822), .B(g7358), .Z(g13120) ) ;
INV     gate8622  (.A(g13120), .Z(II21888) ) ;
INV     gate8623  (.A(II21888), .Z(g15635) ) ;
INV     gate8624  (.A(g12373), .Z(g15638) ) ;
NAND2   gate8625  (.A(g9968), .B(g3834), .Z(g11720) ) ;
INV     gate8626  (.A(g11720), .Z(II21894) ) ;
INV     gate8627  (.A(II21894), .Z(g15641) ) ;
NAND2   gate8628  (.A(g9968), .B(g7488), .Z(g13122) ) ;
INV     gate8629  (.A(g13122), .Z(II21897) ) ;
INV     gate8630  (.A(II21897), .Z(g15644) ) ;
NAND2   gate8631  (.A(g9968), .B(g7426), .Z(g13138) ) ;
INV     gate8632  (.A(g13138), .Z(II21900) ) ;
INV     gate8633  (.A(II21900), .Z(g15647) ) ;
NAND2   gate8634  (.A(g9968), .B(g7426), .Z(g13140) ) ;
INV     gate8635  (.A(g13140), .Z(II21905) ) ;
INV     gate8636  (.A(II21905), .Z(g15652) ) ;
AND2    gate8637  (.A(II20131), .B(II20132), .Z(g13082) ) ;
INV     gate8638  (.A(g13082), .Z(II21908) ) ;
INV     gate8639  (.A(II21908), .Z(g15655) ) ;
INV     gate8640  (.A(g11706), .Z(g15659) ) ;
INV     gate8641  (.A(g12379), .Z(g15665) ) ;
NAND2   gate8642  (.A(g9534), .B(g3366), .Z(g11721) ) ;
INV     gate8643  (.A(g11721), .Z(II21918) ) ;
INV     gate8644  (.A(II21918), .Z(g15667) ) ;
NAND2   gate8645  (.A(g9676), .B(g3522), .Z(g11722) ) ;
INV     gate8646  (.A(g11722), .Z(II21923) ) ;
INV     gate8647  (.A(II21923), .Z(g15672) ) ;
NAND2   gate8648  (.A(g9676), .B(g7162), .Z(g13126) ) ;
INV     gate8649  (.A(g13126), .Z(II21926) ) ;
INV     gate8650  (.A(II21926), .Z(g15675) ) ;
INV     gate8651  (.A(g12382), .Z(g15678) ) ;
INV     gate8652  (.A(g12385), .Z(g15679) ) ;
NAND2   gate8653  (.A(g9822), .B(g3678), .Z(g11723) ) ;
INV     gate8654  (.A(g11723), .Z(II21933) ) ;
INV     gate8655  (.A(II21933), .Z(g15682) ) ;
NAND2   gate8656  (.A(g9822), .B(g7358), .Z(g13128) ) ;
INV     gate8657  (.A(g13128), .Z(II21936) ) ;
INV     gate8658  (.A(II21936), .Z(g15685) ) ;
NAND2   gate8659  (.A(g9822), .B(g7230), .Z(g13142) ) ;
INV     gate8660  (.A(g13142), .Z(II21939) ) ;
INV     gate8661  (.A(II21939), .Z(g15688) ) ;
NAND2   gate8662  (.A(g9822), .B(g3678), .Z(g11724) ) ;
INV     gate8663  (.A(g11724), .Z(II21942) ) ;
INV     gate8664  (.A(II21942), .Z(g15691) ) ;
INV     gate8665  (.A(g12389), .Z(g15698) ) ;
NAND2   gate8666  (.A(g9968), .B(g3834), .Z(g11725) ) ;
INV     gate8667  (.A(g11725), .Z(II21949) ) ;
INV     gate8668  (.A(II21949), .Z(g15701) ) ;
NAND2   gate8669  (.A(g9968), .B(g7488), .Z(g13132) ) ;
INV     gate8670  (.A(g13132), .Z(II21952) ) ;
INV     gate8671  (.A(II21952), .Z(g15704) ) ;
NAND2   gate8672  (.A(g9968), .B(g7426), .Z(g13144) ) ;
INV     gate8673  (.A(g13144), .Z(II21955) ) ;
INV     gate8674  (.A(II21955), .Z(g15707) ) ;
NAND2   gate8675  (.A(g9968), .B(g7488), .Z(g13133) ) ;
INV     gate8676  (.A(g13133), .Z(II21959) ) ;
INV     gate8677  (.A(II21959), .Z(g15711) ) ;
AND2    gate8678  (.A(g10186), .B(g8317), .Z(g13004) ) ;
INV     gate8679  (.A(g13004), .Z(II21962) ) ;
INV     gate8680  (.A(II21962), .Z(g15714) ) ;
INV     gate8681  (.A(g13011), .Z(g15722) ) ;
INV     gate8682  (.A(g12409), .Z(g15724) ) ;
NAND2   gate8683  (.A(g9676), .B(g3522), .Z(g11726) ) ;
INV     gate8684  (.A(g11726), .Z(II21974) ) ;
INV     gate8685  (.A(II21974), .Z(g15726) ) ;
NAND2   gate8686  (.A(g9822), .B(g3678), .Z(g11727) ) ;
INV     gate8687  (.A(g11727), .Z(II21979) ) ;
INV     gate8688  (.A(II21979), .Z(g15731) ) ;
NAND2   gate8689  (.A(g9822), .B(g7358), .Z(g13137) ) ;
INV     gate8690  (.A(g13137), .Z(II21982) ) ;
INV     gate8691  (.A(II21982), .Z(g15734) ) ;
INV     gate8692  (.A(g12412), .Z(g15737) ) ;
INV     gate8693  (.A(g12415), .Z(g15738) ) ;
NAND2   gate8694  (.A(g9968), .B(g3834), .Z(g11728) ) ;
INV     gate8695  (.A(g11728), .Z(II21989) ) ;
INV     gate8696  (.A(II21989), .Z(g15741) ) ;
NAND2   gate8697  (.A(g9968), .B(g7488), .Z(g13139) ) ;
INV     gate8698  (.A(g13139), .Z(II21992) ) ;
INV     gate8699  (.A(II21992), .Z(g15744) ) ;
NAND2   gate8700  (.A(g9968), .B(g7426), .Z(g13146) ) ;
INV     gate8701  (.A(g13146), .Z(II21995) ) ;
INV     gate8702  (.A(II21995), .Z(g15747) ) ;
NAND2   gate8703  (.A(g9968), .B(g3834), .Z(g11729) ) ;
INV     gate8704  (.A(g11729), .Z(II21998) ) ;
INV     gate8705  (.A(II21998), .Z(g15750) ) ;
INV     gate8706  (.A(g13011), .Z(g15762) ) ;
INV     gate8707  (.A(g12421), .Z(g15764) ) ;
NAND2   gate8708  (.A(g9822), .B(g3678), .Z(g11730) ) ;
INV     gate8709  (.A(g11730), .Z(II22014) ) ;
INV     gate8710  (.A(II22014), .Z(g15766) ) ;
NAND2   gate8711  (.A(g9968), .B(g3834), .Z(g11731) ) ;
INV     gate8712  (.A(g11731), .Z(II22019) ) ;
INV     gate8713  (.A(II22019), .Z(g15771) ) ;
NAND2   gate8714  (.A(g9968), .B(g7488), .Z(g13145) ) ;
INV     gate8715  (.A(g13145), .Z(II22022) ) ;
INV     gate8716  (.A(II22022), .Z(g15774) ) ;
NAND2   gate8717  (.A(g8313), .B(g2883), .Z(g11617) ) ;
INV     gate8718  (.A(g11617), .Z(II22025) ) ;
INV     gate8719  (.A(II22025), .Z(g15777) ) ;
INV     gate8720  (.A(g13011), .Z(g15790) ) ;
INV     gate8721  (.A(g12426), .Z(g15792) ) ;
NAND2   gate8722  (.A(g9968), .B(g3834), .Z(g11733) ) ;
INV     gate8723  (.A(g11733), .Z(II22044) ) ;
INV     gate8724  (.A(II22044), .Z(g15794) ) ;
INV     gate8725  (.A(g12909), .Z(g15800) ) ;
INV     gate8726  (.A(g13011), .Z(g15813) ) ;
INV     gate8727  (.A(g13378), .Z(g15859) ) ;
INV     gate8728  (.A(g12909), .Z(II22120) ) ;
INV     gate8729  (.A(II22120), .Z(g15876) ) ;
INV     gate8730  (.A(g11624), .Z(g15880) ) ;
INV     gate8731  (.A(g11600), .Z(g15890) ) ;
INV     gate8732  (.A(g11644), .Z(g15904) ) ;
INV     gate8733  (.A(g11647), .Z(g15913) ) ;
INV     gate8734  (.A(g11630), .Z(g15923) ) ;
INV     gate8735  (.A(g11663), .Z(g15933) ) ;
INV     gate8736  (.A(g11666), .Z(g15942) ) ;
INV     gate8737  (.A(g11653), .Z(g15952) ) ;
INV     gate8738  (.A(g11675), .Z(g15962) ) ;
INV     gate8739  (.A(g11678), .Z(g15971) ) ;
INV     gate8740  (.A(g11687), .Z(g15981) ) ;
NAND2   gate8741  (.A(g2879), .B(g10778), .Z(g12433) ) ;
INV     gate8742  (.A(g12433), .Z(II22163) ) ;
INV     gate8743  (.A(II22163), .Z(g15989) ) ;
INV     gate8744  (.A(g12548), .Z(g15991) ) ;
INV     gate8745  (.A(g12555), .Z(g15994) ) ;
INV     gate8746  (.A(g12561), .Z(g15997) ) ;
INV     gate8747  (.A(g12601), .Z(g16001) ) ;
INV     gate8748  (.A(g12604), .Z(g16002) ) ;
INV     gate8749  (.A(g12608), .Z(g16005) ) ;
INV     gate8750  (.A(g12647), .Z(g16007) ) ;
INV     gate8751  (.A(g12651), .Z(g16011) ) ;
INV     gate8752  (.A(g12654), .Z(g16012) ) ;
INV     gate8753  (.A(g12692), .Z(g16013) ) ;
INV     gate8754  (.A(g12695), .Z(g16014) ) ;
INV     gate8755  (.A(g12699), .Z(g16023) ) ;
INV     gate8756  (.A(g12702), .Z(g16024) ) ;
INV     gate8757  (.A(g12705), .Z(g16025) ) ;
INV     gate8758  (.A(g12708), .Z(g16026) ) ;
INV     gate8759  (.A(g12744), .Z(g16027) ) ;
INV     gate8760  (.A(g12749), .Z(g16034) ) ;
INV     gate8761  (.A(g12752), .Z(g16035) ) ;
INV     gate8762  (.A(g12756), .Z(g16039) ) ;
INV     gate8763  (.A(g12759), .Z(g16040) ) ;
INV     gate8764  (.A(g12762), .Z(g16041) ) ;
INV     gate8765  (.A(g12765), .Z(g16042) ) ;
INV     gate8766  (.A(g12769), .Z(g16043) ) ;
INV     gate8767  (.A(g12772), .Z(g16044) ) ;
INV     gate8768  (.A(g12783), .Z(g16054) ) ;
INV     gate8769  (.A(g12786), .Z(g16055) ) ;
INV     gate8770  (.A(g12791), .Z(g16056) ) ;
INV     gate8771  (.A(g12794), .Z(g16057) ) ;
INV     gate8772  (.A(g12798), .Z(g16061) ) ;
INV     gate8773  (.A(g12801), .Z(g16062) ) ;
INV     gate8774  (.A(g12804), .Z(g16063) ) ;
INV     gate8775  (.A(g12808), .Z(g16064) ) ;
INV     gate8776  (.A(g12811), .Z(g16065) ) ;
NOR3    gate8777  (.A(g9766), .B(g9894), .C(g10013), .Z(g11861) ) ;
INV     gate8778  (.A(g11861), .Z(g16075) ) ;
INV     gate8779  (.A(g12816), .Z(g16088) ) ;
INV     gate8780  (.A(g12822), .Z(g16090) ) ;
INV     gate8781  (.A(g12825), .Z(g16091) ) ;
INV     gate8782  (.A(g12830), .Z(g16092) ) ;
INV     gate8783  (.A(g12833), .Z(g16093) ) ;
INV     gate8784  (.A(g12837), .Z(g16097) ) ;
INV     gate8785  (.A(g12840), .Z(g16098) ) ;
INV     gate8786  (.A(g12844), .Z(g16099) ) ;
NOR3    gate8787  (.A(g9912), .B(g10048), .C(g10122), .Z(g11903) ) ;
INV     gate8788  (.A(g11903), .Z(g16113) ) ;
INV     gate8789  (.A(g12854), .Z(g16126) ) ;
INV     gate8790  (.A(g12860), .Z(g16128) ) ;
INV     gate8791  (.A(g12863), .Z(g16129) ) ;
INV     gate8792  (.A(g12868), .Z(g16130) ) ;
INV     gate8793  (.A(g12871), .Z(g16131) ) ;
INV     gate8794  (.A(g13057), .Z(g16142) ) ;
NOR3    gate8795  (.A(g10434), .B(g10494), .C(g10556), .Z(g12194) ) ;
INV     gate8796  (.A(g12194), .Z(g16154) ) ;
NOR3    gate8797  (.A(g10066), .B(g10157), .C(g10227), .Z(g11953) ) ;
INV     gate8798  (.A(g11953), .Z(g16164) ) ;
INV     gate8799  (.A(g12895), .Z(g16177) ) ;
INV     gate8800  (.A(g12901), .Z(g16179) ) ;
INV     gate8801  (.A(g12904), .Z(g16180) ) ;
INV     gate8802  (.A(g13043), .Z(g16189) ) ;
INV     gate8803  (.A(g13073), .Z(g16201) ) ;
NOR3    gate8804  (.A(g10510), .B(g10568), .C(g10613), .Z(g12249) ) ;
INV     gate8805  (.A(g12249), .Z(g16213) ) ;
NOR3    gate8806  (.A(g10175), .B(g10262), .C(g10329), .Z(g12006) ) ;
INV     gate8807  (.A(g12006), .Z(g16223) ) ;
INV     gate8808  (.A(g12935), .Z(g16236) ) ;
INV     gate8809  (.A(g13033), .Z(g16243) ) ;
INV     gate8810  (.A(g13060), .Z(g16254) ) ;
INV     gate8811  (.A(g13092), .Z(g16266) ) ;
NOR3    gate8812  (.A(g10584), .B(g10625), .C(g10660), .Z(g12292) ) ;
INV     gate8813  (.A(g12292), .Z(g16278) ) ;
INV     gate8814  (.A(g12962), .Z(g16287) ) ;
INV     gate8815  (.A(g13025), .Z(g16293) ) ;
INV     gate8816  (.A(g520), .Z(II22382) ) ;
INV     gate8817  (.A(g13046), .Z(g16302) ) ;
INV     gate8818  (.A(g13076), .Z(g16313) ) ;
INV     gate8819  (.A(g13107), .Z(g16325) ) ;
NOR3    gate8820  (.A(g10641), .B(g10672), .C(g10690), .Z(g12328) ) ;
INV     gate8821  (.A(g12328), .Z(g16337) ) ;
INV     gate8822  (.A(g13036), .Z(g16351) ) ;
INV     gate8823  (.A(g1206), .Z(II22414) ) ;
INV     gate8824  (.A(g13063), .Z(g16360) ) ;
INV     gate8825  (.A(g13095), .Z(g16371) ) ;
INV     gate8826  (.A(g13049), .Z(g16395) ) ;
INV     gate8827  (.A(g1900), .Z(II22444) ) ;
INV     gate8828  (.A(g13079), .Z(g16404) ) ;
INV     gate8829  (.A(g13066), .Z(g16433) ) ;
INV     gate8830  (.A(g2594), .Z(II22475) ) ;
INV     gate8831  (.A(g12017), .Z(g16466) ) ;
INV     gate8832  (.A(g13598), .Z(II22503) ) ;
INV     gate8833  (.A(g13624), .Z(II22506) ) ;
INV     gate8834  (.A(g13610), .Z(II22509) ) ;
INV     gate8835  (.A(g13635), .Z(II22512) ) ;
INV     gate8836  (.A(g13620), .Z(II22515) ) ;
INV     gate8837  (.A(g13647), .Z(II22518) ) ;
INV     gate8838  (.A(g13632), .Z(II22521) ) ;
INV     gate8839  (.A(g13673), .Z(II22524) ) ;
INV     gate8840  (.A(g13469), .Z(II22527) ) ;
INV     gate8841  (.A(g14774), .Z(II22530) ) ;
INV     gate8842  (.A(g14795), .Z(II22533) ) ;
INV     gate8843  (.A(g14829), .Z(II22536) ) ;
INV     gate8844  (.A(g14882), .Z(II22539) ) ;
INV     gate8845  (.A(g14954), .Z(II22542) ) ;
INV     gate8846  (.A(g15018), .Z(II22545) ) ;
INV     gate8847  (.A(g14718), .Z(II22548) ) ;
INV     gate8848  (.A(g14745), .Z(II22551) ) ;
INV     gate8849  (.A(g14765), .Z(II22554) ) ;
INV     gate8850  (.A(g14775), .Z(II22557) ) ;
INV     gate8851  (.A(g14796), .Z(II22560) ) ;
INV     gate8852  (.A(g14830), .Z(II22563) ) ;
INV     gate8853  (.A(g14883), .Z(II22566) ) ;
INV     gate8854  (.A(g14955), .Z(II22569) ) ;
INV     gate8855  (.A(g15019), .Z(II22572) ) ;
INV     gate8856  (.A(g15092), .Z(II22575) ) ;
INV     gate8857  (.A(g14746), .Z(II22578) ) ;
INV     gate8858  (.A(g14766), .Z(II22581) ) ;
INV     gate8859  (.A(g15989), .Z(II22584) ) ;
INV     gate8860  (.A(g14684), .Z(II22587) ) ;
INV     gate8861  (.A(g13863), .Z(II22590) ) ;
INV     gate8862  (.A(g15876), .Z(II22593) ) ;
INV     gate8863  (.A(g14158), .Z(g16501) ) ;
INV     gate8864  (.A(g14966), .Z(II22599) ) ;
INV     gate8865  (.A(II22599), .Z(g16506) ) ;
INV     gate8866  (.A(g14186), .Z(g16507) ) ;
INV     gate8867  (.A(g15080), .Z(II22604) ) ;
INV     gate8868  (.A(II22604), .Z(g16514) ) ;
INV     gate8869  (.A(g14244), .Z(g16515) ) ;
INV     gate8870  (.A(g14273), .Z(g16523) ) ;
INV     gate8871  (.A(g15055), .Z(II22611) ) ;
INV     gate8872  (.A(II22611), .Z(g16528) ) ;
INV     gate8873  (.A(g14301), .Z(g16529) ) ;
INV     gate8874  (.A(g14630), .Z(II22618) ) ;
INV     gate8875  (.A(II22618), .Z(g16540) ) ;
INV     gate8876  (.A(g14347), .Z(g16543) ) ;
INV     gate8877  (.A(g14366), .Z(g16546) ) ;
INV     gate8878  (.A(g14395), .Z(g16554) ) ;
INV     gate8879  (.A(g15151), .Z(II22626) ) ;
INV     gate8880  (.A(II22626), .Z(g16559) ) ;
INV     gate8881  (.A(g14423), .Z(g16560) ) ;
INV     gate8882  (.A(g14650), .Z(II22640) ) ;
INV     gate8883  (.A(II22640), .Z(g16572) ) ;
INV     gate8884  (.A(g14459), .Z(g16575) ) ;
INV     gate8885  (.A(g14478), .Z(g16578) ) ;
INV     gate8886  (.A(g14507), .Z(g16586) ) ;
INV     gate8887  (.A(g14677), .Z(II22651) ) ;
INV     gate8888  (.A(II22651), .Z(g16596) ) ;
INV     gate8889  (.A(g14546), .Z(g16599) ) ;
INV     gate8890  (.A(g14565), .Z(g16602) ) ;
INV     gate8891  (.A(g14657), .Z(II22657) ) ;
INV     gate8892  (.A(II22657), .Z(g16608) ) ;
INV     gate8893  (.A(g14711), .Z(II22663) ) ;
INV     gate8894  (.A(II22663), .Z(g16616) ) ;
INV     gate8895  (.A(g14601), .Z(g16619) ) ;
INV     gate8896  (.A(g14642), .Z(II22667) ) ;
INV     gate8897  (.A(II22667), .Z(g16622) ) ;
INV     gate8898  (.A(g14691), .Z(II22671) ) ;
INV     gate8899  (.A(II22671), .Z(g16626) ) ;
INV     gate8900  (.A(g14630), .Z(II22676) ) ;
INV     gate8901  (.A(II22676), .Z(g16633) ) ;
INV     gate8902  (.A(g14669), .Z(II22679) ) ;
INV     gate8903  (.A(II22679), .Z(g16636) ) ;
INV     gate8904  (.A(g14725), .Z(II22683) ) ;
INV     gate8905  (.A(II22683), .Z(g16640) ) ;
INV     gate8906  (.A(g14650), .Z(II22687) ) ;
INV     gate8907  (.A(II22687), .Z(g16644) ) ;
INV     gate8908  (.A(g14703), .Z(II22690) ) ;
INV     gate8909  (.A(II22690), .Z(g16647) ) ;
INV     gate8910  (.A(g14753), .Z(II22694) ) ;
INV     gate8911  (.A(II22694), .Z(g16651) ) ;
INV     gate8912  (.A(g14677), .Z(II22699) ) ;
INV     gate8913  (.A(II22699), .Z(g16656) ) ;
INV     gate8914  (.A(g14737), .Z(II22702) ) ;
INV     gate8915  (.A(II22702), .Z(g16659) ) ;
INV     gate8916  (.A(g14776), .Z(g16665) ) ;
INV     gate8917  (.A(g14711), .Z(II22715) ) ;
INV     gate8918  (.A(II22715), .Z(g16673) ) ;
INV     gate8919  (.A(g14657), .Z(II22718) ) ;
INV     gate8920  (.A(II22718), .Z(g16676) ) ;
INV     gate8921  (.A(g14797), .Z(g16682) ) ;
INV     gate8922  (.A(g14811), .Z(g16686) ) ;
INV     gate8923  (.A(g14642), .Z(II22726) ) ;
INV     gate8924  (.A(II22726), .Z(g16694) ) ;
INV     gate8925  (.A(g14837), .Z(g16697) ) ;
INV     gate8926  (.A(g14691), .Z(II22730) ) ;
INV     gate8927  (.A(II22730), .Z(g16702) ) ;
INV     gate8928  (.A(g14849), .Z(g16708) ) ;
INV     gate8929  (.A(g14863), .Z(g16712) ) ;
INV     gate8930  (.A(g14630), .Z(II22737) ) ;
INV     gate8931  (.A(II22737), .Z(g16719) ) ;
INV     gate8932  (.A(g14895), .Z(g16722) ) ;
INV     gate8933  (.A(g14669), .Z(II22741) ) ;
INV     gate8934  (.A(II22741), .Z(g16725) ) ;
INV     gate8935  (.A(g14910), .Z(g16728) ) ;
INV     gate8936  (.A(g14725), .Z(II22745) ) ;
INV     gate8937  (.A(II22745), .Z(g16733) ) ;
INV     gate8938  (.A(g14922), .Z(g16739) ) ;
INV     gate8939  (.A(g14936), .Z(g16743) ) ;
NAND2   gate8940  (.A(g13332), .B(g12354), .Z(g15782) ) ;
INV     gate8941  (.A(g15782), .Z(g16749) ) ;
INV     gate8942  (.A(g14657), .Z(II22752) ) ;
INV     gate8943  (.A(II22752), .Z(g16758) ) ;
INV     gate8944  (.A(g14650), .Z(II22755) ) ;
INV     gate8945  (.A(II22755), .Z(g16761) ) ;
INV     gate8946  (.A(g14976), .Z(g16764) ) ;
INV     gate8947  (.A(g14703), .Z(II22759) ) ;
INV     gate8948  (.A(II22759), .Z(g16767) ) ;
INV     gate8949  (.A(g14991), .Z(g16770) ) ;
INV     gate8950  (.A(g14753), .Z(II22763) ) ;
INV     gate8951  (.A(II22763), .Z(g16775) ) ;
INV     gate8952  (.A(g15003), .Z(g16781) ) ;
INV     gate8953  (.A(g14691), .Z(II22768) ) ;
INV     gate8954  (.A(II22768), .Z(g16785) ) ;
INV     gate8955  (.A(g14677), .Z(II22771) ) ;
INV     gate8956  (.A(II22771), .Z(g16788) ) ;
INV     gate8957  (.A(g15065), .Z(g16791) ) ;
INV     gate8958  (.A(g14737), .Z(II22775) ) ;
INV     gate8959  (.A(II22775), .Z(g16794) ) ;
INV     gate8960  (.A(g15080), .Z(g16797) ) ;
NAND2   gate8961  (.A(g13375), .B(g12354), .Z(g15803) ) ;
INV     gate8962  (.A(g15803), .Z(g16804) ) ;
NAND2   gate8963  (.A(g13332), .B(g12392), .Z(g15842) ) ;
INV     gate8964  (.A(g15842), .Z(g16809) ) ;
INV     gate8965  (.A(g13572), .Z(II22783) ) ;
INV     gate8966  (.A(II22783), .Z(g16813) ) ;
INV     gate8967  (.A(g14725), .Z(II22786) ) ;
INV     gate8968  (.A(II22786), .Z(g16814) ) ;
INV     gate8969  (.A(g14711), .Z(II22789) ) ;
INV     gate8970  (.A(II22789), .Z(g16817) ) ;
INV     gate8971  (.A(g15161), .Z(g16820) ) ;
NAND2   gate8972  (.A(g13354), .B(g12392), .Z(g15855) ) ;
INV     gate8973  (.A(g15855), .Z(g16825) ) ;
INV     gate8974  (.A(g14165), .Z(II22797) ) ;
INV     gate8975  (.A(II22797), .Z(g16830) ) ;
INV     gate8976  (.A(g13581), .Z(II22800) ) ;
INV     gate8977  (.A(II22800), .Z(g16831) ) ;
INV     gate8978  (.A(g14753), .Z(II22803) ) ;
INV     gate8979  (.A(II22803), .Z(g16832) ) ;
NAND2   gate8980  (.A(g13024), .B(g12354), .Z(g15818) ) ;
INV     gate8981  (.A(g15818), .Z(g16836) ) ;
NAND2   gate8982  (.A(g13375), .B(g12392), .Z(g15878) ) ;
INV     gate8983  (.A(g15878), .Z(g16840) ) ;
INV     gate8984  (.A(g14280), .Z(II22810) ) ;
INV     gate8985  (.A(II22810), .Z(g16842) ) ;
INV     gate8986  (.A(g13601), .Z(II22813) ) ;
INV     gate8987  (.A(II22813), .Z(g16843) ) ;
NAND2   gate8988  (.A(g13404), .B(g12392), .Z(g15903) ) ;
INV     gate8989  (.A(g15903), .Z(g16846) ) ;
INV     gate8990  (.A(g14402), .Z(II22820) ) ;
INV     gate8991  (.A(II22820), .Z(g16848) ) ;
INV     gate8992  (.A(g13613), .Z(II22823) ) ;
INV     gate8993  (.A(II22823), .Z(g16849) ) ;
INV     gate8994  (.A(g14514), .Z(II22828) ) ;
INV     gate8995  (.A(II22828), .Z(g16852) ) ;
INV     gate8996  (.A(g13571), .Z(II22836) ) ;
INV     gate8997  (.A(II22836), .Z(g16858) ) ;
INV     gate8998  (.A(g13580), .Z(II22842) ) ;
INV     gate8999  (.A(II22842), .Z(g16862) ) ;
INV     gate9000  (.A(g13579), .Z(II22845) ) ;
INV     gate9001  (.A(II22845), .Z(g16863) ) ;
INV     gate9002  (.A(g13589), .Z(g16867) ) ;
INV     gate9003  (.A(g13600), .Z(II22852) ) ;
INV     gate9004  (.A(II22852), .Z(g16877) ) ;
INV     gate9005  (.A(g13588), .Z(II22855) ) ;
INV     gate9006  (.A(II22855), .Z(g16878) ) ;
INV     gate9007  (.A(g14885), .Z(II22860) ) ;
INV     gate9008  (.A(II22860), .Z(g16881) ) ;
INV     gate9009  (.A(g13589), .Z(g16884) ) ;
INV     gate9010  (.A(g13589), .Z(g16895) ) ;
INV     gate9011  (.A(g13612), .Z(II22866) ) ;
INV     gate9012  (.A(II22866), .Z(g16905) ) ;
INV     gate9013  (.A(g13608), .Z(II22869) ) ;
INV     gate9014  (.A(II22869), .Z(g16906) ) ;
INV     gate9015  (.A(g14966), .Z(II22875) ) ;
INV     gate9016  (.A(II22875), .Z(g16910) ) ;
INV     gate9017  (.A(g13589), .Z(g16913) ) ;
INV     gate9018  (.A(g13589), .Z(g16924) ) ;
INV     gate9019  (.A(g13622), .Z(II22881) ) ;
INV     gate9020  (.A(II22881), .Z(g16934) ) ;
INV     gate9021  (.A(g15055), .Z(II22893) ) ;
INV     gate9022  (.A(II22893), .Z(g16940) ) ;
INV     gate9023  (.A(g13589), .Z(g16943) ) ;
INV     gate9024  (.A(g13589), .Z(g16954) ) ;
INV     gate9025  (.A(g15151), .Z(II22912) ) ;
INV     gate9026  (.A(II22912), .Z(g16971) ) ;
INV     gate9027  (.A(g13589), .Z(g16974) ) ;
INV     gate9028  (.A(g14685), .Z(g17029) ) ;
INV     gate9029  (.A(g13519), .Z(g17057) ) ;
INV     gate9030  (.A(g14719), .Z(g17063) ) ;
INV     gate9031  (.A(g13530), .Z(g17092) ) ;
INV     gate9032  (.A(g14747), .Z(g17098) ) ;
INV     gate9033  (.A(g13541), .Z(g17130) ) ;
INV     gate9034  (.A(g14768), .Z(g17136) ) ;
INV     gate9035  (.A(g13552), .Z(g17157) ) ;
INV     gate9036  (.A(g13741), .Z(II23253) ) ;
INV     gate9037  (.A(II23253), .Z(g17189) ) ;
INV     gate9038  (.A(g13741), .Z(II23274) ) ;
INV     gate9039  (.A(II23274), .Z(g17200) ) ;
INV     gate9040  (.A(g13568), .Z(g17203) ) ;
INV     gate9041  (.A(g13741), .Z(II23287) ) ;
INV     gate9042  (.A(II23287), .Z(g17207) ) ;
INV     gate9043  (.A(g13576), .Z(g17208) ) ;
INV     gate9044  (.A(g13741), .Z(II23292) ) ;
INV     gate9045  (.A(II23292), .Z(g17212) ) ;
INV     gate9046  (.A(g13585), .Z(g17214) ) ;
INV     gate9047  (.A(g13605), .Z(g17217) ) ;
NAND2   gate9048  (.A(II22283), .B(II22284), .Z(g16132) ) ;
INV     gate9049  (.A(g16132), .Z(II23309) ) ;
INV     gate9050  (.A(II23309), .Z(g17227) ) ;
NAND2   gate9051  (.A(g12565), .B(g6232), .Z(g15720) ) ;
INV     gate9052  (.A(g15720), .Z(II23314) ) ;
INV     gate9053  (.A(II23314), .Z(g17230) ) ;
NAND2   gate9054  (.A(II22317), .B(II22318), .Z(g16181) ) ;
INV     gate9055  (.A(g16181), .Z(II23317) ) ;
INV     gate9056  (.A(II23317), .Z(g17233) ) ;
NAND2   gate9057  (.A(g12565), .B(g6314), .Z(g15664) ) ;
INV     gate9058  (.A(g15664), .Z(II23323) ) ;
INV     gate9059  (.A(II23323), .Z(g17237) ) ;
NAND2   gate9060  (.A(g12565), .B(g6232), .Z(g15758) ) ;
INV     gate9061  (.A(g15758), .Z(II23326) ) ;
INV     gate9062  (.A(II23326), .Z(g17240) ) ;
NAND2   gate9063  (.A(g12611), .B(g6369), .Z(g15760) ) ;
INV     gate9064  (.A(g15760), .Z(II23329) ) ;
INV     gate9065  (.A(II23329), .Z(g17243) ) ;
NAND2   gate9066  (.A(g12565), .B(g3254), .Z(g16412) ) ;
INV     gate9067  (.A(g16412), .Z(II23335) ) ;
INV     gate9068  (.A(II23335), .Z(g17249) ) ;
NAND2   gate9069  (.A(g12565), .B(g6314), .Z(g15721) ) ;
INV     gate9070  (.A(g15721), .Z(II23338) ) ;
INV     gate9071  (.A(II23338), .Z(g17252) ) ;
NAND2   gate9072  (.A(g12565), .B(g6232), .Z(g15784) ) ;
INV     gate9073  (.A(g15784), .Z(II23341) ) ;
INV     gate9074  (.A(II23341), .Z(g17255) ) ;
AND2    gate9075  (.A(g297), .B(g11770), .Z(g16053) ) ;
INV     gate9076  (.A(g16053), .Z(g17258) ) ;
NAND2   gate9077  (.A(g12611), .B(g6519), .Z(g15723) ) ;
INV     gate9078  (.A(g15723), .Z(II23345) ) ;
INV     gate9079  (.A(II23345), .Z(g17259) ) ;
NAND2   gate9080  (.A(g12611), .B(g6369), .Z(g15786) ) ;
INV     gate9081  (.A(g15786), .Z(II23348) ) ;
INV     gate9082  (.A(II23348), .Z(g17262) ) ;
NAND2   gate9083  (.A(g12657), .B(g6574), .Z(g15788) ) ;
INV     gate9084  (.A(g15788), .Z(II23351) ) ;
INV     gate9085  (.A(II23351), .Z(g17265) ) ;
NAND2   gate9086  (.A(g12565), .B(g3254), .Z(g16442) ) ;
INV     gate9087  (.A(g16442), .Z(II23358) ) ;
INV     gate9088  (.A(II23358), .Z(g17272) ) ;
NAND2   gate9089  (.A(g12565), .B(g6314), .Z(g15759) ) ;
INV     gate9090  (.A(g15759), .Z(II23361) ) ;
INV     gate9091  (.A(II23361), .Z(g17275) ) ;
NAND2   gate9092  (.A(g12565), .B(g6232), .Z(g15805) ) ;
INV     gate9093  (.A(g15805), .Z(II23364) ) ;
INV     gate9094  (.A(II23364), .Z(g17278) ) ;
AND2    gate9095  (.A(g3304), .B(g11783), .Z(g16081) ) ;
INV     gate9096  (.A(g16081), .Z(g17281) ) ;
NAND2   gate9097  (.A(g12611), .B(g3410), .Z(g16446) ) ;
INV     gate9098  (.A(g16446), .Z(II23368) ) ;
INV     gate9099  (.A(II23368), .Z(g17282) ) ;
NAND2   gate9100  (.A(g12611), .B(g6519), .Z(g15761) ) ;
INV     gate9101  (.A(g15761), .Z(II23371) ) ;
INV     gate9102  (.A(II23371), .Z(g17285) ) ;
NAND2   gate9103  (.A(g12611), .B(g6369), .Z(g15807) ) ;
INV     gate9104  (.A(g15807), .Z(II23374) ) ;
INV     gate9105  (.A(II23374), .Z(g17288) ) ;
NAND2   gate9106  (.A(g12657), .B(g6783), .Z(g15763) ) ;
INV     gate9107  (.A(g15763), .Z(II23377) ) ;
INV     gate9108  (.A(II23377), .Z(g17291) ) ;
NAND2   gate9109  (.A(g12657), .B(g6574), .Z(g15809) ) ;
INV     gate9110  (.A(g15809), .Z(II23380) ) ;
INV     gate9111  (.A(II23380), .Z(g17294) ) ;
NAND2   gate9112  (.A(g12711), .B(g6838), .Z(g15811) ) ;
INV     gate9113  (.A(g15811), .Z(II23383) ) ;
INV     gate9114  (.A(II23383), .Z(g17297) ) ;
INV     gate9115  (.A(g13469), .Z(II23386) ) ;
INV     gate9116  (.A(II23386), .Z(g17300) ) ;
NAND2   gate9117  (.A(g12565), .B(g3254), .Z(g13476) ) ;
INV     gate9118  (.A(g13476), .Z(II23392) ) ;
INV     gate9119  (.A(II23392), .Z(g17304) ) ;
NAND2   gate9120  (.A(g12565), .B(g6314), .Z(g15785) ) ;
INV     gate9121  (.A(g15785), .Z(II23395) ) ;
INV     gate9122  (.A(II23395), .Z(g17307) ) ;
NAND2   gate9123  (.A(g12565), .B(g6232), .Z(g15820) ) ;
INV     gate9124  (.A(g15820), .Z(II23398) ) ;
INV     gate9125  (.A(II23398), .Z(g17310) ) ;
AND2    gate9126  (.A(g8277), .B(g11803), .Z(g16109) ) ;
INV     gate9127  (.A(g16109), .Z(g17313) ) ;
AND2    gate9128  (.A(g516), .B(g11804), .Z(g16110) ) ;
INV     gate9129  (.A(g16110), .Z(g17314) ) ;
NAND2   gate9130  (.A(g12611), .B(g3410), .Z(g13478) ) ;
INV     gate9131  (.A(g13478), .Z(II23403) ) ;
INV     gate9132  (.A(II23403), .Z(g17315) ) ;
NAND2   gate9133  (.A(g12611), .B(g6519), .Z(g15787) ) ;
INV     gate9134  (.A(g15787), .Z(II23406) ) ;
INV     gate9135  (.A(II23406), .Z(g17318) ) ;
NAND2   gate9136  (.A(g12611), .B(g6369), .Z(g15822) ) ;
INV     gate9137  (.A(g15822), .Z(II23409) ) ;
INV     gate9138  (.A(II23409), .Z(g17321) ) ;
NAND2   gate9139  (.A(g12657), .B(g3566), .Z(g13482) ) ;
INV     gate9140  (.A(g13482), .Z(II23412) ) ;
INV     gate9141  (.A(II23412), .Z(g17324) ) ;
NAND2   gate9142  (.A(g12657), .B(g6783), .Z(g15789) ) ;
INV     gate9143  (.A(g15789), .Z(II23415) ) ;
INV     gate9144  (.A(II23415), .Z(g17327) ) ;
NAND2   gate9145  (.A(g12657), .B(g6574), .Z(g15824) ) ;
INV     gate9146  (.A(g15824), .Z(II23418) ) ;
INV     gate9147  (.A(II23418), .Z(g17330) ) ;
NAND2   gate9148  (.A(g12711), .B(g7085), .Z(g15791) ) ;
INV     gate9149  (.A(g15791), .Z(II23421) ) ;
INV     gate9150  (.A(II23421), .Z(g17333) ) ;
NAND2   gate9151  (.A(g12711), .B(g6838), .Z(g15826) ) ;
INV     gate9152  (.A(g15826), .Z(II23424) ) ;
INV     gate9153  (.A(II23424), .Z(g17336) ) ;
NAND2   gate9154  (.A(g12565), .B(g3254), .Z(g13494) ) ;
INV     gate9155  (.A(g13494), .Z(II23430) ) ;
INV     gate9156  (.A(II23430), .Z(g17342) ) ;
NAND2   gate9157  (.A(g12565), .B(g6314), .Z(g15806) ) ;
INV     gate9158  (.A(g15806), .Z(II23433) ) ;
INV     gate9159  (.A(II23433), .Z(g17345) ) ;
NAND2   gate9160  (.A(g12565), .B(g6232), .Z(g15832) ) ;
INV     gate9161  (.A(g15832), .Z(II23436) ) ;
INV     gate9162  (.A(II23436), .Z(g17348) ) ;
AND2    gate9163  (.A(g517), .B(g11829), .Z(g16152) ) ;
INV     gate9164  (.A(g16152), .Z(g17351) ) ;
NAND2   gate9165  (.A(g12611), .B(g3410), .Z(g13495) ) ;
INV     gate9166  (.A(g13495), .Z(II23442) ) ;
INV     gate9167  (.A(II23442), .Z(g17354) ) ;
NAND2   gate9168  (.A(g12611), .B(g6519), .Z(g15808) ) ;
INV     gate9169  (.A(g15808), .Z(II23445) ) ;
INV     gate9170  (.A(II23445), .Z(g17357) ) ;
NAND2   gate9171  (.A(g12611), .B(g6369), .Z(g15834) ) ;
INV     gate9172  (.A(g15834), .Z(II23448) ) ;
INV     gate9173  (.A(II23448), .Z(g17360) ) ;
NAND2   gate9174  (.A(g12657), .B(g3566), .Z(g13497) ) ;
INV     gate9175  (.A(g13497), .Z(II23451) ) ;
INV     gate9176  (.A(II23451), .Z(g17363) ) ;
NAND2   gate9177  (.A(g12657), .B(g6783), .Z(g15810) ) ;
INV     gate9178  (.A(g15810), .Z(II23454) ) ;
INV     gate9179  (.A(II23454), .Z(g17366) ) ;
NAND2   gate9180  (.A(g12657), .B(g6574), .Z(g15836) ) ;
INV     gate9181  (.A(g15836), .Z(II23457) ) ;
INV     gate9182  (.A(II23457), .Z(g17369) ) ;
NAND2   gate9183  (.A(g12711), .B(g3722), .Z(g13501) ) ;
INV     gate9184  (.A(g13501), .Z(II23460) ) ;
INV     gate9185  (.A(II23460), .Z(g17372) ) ;
NAND2   gate9186  (.A(g12711), .B(g7085), .Z(g15812) ) ;
INV     gate9187  (.A(g15812), .Z(II23463) ) ;
INV     gate9188  (.A(II23463), .Z(g17375) ) ;
NAND2   gate9189  (.A(g12711), .B(g6838), .Z(g15838) ) ;
INV     gate9190  (.A(g15838), .Z(II23466) ) ;
INV     gate9191  (.A(II23466), .Z(g17378) ) ;
NAND2   gate9192  (.A(g12565), .B(g3254), .Z(g13510) ) ;
INV     gate9193  (.A(g13510), .Z(II23472) ) ;
INV     gate9194  (.A(II23472), .Z(g17384) ) ;
NAND2   gate9195  (.A(g12565), .B(g6314), .Z(g15821) ) ;
INV     gate9196  (.A(g15821), .Z(II23475) ) ;
INV     gate9197  (.A(II23475), .Z(g17387) ) ;
NAND2   gate9198  (.A(g12565), .B(g6232), .Z(g15844) ) ;
INV     gate9199  (.A(g15844), .Z(II23478) ) ;
INV     gate9200  (.A(II23478), .Z(g17390) ) ;
AND2    gate9201  (.A(g518), .B(g11862), .Z(g16197) ) ;
INV     gate9202  (.A(g16197), .Z(g17394) ) ;
NAND2   gate9203  (.A(g12611), .B(g3410), .Z(g13511) ) ;
INV     gate9204  (.A(g13511), .Z(II23487) ) ;
INV     gate9205  (.A(II23487), .Z(g17399) ) ;
NAND2   gate9206  (.A(g12611), .B(g6519), .Z(g15823) ) ;
INV     gate9207  (.A(g15823), .Z(II23490) ) ;
INV     gate9208  (.A(II23490), .Z(g17402) ) ;
NAND2   gate9209  (.A(g12611), .B(g6369), .Z(g15846) ) ;
INV     gate9210  (.A(g15846), .Z(II23493) ) ;
INV     gate9211  (.A(II23493), .Z(g17405) ) ;
NAND2   gate9212  (.A(g12657), .B(g3566), .Z(g13512) ) ;
INV     gate9213  (.A(g13512), .Z(II23498) ) ;
INV     gate9214  (.A(II23498), .Z(g17410) ) ;
NAND2   gate9215  (.A(g12657), .B(g6783), .Z(g15825) ) ;
INV     gate9216  (.A(g15825), .Z(II23501) ) ;
INV     gate9217  (.A(II23501), .Z(g17413) ) ;
NAND2   gate9218  (.A(g12657), .B(g6574), .Z(g15848) ) ;
INV     gate9219  (.A(g15848), .Z(II23504) ) ;
INV     gate9220  (.A(II23504), .Z(g17416) ) ;
NAND2   gate9221  (.A(g12711), .B(g3722), .Z(g13514) ) ;
INV     gate9222  (.A(g13514), .Z(II23507) ) ;
INV     gate9223  (.A(II23507), .Z(g17419) ) ;
NAND2   gate9224  (.A(g12711), .B(g7085), .Z(g15827) ) ;
INV     gate9225  (.A(g15827), .Z(II23510) ) ;
INV     gate9226  (.A(II23510), .Z(g17422) ) ;
NAND2   gate9227  (.A(g12711), .B(g6838), .Z(g15850) ) ;
INV     gate9228  (.A(g15850), .Z(II23513) ) ;
INV     gate9229  (.A(II23513), .Z(g17425) ) ;
NAND2   gate9230  (.A(g12565), .B(g6232), .Z(g15856) ) ;
INV     gate9231  (.A(g15856), .Z(II23518) ) ;
INV     gate9232  (.A(II23518), .Z(g17430) ) ;
NAND2   gate9233  (.A(g12565), .B(g3254), .Z(g13518) ) ;
INV     gate9234  (.A(g13518), .Z(II23521) ) ;
INV     gate9235  (.A(II23521), .Z(g17433) ) ;
NAND2   gate9236  (.A(g12565), .B(g6314), .Z(g15833) ) ;
INV     gate9237  (.A(g15833), .Z(II23524) ) ;
INV     gate9238  (.A(II23524), .Z(g17436) ) ;
NAND2   gate9239  (.A(g12565), .B(g6232), .Z(g15858) ) ;
INV     gate9240  (.A(g15858), .Z(II23527) ) ;
INV     gate9241  (.A(II23527), .Z(g17439) ) ;
INV     gate9242  (.A(g14885), .Z(II23530) ) ;
INV     gate9243  (.A(II23530), .Z(g17442) ) ;
AND2    gate9244  (.A(g519), .B(g11895), .Z(g16250) ) ;
INV     gate9245  (.A(g16250), .Z(g17445) ) ;
NAND2   gate9246  (.A(g12611), .B(g3410), .Z(g13524) ) ;
INV     gate9247  (.A(g13524), .Z(II23539) ) ;
INV     gate9248  (.A(II23539), .Z(g17451) ) ;
NAND2   gate9249  (.A(g12611), .B(g6519), .Z(g15835) ) ;
INV     gate9250  (.A(g15835), .Z(II23542) ) ;
INV     gate9251  (.A(II23542), .Z(g17454) ) ;
NAND2   gate9252  (.A(g12611), .B(g6369), .Z(g15867) ) ;
INV     gate9253  (.A(g15867), .Z(II23545) ) ;
INV     gate9254  (.A(II23545), .Z(g17457) ) ;
NAND2   gate9255  (.A(g12657), .B(g3566), .Z(g13525) ) ;
INV     gate9256  (.A(g13525), .Z(II23553) ) ;
INV     gate9257  (.A(II23553), .Z(g17465) ) ;
NAND2   gate9258  (.A(g12657), .B(g6783), .Z(g15837) ) ;
INV     gate9259  (.A(g15837), .Z(II23556) ) ;
INV     gate9260  (.A(II23556), .Z(g17468) ) ;
NAND2   gate9261  (.A(g12657), .B(g6574), .Z(g15869) ) ;
INV     gate9262  (.A(g15869), .Z(II23559) ) ;
INV     gate9263  (.A(II23559), .Z(g17471) ) ;
NAND2   gate9264  (.A(g12711), .B(g3722), .Z(g13526) ) ;
INV     gate9265  (.A(g13526), .Z(II23564) ) ;
INV     gate9266  (.A(II23564), .Z(g17476) ) ;
NAND2   gate9267  (.A(g12711), .B(g7085), .Z(g15839) ) ;
INV     gate9268  (.A(g15839), .Z(II23567) ) ;
INV     gate9269  (.A(II23567), .Z(g17479) ) ;
NAND2   gate9270  (.A(g12711), .B(g6838), .Z(g15871) ) ;
INV     gate9271  (.A(g15871), .Z(II23570) ) ;
INV     gate9272  (.A(II23570), .Z(g17482) ) ;
NAND2   gate9273  (.A(g12565), .B(g6314), .Z(g15843) ) ;
INV     gate9274  (.A(g15843), .Z(II23575) ) ;
INV     gate9275  (.A(II23575), .Z(g17487) ) ;
NAND2   gate9276  (.A(g12565), .B(g6232), .Z(g15879) ) ;
INV     gate9277  (.A(g15879), .Z(II23578) ) ;
INV     gate9278  (.A(II23578), .Z(g17490) ) ;
NAND2   gate9279  (.A(g12565), .B(g3254), .Z(g13528) ) ;
INV     gate9280  (.A(g13528), .Z(II23581) ) ;
INV     gate9281  (.A(II23581), .Z(g17493) ) ;
NAND2   gate9282  (.A(g12565), .B(g6314), .Z(g15845) ) ;
INV     gate9283  (.A(g15845), .Z(II23584) ) ;
INV     gate9284  (.A(II23584), .Z(g17496) ) ;
AND2    gate9285  (.A(g294), .B(g11932), .Z(g16292) ) ;
INV     gate9286  (.A(g16292), .Z(g17499) ) ;
INV     gate9287  (.A(g14885), .Z(II23588) ) ;
INV     gate9288  (.A(II23588), .Z(g17500) ) ;
INV     gate9289  (.A(g14885), .Z(II23591) ) ;
INV     gate9290  (.A(II23591), .Z(g17503) ) ;
NAND2   gate9291  (.A(g12611), .B(g6369), .Z(g15887) ) ;
INV     gate9292  (.A(g15887), .Z(II23599) ) ;
INV     gate9293  (.A(II23599), .Z(g17511) ) ;
NAND2   gate9294  (.A(g12611), .B(g3410), .Z(g13529) ) ;
INV     gate9295  (.A(g13529), .Z(II23602) ) ;
INV     gate9296  (.A(II23602), .Z(g17514) ) ;
NAND2   gate9297  (.A(g12611), .B(g6519), .Z(g15847) ) ;
INV     gate9298  (.A(g15847), .Z(II23605) ) ;
INV     gate9299  (.A(II23605), .Z(g17517) ) ;
NAND2   gate9300  (.A(g12611), .B(g6369), .Z(g15889) ) ;
INV     gate9301  (.A(g15889), .Z(II23608) ) ;
INV     gate9302  (.A(II23608), .Z(g17520) ) ;
INV     gate9303  (.A(g14966), .Z(II23611) ) ;
INV     gate9304  (.A(II23611), .Z(g17523) ) ;
NAND2   gate9305  (.A(g12657), .B(g3566), .Z(g13535) ) ;
INV     gate9306  (.A(g13535), .Z(II23619) ) ;
INV     gate9307  (.A(II23619), .Z(g17531) ) ;
NAND2   gate9308  (.A(g12657), .B(g6783), .Z(g15849) ) ;
INV     gate9309  (.A(g15849), .Z(II23622) ) ;
INV     gate9310  (.A(II23622), .Z(g17534) ) ;
NAND2   gate9311  (.A(g12657), .B(g6574), .Z(g15898) ) ;
INV     gate9312  (.A(g15898), .Z(II23625) ) ;
INV     gate9313  (.A(II23625), .Z(g17537) ) ;
NAND2   gate9314  (.A(g12711), .B(g3722), .Z(g13536) ) ;
INV     gate9315  (.A(g13536), .Z(II23633) ) ;
INV     gate9316  (.A(II23633), .Z(g17545) ) ;
NAND2   gate9317  (.A(g12711), .B(g7085), .Z(g15851) ) ;
INV     gate9318  (.A(g15851), .Z(II23636) ) ;
INV     gate9319  (.A(II23636), .Z(g17548) ) ;
NAND2   gate9320  (.A(g12711), .B(g6838), .Z(g15900) ) ;
INV     gate9321  (.A(g15900), .Z(II23639) ) ;
INV     gate9322  (.A(II23639), .Z(g17551) ) ;
NAND2   gate9323  (.A(g12565), .B(g3254), .Z(g13537) ) ;
INV     gate9324  (.A(g13537), .Z(II23645) ) ;
INV     gate9325  (.A(II23645), .Z(g17557) ) ;
NAND2   gate9326  (.A(g12565), .B(g6314), .Z(g15857) ) ;
INV     gate9327  (.A(g15857), .Z(II23648) ) ;
INV     gate9328  (.A(II23648), .Z(g17560) ) ;
NAND2   gate9329  (.A(g12565), .B(g3254), .Z(g13538) ) ;
INV     gate9330  (.A(g13538), .Z(II23651) ) ;
INV     gate9331  (.A(II23651), .Z(g17563) ) ;
AND2    gate9332  (.A(g295), .B(g11972), .Z(g16346) ) ;
INV     gate9333  (.A(g16346), .Z(g17566) ) ;
INV     gate9334  (.A(g14831), .Z(II23655) ) ;
INV     gate9335  (.A(II23655), .Z(g17567) ) ;
INV     gate9336  (.A(g14885), .Z(II23658) ) ;
INV     gate9337  (.A(II23658), .Z(g17570) ) ;
NAND2   gate9338  (.A(g12883), .B(g633), .Z(g16085) ) ;
INV     gate9339  (.A(g16085), .Z(II23661) ) ;
INV     gate9340  (.A(II23661), .Z(g17573) ) ;
NAND2   gate9341  (.A(g12611), .B(g6519), .Z(g15866) ) ;
INV     gate9342  (.A(g15866), .Z(II23667) ) ;
INV     gate9343  (.A(II23667), .Z(g17579) ) ;
NAND2   gate9344  (.A(g12611), .B(g6369), .Z(g15912) ) ;
INV     gate9345  (.A(g15912), .Z(II23670) ) ;
INV     gate9346  (.A(II23670), .Z(g17582) ) ;
NAND2   gate9347  (.A(g12611), .B(g3410), .Z(g13539) ) ;
INV     gate9348  (.A(g13539), .Z(II23673) ) ;
INV     gate9349  (.A(II23673), .Z(g17585) ) ;
NAND2   gate9350  (.A(g12611), .B(g6519), .Z(g15868) ) ;
INV     gate9351  (.A(g15868), .Z(II23676) ) ;
INV     gate9352  (.A(II23676), .Z(g17588) ) ;
INV     gate9353  (.A(g14966), .Z(II23679) ) ;
INV     gate9354  (.A(II23679), .Z(g17591) ) ;
INV     gate9355  (.A(g14966), .Z(II23682) ) ;
INV     gate9356  (.A(II23682), .Z(g17594) ) ;
NAND2   gate9357  (.A(g12657), .B(g6574), .Z(g15920) ) ;
INV     gate9358  (.A(g15920), .Z(II23689) ) ;
INV     gate9359  (.A(II23689), .Z(g17601) ) ;
NAND2   gate9360  (.A(g12657), .B(g3566), .Z(g13540) ) ;
INV     gate9361  (.A(g13540), .Z(II23692) ) ;
INV     gate9362  (.A(II23692), .Z(g17604) ) ;
NAND2   gate9363  (.A(g12657), .B(g6783), .Z(g15870) ) ;
INV     gate9364  (.A(g15870), .Z(II23695) ) ;
INV     gate9365  (.A(II23695), .Z(g17607) ) ;
NAND2   gate9366  (.A(g12657), .B(g6574), .Z(g15922) ) ;
INV     gate9367  (.A(g15922), .Z(II23698) ) ;
INV     gate9368  (.A(II23698), .Z(g17610) ) ;
INV     gate9369  (.A(g15055), .Z(II23701) ) ;
INV     gate9370  (.A(II23701), .Z(g17613) ) ;
NAND2   gate9371  (.A(g12711), .B(g3722), .Z(g13546) ) ;
INV     gate9372  (.A(g13546), .Z(II23709) ) ;
INV     gate9373  (.A(II23709), .Z(g17621) ) ;
NAND2   gate9374  (.A(g12711), .B(g7085), .Z(g15872) ) ;
INV     gate9375  (.A(g15872), .Z(II23712) ) ;
INV     gate9376  (.A(II23712), .Z(g17624) ) ;
NAND2   gate9377  (.A(g12711), .B(g6838), .Z(g15931) ) ;
INV     gate9378  (.A(g15931), .Z(II23715) ) ;
INV     gate9379  (.A(II23715), .Z(g17627) ) ;
NAND2   gate9380  (.A(g12565), .B(g3254), .Z(g13547) ) ;
INV     gate9381  (.A(g13547), .Z(II23725) ) ;
INV     gate9382  (.A(II23725), .Z(g17637) ) ;
INV     gate9383  (.A(g13873), .Z(g17640) ) ;
INV     gate9384  (.A(g14337), .Z(II23729) ) ;
INV     gate9385  (.A(II23729), .Z(g17645) ) ;
AND2    gate9386  (.A(g296), .B(g12024), .Z(g16384) ) ;
INV     gate9387  (.A(g16384), .Z(g17648) ) ;
INV     gate9388  (.A(g14831), .Z(II23733) ) ;
INV     gate9389  (.A(II23733), .Z(g17649) ) ;
NAND2   gate9390  (.A(g12611), .B(g3410), .Z(g13548) ) ;
INV     gate9391  (.A(g13548), .Z(II23739) ) ;
INV     gate9392  (.A(II23739), .Z(g17655) ) ;
NAND2   gate9393  (.A(g12611), .B(g6519), .Z(g15888) ) ;
INV     gate9394  (.A(g15888), .Z(II23742) ) ;
INV     gate9395  (.A(II23742), .Z(g17658) ) ;
NAND2   gate9396  (.A(g12611), .B(g3410), .Z(g13549) ) ;
INV     gate9397  (.A(g13549), .Z(II23745) ) ;
INV     gate9398  (.A(II23745), .Z(g17661) ) ;
INV     gate9399  (.A(g14904), .Z(II23748) ) ;
INV     gate9400  (.A(II23748), .Z(g17664) ) ;
INV     gate9401  (.A(g14966), .Z(II23751) ) ;
INV     gate9402  (.A(II23751), .Z(g17667) ) ;
NAND2   gate9403  (.A(g12923), .B(g1319), .Z(g16123) ) ;
INV     gate9404  (.A(g16123), .Z(II23754) ) ;
INV     gate9405  (.A(II23754), .Z(g17670) ) ;
NAND2   gate9406  (.A(g12657), .B(g6783), .Z(g15897) ) ;
INV     gate9407  (.A(g15897), .Z(II23760) ) ;
INV     gate9408  (.A(II23760), .Z(g17676) ) ;
NAND2   gate9409  (.A(g12657), .B(g6574), .Z(g15941) ) ;
INV     gate9410  (.A(g15941), .Z(II23763) ) ;
INV     gate9411  (.A(II23763), .Z(g17679) ) ;
NAND2   gate9412  (.A(g12657), .B(g3566), .Z(g13550) ) ;
INV     gate9413  (.A(g13550), .Z(II23766) ) ;
INV     gate9414  (.A(II23766), .Z(g17682) ) ;
NAND2   gate9415  (.A(g12657), .B(g6783), .Z(g15899) ) ;
INV     gate9416  (.A(g15899), .Z(II23769) ) ;
INV     gate9417  (.A(II23769), .Z(g17685) ) ;
INV     gate9418  (.A(g15055), .Z(II23772) ) ;
INV     gate9419  (.A(II23772), .Z(g17688) ) ;
INV     gate9420  (.A(g15055), .Z(II23775) ) ;
INV     gate9421  (.A(II23775), .Z(g17691) ) ;
NAND2   gate9422  (.A(g12711), .B(g6838), .Z(g15949) ) ;
INV     gate9423  (.A(g15949), .Z(II23782) ) ;
INV     gate9424  (.A(II23782), .Z(g17698) ) ;
NAND2   gate9425  (.A(g12711), .B(g3722), .Z(g13551) ) ;
INV     gate9426  (.A(g13551), .Z(II23785) ) ;
INV     gate9427  (.A(II23785), .Z(g17701) ) ;
NAND2   gate9428  (.A(g12711), .B(g7085), .Z(g15901) ) ;
INV     gate9429  (.A(g15901), .Z(II23788) ) ;
INV     gate9430  (.A(II23788), .Z(g17704) ) ;
NAND2   gate9431  (.A(g12711), .B(g6838), .Z(g15951) ) ;
INV     gate9432  (.A(g15951), .Z(II23791) ) ;
INV     gate9433  (.A(II23791), .Z(g17707) ) ;
INV     gate9434  (.A(g15151), .Z(II23794) ) ;
INV     gate9435  (.A(II23794), .Z(g17710) ) ;
NAND2   gate9436  (.A(g13310), .B(g12354), .Z(g15853) ) ;
INV     gate9437  (.A(g15853), .Z(g17720) ) ;
INV     gate9438  (.A(g13886), .Z(g17724) ) ;
NAND2   gate9439  (.A(g12611), .B(g3410), .Z(g13557) ) ;
INV     gate9440  (.A(g13557), .Z(II23817) ) ;
INV     gate9441  (.A(II23817), .Z(g17738) ) ;
INV     gate9442  (.A(g13895), .Z(g17741) ) ;
INV     gate9443  (.A(g14337), .Z(II23821) ) ;
INV     gate9444  (.A(II23821), .Z(g17746) ) ;
INV     gate9445  (.A(g14904), .Z(II23824) ) ;
INV     gate9446  (.A(II23824), .Z(g17749) ) ;
NAND2   gate9447  (.A(g12657), .B(g3566), .Z(g13558) ) ;
INV     gate9448  (.A(g13558), .Z(II23830) ) ;
INV     gate9449  (.A(II23830), .Z(g17755) ) ;
NAND2   gate9450  (.A(g12657), .B(g6783), .Z(g15921) ) ;
INV     gate9451  (.A(g15921), .Z(II23833) ) ;
INV     gate9452  (.A(II23833), .Z(g17758) ) ;
NAND2   gate9453  (.A(g12657), .B(g3566), .Z(g13559) ) ;
INV     gate9454  (.A(g13559), .Z(II23836) ) ;
INV     gate9455  (.A(II23836), .Z(g17761) ) ;
INV     gate9456  (.A(g14985), .Z(II23839) ) ;
INV     gate9457  (.A(II23839), .Z(g17764) ) ;
INV     gate9458  (.A(g15055), .Z(II23842) ) ;
INV     gate9459  (.A(II23842), .Z(g17767) ) ;
NAND2   gate9460  (.A(g12952), .B(g2013), .Z(g16174) ) ;
INV     gate9461  (.A(g16174), .Z(II23845) ) ;
INV     gate9462  (.A(II23845), .Z(g17770) ) ;
NAND2   gate9463  (.A(g12711), .B(g7085), .Z(g15930) ) ;
INV     gate9464  (.A(g15930), .Z(II23851) ) ;
INV     gate9465  (.A(II23851), .Z(g17776) ) ;
NAND2   gate9466  (.A(g12711), .B(g6838), .Z(g15970) ) ;
INV     gate9467  (.A(g15970), .Z(II23854) ) ;
INV     gate9468  (.A(II23854), .Z(g17779) ) ;
NAND2   gate9469  (.A(g12711), .B(g3722), .Z(g13560) ) ;
INV     gate9470  (.A(g13560), .Z(II23857) ) ;
INV     gate9471  (.A(II23857), .Z(g17782) ) ;
NAND2   gate9472  (.A(g12711), .B(g7085), .Z(g15932) ) ;
INV     gate9473  (.A(g15932), .Z(II23860) ) ;
INV     gate9474  (.A(II23860), .Z(g17785) ) ;
INV     gate9475  (.A(g15151), .Z(II23863) ) ;
INV     gate9476  (.A(II23863), .Z(g17788) ) ;
INV     gate9477  (.A(g15151), .Z(II23866) ) ;
INV     gate9478  (.A(II23866), .Z(g17791) ) ;
NOR2    gate9479  (.A(g13305), .B(g7143), .Z(g15797) ) ;
INV     gate9480  (.A(g15797), .Z(II23874) ) ;
INV     gate9481  (.A(II23874), .Z(g17799) ) ;
INV     gate9482  (.A(g13907), .Z(g17802) ) ;
INV     gate9483  (.A(g14685), .Z(II23888) ) ;
INV     gate9484  (.A(II23888), .Z(g17815) ) ;
INV     gate9485  (.A(g13927), .Z(g17825) ) ;
NAND2   gate9486  (.A(g12657), .B(g3566), .Z(g13561) ) ;
INV     gate9487  (.A(g13561), .Z(II23904) ) ;
INV     gate9488  (.A(II23904), .Z(g17839) ) ;
INV     gate9489  (.A(g13936), .Z(g17842) ) ;
INV     gate9490  (.A(g14337), .Z(II23908) ) ;
INV     gate9491  (.A(II23908), .Z(g17847) ) ;
INV     gate9492  (.A(g14985), .Z(II23911) ) ;
INV     gate9493  (.A(II23911), .Z(g17850) ) ;
NAND2   gate9494  (.A(g12711), .B(g3722), .Z(g13562) ) ;
INV     gate9495  (.A(g13562), .Z(II23917) ) ;
INV     gate9496  (.A(II23917), .Z(g17856) ) ;
NAND2   gate9497  (.A(g12711), .B(g7085), .Z(g15950) ) ;
INV     gate9498  (.A(g15950), .Z(II23920) ) ;
INV     gate9499  (.A(II23920), .Z(g17859) ) ;
NAND2   gate9500  (.A(g12711), .B(g3722), .Z(g13563) ) ;
INV     gate9501  (.A(g13563), .Z(II23923) ) ;
INV     gate9502  (.A(II23923), .Z(g17862) ) ;
INV     gate9503  (.A(g15074), .Z(II23926) ) ;
INV     gate9504  (.A(II23926), .Z(g17865) ) ;
INV     gate9505  (.A(g15151), .Z(II23929) ) ;
INV     gate9506  (.A(II23929), .Z(g17868) ) ;
NAND2   gate9507  (.A(g12981), .B(g2707), .Z(g16233) ) ;
INV     gate9508  (.A(g16233), .Z(II23932) ) ;
INV     gate9509  (.A(II23932), .Z(g17871) ) ;
NAND2   gate9510  (.A(g13310), .B(g12392), .Z(g15830) ) ;
INV     gate9511  (.A(g15830), .Z(g17878) ) ;
INV     gate9512  (.A(g13946), .Z(g17882) ) ;
INV     gate9513  (.A(g13954), .Z(g17892) ) ;
INV     gate9514  (.A(g14165), .Z(g17893) ) ;
INV     gate9515  (.A(g16154), .Z(II23954) ) ;
INV     gate9516  (.A(II23954), .Z(g17903) ) ;
INV     gate9517  (.A(g13963), .Z(g17914) ) ;
INV     gate9518  (.A(g14719), .Z(II23976) ) ;
INV     gate9519  (.A(II23976), .Z(g17927) ) ;
INV     gate9520  (.A(g13983), .Z(g17937) ) ;
NAND2   gate9521  (.A(g12711), .B(g3722), .Z(g13564) ) ;
INV     gate9522  (.A(g13564), .Z(II23992) ) ;
INV     gate9523  (.A(II23992), .Z(g17951) ) ;
INV     gate9524  (.A(g13992), .Z(g17954) ) ;
INV     gate9525  (.A(g14337), .Z(II23996) ) ;
INV     gate9526  (.A(II23996), .Z(g17959) ) ;
INV     gate9527  (.A(g15074), .Z(II23999) ) ;
INV     gate9528  (.A(II23999), .Z(g17962) ) ;
NAND2   gate9529  (.A(g13331), .B(g12392), .Z(g15841) ) ;
INV     gate9530  (.A(g15841), .Z(g17969) ) ;
INV     gate9531  (.A(g14001), .Z(g17974) ) ;
INV     gate9532  (.A(g14008), .Z(g17984) ) ;
INV     gate9533  (.A(g14685), .Z(g17988) ) ;
INV     gate9534  (.A(g14450), .Z(g17991) ) ;
INV     gate9535  (.A(g14016), .Z(g17993) ) ;
INV     gate9536  (.A(g14024), .Z(g18003) ) ;
INV     gate9537  (.A(g14280), .Z(g18004) ) ;
INV     gate9538  (.A(g16213), .Z(II24049) ) ;
INV     gate9539  (.A(II24049), .Z(g18014) ) ;
INV     gate9540  (.A(g14033), .Z(g18025) ) ;
INV     gate9541  (.A(g14747), .Z(II24071) ) ;
INV     gate9542  (.A(II24071), .Z(g18038) ) ;
INV     gate9543  (.A(g14053), .Z(g18048) ) ;
NAND2   gate9544  (.A(g13401), .B(g12354), .Z(g15660) ) ;
INV     gate9545  (.A(g15660), .Z(g18063) ) ;
NAND2   gate9546  (.A(g13353), .B(g12392), .Z(g15854) ) ;
INV     gate9547  (.A(g15854), .Z(g18070) ) ;
INV     gate9548  (.A(g14062), .Z(g18074) ) ;
INV     gate9549  (.A(g14068), .Z(g18084) ) ;
INV     gate9550  (.A(g14355), .Z(g18089) ) ;
INV     gate9551  (.A(g14092), .Z(g18091) ) ;
INV     gate9552  (.A(g14099), .Z(g18101) ) ;
INV     gate9553  (.A(g14719), .Z(g18105) ) ;
INV     gate9554  (.A(g14537), .Z(g18108) ) ;
INV     gate9555  (.A(g14107), .Z(g18110) ) ;
INV     gate9556  (.A(g14115), .Z(g18120) ) ;
INV     gate9557  (.A(g14402), .Z(g18121) ) ;
INV     gate9558  (.A(g16278), .Z(II24144) ) ;
INV     gate9559  (.A(II24144), .Z(g18131) ) ;
INV     gate9560  (.A(g14124), .Z(g18142) ) ;
INV     gate9561  (.A(g14768), .Z(II24166) ) ;
INV     gate9562  (.A(II24166), .Z(g18155) ) ;
NAND2   gate9563  (.A(g13082), .B(g2912), .Z(g16439) ) ;
INV     gate9564  (.A(g16439), .Z(II24171) ) ;
INV     gate9565  (.A(II24171), .Z(g18166) ) ;
NAND2   gate9566  (.A(g13374), .B(g12392), .Z(g15877) ) ;
INV     gate9567  (.A(g15877), .Z(g18170) ) ;
INV     gate9568  (.A(g14148), .Z(g18174) ) ;
INV     gate9569  (.A(g14153), .Z(g18179) ) ;
INV     gate9570  (.A(g14252), .Z(g18188) ) ;
INV     gate9571  (.A(g14177), .Z(g18190) ) ;
INV     gate9572  (.A(g14183), .Z(g18200) ) ;
INV     gate9573  (.A(g14467), .Z(g18205) ) ;
INV     gate9574  (.A(g14207), .Z(g18207) ) ;
INV     gate9575  (.A(g14214), .Z(g18217) ) ;
INV     gate9576  (.A(g14747), .Z(g18221) ) ;
INV     gate9577  (.A(g14592), .Z(g18224) ) ;
INV     gate9578  (.A(g14222), .Z(g18226) ) ;
INV     gate9579  (.A(g14230), .Z(g18236) ) ;
INV     gate9580  (.A(g14514), .Z(g18237) ) ;
INV     gate9581  (.A(g16337), .Z(II24247) ) ;
INV     gate9582  (.A(II24247), .Z(g18247) ) ;
NAND2   gate9583  (.A(g13004), .B(g3018), .Z(g16463) ) ;
INV     gate9584  (.A(g16463), .Z(II24258) ) ;
INV     gate9585  (.A(II24258), .Z(g18258) ) ;
NAND2   gate9586  (.A(g13401), .B(g12392), .Z(g15719) ) ;
INV     gate9587  (.A(g15719), .Z(g18261) ) ;
INV     gate9588  (.A(g14238), .Z(g18265) ) ;
INV     gate9589  (.A(g14171), .Z(g18275) ) ;
NAND2   gate9590  (.A(g12886), .B(g6678), .Z(g15992) ) ;
INV     gate9591  (.A(g15992), .Z(II24285) ) ;
INV     gate9592  (.A(II24285), .Z(g18278) ) ;
INV     gate9593  (.A(g14263), .Z(g18281) ) ;
INV     gate9594  (.A(g14268), .Z(g18286) ) ;
INV     gate9595  (.A(g14374), .Z(g18295) ) ;
INV     gate9596  (.A(g14292), .Z(g18297) ) ;
INV     gate9597  (.A(g14298), .Z(g18307) ) ;
INV     gate9598  (.A(g14554), .Z(g18312) ) ;
INV     gate9599  (.A(g14322), .Z(g18314) ) ;
INV     gate9600  (.A(g14329), .Z(g18324) ) ;
INV     gate9601  (.A(g14768), .Z(g18328) ) ;
INV     gate9602  (.A(g14626), .Z(g18331) ) ;
NOR2    gate9603  (.A(g11617), .B(g7562), .Z(g15873) ) ;
INV     gate9604  (.A(g15873), .Z(II24346) ) ;
INV     gate9605  (.A(II24346), .Z(g18334) ) ;
NAND2   gate9606  (.A(g11622), .B(g12392), .Z(g15757) ) ;
INV     gate9607  (.A(g15757), .Z(g18337) ) ;
INV     gate9608  (.A(g14342), .Z(g18341) ) ;
INV     gate9609  (.A(g13741), .Z(g18351) ) ;
INV     gate9610  (.A(g13918), .Z(g18353) ) ;
NAND2   gate9611  (.A(g12886), .B(g6912), .Z(g15990) ) ;
INV     gate9612  (.A(g15990), .Z(II24368) ) ;
INV     gate9613  (.A(II24368), .Z(g18355) ) ;
INV     gate9614  (.A(g14360), .Z(g18358) ) ;
INV     gate9615  (.A(g14286), .Z(g18368) ) ;
NAND2   gate9616  (.A(g12926), .B(g6980), .Z(g15995) ) ;
INV     gate9617  (.A(g15995), .Z(II24394) ) ;
INV     gate9618  (.A(II24394), .Z(g18371) ) ;
INV     gate9619  (.A(g14385), .Z(g18374) ) ;
INV     gate9620  (.A(g14390), .Z(g18379) ) ;
INV     gate9621  (.A(g14486), .Z(g18388) ) ;
INV     gate9622  (.A(g14414), .Z(g18390) ) ;
INV     gate9623  (.A(g14420), .Z(g18400) ) ;
INV     gate9624  (.A(g14609), .Z(g18405) ) ;
NOR2    gate9625  (.A(g2814), .B(g13082), .Z(g15959) ) ;
INV     gate9626  (.A(g15959), .Z(g18407) ) ;
NAND2   gate9627  (.A(g13286), .B(g12354), .Z(g15718) ) ;
INV     gate9628  (.A(g15718), .Z(g18414) ) ;
NAND2   gate9629  (.A(g11643), .B(g12392), .Z(g15783) ) ;
INV     gate9630  (.A(g15783), .Z(g18415) ) ;
INV     gate9631  (.A(g14831), .Z(g18429) ) ;
NAND2   gate9632  (.A(g12886), .B(g3366), .Z(g13599) ) ;
INV     gate9633  (.A(g13599), .Z(II24459) ) ;
INV     gate9634  (.A(II24459), .Z(g18432) ) ;
INV     gate9635  (.A(g14359), .Z(g18435) ) ;
INV     gate9636  (.A(g14454), .Z(g18436) ) ;
INV     gate9637  (.A(g13741), .Z(g18446) ) ;
INV     gate9638  (.A(g13974), .Z(g18448) ) ;
NAND2   gate9639  (.A(g12926), .B(g7162), .Z(g15993) ) ;
INV     gate9640  (.A(g15993), .Z(II24481) ) ;
INV     gate9641  (.A(II24481), .Z(g18450) ) ;
INV     gate9642  (.A(g14472), .Z(g18453) ) ;
INV     gate9643  (.A(g14408), .Z(g18463) ) ;
NAND2   gate9644  (.A(g12955), .B(g7230), .Z(g15999) ) ;
INV     gate9645  (.A(g15999), .Z(II24507) ) ;
INV     gate9646  (.A(II24507), .Z(g18466) ) ;
INV     gate9647  (.A(g14497), .Z(g18469) ) ;
INV     gate9648  (.A(g14502), .Z(g18474) ) ;
INV     gate9649  (.A(g14573), .Z(g18483) ) ;
NAND2   gate9650  (.A(g13313), .B(g12354), .Z(g15756) ) ;
INV     gate9651  (.A(g15756), .Z(g18485) ) ;
NAND2   gate9652  (.A(g11660), .B(g12392), .Z(g15804) ) ;
INV     gate9653  (.A(g15804), .Z(g18486) ) ;
INV     gate9654  (.A(g13565), .Z(g18490) ) ;
INV     gate9655  (.A(g14904), .Z(g18502) ) ;
NAND2   gate9656  (.A(g12926), .B(g3522), .Z(g13611) ) ;
INV     gate9657  (.A(g13611), .Z(II24560) ) ;
INV     gate9658  (.A(II24560), .Z(g18505) ) ;
INV     gate9659  (.A(g14471), .Z(g18508) ) ;
INV     gate9660  (.A(g14541), .Z(g18509) ) ;
INV     gate9661  (.A(g13741), .Z(g18519) ) ;
INV     gate9662  (.A(g14044), .Z(g18521) ) ;
NAND2   gate9663  (.A(g12955), .B(g7358), .Z(g15996) ) ;
INV     gate9664  (.A(g15996), .Z(II24582) ) ;
INV     gate9665  (.A(II24582), .Z(g18523) ) ;
INV     gate9666  (.A(g14559), .Z(g18526) ) ;
INV     gate9667  (.A(g14520), .Z(g18536) ) ;
NAND2   gate9668  (.A(g12984), .B(g7426), .Z(g16006) ) ;
INV     gate9669  (.A(g16006), .Z(II24608) ) ;
INV     gate9670  (.A(II24608), .Z(g18539) ) ;
NAND2   gate9671  (.A(g13286), .B(g12392), .Z(g15819) ) ;
INV     gate9672  (.A(g15819), .Z(g18543) ) ;
INV     gate9673  (.A(g16154), .Z(g18552) ) ;
INV     gate9674  (.A(g13573), .Z(g18554) ) ;
INV     gate9675  (.A(g14985), .Z(g18566) ) ;
NAND2   gate9676  (.A(g12955), .B(g3678), .Z(g13621) ) ;
INV     gate9677  (.A(g13621), .Z(II24662) ) ;
INV     gate9678  (.A(II24662), .Z(g18569) ) ;
INV     gate9679  (.A(g14558), .Z(g18572) ) ;
INV     gate9680  (.A(g14596), .Z(g18573) ) ;
INV     gate9681  (.A(g13741), .Z(g18583) ) ;
INV     gate9682  (.A(g14135), .Z(g18585) ) ;
NAND2   gate9683  (.A(g12984), .B(g7488), .Z(g16000) ) ;
INV     gate9684  (.A(g16000), .Z(II24684) ) ;
INV     gate9685  (.A(II24684), .Z(g18587) ) ;
NAND2   gate9686  (.A(g13313), .B(g12392), .Z(g15831) ) ;
INV     gate9687  (.A(g15831), .Z(g18593) ) ;
INV     gate9688  (.A(g16213), .Z(g18602) ) ;
INV     gate9689  (.A(g13582), .Z(g18604) ) ;
INV     gate9690  (.A(g15074), .Z(g18616) ) ;
NAND2   gate9691  (.A(g12984), .B(g3834), .Z(g13633) ) ;
INV     gate9692  (.A(g13633), .Z(II24732) ) ;
INV     gate9693  (.A(II24732), .Z(g18619) ) ;
INV     gate9694  (.A(g14613), .Z(g18622) ) ;
INV     gate9695  (.A(g16278), .Z(g18634) ) ;
INV     gate9696  (.A(g13602), .Z(g18636) ) ;
INV     gate9697  (.A(g16337), .Z(g18643) ) ;
NAND2   gate9698  (.A(g12377), .B(g12407), .Z(g16341) ) ;
INV     gate9699  (.A(g16341), .Z(g18646) ) ;
INV     gate9700  (.A(g14776), .Z(g18656) ) ;
INV     gate9701  (.A(g14797), .Z(g18670) ) ;
INV     gate9702  (.A(g14811), .Z(g18679) ) ;
INV     gate9703  (.A(g14885), .Z(g18691) ) ;
INV     gate9704  (.A(g14837), .Z(g18692) ) ;
INV     gate9705  (.A(g14849), .Z(g18699) ) ;
INV     gate9706  (.A(g14863), .Z(g18708) ) ;
INV     gate9707  (.A(g14895), .Z(g18720) ) ;
AND2    gate9708  (.A(g548), .B(g12748), .Z(g13865) ) ;
INV     gate9709  (.A(g13865), .Z(g18725) ) ;
INV     gate9710  (.A(g14966), .Z(g18727) ) ;
INV     gate9711  (.A(g14910), .Z(g18728) ) ;
INV     gate9712  (.A(g14922), .Z(g18735) ) ;
INV     gate9713  (.A(g14936), .Z(g18744) ) ;
INV     gate9714  (.A(g14960), .Z(g18756) ) ;
INV     gate9715  (.A(g14963), .Z(g18757) ) ;
INV     gate9716  (.A(g14976), .Z(g18758) ) ;
INV     gate9717  (.A(g15055), .Z(g18764) ) ;
INV     gate9718  (.A(g14991), .Z(g18765) ) ;
INV     gate9719  (.A(g15003), .Z(g18772) ) ;
INV     gate9720  (.A(g15034), .Z(g18783) ) ;
INV     gate9721  (.A(g15037), .Z(g18784) ) ;
INV     gate9722  (.A(g15040), .Z(g18785) ) ;
INV     gate9723  (.A(g15043), .Z(g18786) ) ;
INV     gate9724  (.A(g15049), .Z(g18787) ) ;
INV     gate9725  (.A(g15052), .Z(g18788) ) ;
INV     gate9726  (.A(g15065), .Z(g18789) ) ;
INV     gate9727  (.A(g15151), .Z(g18795) ) ;
INV     gate9728  (.A(g15080), .Z(g18796) ) ;
INV     gate9729  (.A(g15106), .Z(g18805) ) ;
INV     gate9730  (.A(g15109), .Z(g18806) ) ;
INV     gate9731  (.A(g15112), .Z(g18807) ) ;
INV     gate9732  (.A(g15115), .Z(g18808) ) ;
INV     gate9733  (.A(g15130), .Z(g18809) ) ;
INV     gate9734  (.A(g15133), .Z(g18810) ) ;
INV     gate9735  (.A(g15136), .Z(g18811) ) ;
INV     gate9736  (.A(g15139), .Z(g18812) ) ;
INV     gate9737  (.A(g15145), .Z(g18813) ) ;
INV     gate9738  (.A(g15148), .Z(g18814) ) ;
INV     gate9739  (.A(g15161), .Z(g18815) ) ;
INV     gate9740  (.A(g15179), .Z(g18822) ) ;
INV     gate9741  (.A(g15182), .Z(g18823) ) ;
INV     gate9742  (.A(g15185), .Z(g18824) ) ;
INV     gate9743  (.A(g15198), .Z(g18825) ) ;
INV     gate9744  (.A(g15201), .Z(g18826) ) ;
INV     gate9745  (.A(g15204), .Z(g18827) ) ;
INV     gate9746  (.A(g15207), .Z(g18828) ) ;
INV     gate9747  (.A(g15222), .Z(g18829) ) ;
INV     gate9748  (.A(g15225), .Z(g18830) ) ;
INV     gate9749  (.A(g15228), .Z(g18831) ) ;
INV     gate9750  (.A(g15231), .Z(g18832) ) ;
INV     gate9751  (.A(g15237), .Z(g18833) ) ;
INV     gate9752  (.A(g15240), .Z(g18834) ) ;
INV     gate9753  (.A(g15248), .Z(g18838) ) ;
INV     gate9754  (.A(g15251), .Z(g18839) ) ;
INV     gate9755  (.A(g15254), .Z(g18840) ) ;
INV     gate9756  (.A(g15265), .Z(g18841) ) ;
INV     gate9757  (.A(g15268), .Z(g18842) ) ;
INV     gate9758  (.A(g15271), .Z(g18843) ) ;
INV     gate9759  (.A(g15284), .Z(g18844) ) ;
INV     gate9760  (.A(g15287), .Z(g18845) ) ;
INV     gate9761  (.A(g15290), .Z(g18846) ) ;
INV     gate9762  (.A(g15293), .Z(g18847) ) ;
INV     gate9763  (.A(g15308), .Z(g18848) ) ;
INV     gate9764  (.A(g15311), .Z(g18849) ) ;
INV     gate9765  (.A(g15314), .Z(g18850) ) ;
INV     gate9766  (.A(g15317), .Z(g18851) ) ;
INV     gate9767  (.A(g15326), .Z(g18853) ) ;
INV     gate9768  (.A(g15329), .Z(g18854) ) ;
INV     gate9769  (.A(g15332), .Z(g18855) ) ;
INV     gate9770  (.A(g15340), .Z(g18856) ) ;
INV     gate9771  (.A(g15343), .Z(g18857) ) ;
INV     gate9772  (.A(g15346), .Z(g18858) ) ;
INV     gate9773  (.A(g15357), .Z(g18859) ) ;
INV     gate9774  (.A(g15360), .Z(g18860) ) ;
INV     gate9775  (.A(g15363), .Z(g18861) ) ;
INV     gate9776  (.A(g15376), .Z(g18862) ) ;
INV     gate9777  (.A(g15379), .Z(g18863) ) ;
INV     gate9778  (.A(g15382), .Z(g18864) ) ;
INV     gate9779  (.A(g15385), .Z(g18865) ) ;
INV     gate9780  (.A(g14797), .Z(II24894) ) ;
INV     gate9781  (.A(II24894), .Z(g18869) ) ;
INV     gate9782  (.A(g15393), .Z(g18870) ) ;
INV     gate9783  (.A(g15396), .Z(g18871) ) ;
INV     gate9784  (.A(g15399), .Z(g18872) ) ;
INV     gate9785  (.A(g15404), .Z(g18873) ) ;
INV     gate9786  (.A(g15412), .Z(g18874) ) ;
INV     gate9787  (.A(g15415), .Z(g18875) ) ;
INV     gate9788  (.A(g15418), .Z(g18876) ) ;
INV     gate9789  (.A(g15426), .Z(g18877) ) ;
INV     gate9790  (.A(g15429), .Z(g18878) ) ;
INV     gate9791  (.A(g15432), .Z(g18879) ) ;
INV     gate9792  (.A(g15443), .Z(g18880) ) ;
INV     gate9793  (.A(g15446), .Z(g18881) ) ;
INV     gate9794  (.A(g15449), .Z(g18882) ) ;
INV     gate9795  (.A(g13469), .Z(g18884) ) ;
INV     gate9796  (.A(g15800), .Z(II24913) ) ;
INV     gate9797  (.A(II24913), .Z(g18886) ) ;
INV     gate9798  (.A(g14776), .Z(II24916) ) ;
INV     gate9799  (.A(II24916), .Z(g18890) ) ;
INV     gate9800  (.A(g15461), .Z(g18891) ) ;
INV     gate9801  (.A(g15464), .Z(g18892) ) ;
INV     gate9802  (.A(g15467), .Z(g18893) ) ;
INV     gate9803  (.A(g15471), .Z(g18894) ) ;
INV     gate9804  (.A(g14849), .Z(II24923) ) ;
INV     gate9805  (.A(II24923), .Z(g18895) ) ;
INV     gate9806  (.A(g15477), .Z(g18896) ) ;
INV     gate9807  (.A(g15480), .Z(g18897) ) ;
INV     gate9808  (.A(g15483), .Z(g18898) ) ;
INV     gate9809  (.A(g15488), .Z(g18899) ) ;
INV     gate9810  (.A(g15496), .Z(g18900) ) ;
INV     gate9811  (.A(g15499), .Z(g18901) ) ;
INV     gate9812  (.A(g15502), .Z(g18902) ) ;
INV     gate9813  (.A(g15510), .Z(g18903) ) ;
INV     gate9814  (.A(g15513), .Z(g18904) ) ;
INV     gate9815  (.A(g15516), .Z(g18905) ) ;
INV     gate9816  (.A(g15521), .Z(g18908) ) ;
INV     gate9817  (.A(g15528), .Z(g18909) ) ;
INV     gate9818  (.A(g15531), .Z(g18910) ) ;
INV     gate9819  (.A(g15534), .Z(g18911) ) ;
INV     gate9820  (.A(g15537), .Z(g18912) ) ;
INV     gate9821  (.A(g14811), .Z(II24943) ) ;
INV     gate9822  (.A(II24943), .Z(g18913) ) ;
INV     gate9823  (.A(g15547), .Z(g18914) ) ;
INV     gate9824  (.A(g15550), .Z(g18915) ) ;
INV     gate9825  (.A(g15553), .Z(g18916) ) ;
INV     gate9826  (.A(g15557), .Z(g18917) ) ;
INV     gate9827  (.A(g14922), .Z(II24950) ) ;
INV     gate9828  (.A(II24950), .Z(g18918) ) ;
INV     gate9829  (.A(g15563), .Z(g18919) ) ;
INV     gate9830  (.A(g15566), .Z(g18920) ) ;
INV     gate9831  (.A(g15569), .Z(g18921) ) ;
INV     gate9832  (.A(g15574), .Z(g18922) ) ;
INV     gate9833  (.A(g15582), .Z(g18923) ) ;
INV     gate9834  (.A(g15585), .Z(g18924) ) ;
INV     gate9835  (.A(g15588), .Z(g18925) ) ;
INV     gate9836  (.A(g15596), .Z(g18926) ) ;
INV     gate9837  (.A(g15599), .Z(g18927) ) ;
INV     gate9838  (.A(g15606), .Z(g18928) ) ;
INV     gate9839  (.A(g15609), .Z(g18929) ) ;
INV     gate9840  (.A(g15612), .Z(g18930) ) ;
INV     gate9841  (.A(g15615), .Z(g18931) ) ;
INV     gate9842  (.A(g14863), .Z(II24966) ) ;
INV     gate9843  (.A(II24966), .Z(g18932) ) ;
INV     gate9844  (.A(g15625), .Z(g18933) ) ;
INV     gate9845  (.A(g15628), .Z(g18934) ) ;
INV     gate9846  (.A(g15631), .Z(g18935) ) ;
INV     gate9847  (.A(g15635), .Z(g18936) ) ;
INV     gate9848  (.A(g15003), .Z(II24973) ) ;
INV     gate9849  (.A(II24973), .Z(g18937) ) ;
INV     gate9850  (.A(g15641), .Z(g18938) ) ;
INV     gate9851  (.A(g15644), .Z(g18939) ) ;
INV     gate9852  (.A(g15647), .Z(g18940) ) ;
INV     gate9853  (.A(g15652), .Z(g18941) ) ;
INV     gate9854  (.A(g15655), .Z(g18943) ) ;
INV     gate9855  (.A(g14347), .Z(II24982) ) ;
INV     gate9856  (.A(II24982), .Z(g18944) ) ;
INV     gate9857  (.A(g15667), .Z(g18945) ) ;
INV     gate9858  (.A(g15672), .Z(g18946) ) ;
INV     gate9859  (.A(g15675), .Z(g18947) ) ;
INV     gate9860  (.A(g15682), .Z(g18948) ) ;
INV     gate9861  (.A(g15685), .Z(g18949) ) ;
INV     gate9862  (.A(g15688), .Z(g18950) ) ;
INV     gate9863  (.A(g15691), .Z(g18951) ) ;
INV     gate9864  (.A(g14936), .Z(II24992) ) ;
INV     gate9865  (.A(II24992), .Z(g18952) ) ;
INV     gate9866  (.A(g15701), .Z(g18953) ) ;
INV     gate9867  (.A(g15704), .Z(g18954) ) ;
INV     gate9868  (.A(g15707), .Z(g18955) ) ;
INV     gate9869  (.A(g15711), .Z(g18956) ) ;
INV     gate9870  (.A(g15714), .Z(g18958) ) ;
INV     gate9871  (.A(g14244), .Z(II25001) ) ;
INV     gate9872  (.A(II25001), .Z(g18959) ) ;
INV     gate9873  (.A(g14459), .Z(II25004) ) ;
INV     gate9874  (.A(II25004), .Z(g18960) ) ;
INV     gate9875  (.A(g15726), .Z(g18961) ) ;
INV     gate9876  (.A(g15731), .Z(g18962) ) ;
INV     gate9877  (.A(g15734), .Z(g18963) ) ;
INV     gate9878  (.A(g15741), .Z(g18964) ) ;
INV     gate9879  (.A(g15744), .Z(g18965) ) ;
INV     gate9880  (.A(g15747), .Z(g18966) ) ;
INV     gate9881  (.A(g15750), .Z(g18967) ) ;
INV     gate9882  (.A(g14158), .Z(II25015) ) ;
INV     gate9883  (.A(II25015), .Z(g18969) ) ;
INV     gate9884  (.A(g14366), .Z(II25018) ) ;
INV     gate9885  (.A(II25018), .Z(g18970) ) ;
INV     gate9886  (.A(g14546), .Z(II25021) ) ;
INV     gate9887  (.A(II25021), .Z(g18971) ) ;
INV     gate9888  (.A(g15766), .Z(g18972) ) ;
INV     gate9889  (.A(g15771), .Z(g18973) ) ;
INV     gate9890  (.A(g15774), .Z(g18974) ) ;
INV     gate9891  (.A(g15777), .Z(g18976) ) ;
INV     gate9892  (.A(g14071), .Z(II25037) ) ;
INV     gate9893  (.A(II25037), .Z(g18981) ) ;
INV     gate9894  (.A(g14895), .Z(II25041) ) ;
INV     gate9895  (.A(II25041), .Z(g18983) ) ;
INV     gate9896  (.A(g14273), .Z(II25044) ) ;
INV     gate9897  (.A(II25044), .Z(g18984) ) ;
INV     gate9898  (.A(g14478), .Z(II25047) ) ;
INV     gate9899  (.A(II25047), .Z(g18985) ) ;
INV     gate9900  (.A(g14601), .Z(II25050) ) ;
INV     gate9901  (.A(II25050), .Z(g18986) ) ;
INV     gate9902  (.A(g15794), .Z(g18987) ) ;
INV     gate9903  (.A(g14837), .Z(II25054) ) ;
INV     gate9904  (.A(II25054), .Z(g18988) ) ;
INV     gate9905  (.A(g14186), .Z(II25057) ) ;
INV     gate9906  (.A(II25057), .Z(g18989) ) ;
INV     gate9907  (.A(g14976), .Z(II25061) ) ;
INV     gate9908  (.A(II25061), .Z(g18991) ) ;
INV     gate9909  (.A(g14395), .Z(II25064) ) ;
INV     gate9910  (.A(II25064), .Z(g18992) ) ;
INV     gate9911  (.A(g14565), .Z(II25067) ) ;
INV     gate9912  (.A(II25067), .Z(g18993) ) ;
INV     gate9913  (.A(g14910), .Z(II25071) ) ;
INV     gate9914  (.A(II25071), .Z(g18995) ) ;
INV     gate9915  (.A(g14301), .Z(II25074) ) ;
INV     gate9916  (.A(II25074), .Z(g18996) ) ;
INV     gate9917  (.A(g15065), .Z(II25078) ) ;
INV     gate9918  (.A(II25078), .Z(g18998) ) ;
INV     gate9919  (.A(g14507), .Z(II25081) ) ;
INV     gate9920  (.A(II25081), .Z(g18999) ) ;
INV     gate9921  (.A(g14885), .Z(II25084) ) ;
INV     gate9922  (.A(II25084), .Z(g19000) ) ;
INV     gate9923  (.A(g14071), .Z(g19001) ) ;
INV     gate9924  (.A(g14991), .Z(II25089) ) ;
INV     gate9925  (.A(II25089), .Z(g19008) ) ;
INV     gate9926  (.A(g14423), .Z(II25092) ) ;
INV     gate9927  (.A(II25092), .Z(g19009) ) ;
INV     gate9928  (.A(g15161), .Z(II25096) ) ;
INV     gate9929  (.A(II25096), .Z(g19011) ) ;
INV     gate9930  (.A(g19000), .Z(II25099) ) ;
INV     gate9931  (.A(g18944), .Z(II25102) ) ;
INV     gate9932  (.A(g18959), .Z(II25105) ) ;
INV     gate9933  (.A(g18969), .Z(II25108) ) ;
INV     gate9934  (.A(g18981), .Z(II25111) ) ;
INV     gate9935  (.A(g18983), .Z(II25114) ) ;
INV     gate9936  (.A(g18988), .Z(II25117) ) ;
INV     gate9937  (.A(g18869), .Z(II25120) ) ;
INV     gate9938  (.A(g18890), .Z(II25123) ) ;
INV     gate9939  (.A(g16858), .Z(II25126) ) ;
INV     gate9940  (.A(g16813), .Z(II25129) ) ;
INV     gate9941  (.A(g16862), .Z(II25132) ) ;
INV     gate9942  (.A(g16506), .Z(II25135) ) ;
INV     gate9943  (.A(g18960), .Z(II25138) ) ;
INV     gate9944  (.A(g18970), .Z(II25141) ) ;
INV     gate9945  (.A(g18984), .Z(II25144) ) ;
INV     gate9946  (.A(g18989), .Z(II25147) ) ;
INV     gate9947  (.A(g18991), .Z(II25150) ) ;
INV     gate9948  (.A(g18995), .Z(II25153) ) ;
INV     gate9949  (.A(g18895), .Z(II25156) ) ;
INV     gate9950  (.A(g18913), .Z(II25159) ) ;
INV     gate9951  (.A(g16863), .Z(II25162) ) ;
INV     gate9952  (.A(g16831), .Z(II25165) ) ;
INV     gate9953  (.A(g16877), .Z(II25168) ) ;
INV     gate9954  (.A(g16528), .Z(II25171) ) ;
INV     gate9955  (.A(g18971), .Z(II25174) ) ;
INV     gate9956  (.A(g18985), .Z(II25177) ) ;
INV     gate9957  (.A(g18992), .Z(II25180) ) ;
INV     gate9958  (.A(g18996), .Z(II25183) ) ;
INV     gate9959  (.A(g18998), .Z(II25186) ) ;
INV     gate9960  (.A(g19008), .Z(II25189) ) ;
INV     gate9961  (.A(g18918), .Z(II25192) ) ;
INV     gate9962  (.A(g18932), .Z(II25195) ) ;
INV     gate9963  (.A(g16878), .Z(II25198) ) ;
INV     gate9964  (.A(g16843), .Z(II25201) ) ;
INV     gate9965  (.A(g16905), .Z(II25204) ) ;
INV     gate9966  (.A(g16559), .Z(II25207) ) ;
INV     gate9967  (.A(g18986), .Z(II25210) ) ;
INV     gate9968  (.A(g18993), .Z(II25213) ) ;
INV     gate9969  (.A(g18999), .Z(II25216) ) ;
INV     gate9970  (.A(g19009), .Z(II25219) ) ;
INV     gate9971  (.A(g19011), .Z(II25222) ) ;
INV     gate9972  (.A(g16514), .Z(II25225) ) ;
INV     gate9973  (.A(g18937), .Z(II25228) ) ;
INV     gate9974  (.A(g18952), .Z(II25231) ) ;
INV     gate9975  (.A(g16906), .Z(II25234) ) ;
INV     gate9976  (.A(g16849), .Z(II25237) ) ;
INV     gate9977  (.A(g16934), .Z(II25240) ) ;
INV     gate9978  (.A(g17227), .Z(II25243) ) ;
INV     gate9979  (.A(g17233), .Z(II25246) ) ;
INV     gate9980  (.A(g17300), .Z(II25249) ) ;
NOR3    gate9981  (.A(g14725), .B(g15942), .C(g14677), .Z(g17124) ) ;
INV     gate9982  (.A(g17124), .Z(II25253) ) ;
INV     gate9983  (.A(II25253), .Z(g19064) ) ;
INV     gate9984  (.A(g18583), .Z(g19070) ) ;
INV     gate9985  (.A(g16974), .Z(II25258) ) ;
INV     gate9986  (.A(II25258), .Z(g19075) ) ;
INV     gate9987  (.A(g18619), .Z(g19078) ) ;
NOR3    gate9988  (.A(g14753), .B(g15971), .C(g14711), .Z(g17151) ) ;
INV     gate9989  (.A(g17151), .Z(II25264) ) ;
INV     gate9990  (.A(II25264), .Z(g19081) ) ;
NOR3    gate9991  (.A(g14657), .B(g15880), .C(g14630), .Z(g17051) ) ;
INV     gate9992  (.A(g17051), .Z(II25272) ) ;
INV     gate9993  (.A(II25272), .Z(g19091) ) ;
NAND2   gate9994  (.A(II25031), .B(II25032), .Z(g18980) ) ;
INV     gate9995  (.A(g18980), .Z(g19096) ) ;
NOR3    gate9996  (.A(g14691), .B(g15913), .C(g14650), .Z(g17086) ) ;
INV     gate9997  (.A(g17086), .Z(II25283) ) ;
INV     gate9998  (.A(II25283), .Z(g19098) ) ;
INV     gate9999  (.A(g17124), .Z(II25294) ) ;
INV     gate10000  (.A(II25294), .Z(g19105) ) ;
INV     gate10001  (.A(g17151), .Z(II25303) ) ;
INV     gate10002  (.A(II25303), .Z(g19110) ) ;
INV     gate10003  (.A(g16867), .Z(II25308) ) ;
INV     gate10004  (.A(II25308), .Z(g19113) ) ;
INV     gate10005  (.A(g16895), .Z(II25315) ) ;
INV     gate10006  (.A(II25315), .Z(g19118) ) ;
INV     gate10007  (.A(g16924), .Z(II25320) ) ;
INV     gate10008  (.A(II25320), .Z(g19125) ) ;
INV     gate10009  (.A(g16954), .Z(II25325) ) ;
INV     gate10010  (.A(II25325), .Z(g19132) ) ;
INV     gate10011  (.A(g17645), .Z(II25334) ) ;
INV     gate10012  (.A(II25334), .Z(g19145) ) ;
INV     gate10013  (.A(g17746), .Z(II25338) ) ;
INV     gate10014  (.A(II25338), .Z(g19147) ) ;
INV     gate10015  (.A(g17847), .Z(II25344) ) ;
INV     gate10016  (.A(II25344), .Z(g19151) ) ;
INV     gate10017  (.A(g17959), .Z(II25351) ) ;
INV     gate10018  (.A(II25351), .Z(g19156) ) ;
NOR2    gate10019  (.A(g13623), .B(g13634), .Z(g18669) ) ;
INV     gate10020  (.A(g18669), .Z(II25355) ) ;
INV     gate10021  (.A(II25355), .Z(g19158) ) ;
NOR2    gate10022  (.A(g13625), .B(g11771), .Z(g18678) ) ;
INV     gate10023  (.A(g18678), .Z(II25358) ) ;
INV     gate10024  (.A(II25358), .Z(g19159) ) ;
NOR2    gate10025  (.A(g13636), .B(g11788), .Z(g18707) ) ;
INV     gate10026  (.A(g18707), .Z(II25365) ) ;
INV     gate10027  (.A(II25365), .Z(g19164) ) ;
NOR2    gate10028  (.A(g13643), .B(g13656), .Z(g18719) ) ;
INV     gate10029  (.A(g18719), .Z(II25371) ) ;
INV     gate10030  (.A(II25371), .Z(g19168) ) ;
NOR2    gate10031  (.A(g13645), .B(g11805), .Z(g18726) ) ;
INV     gate10032  (.A(g18726), .Z(II25374) ) ;
INV     gate10033  (.A(II25374), .Z(g19169) ) ;
NOR2    gate10034  (.A(g13648), .B(g11814), .Z(g18743) ) ;
INV     gate10035  (.A(g18743), .Z(II25377) ) ;
INV     gate10036  (.A(II25377), .Z(g19170) ) ;
NOR2    gate10037  (.A(g13871), .B(g12274), .Z(g18755) ) ;
INV     gate10038  (.A(g18755), .Z(II25383) ) ;
INV     gate10039  (.A(II25383), .Z(g19174) ) ;
NOR2    gate10040  (.A(g13671), .B(g11838), .Z(g18763) ) ;
INV     gate10041  (.A(g18763), .Z(II25386) ) ;
INV     gate10042  (.A(II25386), .Z(g19175) ) ;
NOR2    gate10043  (.A(g13674), .B(g11847), .Z(g18780) ) ;
INV     gate10044  (.A(g18780), .Z(II25389) ) ;
INV     gate10045  (.A(II25389), .Z(g19176) ) ;
NOR2    gate10046  (.A(g13676), .B(g13705), .Z(g18782) ) ;
INV     gate10047  (.A(g18782), .Z(II25395) ) ;
INV     gate10048  (.A(II25395), .Z(g19180) ) ;
NOR2    gate10049  (.A(g13701), .B(g11880), .Z(g18794) ) ;
INV     gate10050  (.A(g18794), .Z(II25399) ) ;
INV     gate10051  (.A(II25399), .Z(g19182) ) ;
NOR2    gate10052  (.A(g13740), .B(g11926), .Z(g18821) ) ;
INV     gate10053  (.A(g18821), .Z(II25402) ) ;
INV     gate10054  (.A(II25402), .Z(g19183) ) ;
NOR2    gate10055  (.A(g13905), .B(g12331), .Z(g18804) ) ;
INV     gate10056  (.A(g18804), .Z(II25406) ) ;
INV     gate10057  (.A(II25406), .Z(g19185) ) ;
NOR2    gate10058  (.A(g13738), .B(g11922), .Z(g18820) ) ;
INV     gate10059  (.A(g18820), .Z(II25412) ) ;
INV     gate10060  (.A(II25412), .Z(g19189) ) ;
NOR2    gate10061  (.A(g13788), .B(g11966), .Z(g18835) ) ;
INV     gate10062  (.A(g18835), .Z(II25415) ) ;
INV     gate10063  (.A(II25415), .Z(g19190) ) ;
NOR2    gate10064  (.A(g13815), .B(g12012), .Z(g18852) ) ;
INV     gate10065  (.A(g18852), .Z(II25423) ) ;
INV     gate10066  (.A(II25423), .Z(g19196) ) ;
NOR2    gate10067  (.A(g13789), .B(g11967), .Z(g18836) ) ;
INV     gate10068  (.A(g18836), .Z(II25426) ) ;
INV     gate10069  (.A(II25426), .Z(g19197) ) ;
NOR2    gate10070  (.A(g13944), .B(g12353), .Z(g18975) ) ;
INV     gate10071  (.A(g18975), .Z(II25429) ) ;
INV     gate10072  (.A(II25429), .Z(g19198) ) ;
NOR2    gate10073  (.A(g13998), .B(g12376), .Z(g18837) ) ;
INV     gate10074  (.A(g18837), .Z(II25432) ) ;
INV     gate10075  (.A(II25432), .Z(g19199) ) ;
NOR2    gate10076  (.A(g13834), .B(g12069), .Z(g18866) ) ;
INV     gate10077  (.A(g18866), .Z(II25442) ) ;
INV     gate10078  (.A(II25442), .Z(g19207) ) ;
NOR2    gate10079  (.A(g13904), .B(g12330), .Z(g18968) ) ;
INV     gate10080  (.A(g18968), .Z(II25445) ) ;
INV     gate10081  (.A(II25445), .Z(g19208) ) ;
NOR2    gate10082  (.A(g13846), .B(g12128), .Z(g18883) ) ;
INV     gate10083  (.A(g18883), .Z(II25456) ) ;
INV     gate10084  (.A(II25456), .Z(g19217) ) ;
NOR2    gate10085  (.A(g13835), .B(g12070), .Z(g18867) ) ;
INV     gate10086  (.A(g18867), .Z(II25459) ) ;
INV     gate10087  (.A(II25459), .Z(g19218) ) ;
NOR2    gate10088  (.A(g14143), .B(g12419), .Z(g18868) ) ;
INV     gate10089  (.A(g18868), .Z(II25463) ) ;
INV     gate10090  (.A(II25463), .Z(g19220) ) ;
NOR2    gate10091  (.A(g13847), .B(g12129), .Z(g18885) ) ;
INV     gate10092  (.A(g18885), .Z(II25474) ) ;
INV     gate10093  (.A(II25474), .Z(g19229) ) ;
NOR2    gate10094  (.A(g13655), .B(g11816), .Z(g18754) ) ;
INV     gate10095  (.A(g18754), .Z(II25486) ) ;
INV     gate10096  (.A(II25486), .Z(g19237) ) ;
NOR2    gate10097  (.A(g13855), .B(g12186), .Z(g18906) ) ;
INV     gate10098  (.A(g18906), .Z(II25489) ) ;
INV     gate10099  (.A(II25489), .Z(g19238) ) ;
NOR2    gate10100  (.A(g14336), .B(g12429), .Z(g18907) ) ;
INV     gate10101  (.A(g18907), .Z(II25492) ) ;
INV     gate10102  (.A(II25492), .Z(g19239) ) ;
NOR2    gate10103  (.A(g13675), .B(g11851), .Z(g18781) ) ;
INV     gate10104  (.A(g18781), .Z(II25506) ) ;
INV     gate10105  (.A(II25506), .Z(g19247) ) ;
NAND2   gate10106  (.A(II24612), .B(II24613), .Z(g18542) ) ;
INV     gate10107  (.A(g18542), .Z(II25510) ) ;
INV     gate10108  (.A(II25510), .Z(g19249) ) ;
INV     gate10109  (.A(g16540), .Z(g19251) ) ;
NOR2    gate10110  (.A(g13704), .B(g11885), .Z(g18803) ) ;
INV     gate10111  (.A(g18803), .Z(II25525) ) ;
INV     gate10112  (.A(II25525), .Z(g19258) ) ;
NOR2    gate10113  (.A(g13870), .B(g12273), .Z(g18942) ) ;
INV     gate10114  (.A(g18942), .Z(II25528) ) ;
INV     gate10115  (.A(II25528), .Z(g19259) ) ;
INV     gate10116  (.A(g16572), .Z(g19265) ) ;
NOR2    gate10117  (.A(g13884), .B(g12307), .Z(g18957) ) ;
INV     gate10118  (.A(g18957), .Z(II25557) ) ;
INV     gate10119  (.A(II25557), .Z(g19270) ) ;
NOR2    gate10120  (.A(g7949), .B(g14144), .Z(g17186) ) ;
INV     gate10121  (.A(g17186), .Z(II25567) ) ;
INV     gate10122  (.A(II25567), .Z(g19272) ) ;
INV     gate10123  (.A(g16596), .Z(g19280) ) ;
INV     gate10124  (.A(g16608), .Z(g19287) ) ;
NOR2    gate10125  (.A(g8000), .B(g14259), .Z(g17197) ) ;
INV     gate10126  (.A(g17197), .Z(II25612) ) ;
INV     gate10127  (.A(II25612), .Z(g19291) ) ;
INV     gate10128  (.A(g16616), .Z(g19299) ) ;
INV     gate10129  (.A(g16622), .Z(g19301) ) ;
NOR3    gate10130  (.A(g15904), .B(g15880), .C(g15859), .Z(g17025) ) ;
INV     gate10131  (.A(g17025), .Z(g19302) ) ;
INV     gate10132  (.A(g16626), .Z(g19305) ) ;
NOR2    gate10133  (.A(g8075), .B(g14381), .Z(g17204) ) ;
INV     gate10134  (.A(g17204), .Z(II25660) ) ;
INV     gate10135  (.A(II25660), .Z(g19309) ) ;
INV     gate10136  (.A(g16633), .Z(g19319) ) ;
INV     gate10137  (.A(g16636), .Z(g19322) ) ;
NOR3    gate10138  (.A(g15933), .B(g15913), .C(g15890), .Z(g17059) ) ;
INV     gate10139  (.A(g17059), .Z(g19323) ) ;
INV     gate10140  (.A(g16640), .Z(g19326) ) ;
NOR2    gate10141  (.A(g8160), .B(g14493), .Z(g17209) ) ;
INV     gate10142  (.A(g17209), .Z(II25717) ) ;
INV     gate10143  (.A(II25717), .Z(g19330) ) ;
NAND2   gate10144  (.A(g13915), .B(g13893), .Z(g17118) ) ;
INV     gate10145  (.A(g17118), .Z(II25728) ) ;
INV     gate10146  (.A(II25728), .Z(g19335) ) ;
INV     gate10147  (.A(g16644), .Z(g19346) ) ;
INV     gate10148  (.A(g16647), .Z(g19349) ) ;
NOR3    gate10149  (.A(g15962), .B(g15942), .C(g15923), .Z(g17094) ) ;
INV     gate10150  (.A(g17094), .Z(g19350) ) ;
INV     gate10151  (.A(g16651), .Z(g19353) ) ;
NAND2   gate10152  (.A(g13957), .B(g13915), .Z(g17139) ) ;
INV     gate10153  (.A(g17139), .Z(II25768) ) ;
INV     gate10154  (.A(II25768), .Z(g19358) ) ;
NAND2   gate10155  (.A(g13971), .B(g13934), .Z(g17145) ) ;
INV     gate10156  (.A(g17145), .Z(II25778) ) ;
INV     gate10157  (.A(II25778), .Z(g19369) ) ;
INV     gate10158  (.A(g16656), .Z(g19380) ) ;
INV     gate10159  (.A(g16659), .Z(g19383) ) ;
NOR3    gate10160  (.A(g15981), .B(g15971), .C(g15952), .Z(g17132) ) ;
INV     gate10161  (.A(g17132), .Z(g19384) ) ;
NOR3    gate10162  (.A(g15904), .B(g15880), .C(g15859), .Z(g16567) ) ;
INV     gate10163  (.A(g16567), .Z(g19387) ) ;
INV     gate10164  (.A(g17139), .Z(g19388) ) ;
NAND2   gate10165  (.A(g14027), .B(g13971), .Z(g17162) ) ;
INV     gate10166  (.A(g17162), .Z(II25816) ) ;
INV     gate10167  (.A(II25816), .Z(g19390) ) ;
NAND2   gate10168  (.A(g14041), .B(g13990), .Z(g17168) ) ;
INV     gate10169  (.A(g17168), .Z(II25826) ) ;
INV     gate10170  (.A(II25826), .Z(g19401) ) ;
INV     gate10171  (.A(g16673), .Z(g19412) ) ;
INV     gate10172  (.A(g16676), .Z(g19415) ) ;
NOR3    gate10173  (.A(g15933), .B(g15913), .C(g15890), .Z(g16591) ) ;
INV     gate10174  (.A(g16591), .Z(g19417) ) ;
INV     gate10175  (.A(g17162), .Z(g19418) ) ;
NAND2   gate10176  (.A(g14118), .B(g14041), .Z(g17177) ) ;
INV     gate10177  (.A(g17177), .Z(II25862) ) ;
INV     gate10178  (.A(II25862), .Z(g19420) ) ;
NAND2   gate10179  (.A(g14132), .B(g14060), .Z(g17183) ) ;
INV     gate10180  (.A(g17183), .Z(II25872) ) ;
INV     gate10181  (.A(II25872), .Z(g19431) ) ;
NOR2    gate10182  (.A(g4326), .B(g14442), .Z(g17213) ) ;
INV     gate10183  (.A(g17213), .Z(g19441) ) ;
NAND2   gate10184  (.A(g14641), .B(g9636), .Z(g17985) ) ;
INV     gate10185  (.A(g17985), .Z(g19444) ) ;
INV     gate10186  (.A(g16694), .Z(g19448) ) ;
INV     gate10187  (.A(g16702), .Z(g19452) ) ;
NOR3    gate10188  (.A(g15962), .B(g15942), .C(g15923), .Z(g16611) ) ;
INV     gate10189  (.A(g16611), .Z(g19454) ) ;
INV     gate10190  (.A(g17177), .Z(g19455) ) ;
NAND2   gate10191  (.A(g14233), .B(g14132), .Z(g17194) ) ;
INV     gate10192  (.A(g17194), .Z(II25904) ) ;
INV     gate10193  (.A(II25904), .Z(g19457) ) ;
INV     gate10194  (.A(g16719), .Z(g19467) ) ;
NOR2    gate10195  (.A(g4495), .B(g14529), .Z(g17216) ) ;
INV     gate10196  (.A(g17216), .Z(g19468) ) ;
NAND2   gate10197  (.A(g14668), .B(g9782), .Z(g18102) ) ;
INV     gate10198  (.A(g18102), .Z(g19471) ) ;
INV     gate10199  (.A(g16725), .Z(g19475) ) ;
INV     gate10200  (.A(g16733), .Z(g19479) ) ;
NOR3    gate10201  (.A(g15981), .B(g15971), .C(g15952), .Z(g16629) ) ;
INV     gate10202  (.A(g16629), .Z(g19481) ) ;
INV     gate10203  (.A(g17194), .Z(g19482) ) ;
INV     gate10204  (.A(g16758), .Z(g19483) ) ;
INV     gate10205  (.A(g16867), .Z(g19484) ) ;
INV     gate10206  (.A(g16761), .Z(g19490) ) ;
NOR2    gate10207  (.A(g4671), .B(g14584), .Z(g17219) ) ;
INV     gate10208  (.A(g17219), .Z(g19491) ) ;
NAND2   gate10209  (.A(g14702), .B(g9928), .Z(g18218) ) ;
INV     gate10210  (.A(g18218), .Z(g19494) ) ;
INV     gate10211  (.A(g16767), .Z(g19498) ) ;
INV     gate10212  (.A(g16775), .Z(g19502) ) ;
INV     gate10213  (.A(g16785), .Z(g19504) ) ;
INV     gate10214  (.A(g16895), .Z(g19505) ) ;
INV     gate10215  (.A(g16788), .Z(g19511) ) ;
NOR2    gate10216  (.A(g4848), .B(g14618), .Z(g17221) ) ;
INV     gate10217  (.A(g17221), .Z(g19512) ) ;
NAND2   gate10218  (.A(g14736), .B(g10082), .Z(g18325) ) ;
INV     gate10219  (.A(g18325), .Z(g19515) ) ;
INV     gate10220  (.A(g16794), .Z(g19519) ) ;
INV     gate10221  (.A(g16814), .Z(g19523) ) ;
INV     gate10222  (.A(g16924), .Z(g19524) ) ;
INV     gate10223  (.A(g16817), .Z(g19530) ) ;
INV     gate10224  (.A(g16832), .Z(g19533) ) ;
INV     gate10225  (.A(g16954), .Z(g19534) ) ;
NOR2    gate10226  (.A(g14690), .B(g12477), .Z(g16654) ) ;
INV     gate10227  (.A(g16654), .Z(II25966) ) ;
INV     gate10228  (.A(II25966), .Z(g19543) ) ;
NOR2    gate10229  (.A(g14724), .B(g12494), .Z(g16671) ) ;
INV     gate10230  (.A(g16671), .Z(II25971) ) ;
INV     gate10231  (.A(II25971), .Z(g19546) ) ;
NOR2    gate10232  (.A(g14752), .B(g12514), .Z(g16692) ) ;
INV     gate10233  (.A(g16692), .Z(II25977) ) ;
INV     gate10234  (.A(II25977), .Z(g19550) ) ;
NOR2    gate10235  (.A(g14773), .B(g12531), .Z(g16718) ) ;
INV     gate10236  (.A(g16718), .Z(II25985) ) ;
INV     gate10237  (.A(II25985), .Z(g19556) ) ;
NOR2    gate10238  (.A(g15828), .B(g13031), .Z(g16860) ) ;
INV     gate10239  (.A(g16860), .Z(II25994) ) ;
INV     gate10240  (.A(II25994), .Z(g19563) ) ;
NOR2    gate10241  (.A(g15840), .B(g13042), .Z(g16866) ) ;
INV     gate10242  (.A(g16866), .Z(II26006) ) ;
INV     gate10243  (.A(II26006), .Z(g19573) ) ;
INV     gate10244  (.A(g16881), .Z(g19577) ) ;
INV     gate10245  (.A(g16884), .Z(g19578) ) ;
NOR2    gate10246  (.A(g15593), .B(g12908), .Z(g16803) ) ;
INV     gate10247  (.A(g16803), .Z(II26025) ) ;
INV     gate10248  (.A(II26025), .Z(g19595) ) ;
NAND2   gate10249  (.A(II22631), .B(II22632), .Z(g16566) ) ;
INV     gate10250  (.A(g16566), .Z(II26028) ) ;
INV     gate10251  (.A(II26028), .Z(g19596) ) ;
INV     gate10252  (.A(g16910), .Z(g19607) ) ;
INV     gate10253  (.A(g16913), .Z(g19608) ) ;
NOR2    gate10254  (.A(g15658), .B(g12938), .Z(g16824) ) ;
INV     gate10255  (.A(g16824), .Z(II26051) ) ;
INV     gate10256  (.A(II26051), .Z(g19622) ) ;
INV     gate10257  (.A(g16940), .Z(g19640) ) ;
INV     gate10258  (.A(g16943), .Z(g19641) ) ;
NOR2    gate10259  (.A(g15717), .B(g12966), .Z(g16835) ) ;
INV     gate10260  (.A(g16835), .Z(II26078) ) ;
INV     gate10261  (.A(II26078), .Z(g19652) ) ;
NOR2    gate10262  (.A(g16085), .B(g6363), .Z(g18085) ) ;
INV     gate10263  (.A(g18085), .Z(II26085) ) ;
INV     gate10264  (.A(II26085), .Z(g19657) ) ;
INV     gate10265  (.A(g16971), .Z(g19680) ) ;
INV     gate10266  (.A(g16974), .Z(g19681) ) ;
NOR2    gate10267  (.A(g15754), .B(g12989), .Z(g16844) ) ;
INV     gate10268  (.A(g16844), .Z(II26112) ) ;
INV     gate10269  (.A(II26112), .Z(g19689) ) ;
NOR2    gate10270  (.A(g15755), .B(g12990), .Z(g16845) ) ;
INV     gate10271  (.A(g16845), .Z(II26115) ) ;
INV     gate10272  (.A(II26115), .Z(g19690) ) ;
INV     gate10273  (.A(g17503), .Z(II26123) ) ;
INV     gate10274  (.A(II26123), .Z(g19696) ) ;
NOR2    gate10275  (.A(g16123), .B(g6568), .Z(g18201) ) ;
INV     gate10276  (.A(g18201), .Z(II26134) ) ;
INV     gate10277  (.A(II26134), .Z(g19705) ) ;
NOR2    gate10278  (.A(g15781), .B(g13000), .Z(g16851) ) ;
INV     gate10279  (.A(g16851), .Z(II26154) ) ;
INV     gate10280  (.A(II26154), .Z(g19725) ) ;
INV     gate10281  (.A(g17594), .Z(II26171) ) ;
INV     gate10282  (.A(II26171), .Z(g19740) ) ;
NOR2    gate10283  (.A(g16174), .B(g6832), .Z(g18308) ) ;
INV     gate10284  (.A(g18308), .Z(II26182) ) ;
INV     gate10285  (.A(II26182), .Z(g19749) ) ;
NOR2    gate10286  (.A(g15801), .B(g13009), .Z(g16853) ) ;
INV     gate10287  (.A(g16853), .Z(II26195) ) ;
INV     gate10288  (.A(II26195), .Z(g19762) ) ;
NOR2    gate10289  (.A(g15802), .B(g13010), .Z(g16854) ) ;
INV     gate10290  (.A(g16854), .Z(II26198) ) ;
INV     gate10291  (.A(II26198), .Z(g19763) ) ;
INV     gate10292  (.A(g17691), .Z(II26220) ) ;
INV     gate10293  (.A(II26220), .Z(g19783) ) ;
NOR2    gate10294  (.A(g16233), .B(g7134), .Z(g18401) ) ;
INV     gate10295  (.A(g18401), .Z(II26231) ) ;
INV     gate10296  (.A(II26231), .Z(g19792) ) ;
NOR2    gate10297  (.A(g15817), .B(g13023), .Z(g16857) ) ;
INV     gate10298  (.A(g16857), .Z(II26237) ) ;
INV     gate10299  (.A(II26237), .Z(g19798) ) ;
INV     gate10300  (.A(g17791), .Z(II26266) ) ;
INV     gate10301  (.A(II26266), .Z(g19825) ) ;
INV     gate10302  (.A(g18886), .Z(g19830) ) ;
NOR2    gate10303  (.A(g15829), .B(g13032), .Z(g16861) ) ;
INV     gate10304  (.A(g16861), .Z(II26276) ) ;
INV     gate10305  (.A(II26276), .Z(g19838) ) ;
NAND2   gate10306  (.A(g15797), .B(g3006), .Z(g18977) ) ;
INV     gate10307  (.A(g18977), .Z(II26334) ) ;
INV     gate10308  (.A(II26334), .Z(g19890) ) ;
NOR2    gate10309  (.A(g15852), .B(g13056), .Z(g16880) ) ;
INV     gate10310  (.A(g16880), .Z(II26337) ) ;
INV     gate10311  (.A(II26337), .Z(g19893) ) ;
INV     gate10312  (.A(g17025), .Z(II26340) ) ;
INV     gate10313  (.A(II26340), .Z(g19894) ) ;
NOR2    gate10314  (.A(g16463), .B(g7549), .Z(g18626) ) ;
INV     gate10315  (.A(g18626), .Z(II26365) ) ;
INV     gate10316  (.A(II26365), .Z(g19915) ) ;
INV     gate10317  (.A(g18646), .Z(g19918) ) ;
INV     gate10318  (.A(g17059), .Z(II26369) ) ;
INV     gate10319  (.A(II26369), .Z(g19919) ) ;
NOR2    gate10320  (.A(g14249), .B(g16082), .Z(g18548) ) ;
INV     gate10321  (.A(g18548), .Z(g19933) ) ;
INV     gate10322  (.A(g17094), .Z(II26388) ) ;
INV     gate10323  (.A(II26388), .Z(g19934) ) ;
NOR3    gate10324  (.A(g14657), .B(g14642), .C(g15859), .Z(g17012) ) ;
INV     gate10325  (.A(g17012), .Z(II26401) ) ;
INV     gate10326  (.A(II26401), .Z(g19945) ) ;
NOR2    gate10327  (.A(g14352), .B(g16020), .Z(g17896) ) ;
INV     gate10328  (.A(g17896), .Z(g19948) ) ;
NOR2    gate10329  (.A(g14371), .B(g16120), .Z(g18598) ) ;
INV     gate10330  (.A(g18598), .Z(g19950) ) ;
INV     gate10331  (.A(g17132), .Z(II26407) ) ;
INV     gate10332  (.A(II26407), .Z(g19951) ) ;
NOR3    gate10333  (.A(g15904), .B(g14642), .C(g15859), .Z(g16643) ) ;
INV     gate10334  (.A(g16643), .Z(II26413) ) ;
INV     gate10335  (.A(II26413), .Z(g19957) ) ;
NOR3    gate10336  (.A(g14691), .B(g14669), .C(g15890), .Z(g17042) ) ;
INV     gate10337  (.A(g17042), .Z(II26420) ) ;
INV     gate10338  (.A(II26420), .Z(g19972) ) ;
NOR2    gate10339  (.A(g14464), .B(g16036), .Z(g18007) ) ;
INV     gate10340  (.A(g18007), .Z(g19975) ) ;
NOR2    gate10341  (.A(g14483), .B(g16171), .Z(g18630) ) ;
INV     gate10342  (.A(g18630), .Z(g19977) ) ;
NAND2   gate10343  (.A(g15873), .B(g2896), .Z(g16536) ) ;
INV     gate10344  (.A(g16536), .Z(II26426) ) ;
INV     gate10345  (.A(II26426), .Z(g19978) ) ;
NOR3    gate10346  (.A(g15933), .B(g14669), .C(g15890), .Z(g16655) ) ;
INV     gate10347  (.A(g16655), .Z(II26437) ) ;
INV     gate10348  (.A(II26437), .Z(g19987) ) ;
NOR3    gate10349  (.A(g14725), .B(g14703), .C(g15923), .Z(g17076) ) ;
INV     gate10350  (.A(g17076), .Z(II26444) ) ;
INV     gate10351  (.A(II26444), .Z(g20002) ) ;
NOR2    gate10352  (.A(g14551), .B(g16058), .Z(g18124) ) ;
INV     gate10353  (.A(g18124), .Z(g20005) ) ;
NOR2    gate10354  (.A(g14570), .B(g16230), .Z(g18639) ) ;
INV     gate10355  (.A(g18639), .Z(g20007) ) ;
INV     gate10356  (.A(g17985), .Z(II26458) ) ;
INV     gate10357  (.A(II26458), .Z(g20016) ) ;
NOR3    gate10358  (.A(g15962), .B(g14703), .C(g15923), .Z(g16672) ) ;
INV     gate10359  (.A(g16672), .Z(II26469) ) ;
INV     gate10360  (.A(II26469), .Z(g20025) ) ;
NOR3    gate10361  (.A(g14753), .B(g14737), .C(g15952), .Z(g17111) ) ;
INV     gate10362  (.A(g17111), .Z(II26476) ) ;
INV     gate10363  (.A(II26476), .Z(g20040) ) ;
NOR2    gate10364  (.A(g14606), .B(g16094), .Z(g18240) ) ;
INV     gate10365  (.A(g18240), .Z(g20043) ) ;
NOR2    gate10366  (.A(g16439), .B(g7522), .Z(g18590) ) ;
INV     gate10367  (.A(g18590), .Z(II26481) ) ;
INV     gate10368  (.A(II26481), .Z(g20045) ) ;
INV     gate10369  (.A(g18102), .Z(II26494) ) ;
INV     gate10370  (.A(II26494), .Z(g20058) ) ;
NOR3    gate10371  (.A(g15981), .B(g14737), .C(g15952), .Z(g16693) ) ;
INV     gate10372  (.A(g16693), .Z(II26505) ) ;
INV     gate10373  (.A(II26505), .Z(g20067) ) ;
NOR2    gate10374  (.A(g13469), .B(g3897), .Z(g16802) ) ;
INV     gate10375  (.A(g16802), .Z(II26512) ) ;
INV     gate10376  (.A(II26512), .Z(g20082) ) ;
NAND2   gate10377  (.A(II24006), .B(II24007), .Z(g17968) ) ;
INV     gate10378  (.A(g17968), .Z(g20083) ) ;
INV     gate10379  (.A(g18218), .Z(II26535) ) ;
INV     gate10380  (.A(II26535), .Z(g20099) ) ;
NOR2    gate10381  (.A(g5362), .B(g13469), .Z(g16823) ) ;
INV     gate10382  (.A(g16823), .Z(II26545) ) ;
INV     gate10383  (.A(II26545), .Z(g20105) ) ;
INV     gate10384  (.A(g18325), .Z(II26574) ) ;
INV     gate10385  (.A(II26574), .Z(g20124) ) ;
NOR2    gate10386  (.A(g15902), .B(g2814), .Z(g18623) ) ;
INV     gate10387  (.A(g18623), .Z(g20127) ) ;
INV     gate10388  (.A(g16830), .Z(g20140) ) ;
OR2     gate10389  (.A(g11623), .B(g15659), .Z(g17973) ) ;
INV     gate10390  (.A(g17973), .Z(g20163) ) ;
INV     gate10391  (.A(g17645), .Z(II26612) ) ;
INV     gate10392  (.A(II26612), .Z(g20164) ) ;
INV     gate10393  (.A(g16842), .Z(g20178) ) ;
INV     gate10394  (.A(g18691), .Z(g20193) ) ;
INV     gate10395  (.A(g17746), .Z(II26642) ) ;
INV     gate10396  (.A(II26642), .Z(g20198) ) ;
INV     gate10397  (.A(g16848), .Z(g20212) ) ;
INV     gate10398  (.A(g18727), .Z(g20223) ) ;
INV     gate10399  (.A(g17847), .Z(II26664) ) ;
INV     gate10400  (.A(II26664), .Z(g20228) ) ;
INV     gate10401  (.A(g16852), .Z(g20242) ) ;
INV     gate10402  (.A(g18764), .Z(g20250) ) ;
INV     gate10403  (.A(g17959), .Z(II26679) ) ;
INV     gate10404  (.A(II26679), .Z(g20255) ) ;
INV     gate10405  (.A(g17230), .Z(g20269) ) ;
INV     gate10406  (.A(g18795), .Z(g20273) ) ;
INV     gate10407  (.A(g17237), .Z(g20278) ) ;
INV     gate10408  (.A(g17240), .Z(g20279) ) ;
INV     gate10409  (.A(g17243), .Z(g20281) ) ;
INV     gate10410  (.A(g17249), .Z(g20286) ) ;
INV     gate10411  (.A(g17252), .Z(g20287) ) ;
INV     gate10412  (.A(g17255), .Z(g20288) ) ;
INV     gate10413  (.A(g17259), .Z(g20289) ) ;
INV     gate10414  (.A(g17262), .Z(g20290) ) ;
INV     gate10415  (.A(g17265), .Z(g20292) ) ;
INV     gate10416  (.A(g17720), .Z(II26714) ) ;
INV     gate10417  (.A(II26714), .Z(g20295) ) ;
INV     gate10418  (.A(g17272), .Z(g20296) ) ;
INV     gate10419  (.A(g17275), .Z(g20297) ) ;
INV     gate10420  (.A(g17278), .Z(g20298) ) ;
INV     gate10421  (.A(g17282), .Z(g20302) ) ;
INV     gate10422  (.A(g17285), .Z(g20303) ) ;
INV     gate10423  (.A(g17288), .Z(g20304) ) ;
INV     gate10424  (.A(g17291), .Z(g20305) ) ;
INV     gate10425  (.A(g17294), .Z(g20306) ) ;
INV     gate10426  (.A(g17297), .Z(g20308) ) ;
INV     gate10427  (.A(g17304), .Z(g20311) ) ;
INV     gate10428  (.A(g17307), .Z(g20312) ) ;
INV     gate10429  (.A(g17310), .Z(g20313) ) ;
INV     gate10430  (.A(g17315), .Z(g20315) ) ;
INV     gate10431  (.A(g17318), .Z(g20316) ) ;
INV     gate10432  (.A(g17321), .Z(g20317) ) ;
INV     gate10433  (.A(g17324), .Z(g20321) ) ;
INV     gate10434  (.A(g17327), .Z(g20322) ) ;
INV     gate10435  (.A(g17330), .Z(g20323) ) ;
INV     gate10436  (.A(g17333), .Z(g20324) ) ;
INV     gate10437  (.A(g17336), .Z(g20325) ) ;
INV     gate10438  (.A(g17342), .Z(g20327) ) ;
INV     gate10439  (.A(g17345), .Z(g20328) ) ;
INV     gate10440  (.A(g17348), .Z(g20329) ) ;
INV     gate10441  (.A(g17354), .Z(g20330) ) ;
INV     gate10442  (.A(g17357), .Z(g20331) ) ;
INV     gate10443  (.A(g17360), .Z(g20332) ) ;
INV     gate10444  (.A(g17363), .Z(g20334) ) ;
INV     gate10445  (.A(g17366), .Z(g20335) ) ;
INV     gate10446  (.A(g17369), .Z(g20336) ) ;
INV     gate10447  (.A(g17372), .Z(g20340) ) ;
INV     gate10448  (.A(g17375), .Z(g20341) ) ;
INV     gate10449  (.A(g17378), .Z(g20342) ) ;
INV     gate10450  (.A(g17384), .Z(g20344) ) ;
INV     gate10451  (.A(g17387), .Z(g20345) ) ;
INV     gate10452  (.A(g17390), .Z(g20346) ) ;
INV     gate10453  (.A(g17399), .Z(g20347) ) ;
INV     gate10454  (.A(g17402), .Z(g20348) ) ;
INV     gate10455  (.A(g17405), .Z(g20349) ) ;
INV     gate10456  (.A(g17410), .Z(g20350) ) ;
INV     gate10457  (.A(g17413), .Z(g20351) ) ;
INV     gate10458  (.A(g17416), .Z(g20352) ) ;
INV     gate10459  (.A(g17419), .Z(g20354) ) ;
INV     gate10460  (.A(g17422), .Z(g20355) ) ;
INV     gate10461  (.A(g17425), .Z(g20356) ) ;
NOR2    gate10462  (.A(g15998), .B(g16003), .Z(g17222) ) ;
INV     gate10463  (.A(g17222), .Z(II26777) ) ;
INV     gate10464  (.A(II26777), .Z(g20360) ) ;
INV     gate10465  (.A(g17430), .Z(g20361) ) ;
INV     gate10466  (.A(g17433), .Z(g20362) ) ;
INV     gate10467  (.A(g17436), .Z(g20363) ) ;
INV     gate10468  (.A(g17439), .Z(g20364) ) ;
INV     gate10469  (.A(g17442), .Z(g20365) ) ;
INV     gate10470  (.A(g17451), .Z(g20366) ) ;
INV     gate10471  (.A(g17454), .Z(g20367) ) ;
INV     gate10472  (.A(g17457), .Z(g20368) ) ;
INV     gate10473  (.A(g17465), .Z(g20369) ) ;
INV     gate10474  (.A(g17468), .Z(g20370) ) ;
INV     gate10475  (.A(g17471), .Z(g20371) ) ;
INV     gate10476  (.A(g17476), .Z(g20372) ) ;
INV     gate10477  (.A(g17479), .Z(g20373) ) ;
INV     gate10478  (.A(g17482), .Z(g20374) ) ;
NOR2    gate10479  (.A(g16004), .B(g16009), .Z(g17224) ) ;
INV     gate10480  (.A(g17224), .Z(II26796) ) ;
INV     gate10481  (.A(II26796), .Z(g20377) ) ;
INV     gate10482  (.A(g17487), .Z(g20378) ) ;
INV     gate10483  (.A(g17490), .Z(g20379) ) ;
INV     gate10484  (.A(g17493), .Z(g20380) ) ;
INV     gate10485  (.A(g17496), .Z(g20381) ) ;
INV     gate10486  (.A(g17500), .Z(g20382) ) ;
INV     gate10487  (.A(g17503), .Z(g20383) ) ;
INV     gate10488  (.A(g17511), .Z(g20384) ) ;
INV     gate10489  (.A(g17514), .Z(g20385) ) ;
INV     gate10490  (.A(g17517), .Z(g20386) ) ;
INV     gate10491  (.A(g17520), .Z(g20387) ) ;
INV     gate10492  (.A(g17523), .Z(g20388) ) ;
INV     gate10493  (.A(g17531), .Z(g20389) ) ;
INV     gate10494  (.A(g17534), .Z(g20390) ) ;
INV     gate10495  (.A(g17537), .Z(g20391) ) ;
INV     gate10496  (.A(g17545), .Z(g20392) ) ;
INV     gate10497  (.A(g17548), .Z(g20393) ) ;
INV     gate10498  (.A(g17551), .Z(g20394) ) ;
NOR2    gate10499  (.A(g16008), .B(g16015), .Z(g17225) ) ;
INV     gate10500  (.A(g17225), .Z(II26816) ) ;
INV     gate10501  (.A(II26816), .Z(g20395) ) ;
NOR2    gate10502  (.A(g16010), .B(g16017), .Z(g17226) ) ;
INV     gate10503  (.A(g17226), .Z(II26819) ) ;
INV     gate10504  (.A(II26819), .Z(g20396) ) ;
INV     gate10505  (.A(g17557), .Z(g20397) ) ;
INV     gate10506  (.A(g17560), .Z(g20398) ) ;
INV     gate10507  (.A(g17563), .Z(g20399) ) ;
INV     gate10508  (.A(g17567), .Z(g20400) ) ;
INV     gate10509  (.A(g17570), .Z(g20401) ) ;
INV     gate10510  (.A(g17573), .Z(g20402) ) ;
INV     gate10511  (.A(g17579), .Z(g20403) ) ;
INV     gate10512  (.A(g17582), .Z(g20404) ) ;
INV     gate10513  (.A(g17585), .Z(g20405) ) ;
INV     gate10514  (.A(g17588), .Z(g20406) ) ;
INV     gate10515  (.A(g17591), .Z(g20407) ) ;
INV     gate10516  (.A(g17594), .Z(g20408) ) ;
INV     gate10517  (.A(g17601), .Z(g20409) ) ;
INV     gate10518  (.A(g17604), .Z(g20410) ) ;
INV     gate10519  (.A(g17607), .Z(g20411) ) ;
INV     gate10520  (.A(g17610), .Z(g20412) ) ;
INV     gate10521  (.A(g17613), .Z(g20413) ) ;
INV     gate10522  (.A(g17621), .Z(g20414) ) ;
INV     gate10523  (.A(g17624), .Z(g20415) ) ;
INV     gate10524  (.A(g17627), .Z(g20416) ) ;
NOR2    gate10525  (.A(g16016), .B(g16029), .Z(g17228) ) ;
INV     gate10526  (.A(g17228), .Z(II26843) ) ;
INV     gate10527  (.A(II26843), .Z(g20418) ) ;
NOR2    gate10528  (.A(g16019), .B(g16032), .Z(g17229) ) ;
INV     gate10529  (.A(g17229), .Z(II26846) ) ;
INV     gate10530  (.A(II26846), .Z(g20419) ) ;
INV     gate10531  (.A(g17637), .Z(g20420) ) ;
INV     gate10532  (.A(g17649), .Z(g20421) ) ;
INV     gate10533  (.A(g17655), .Z(g20422) ) ;
INV     gate10534  (.A(g17658), .Z(g20423) ) ;
INV     gate10535  (.A(g17661), .Z(g20424) ) ;
INV     gate10536  (.A(g17664), .Z(g20425) ) ;
INV     gate10537  (.A(g17667), .Z(g20426) ) ;
INV     gate10538  (.A(g17670), .Z(g20427) ) ;
INV     gate10539  (.A(g17676), .Z(g20428) ) ;
INV     gate10540  (.A(g17679), .Z(g20429) ) ;
INV     gate10541  (.A(g17682), .Z(g20430) ) ;
INV     gate10542  (.A(g17685), .Z(g20431) ) ;
INV     gate10543  (.A(g17688), .Z(g20432) ) ;
INV     gate10544  (.A(g17691), .Z(g20433) ) ;
INV     gate10545  (.A(g17698), .Z(g20434) ) ;
INV     gate10546  (.A(g17701), .Z(g20435) ) ;
INV     gate10547  (.A(g17704), .Z(g20436) ) ;
INV     gate10548  (.A(g17707), .Z(g20437) ) ;
INV     gate10549  (.A(g17710), .Z(g20438) ) ;
NOR2    gate10550  (.A(g16028), .B(g16045), .Z(g17234) ) ;
INV     gate10551  (.A(g17234), .Z(II26868) ) ;
INV     gate10552  (.A(II26868), .Z(g20439) ) ;
NOR2    gate10553  (.A(g16030), .B(g16047), .Z(g17235) ) ;
INV     gate10554  (.A(g17235), .Z(II26871) ) ;
INV     gate10555  (.A(II26871), .Z(g20440) ) ;
NOR2    gate10556  (.A(g16033), .B(g16051), .Z(g17236) ) ;
INV     gate10557  (.A(g17236), .Z(II26874) ) ;
INV     gate10558  (.A(II26874), .Z(g20441) ) ;
INV     gate10559  (.A(g17738), .Z(g20442) ) ;
INV     gate10560  (.A(g17749), .Z(g20443) ) ;
INV     gate10561  (.A(g17755), .Z(g20444) ) ;
INV     gate10562  (.A(g17758), .Z(g20445) ) ;
INV     gate10563  (.A(g17761), .Z(g20446) ) ;
INV     gate10564  (.A(g17764), .Z(g20447) ) ;
INV     gate10565  (.A(g17767), .Z(g20448) ) ;
INV     gate10566  (.A(g17770), .Z(g20449) ) ;
INV     gate10567  (.A(g17776), .Z(g20450) ) ;
INV     gate10568  (.A(g17779), .Z(g20451) ) ;
INV     gate10569  (.A(g17782), .Z(g20452) ) ;
INV     gate10570  (.A(g17785), .Z(g20453) ) ;
INV     gate10571  (.A(g17788), .Z(g20454) ) ;
INV     gate10572  (.A(g17791), .Z(g20455) ) ;
INV     gate10573  (.A(g17799), .Z(g20456) ) ;
NOR2    gate10574  (.A(g16046), .B(g16066), .Z(g17246) ) ;
INV     gate10575  (.A(g17246), .Z(II26892) ) ;
INV     gate10576  (.A(II26892), .Z(g20457) ) ;
NOR2    gate10577  (.A(g16050), .B(g16070), .Z(g17247) ) ;
INV     gate10578  (.A(g17247), .Z(II26895) ) ;
INV     gate10579  (.A(II26895), .Z(g20458) ) ;
NOR2    gate10580  (.A(g16052), .B(g16072), .Z(g17248) ) ;
INV     gate10581  (.A(g17248), .Z(II26898) ) ;
INV     gate10582  (.A(II26898), .Z(g20459) ) ;
INV     gate10583  (.A(g17839), .Z(g20461) ) ;
INV     gate10584  (.A(g17850), .Z(g20462) ) ;
INV     gate10585  (.A(g17856), .Z(g20463) ) ;
INV     gate10586  (.A(g17859), .Z(g20464) ) ;
INV     gate10587  (.A(g17862), .Z(g20465) ) ;
INV     gate10588  (.A(g17865), .Z(g20466) ) ;
INV     gate10589  (.A(g17868), .Z(g20467) ) ;
INV     gate10590  (.A(g17871), .Z(g20468) ) ;
NOR2    gate10591  (.A(g16067), .B(g16100), .Z(g17269) ) ;
INV     gate10592  (.A(g17269), .Z(II26910) ) ;
INV     gate10593  (.A(II26910), .Z(g20469) ) ;
NOR2    gate10594  (.A(g16071), .B(g16104), .Z(g17270) ) ;
INV     gate10595  (.A(g17270), .Z(II26913) ) ;
INV     gate10596  (.A(II26913), .Z(g20470) ) ;
NOR2    gate10597  (.A(g16073), .B(g16106), .Z(g17271) ) ;
INV     gate10598  (.A(g17271), .Z(II26916) ) ;
INV     gate10599  (.A(II26916), .Z(g20471) ) ;
INV     gate10600  (.A(g17951), .Z(g20476) ) ;
INV     gate10601  (.A(g17962), .Z(g20477) ) ;
NOR2    gate10602  (.A(g16103), .B(g16135), .Z(g17302) ) ;
INV     gate10603  (.A(g17302), .Z(II26923) ) ;
INV     gate10604  (.A(II26923), .Z(g20478) ) ;
NOR2    gate10605  (.A(g16105), .B(g16137), .Z(g17303) ) ;
INV     gate10606  (.A(g17303), .Z(II26926) ) ;
INV     gate10607  (.A(II26926), .Z(g20479) ) ;
NOR2    gate10608  (.A(g16136), .B(g16183), .Z(g17340) ) ;
INV     gate10609  (.A(g17340), .Z(II26931) ) ;
INV     gate10610  (.A(II26931), .Z(g20484) ) ;
NOR2    gate10611  (.A(g16138), .B(g16185), .Z(g17341) ) ;
INV     gate10612  (.A(g17341), .Z(II26934) ) ;
INV     gate10613  (.A(II26934), .Z(g20485) ) ;
INV     gate10614  (.A(g18166), .Z(g20490) ) ;
NOR2    gate10615  (.A(g16184), .B(g16238), .Z(g17383) ) ;
INV     gate10616  (.A(g17383), .Z(II26940) ) ;
INV     gate10617  (.A(II26940), .Z(g20491) ) ;
INV     gate10618  (.A(g18258), .Z(g20496) ) ;
NOR2    gate10619  (.A(g16239), .B(g16288), .Z(g17429) ) ;
INV     gate10620  (.A(g17429), .Z(II26947) ) ;
INV     gate10621  (.A(II26947), .Z(g20498) ) ;
INV     gate10622  (.A(g18278), .Z(g20500) ) ;
INV     gate10623  (.A(g18334), .Z(g20501) ) ;
INV     gate10624  (.A(g18355), .Z(g20504) ) ;
INV     gate10625  (.A(g18371), .Z(g20505) ) ;
INV     gate10626  (.A(g18351), .Z(g20507) ) ;
INV     gate10627  (.A(g16884), .Z(II26960) ) ;
INV     gate10628  (.A(II26960), .Z(g20513) ) ;
INV     gate10629  (.A(g18432), .Z(g20516) ) ;
INV     gate10630  (.A(g18450), .Z(g20517) ) ;
INV     gate10631  (.A(g18466), .Z(g20518) ) ;
INV     gate10632  (.A(g17051), .Z(II26966) ) ;
INV     gate10633  (.A(II26966), .Z(g20519) ) ;
INV     gate10634  (.A(g18446), .Z(g20526) ) ;
INV     gate10635  (.A(g16913), .Z(II26972) ) ;
INV     gate10636  (.A(II26972), .Z(g20531) ) ;
INV     gate10637  (.A(g18505), .Z(g20534) ) ;
INV     gate10638  (.A(g18523), .Z(g20535) ) ;
INV     gate10639  (.A(g18539), .Z(g20536) ) ;
INV     gate10640  (.A(g17086), .Z(II26980) ) ;
INV     gate10641  (.A(II26980), .Z(g20539) ) ;
INV     gate10642  (.A(g18519), .Z(g20545) ) ;
INV     gate10643  (.A(g16943), .Z(II26985) ) ;
INV     gate10644  (.A(II26985), .Z(g20550) ) ;
INV     gate10645  (.A(g18569), .Z(g20553) ) ;
INV     gate10646  (.A(g18587), .Z(g20554) ) ;
INV     gate10647  (.A(g19145), .Z(II26990) ) ;
INV     gate10648  (.A(g19159), .Z(II26993) ) ;
INV     gate10649  (.A(g19169), .Z(II26996) ) ;
INV     gate10650  (.A(g19543), .Z(II26999) ) ;
INV     gate10651  (.A(g19147), .Z(II27002) ) ;
INV     gate10652  (.A(g19164), .Z(II27005) ) ;
INV     gate10653  (.A(g19175), .Z(II27008) ) ;
INV     gate10654  (.A(g19546), .Z(II27011) ) ;
INV     gate10655  (.A(g19151), .Z(II27014) ) ;
INV     gate10656  (.A(g19170), .Z(II27017) ) ;
INV     gate10657  (.A(g19182), .Z(II27020) ) ;
INV     gate10658  (.A(g19550), .Z(II27023) ) ;
INV     gate10659  (.A(g19156), .Z(II27026) ) ;
INV     gate10660  (.A(g19176), .Z(II27029) ) ;
INV     gate10661  (.A(g19189), .Z(II27032) ) ;
INV     gate10662  (.A(g19556), .Z(II27035) ) ;
INV     gate10663  (.A(g20082), .Z(II27038) ) ;
INV     gate10664  (.A(g19237), .Z(II27041) ) ;
INV     gate10665  (.A(g19247), .Z(II27044) ) ;
INV     gate10666  (.A(g19258), .Z(II27047) ) ;
INV     gate10667  (.A(g19183), .Z(II27050) ) ;
INV     gate10668  (.A(g19190), .Z(II27053) ) ;
INV     gate10669  (.A(g19196), .Z(II27056) ) ;
INV     gate10670  (.A(g19207), .Z(II27059) ) ;
INV     gate10671  (.A(g19217), .Z(II27062) ) ;
INV     gate10672  (.A(g19270), .Z(II27065) ) ;
INV     gate10673  (.A(g19197), .Z(II27068) ) ;
INV     gate10674  (.A(g19218), .Z(II27071) ) ;
INV     gate10675  (.A(g19238), .Z(II27074) ) ;
INV     gate10676  (.A(g19259), .Z(II27077) ) ;
INV     gate10677  (.A(g19198), .Z(II27080) ) ;
INV     gate10678  (.A(g19208), .Z(II27083) ) ;
INV     gate10679  (.A(g19229), .Z(II27086) ) ;
INV     gate10680  (.A(g20105), .Z(II27089) ) ;
INV     gate10681  (.A(g19174), .Z(II27092) ) ;
INV     gate10682  (.A(g19185), .Z(II27095) ) ;
INV     gate10683  (.A(g19199), .Z(II27098) ) ;
INV     gate10684  (.A(g19220), .Z(II27101) ) ;
INV     gate10685  (.A(g19239), .Z(II27104) ) ;
INV     gate10686  (.A(g19249), .Z(II27107) ) ;
INV     gate10687  (.A(g19622), .Z(II27110) ) ;
INV     gate10688  (.A(g19689), .Z(II27113) ) ;
INV     gate10689  (.A(g19762), .Z(II27116) ) ;
INV     gate10690  (.A(g19563), .Z(II27119) ) ;
INV     gate10691  (.A(g19595), .Z(II27122) ) ;
INV     gate10692  (.A(g19652), .Z(II27125) ) ;
INV     gate10693  (.A(g19725), .Z(II27128) ) ;
INV     gate10694  (.A(g19798), .Z(II27131) ) ;
INV     gate10695  (.A(g19573), .Z(II27134) ) ;
INV     gate10696  (.A(g19596), .Z(II27137) ) ;
INV     gate10697  (.A(g19690), .Z(II27140) ) ;
INV     gate10698  (.A(g19763), .Z(II27143) ) ;
INV     gate10699  (.A(g19838), .Z(II27146) ) ;
INV     gate10700  (.A(g19893), .Z(II27149) ) ;
INV     gate10701  (.A(g20360), .Z(II27152) ) ;
INV     gate10702  (.A(g20395), .Z(II27155) ) ;
INV     gate10703  (.A(g20439), .Z(II27158) ) ;
INV     gate10704  (.A(g20377), .Z(II27161) ) ;
INV     gate10705  (.A(g20418), .Z(II27164) ) ;
INV     gate10706  (.A(g20457), .Z(II27167) ) ;
INV     gate10707  (.A(g20396), .Z(II27170) ) ;
INV     gate10708  (.A(g20440), .Z(II27173) ) ;
INV     gate10709  (.A(g20469), .Z(II27176) ) ;
INV     gate10710  (.A(g20419), .Z(II27179) ) ;
INV     gate10711  (.A(g20458), .Z(II27182) ) ;
INV     gate10712  (.A(g20478), .Z(II27185) ) ;
INV     gate10713  (.A(g20441), .Z(II27188) ) ;
INV     gate10714  (.A(g20470), .Z(II27191) ) ;
INV     gate10715  (.A(g20484), .Z(II27194) ) ;
INV     gate10716  (.A(g20459), .Z(II27197) ) ;
INV     gate10717  (.A(g20479), .Z(II27200) ) ;
INV     gate10718  (.A(g20491), .Z(II27203) ) ;
INV     gate10719  (.A(g20471), .Z(II27206) ) ;
INV     gate10720  (.A(g20485), .Z(II27209) ) ;
INV     gate10721  (.A(g20498), .Z(II27212) ) ;
INV     gate10722  (.A(g19158), .Z(II27215) ) ;
INV     gate10723  (.A(g19168), .Z(II27218) ) ;
INV     gate10724  (.A(g19180), .Z(II27221) ) ;
INV     gate10725  (.A(g19358), .Z(II27225) ) ;
INV     gate10726  (.A(II27225), .Z(g20634) ) ;
INV     gate10727  (.A(g19390), .Z(II27228) ) ;
INV     gate10728  (.A(II27228), .Z(g20637) ) ;
INV     gate10729  (.A(g19401), .Z(II27232) ) ;
INV     gate10730  (.A(II27232), .Z(g20641) ) ;
INV     gate10731  (.A(g19420), .Z(II27235) ) ;
INV     gate10732  (.A(II27235), .Z(g20644) ) ;
INV     gate10733  (.A(g19335), .Z(II27240) ) ;
INV     gate10734  (.A(II27240), .Z(g20649) ) ;
INV     gate10735  (.A(g19335), .Z(II27243) ) ;
INV     gate10736  (.A(II27243), .Z(g20652) ) ;
INV     gate10737  (.A(g19335), .Z(II27246) ) ;
INV     gate10738  (.A(II27246), .Z(g20655) ) ;
INV     gate10739  (.A(g19390), .Z(II27250) ) ;
INV     gate10740  (.A(II27250), .Z(g20659) ) ;
INV     gate10741  (.A(g19420), .Z(II27253) ) ;
INV     gate10742  (.A(II27253), .Z(g20662) ) ;
INV     gate10743  (.A(g19431), .Z(II27257) ) ;
INV     gate10744  (.A(II27257), .Z(g20666) ) ;
INV     gate10745  (.A(g19457), .Z(II27260) ) ;
INV     gate10746  (.A(II27260), .Z(g20669) ) ;
INV     gate10747  (.A(g19358), .Z(II27264) ) ;
INV     gate10748  (.A(II27264), .Z(g20673) ) ;
INV     gate10749  (.A(g19358), .Z(II27267) ) ;
INV     gate10750  (.A(II27267), .Z(g20676) ) ;
INV     gate10751  (.A(g19335), .Z(II27270) ) ;
INV     gate10752  (.A(II27270), .Z(g20679) ) ;
INV     gate10753  (.A(g19369), .Z(II27275) ) ;
INV     gate10754  (.A(II27275), .Z(g20684) ) ;
INV     gate10755  (.A(g19369), .Z(II27278) ) ;
INV     gate10756  (.A(II27278), .Z(g20687) ) ;
INV     gate10757  (.A(g19369), .Z(II27281) ) ;
INV     gate10758  (.A(II27281), .Z(g20690) ) ;
INV     gate10759  (.A(g19420), .Z(II27285) ) ;
INV     gate10760  (.A(II27285), .Z(g20694) ) ;
INV     gate10761  (.A(g19457), .Z(II27288) ) ;
INV     gate10762  (.A(II27288), .Z(g20697) ) ;
INV     gate10763  (.A(g19335), .Z(II27293) ) ;
INV     gate10764  (.A(II27293), .Z(g20704) ) ;
INV     gate10765  (.A(g19390), .Z(II27297) ) ;
INV     gate10766  (.A(II27297), .Z(g20708) ) ;
INV     gate10767  (.A(g19390), .Z(II27300) ) ;
INV     gate10768  (.A(II27300), .Z(g20711) ) ;
INV     gate10769  (.A(g19369), .Z(II27303) ) ;
INV     gate10770  (.A(II27303), .Z(g20714) ) ;
INV     gate10771  (.A(g19401), .Z(II27308) ) ;
INV     gate10772  (.A(II27308), .Z(g20719) ) ;
INV     gate10773  (.A(g19401), .Z(II27311) ) ;
INV     gate10774  (.A(II27311), .Z(g20722) ) ;
INV     gate10775  (.A(g19401), .Z(II27314) ) ;
INV     gate10776  (.A(II27314), .Z(g20725) ) ;
INV     gate10777  (.A(g19457), .Z(II27318) ) ;
INV     gate10778  (.A(II27318), .Z(g20729) ) ;
INV     gate10779  (.A(g19335), .Z(II27321) ) ;
INV     gate10780  (.A(II27321), .Z(g20732) ) ;
INV     gate10781  (.A(g19358), .Z(II27324) ) ;
INV     gate10782  (.A(II27324), .Z(g20735) ) ;
INV     gate10783  (.A(g19369), .Z(II27328) ) ;
INV     gate10784  (.A(II27328), .Z(g20739) ) ;
INV     gate10785  (.A(g19420), .Z(II27332) ) ;
INV     gate10786  (.A(II27332), .Z(g20743) ) ;
INV     gate10787  (.A(g19420), .Z(II27335) ) ;
INV     gate10788  (.A(II27335), .Z(g20746) ) ;
INV     gate10789  (.A(g19401), .Z(II27338) ) ;
INV     gate10790  (.A(II27338), .Z(g20749) ) ;
INV     gate10791  (.A(g19431), .Z(II27343) ) ;
INV     gate10792  (.A(II27343), .Z(g20754) ) ;
INV     gate10793  (.A(g19431), .Z(II27346) ) ;
INV     gate10794  (.A(II27346), .Z(g20757) ) ;
INV     gate10795  (.A(g19431), .Z(II27349) ) ;
INV     gate10796  (.A(II27349), .Z(g20760) ) ;
INV     gate10797  (.A(g19358), .Z(II27352) ) ;
INV     gate10798  (.A(II27352), .Z(g20763) ) ;
INV     gate10799  (.A(g19335), .Z(II27355) ) ;
INV     gate10800  (.A(II27355), .Z(g20766) ) ;
INV     gate10801  (.A(g19369), .Z(II27358) ) ;
INV     gate10802  (.A(II27358), .Z(g20769) ) ;
INV     gate10803  (.A(g19390), .Z(II27361) ) ;
INV     gate10804  (.A(II27361), .Z(g20772) ) ;
INV     gate10805  (.A(g19401), .Z(II27365) ) ;
INV     gate10806  (.A(II27365), .Z(g20776) ) ;
INV     gate10807  (.A(g19457), .Z(II27369) ) ;
INV     gate10808  (.A(II27369), .Z(g20780) ) ;
INV     gate10809  (.A(g19457), .Z(II27372) ) ;
INV     gate10810  (.A(II27372), .Z(g20783) ) ;
INV     gate10811  (.A(g19431), .Z(II27375) ) ;
INV     gate10812  (.A(II27375), .Z(g20786) ) ;
INV     gate10813  (.A(g19358), .Z(II27379) ) ;
INV     gate10814  (.A(II27379), .Z(g20790) ) ;
INV     gate10815  (.A(g19390), .Z(II27382) ) ;
INV     gate10816  (.A(II27382), .Z(g20793) ) ;
INV     gate10817  (.A(g19369), .Z(II27385) ) ;
INV     gate10818  (.A(II27385), .Z(g20796) ) ;
INV     gate10819  (.A(g19401), .Z(II27388) ) ;
INV     gate10820  (.A(II27388), .Z(g20799) ) ;
INV     gate10821  (.A(g19420), .Z(II27391) ) ;
INV     gate10822  (.A(II27391), .Z(g20802) ) ;
INV     gate10823  (.A(g19431), .Z(II27395) ) ;
INV     gate10824  (.A(II27395), .Z(g20806) ) ;
INV     gate10825  (.A(g19390), .Z(II27399) ) ;
INV     gate10826  (.A(II27399), .Z(g20810) ) ;
INV     gate10827  (.A(g19420), .Z(II27402) ) ;
INV     gate10828  (.A(II27402), .Z(g20813) ) ;
INV     gate10829  (.A(g19401), .Z(II27405) ) ;
INV     gate10830  (.A(II27405), .Z(g20816) ) ;
INV     gate10831  (.A(g19431), .Z(II27408) ) ;
INV     gate10832  (.A(II27408), .Z(g20819) ) ;
INV     gate10833  (.A(g19457), .Z(II27411) ) ;
INV     gate10834  (.A(II27411), .Z(g20822) ) ;
INV     gate10835  (.A(g19420), .Z(II27416) ) ;
INV     gate10836  (.A(II27416), .Z(g20827) ) ;
INV     gate10837  (.A(g19457), .Z(II27419) ) ;
INV     gate10838  (.A(II27419), .Z(g20830) ) ;
INV     gate10839  (.A(g19431), .Z(II27422) ) ;
INV     gate10840  (.A(II27422), .Z(g20833) ) ;
INV     gate10841  (.A(g19457), .Z(II27426) ) ;
INV     gate10842  (.A(II27426), .Z(g20837) ) ;
INV     gate10843  (.A(g19441), .Z(g20842) ) ;
INV     gate10844  (.A(g19468), .Z(g20850) ) ;
INV     gate10845  (.A(g19491), .Z(g20858) ) ;
INV     gate10846  (.A(g19512), .Z(g20866) ) ;
NAND2   gate10847  (.A(g16607), .B(g9636), .Z(g19865) ) ;
INV     gate10848  (.A(g19865), .Z(g20885) ) ;
NAND2   gate10849  (.A(g16625), .B(g9782), .Z(g19896) ) ;
INV     gate10850  (.A(g19896), .Z(g20904) ) ;
NAND2   gate10851  (.A(g16639), .B(g9928), .Z(g19921) ) ;
INV     gate10852  (.A(g19921), .Z(g20928) ) ;
NOR2    gate10853  (.A(g16850), .B(g13654), .Z(g20310) ) ;
INV     gate10854  (.A(g20310), .Z(II27488) ) ;
INV     gate10855  (.A(II27488), .Z(g20942) ) ;
NOR2    gate10856  (.A(g13646), .B(g16855), .Z(g20314) ) ;
INV     gate10857  (.A(g20314), .Z(II27491) ) ;
INV     gate10858  (.A(II27491), .Z(g20943) ) ;
NAND2   gate10859  (.A(g16650), .B(g10082), .Z(g19936) ) ;
INV     gate10860  (.A(g19936), .Z(g20956) ) ;
NOR2    gate10861  (.A(g13672), .B(g16859), .Z(g20333) ) ;
INV     gate10862  (.A(g20333), .Z(II27516) ) ;
INV     gate10863  (.A(II27516), .Z(g20971) ) ;
NOR2    gate10864  (.A(g16856), .B(g13703), .Z(g20343) ) ;
INV     gate10865  (.A(g20343), .Z(II27531) ) ;
INV     gate10866  (.A(II27531), .Z(g20984) ) ;
INV     gate10867  (.A(g20083), .Z(II27534) ) ;
INV     gate10868  (.A(II27534), .Z(g20985) ) ;
INV     gate10869  (.A(g19957), .Z(II27537) ) ;
INV     gate10870  (.A(II27537), .Z(g20986) ) ;
NOR2    gate10871  (.A(g13702), .B(g16864), .Z(g20353) ) ;
INV     gate10872  (.A(g20353), .Z(II27549) ) ;
INV     gate10873  (.A(II27549), .Z(g20998) ) ;
INV     gate10874  (.A(g19987), .Z(II27565) ) ;
INV     gate10875  (.A(II27565), .Z(g21012) ) ;
NOR2    gate10876  (.A(g13739), .B(g16879), .Z(g20375) ) ;
INV     gate10877  (.A(g20375), .Z(II27577) ) ;
INV     gate10878  (.A(II27577), .Z(g21024) ) ;
NOR2    gate10879  (.A(g16865), .B(g13787), .Z(g20376) ) ;
INV     gate10880  (.A(g20376), .Z(II27585) ) ;
INV     gate10881  (.A(II27585), .Z(g21030) ) ;
INV     gate10882  (.A(g20025), .Z(II27593) ) ;
INV     gate10883  (.A(II27593), .Z(g21036) ) ;
INV     gate10884  (.A(g20513), .Z(g21050) ) ;
INV     gate10885  (.A(g20067), .Z(II27614) ) ;
INV     gate10886  (.A(II27614), .Z(g21057) ) ;
NOR2    gate10887  (.A(g16907), .B(g13833), .Z(g20417) ) ;
INV     gate10888  (.A(g20417), .Z(II27621) ) ;
INV     gate10889  (.A(II27621), .Z(g21064) ) ;
INV     gate10890  (.A(g20519), .Z(g21066) ) ;
INV     gate10891  (.A(g20531), .Z(g21069) ) ;
INV     gate10892  (.A(g20539), .Z(g21076) ) ;
INV     gate10893  (.A(g20550), .Z(g21079) ) ;
INV     gate10894  (.A(g20507), .Z(II27646) ) ;
INV     gate10895  (.A(II27646), .Z(g21087) ) ;
INV     gate10896  (.A(g19064), .Z(g21090) ) ;
INV     gate10897  (.A(g19075), .Z(g21093) ) ;
INV     gate10898  (.A(g20526), .Z(II27658) ) ;
INV     gate10899  (.A(II27658), .Z(g21099) ) ;
INV     gate10900  (.A(g19081), .Z(g21102) ) ;
INV     gate10901  (.A(g20507), .Z(II27667) ) ;
INV     gate10902  (.A(II27667), .Z(g21108) ) ;
INV     gate10903  (.A(g20545), .Z(II27672) ) ;
INV     gate10904  (.A(II27672), .Z(g21113) ) ;
INV     gate10905  (.A(g20526), .Z(II27684) ) ;
INV     gate10906  (.A(II27684), .Z(g21125) ) ;
INV     gate10907  (.A(g19070), .Z(II27689) ) ;
INV     gate10908  (.A(II27689), .Z(g21130) ) ;
INV     gate10909  (.A(g20545), .Z(II27705) ) ;
INV     gate10910  (.A(II27705), .Z(g21144) ) ;
INV     gate10911  (.A(g19070), .Z(II27727) ) ;
INV     gate10912  (.A(II27727), .Z(g21164) ) ;
NAND2   gate10913  (.A(g17186), .B(g92), .Z(g19954) ) ;
INV     gate10914  (.A(g19954), .Z(II27749) ) ;
INV     gate10915  (.A(II27749), .Z(g21184) ) ;
INV     gate10916  (.A(g19113), .Z(g21187) ) ;
NAND2   gate10917  (.A(g17197), .B(g780), .Z(g19984) ) ;
INV     gate10918  (.A(g19984), .Z(II27766) ) ;
INV     gate10919  (.A(II27766), .Z(g21199) ) ;
INV     gate10920  (.A(g19118), .Z(g21202) ) ;
NAND2   gate10921  (.A(g17204), .B(g1466), .Z(g20022) ) ;
INV     gate10922  (.A(g20022), .Z(II27779) ) ;
INV     gate10923  (.A(II27779), .Z(g21214) ) ;
INV     gate10924  (.A(g19125), .Z(g21217) ) ;
NAND2   gate10925  (.A(g17209), .B(g2160), .Z(g20064) ) ;
INV     gate10926  (.A(g20064), .Z(II27785) ) ;
INV     gate10927  (.A(II27785), .Z(g21222) ) ;
INV     gate10928  (.A(g19132), .Z(g21225) ) ;
INV     gate10929  (.A(g19945), .Z(g21241) ) ;
INV     gate10930  (.A(g19972), .Z(g21249) ) ;
INV     gate10931  (.A(g20002), .Z(g21258) ) ;
INV     gate10932  (.A(g20040), .Z(g21266) ) ;
INV     gate10933  (.A(g19865), .Z(II27822) ) ;
INV     gate10934  (.A(II27822), .Z(g21271) ) ;
INV     gate10935  (.A(g19896), .Z(II27827) ) ;
INV     gate10936  (.A(II27827), .Z(g21278) ) ;
INV     gate10937  (.A(g19921), .Z(II27832) ) ;
INV     gate10938  (.A(II27832), .Z(g21285) ) ;
INV     gate10939  (.A(g19936), .Z(II27838) ) ;
INV     gate10940  (.A(II27838), .Z(g21293) ) ;
NOR2    gate10941  (.A(g17268), .B(g14884), .Z(g19144) ) ;
INV     gate10942  (.A(g19144), .Z(II27868) ) ;
INV     gate10943  (.A(II27868), .Z(g21327) ) ;
NOR2    gate10944  (.A(g17339), .B(g15020), .Z(g19149) ) ;
INV     gate10945  (.A(g19149), .Z(II27897) ) ;
INV     gate10946  (.A(II27897), .Z(g21358) ) ;
INV     gate10947  (.A(g19096), .Z(II27900) ) ;
INV     gate10948  (.A(II27900), .Z(g21359) ) ;
NOR2    gate10949  (.A(g17381), .B(g15093), .Z(g19153) ) ;
INV     gate10950  (.A(g19153), .Z(II27917) ) ;
INV     gate10951  (.A(II27917), .Z(g21376) ) ;
NOR2    gate10952  (.A(g17382), .B(g15094), .Z(g19154) ) ;
INV     gate10953  (.A(g19154), .Z(II27920) ) ;
INV     gate10954  (.A(II27920), .Z(g21377) ) ;
INV     gate10955  (.A(g19957), .Z(II27927) ) ;
INV     gate10956  (.A(II27927), .Z(g21382) ) ;
NOR2    gate10957  (.A(g17428), .B(g15171), .Z(g19157) ) ;
INV     gate10958  (.A(g19157), .Z(II27942) ) ;
INV     gate10959  (.A(II27942), .Z(g21399) ) ;
INV     gate10960  (.A(g19918), .Z(g21400) ) ;
INV     gate10961  (.A(g19957), .Z(II27949) ) ;
INV     gate10962  (.A(II27949), .Z(g21404) ) ;
INV     gate10963  (.A(g19987), .Z(II27958) ) ;
INV     gate10964  (.A(II27958), .Z(g21415) ) ;
NOR2    gate10965  (.A(g17485), .B(g15243), .Z(g19162) ) ;
INV     gate10966  (.A(g19162), .Z(II27969) ) ;
INV     gate10967  (.A(II27969), .Z(g21426) ) ;
NOR2    gate10968  (.A(g17486), .B(g15244), .Z(g19163) ) ;
INV     gate10969  (.A(g19163), .Z(II27972) ) ;
INV     gate10970  (.A(II27972), .Z(g21427) ) ;
INV     gate10971  (.A(g19957), .Z(II27976) ) ;
INV     gate10972  (.A(II27976), .Z(g21429) ) ;
INV     gate10973  (.A(g19987), .Z(II27984) ) ;
INV     gate10974  (.A(II27984), .Z(g21441) ) ;
INV     gate10975  (.A(g20025), .Z(II27992) ) ;
INV     gate10976  (.A(II27992), .Z(g21449) ) ;
NOR2    gate10977  (.A(g17556), .B(g15320), .Z(g19167) ) ;
INV     gate10978  (.A(g19167), .Z(II28000) ) ;
INV     gate10979  (.A(II28000), .Z(g21457) ) ;
INV     gate10980  (.A(g19957), .Z(II28003) ) ;
INV     gate10981  (.A(II28003), .Z(g21458) ) ;
INV     gate10982  (.A(g19957), .Z(g21461) ) ;
NAND2   gate10983  (.A(g18085), .B(g646), .Z(g20473) ) ;
INV     gate10984  (.A(g20473), .Z(II28009) ) ;
INV     gate10985  (.A(II28009), .Z(g21473) ) ;
INV     gate10986  (.A(g19987), .Z(II28013) ) ;
INV     gate10987  (.A(II28013), .Z(g21477) ) ;
INV     gate10988  (.A(g20025), .Z(II28019) ) ;
INV     gate10989  (.A(II28019), .Z(g21483) ) ;
INV     gate10990  (.A(g20067), .Z(II28027) ) ;
INV     gate10991  (.A(II28027), .Z(g21491) ) ;
NOR2    gate10992  (.A(g17635), .B(g15388), .Z(g19172) ) ;
INV     gate10993  (.A(g19172), .Z(II28031) ) ;
INV     gate10994  (.A(II28031), .Z(g21495) ) ;
NOR2    gate10995  (.A(g17636), .B(g15389), .Z(g19173) ) ;
INV     gate10996  (.A(g19173), .Z(II28034) ) ;
INV     gate10997  (.A(II28034), .Z(g21496) ) ;
INV     gate10998  (.A(g19957), .Z(II28038) ) ;
INV     gate10999  (.A(II28038), .Z(g21498) ) ;
INV     gate11000  (.A(g19987), .Z(II28043) ) ;
INV     gate11001  (.A(II28043), .Z(g21505) ) ;
INV     gate11002  (.A(g19987), .Z(g21508) ) ;
NAND2   gate11003  (.A(g18201), .B(g1332), .Z(g20481) ) ;
INV     gate11004  (.A(g20481), .Z(II28047) ) ;
INV     gate11005  (.A(II28047), .Z(g21514) ) ;
INV     gate11006  (.A(g20025), .Z(II28051) ) ;
INV     gate11007  (.A(II28051), .Z(g21518) ) ;
INV     gate11008  (.A(g20067), .Z(II28057) ) ;
INV     gate11009  (.A(II28057), .Z(g21524) ) ;
NOR2    gate11010  (.A(g17718), .B(g15452), .Z(g19178) ) ;
INV     gate11011  (.A(g19178), .Z(II28061) ) ;
INV     gate11012  (.A(II28061), .Z(g21528) ) ;
INV     gate11013  (.A(g19272), .Z(g21529) ) ;
INV     gate11014  (.A(g19957), .Z(II28065) ) ;
INV     gate11015  (.A(II28065), .Z(g21530) ) ;
INV     gate11016  (.A(g19987), .Z(II28072) ) ;
INV     gate11017  (.A(II28072), .Z(g21537) ) ;
INV     gate11018  (.A(g20025), .Z(II28076) ) ;
INV     gate11019  (.A(II28076), .Z(g21541) ) ;
INV     gate11020  (.A(g20025), .Z(g21544) ) ;
NAND2   gate11021  (.A(g18308), .B(g2026), .Z(g20487) ) ;
INV     gate11022  (.A(g20487), .Z(II28080) ) ;
INV     gate11023  (.A(II28080), .Z(g21550) ) ;
INV     gate11024  (.A(g20067), .Z(II28084) ) ;
INV     gate11025  (.A(II28084), .Z(g21554) ) ;
NOR2    gate11026  (.A(g17798), .B(g15520), .Z(g19184) ) ;
INV     gate11027  (.A(g19184), .Z(II28087) ) ;
INV     gate11028  (.A(II28087), .Z(g21557) ) ;
NOR2    gate11029  (.A(g18977), .B(g7338), .Z(g20008) ) ;
INV     gate11030  (.A(g20008), .Z(II28090) ) ;
INV     gate11031  (.A(II28090), .Z(g21558) ) ;
INV     gate11032  (.A(g19957), .Z(II28093) ) ;
INV     gate11033  (.A(II28093), .Z(g21561) ) ;
INV     gate11034  (.A(g19291), .Z(g21565) ) ;
INV     gate11035  (.A(g19987), .Z(II28100) ) ;
INV     gate11036  (.A(II28100), .Z(g21566) ) ;
INV     gate11037  (.A(g20025), .Z(II28107) ) ;
INV     gate11038  (.A(II28107), .Z(g21573) ) ;
INV     gate11039  (.A(g20067), .Z(II28111) ) ;
INV     gate11040  (.A(II28111), .Z(g21577) ) ;
INV     gate11041  (.A(g20067), .Z(g21580) ) ;
NAND2   gate11042  (.A(g18401), .B(g2720), .Z(g20493) ) ;
INV     gate11043  (.A(g20493), .Z(II28115) ) ;
INV     gate11044  (.A(II28115), .Z(g21586) ) ;
INV     gate11045  (.A(g19957), .Z(II28119) ) ;
INV     gate11046  (.A(II28119), .Z(g21590) ) ;
INV     gate11047  (.A(g19987), .Z(II28123) ) ;
INV     gate11048  (.A(II28123), .Z(g21594) ) ;
INV     gate11049  (.A(g19309), .Z(g21598) ) ;
INV     gate11050  (.A(g20025), .Z(II28130) ) ;
INV     gate11051  (.A(II28130), .Z(g21599) ) ;
INV     gate11052  (.A(g20067), .Z(II28137) ) ;
INV     gate11053  (.A(II28137), .Z(g21606) ) ;
INV     gate11054  (.A(g19957), .Z(II28143) ) ;
INV     gate11055  (.A(II28143), .Z(g21612) ) ;
INV     gate11056  (.A(g19987), .Z(II28148) ) ;
INV     gate11057  (.A(II28148), .Z(g21619) ) ;
INV     gate11058  (.A(g20025), .Z(II28152) ) ;
INV     gate11059  (.A(II28152), .Z(g21623) ) ;
INV     gate11060  (.A(g19330), .Z(g21627) ) ;
INV     gate11061  (.A(g20067), .Z(II28159) ) ;
INV     gate11062  (.A(II28159), .Z(g21628) ) ;
INV     gate11063  (.A(g19987), .Z(II28169) ) ;
INV     gate11064  (.A(II28169), .Z(g21640) ) ;
INV     gate11065  (.A(g20025), .Z(II28174) ) ;
INV     gate11066  (.A(II28174), .Z(g21647) ) ;
INV     gate11067  (.A(g20067), .Z(II28178) ) ;
INV     gate11068  (.A(II28178), .Z(g21651) ) ;
NAND2   gate11069  (.A(g18590), .B(g2924), .Z(g19103) ) ;
INV     gate11070  (.A(g19103), .Z(II28184) ) ;
INV     gate11071  (.A(II28184), .Z(g21655) ) ;
INV     gate11072  (.A(g19091), .Z(g21661) ) ;
INV     gate11073  (.A(g20025), .Z(II28201) ) ;
INV     gate11074  (.A(II28201), .Z(g21671) ) ;
INV     gate11075  (.A(g20067), .Z(II28206) ) ;
INV     gate11076  (.A(II28206), .Z(g21678) ) ;
NAND2   gate11077  (.A(g18626), .B(g3036), .Z(g20537) ) ;
INV     gate11078  (.A(g20537), .Z(II28210) ) ;
INV     gate11079  (.A(II28210), .Z(g21682) ) ;
INV     gate11080  (.A(g19098), .Z(g21690) ) ;
INV     gate11081  (.A(g20067), .Z(II28229) ) ;
INV     gate11082  (.A(II28229), .Z(g21700) ) ;
NOR2    gate11083  (.A(g16536), .B(g7583), .Z(g20153) ) ;
INV     gate11084  (.A(g20153), .Z(II28235) ) ;
INV     gate11085  (.A(II28235), .Z(g21708) ) ;
INV     gate11086  (.A(g19894), .Z(g21716) ) ;
INV     gate11087  (.A(g19105), .Z(g21726) ) ;
INV     gate11088  (.A(g19919), .Z(g21742) ) ;
INV     gate11089  (.A(g19110), .Z(g21752) ) ;
INV     gate11090  (.A(g19934), .Z(g21766) ) ;
INV     gate11091  (.A(g19951), .Z(g21782) ) ;
NAND2   gate11092  (.A(g5378), .B(g18884), .Z(g19152) ) ;
INV     gate11093  (.A(g19152), .Z(II28314) ) ;
INV     gate11094  (.A(II28314), .Z(g21795) ) ;
NAND2   gate11095  (.A(g5410), .B(g18886), .Z(g20497) ) ;
INV     gate11096  (.A(g20497), .Z(II28357) ) ;
INV     gate11097  (.A(II28357), .Z(g21824) ) ;
INV     gate11098  (.A(g20163), .Z(II28360) ) ;
INV     gate11099  (.A(II28360), .Z(g21825) ) ;
INV     gate11100  (.A(g19657), .Z(g21861) ) ;
INV     gate11101  (.A(g19705), .Z(g21867) ) ;
INV     gate11102  (.A(g19749), .Z(g21872) ) ;
INV     gate11103  (.A(g19792), .Z(g21876) ) ;
INV     gate11104  (.A(g19890), .Z(g21883) ) ;
INV     gate11105  (.A(g19915), .Z(g21886) ) ;
INV     gate11106  (.A(g19945), .Z(g21895) ) ;
INV     gate11107  (.A(g19978), .Z(g21902) ) ;
INV     gate11108  (.A(g19972), .Z(g21907) ) ;
INV     gate11109  (.A(g19335), .Z(II28432) ) ;
INV     gate11110  (.A(II28432), .Z(g21914) ) ;
INV     gate11111  (.A(g19358), .Z(II28435) ) ;
INV     gate11112  (.A(II28435), .Z(g21917) ) ;
INV     gate11113  (.A(g20002), .Z(g21921) ) ;
INV     gate11114  (.A(g20045), .Z(g21927) ) ;
INV     gate11115  (.A(g19358), .Z(II28443) ) ;
INV     gate11116  (.A(II28443), .Z(g21928) ) ;
INV     gate11117  (.A(g19369), .Z(II28447) ) ;
INV     gate11118  (.A(II28447), .Z(g21932) ) ;
INV     gate11119  (.A(g19390), .Z(II28450) ) ;
INV     gate11120  (.A(II28450), .Z(g21935) ) ;
INV     gate11121  (.A(g20040), .Z(g21939) ) ;
INV     gate11122  (.A(g20943), .Z(II28455) ) ;
INV     gate11123  (.A(g20971), .Z(II28458) ) ;
INV     gate11124  (.A(g20998), .Z(II28461) ) ;
INV     gate11125  (.A(g21024), .Z(II28464) ) ;
INV     gate11126  (.A(g20942), .Z(II28467) ) ;
INV     gate11127  (.A(g20984), .Z(II28470) ) ;
INV     gate11128  (.A(g21030), .Z(II28473) ) ;
INV     gate11129  (.A(g21064), .Z(II28476) ) ;
INV     gate11130  (.A(g21795), .Z(II28479) ) ;
INV     gate11131  (.A(g21376), .Z(II28482) ) ;
INV     gate11132  (.A(g21426), .Z(II28485) ) ;
INV     gate11133  (.A(g21495), .Z(II28488) ) ;
INV     gate11134  (.A(g21327), .Z(II28491) ) ;
INV     gate11135  (.A(g21358), .Z(II28494) ) ;
INV     gate11136  (.A(g21399), .Z(II28497) ) ;
INV     gate11137  (.A(g21457), .Z(II28500) ) ;
INV     gate11138  (.A(g21528), .Z(II28503) ) ;
INV     gate11139  (.A(g21377), .Z(II28506) ) ;
INV     gate11140  (.A(g21427), .Z(II28509) ) ;
INV     gate11141  (.A(g21496), .Z(II28512) ) ;
INV     gate11142  (.A(g21557), .Z(II28515) ) ;
INV     gate11143  (.A(g20985), .Z(II28518) ) ;
INV     gate11144  (.A(g21824), .Z(II28521) ) ;
INV     gate11145  (.A(g21359), .Z(II28524) ) ;
NOR2    gate11146  (.A(g20499), .B(g13316), .Z(g21407) ) ;
INV     gate11147  (.A(g21407), .Z(II28527) ) ;
INV     gate11148  (.A(II28527), .Z(g21967) ) ;
NOR2    gate11149  (.A(g20506), .B(g13355), .Z(g21467) ) ;
INV     gate11150  (.A(g21467), .Z(II28541) ) ;
INV     gate11151  (.A(II28541), .Z(g21982) ) ;
NOR2    gate11152  (.A(g20502), .B(g13335), .Z(g21432) ) ;
INV     gate11153  (.A(g21432), .Z(II28550) ) ;
INV     gate11154  (.A(II28550), .Z(g21995) ) ;
INV     gate11155  (.A(g21407), .Z(II28557) ) ;
INV     gate11156  (.A(II28557), .Z(g22003) ) ;
NOR2    gate11157  (.A(g20492), .B(g13289), .Z(g21385) ) ;
INV     gate11158  (.A(g21385), .Z(II28564) ) ;
INV     gate11159  (.A(II28564), .Z(g22014) ) ;
NOR2    gate11160  (.A(g13609), .B(g19150), .Z(g21842) ) ;
INV     gate11161  (.A(g21842), .Z(II28628) ) ;
INV     gate11162  (.A(II28628), .Z(g22082) ) ;
NOR2    gate11163  (.A(g13619), .B(g19155), .Z(g21843) ) ;
INV     gate11164  (.A(g21843), .Z(II28649) ) ;
INV     gate11165  (.A(II28649), .Z(g22107) ) ;
NOR2    gate11166  (.A(g13631), .B(g19161), .Z(g21845) ) ;
INV     gate11167  (.A(g21845), .Z(II28671) ) ;
INV     gate11168  (.A(II28671), .Z(g22133) ) ;
NOR2    gate11169  (.A(g13642), .B(g19166), .Z(g21847) ) ;
INV     gate11170  (.A(g21847), .Z(II28693) ) ;
INV     gate11171  (.A(II28693), .Z(g22156) ) ;
NOR2    gate11172  (.A(g19252), .B(g8842), .Z(g21851) ) ;
INV     gate11173  (.A(g21851), .Z(II28712) ) ;
INV     gate11174  (.A(II28712), .Z(g22176) ) ;
INV     gate11175  (.A(g21914), .Z(g22212) ) ;
INV     gate11176  (.A(g21917), .Z(g22213) ) ;
INV     gate11177  (.A(g21928), .Z(g22217) ) ;
NOR2    gate11178  (.A(g20472), .B(g16153), .Z(g21331) ) ;
INV     gate11179  (.A(g21331), .Z(II28781) ) ;
INV     gate11180  (.A(II28781), .Z(g22219) ) ;
INV     gate11181  (.A(g21932), .Z(g22221) ) ;
INV     gate11182  (.A(g21935), .Z(g22222) ) ;
NOR2    gate11183  (.A(g16964), .B(g19228), .Z(g21878) ) ;
INV     gate11184  (.A(g21878), .Z(II28789) ) ;
INV     gate11185  (.A(II28789), .Z(g22225) ) ;
NOR2    gate11186  (.A(g13854), .B(g19236), .Z(g21880) ) ;
INV     gate11187  (.A(g21880), .Z(II28792) ) ;
INV     gate11188  (.A(II28792), .Z(g22226) ) ;
INV     gate11189  (.A(g20634), .Z(g22230) ) ;
NOR2    gate11190  (.A(g20460), .B(g16111), .Z(g21316) ) ;
INV     gate11191  (.A(g21316), .Z(II28800) ) ;
INV     gate11192  (.A(II28800), .Z(g22232) ) ;
INV     gate11193  (.A(g20637), .Z(g22233) ) ;
INV     gate11194  (.A(g20641), .Z(g22236) ) ;
INV     gate11195  (.A(g20644), .Z(g22237) ) ;
INV     gate11196  (.A(g20649), .Z(g22239) ) ;
INV     gate11197  (.A(g20652), .Z(g22240) ) ;
INV     gate11198  (.A(g20655), .Z(g22241) ) ;
NOR2    gate11199  (.A(g20525), .B(g16445), .Z(g21502) ) ;
INV     gate11200  (.A(g21502), .Z(II28813) ) ;
INV     gate11201  (.A(II28813), .Z(g22243) ) ;
INV     gate11202  (.A(g20659), .Z(g22246) ) ;
INV     gate11203  (.A(g20662), .Z(g22248) ) ;
INV     gate11204  (.A(g20666), .Z(g22251) ) ;
INV     gate11205  (.A(g20669), .Z(g22252) ) ;
NOR2    gate11206  (.A(g13862), .B(g19248), .Z(g21882) ) ;
INV     gate11207  (.A(g21882), .Z(II28825) ) ;
INV     gate11208  (.A(II28825), .Z(g22253) ) ;
INV     gate11209  (.A(g20673), .Z(g22256) ) ;
INV     gate11210  (.A(g20676), .Z(g22257) ) ;
INV     gate11211  (.A(g20679), .Z(g22258) ) ;
NOR2    gate11212  (.A(g20512), .B(g16417), .Z(g21470) ) ;
INV     gate11213  (.A(g21470), .Z(II28833) ) ;
INV     gate11214  (.A(II28833), .Z(g22259) ) ;
INV     gate11215  (.A(g20684), .Z(g22260) ) ;
INV     gate11216  (.A(g20687), .Z(g22261) ) ;
INV     gate11217  (.A(g20690), .Z(g22262) ) ;
INV     gate11218  (.A(g20694), .Z(g22266) ) ;
INV     gate11219  (.A(g20697), .Z(g22268) ) ;
INV     gate11220  (.A(g20704), .Z(g22271) ) ;
INV     gate11221  (.A(g20708), .Z(g22274) ) ;
INV     gate11222  (.A(g20711), .Z(g22275) ) ;
INV     gate11223  (.A(g20714), .Z(g22276) ) ;
INV     gate11224  (.A(g20719), .Z(g22277) ) ;
INV     gate11225  (.A(g20722), .Z(g22278) ) ;
INV     gate11226  (.A(g20725), .Z(g22279) ) ;
INV     gate11227  (.A(g20729), .Z(g22283) ) ;
INV     gate11228  (.A(g20732), .Z(g22286) ) ;
INV     gate11229  (.A(g20735), .Z(g22287) ) ;
INV     gate11230  (.A(g20739), .Z(g22290) ) ;
INV     gate11231  (.A(g20743), .Z(g22293) ) ;
INV     gate11232  (.A(g20746), .Z(g22294) ) ;
INV     gate11233  (.A(g20749), .Z(g22295) ) ;
INV     gate11234  (.A(g20754), .Z(g22296) ) ;
INV     gate11235  (.A(g20757), .Z(g22297) ) ;
INV     gate11236  (.A(g20760), .Z(g22298) ) ;
NOR2    gate11237  (.A(g19954), .B(g5890), .Z(g21238) ) ;
INV     gate11238  (.A(g21238), .Z(II28876) ) ;
INV     gate11239  (.A(II28876), .Z(g22300) ) ;
INV     gate11240  (.A(g20763), .Z(g22303) ) ;
INV     gate11241  (.A(g20766), .Z(g22304) ) ;
INV     gate11242  (.A(g20769), .Z(g22306) ) ;
INV     gate11243  (.A(g20772), .Z(g22307) ) ;
INV     gate11244  (.A(g20776), .Z(g22310) ) ;
INV     gate11245  (.A(g20780), .Z(g22313) ) ;
INV     gate11246  (.A(g20783), .Z(g22314) ) ;
INV     gate11247  (.A(g20786), .Z(g22315) ) ;
NOR2    gate11248  (.A(g20015), .B(g19981), .Z(g21149) ) ;
INV     gate11249  (.A(g21149), .Z(g22316) ) ;
INV     gate11250  (.A(g20790), .Z(g22318) ) ;
NOR2    gate11251  (.A(g19388), .B(g17118), .Z(g21228) ) ;
INV     gate11252  (.A(g21228), .Z(g22319) ) ;
NOR2    gate11253  (.A(g19984), .B(g5929), .Z(g21246) ) ;
INV     gate11254  (.A(g21246), .Z(II28896) ) ;
INV     gate11255  (.A(II28896), .Z(g22328) ) ;
INV     gate11256  (.A(g20793), .Z(g22331) ) ;
INV     gate11257  (.A(g20796), .Z(g22332) ) ;
INV     gate11258  (.A(g20799), .Z(g22334) ) ;
INV     gate11259  (.A(g20802), .Z(g22335) ) ;
INV     gate11260  (.A(g20806), .Z(g22338) ) ;
NOR2    gate11261  (.A(g20057), .B(g20019), .Z(g21169) ) ;
INV     gate11262  (.A(g21169), .Z(g22341) ) ;
INV     gate11263  (.A(g20810), .Z(g22343) ) ;
NOR2    gate11264  (.A(g19418), .B(g17145), .Z(g21233) ) ;
INV     gate11265  (.A(g21233), .Z(g22344) ) ;
NOR2    gate11266  (.A(g20022), .B(g5963), .Z(g21255) ) ;
INV     gate11267  (.A(g21255), .Z(II28913) ) ;
INV     gate11268  (.A(II28913), .Z(g22353) ) ;
INV     gate11269  (.A(g20813), .Z(g22356) ) ;
INV     gate11270  (.A(g20816), .Z(g22357) ) ;
INV     gate11271  (.A(g20819), .Z(g22359) ) ;
INV     gate11272  (.A(g20822), .Z(g22360) ) ;
NOR2    gate11273  (.A(g20098), .B(g20061), .Z(g21189) ) ;
INV     gate11274  (.A(g21189), .Z(g22364) ) ;
INV     gate11275  (.A(g20827), .Z(g22366) ) ;
NOR2    gate11276  (.A(g19455), .B(g17168), .Z(g21242) ) ;
INV     gate11277  (.A(g21242), .Z(g22367) ) ;
NOR2    gate11278  (.A(g20064), .B(g5992), .Z(g21263) ) ;
INV     gate11279  (.A(g21263), .Z(II28928) ) ;
INV     gate11280  (.A(II28928), .Z(g22376) ) ;
INV     gate11281  (.A(g20830), .Z(g22379) ) ;
INV     gate11282  (.A(g20833), .Z(g22380) ) ;
NOR2    gate11283  (.A(g20123), .B(g20102), .Z(g21204) ) ;
INV     gate11284  (.A(g21204), .Z(g22384) ) ;
INV     gate11285  (.A(g20837), .Z(g22386) ) ;
NOR2    gate11286  (.A(g19482), .B(g17183), .Z(g21250) ) ;
INV     gate11287  (.A(g21250), .Z(g22387) ) ;
AND4    gate11288  (.A(g17724), .B(g18179), .C(g19799), .D(II28068), .Z(g21533) ) ;
INV     gate11289  (.A(g21533), .Z(g22401) ) ;
AND4    gate11290  (.A(g17825), .B(g18286), .C(g19843), .D(II28103), .Z(g21569) ) ;
INV     gate11291  (.A(g21569), .Z(g22402) ) ;
AND4    gate11292  (.A(g17937), .B(g18379), .C(g19876), .D(II28133), .Z(g21602) ) ;
INV     gate11293  (.A(g21602), .Z(g22403) ) ;
AND4    gate11294  (.A(g18048), .B(g18474), .C(g19907), .D(II28162), .Z(g21631) ) ;
INV     gate11295  (.A(g21631), .Z(g22404) ) ;
NAND2   gate11296  (.A(g20164), .B(g6232), .Z(g21685) ) ;
INV     gate11297  (.A(g21685), .Z(II28949) ) ;
INV     gate11298  (.A(II28949), .Z(g22405) ) ;
INV     gate11299  (.A(g20986), .Z(g22408) ) ;
NAND2   gate11300  (.A(g20164), .B(g6314), .Z(g21659) ) ;
INV     gate11301  (.A(g21659), .Z(II28953) ) ;
INV     gate11302  (.A(II28953), .Z(g22409) ) ;
NAND2   gate11303  (.A(g20164), .B(g6232), .Z(g21714) ) ;
INV     gate11304  (.A(g21714), .Z(II28956) ) ;
INV     gate11305  (.A(II28956), .Z(g22412) ) ;
NOR2    gate11306  (.A(g20473), .B(g6513), .Z(g21636) ) ;
INV     gate11307  (.A(g21636), .Z(II28959) ) ;
INV     gate11308  (.A(II28959), .Z(g22415) ) ;
NAND2   gate11309  (.A(g20198), .B(g6369), .Z(g21721) ) ;
INV     gate11310  (.A(g21721), .Z(II28962) ) ;
INV     gate11311  (.A(II28962), .Z(g22418) ) ;
INV     gate11312  (.A(g21012), .Z(g22421) ) ;
NAND2   gate11313  (.A(g20164), .B(g3254), .Z(g20633) ) ;
INV     gate11314  (.A(g20633), .Z(II28966) ) ;
INV     gate11315  (.A(II28966), .Z(g22422) ) ;
NAND2   gate11316  (.A(g20164), .B(g6314), .Z(g21686) ) ;
INV     gate11317  (.A(g21686), .Z(II28969) ) ;
INV     gate11318  (.A(II28969), .Z(g22425) ) ;
NAND2   gate11319  (.A(g20164), .B(g6232), .Z(g21736) ) ;
INV     gate11320  (.A(g21736), .Z(II28972) ) ;
INV     gate11321  (.A(II28972), .Z(g22428) ) ;
NAND2   gate11322  (.A(g20198), .B(g6519), .Z(g21688) ) ;
INV     gate11323  (.A(g21688), .Z(II28975) ) ;
INV     gate11324  (.A(II28975), .Z(g22431) ) ;
NAND2   gate11325  (.A(g20198), .B(g6369), .Z(g21740) ) ;
INV     gate11326  (.A(g21740), .Z(II28978) ) ;
INV     gate11327  (.A(II28978), .Z(g22434) ) ;
NOR2    gate11328  (.A(g20481), .B(g6777), .Z(g21667) ) ;
INV     gate11329  (.A(g21667), .Z(II28981) ) ;
INV     gate11330  (.A(II28981), .Z(g22437) ) ;
NAND2   gate11331  (.A(g20228), .B(g6574), .Z(g21747) ) ;
INV     gate11332  (.A(g21747), .Z(II28984) ) ;
INV     gate11333  (.A(II28984), .Z(g22440) ) ;
INV     gate11334  (.A(g21036), .Z(g22443) ) ;
NOR2    gate11335  (.A(g17301), .B(g19594), .Z(g20874) ) ;
INV     gate11336  (.A(g20874), .Z(II28988) ) ;
INV     gate11337  (.A(II28988), .Z(g22444) ) ;
NAND2   gate11338  (.A(g20164), .B(g3254), .Z(g20648) ) ;
INV     gate11339  (.A(g20648), .Z(II28991) ) ;
INV     gate11340  (.A(II28991), .Z(g22445) ) ;
NAND2   gate11341  (.A(g20164), .B(g6314), .Z(g21715) ) ;
INV     gate11342  (.A(g21715), .Z(II28994) ) ;
INV     gate11343  (.A(II28994), .Z(g22448) ) ;
NAND2   gate11344  (.A(g20164), .B(g6232), .Z(g21759) ) ;
INV     gate11345  (.A(g21759), .Z(II28997) ) ;
INV     gate11346  (.A(II28997), .Z(g22451) ) ;
NAND2   gate11347  (.A(g20198), .B(g3410), .Z(g20658) ) ;
INV     gate11348  (.A(g20658), .Z(II29001) ) ;
INV     gate11349  (.A(II29001), .Z(g22455) ) ;
NAND2   gate11350  (.A(g20198), .B(g6519), .Z(g21722) ) ;
INV     gate11351  (.A(g21722), .Z(II29004) ) ;
INV     gate11352  (.A(II29004), .Z(g22458) ) ;
NAND2   gate11353  (.A(g20198), .B(g6369), .Z(g21760) ) ;
INV     gate11354  (.A(g21760), .Z(II29007) ) ;
INV     gate11355  (.A(II29007), .Z(g22461) ) ;
NAND2   gate11356  (.A(g20228), .B(g6783), .Z(g21724) ) ;
INV     gate11357  (.A(g21724), .Z(II29010) ) ;
INV     gate11358  (.A(II29010), .Z(g22464) ) ;
NAND2   gate11359  (.A(g20228), .B(g6574), .Z(g21764) ) ;
INV     gate11360  (.A(g21764), .Z(II29013) ) ;
INV     gate11361  (.A(II29013), .Z(g22467) ) ;
NOR2    gate11362  (.A(g20487), .B(g7079), .Z(g21696) ) ;
INV     gate11363  (.A(g21696), .Z(II29016) ) ;
INV     gate11364  (.A(II29016), .Z(g22470) ) ;
NAND2   gate11365  (.A(g20255), .B(g6838), .Z(g21771) ) ;
INV     gate11366  (.A(g21771), .Z(II29019) ) ;
INV     gate11367  (.A(II29019), .Z(g22473) ) ;
INV     gate11368  (.A(g21057), .Z(g22476) ) ;
NAND2   gate11369  (.A(g20164), .B(g3254), .Z(g20672) ) ;
INV     gate11370  (.A(g20672), .Z(II29023) ) ;
INV     gate11371  (.A(II29023), .Z(g22477) ) ;
NAND2   gate11372  (.A(g20164), .B(g6314), .Z(g21737) ) ;
INV     gate11373  (.A(g21737), .Z(II29026) ) ;
INV     gate11374  (.A(II29026), .Z(g22480) ) ;
NAND2   gate11375  (.A(g20198), .B(g3410), .Z(g20683) ) ;
INV     gate11376  (.A(g20683), .Z(II29030) ) ;
INV     gate11377  (.A(II29030), .Z(g22484) ) ;
NAND2   gate11378  (.A(g20198), .B(g6519), .Z(g21741) ) ;
INV     gate11379  (.A(g21741), .Z(II29033) ) ;
INV     gate11380  (.A(II29033), .Z(g22487) ) ;
NAND2   gate11381  (.A(g20198), .B(g6369), .Z(g21775) ) ;
INV     gate11382  (.A(g21775), .Z(II29036) ) ;
INV     gate11383  (.A(II29036), .Z(g22490) ) ;
NAND2   gate11384  (.A(g20228), .B(g3566), .Z(g20693) ) ;
INV     gate11385  (.A(g20693), .Z(II29040) ) ;
INV     gate11386  (.A(II29040), .Z(g22494) ) ;
NAND2   gate11387  (.A(g20228), .B(g6783), .Z(g21748) ) ;
INV     gate11388  (.A(g21748), .Z(II29043) ) ;
INV     gate11389  (.A(II29043), .Z(g22497) ) ;
NAND2   gate11390  (.A(g20228), .B(g6574), .Z(g21776) ) ;
INV     gate11391  (.A(g21776), .Z(II29046) ) ;
INV     gate11392  (.A(II29046), .Z(g22500) ) ;
NAND2   gate11393  (.A(g20255), .B(g7085), .Z(g21750) ) ;
INV     gate11394  (.A(g21750), .Z(II29049) ) ;
INV     gate11395  (.A(II29049), .Z(g22503) ) ;
NAND2   gate11396  (.A(g20255), .B(g6838), .Z(g21780) ) ;
INV     gate11397  (.A(g21780), .Z(II29052) ) ;
INV     gate11398  (.A(II29052), .Z(g22506) ) ;
NOR2    gate11399  (.A(g20493), .B(g7329), .Z(g21732) ) ;
INV     gate11400  (.A(g21732), .Z(II29055) ) ;
INV     gate11401  (.A(II29055), .Z(g22509) ) ;
NAND2   gate11402  (.A(g20164), .B(g3254), .Z(g20703) ) ;
INV     gate11403  (.A(g20703), .Z(II29058) ) ;
INV     gate11404  (.A(II29058), .Z(g22512) ) ;
NOR2    gate11405  (.A(g19584), .B(g17352), .Z(g20875) ) ;
INV     gate11406  (.A(g20875), .Z(II29064) ) ;
INV     gate11407  (.A(II29064), .Z(g22518) ) ;
NOR2    gate11408  (.A(g19585), .B(g17353), .Z(g20876) ) ;
INV     gate11409  (.A(g20876), .Z(II29067) ) ;
INV     gate11410  (.A(II29067), .Z(g22519) ) ;
NAND2   gate11411  (.A(g20198), .B(g3410), .Z(g20707) ) ;
INV     gate11412  (.A(g20707), .Z(II29070) ) ;
INV     gate11413  (.A(II29070), .Z(g22520) ) ;
NAND2   gate11414  (.A(g20198), .B(g6519), .Z(g21761) ) ;
INV     gate11415  (.A(g21761), .Z(II29073) ) ;
INV     gate11416  (.A(II29073), .Z(g22523) ) ;
NAND2   gate11417  (.A(g20228), .B(g3566), .Z(g20718) ) ;
INV     gate11418  (.A(g20718), .Z(II29077) ) ;
INV     gate11419  (.A(II29077), .Z(g22527) ) ;
NAND2   gate11420  (.A(g20228), .B(g6783), .Z(g21765) ) ;
INV     gate11421  (.A(g21765), .Z(II29080) ) ;
INV     gate11422  (.A(II29080), .Z(g22530) ) ;
NAND2   gate11423  (.A(g20228), .B(g6574), .Z(g21790) ) ;
INV     gate11424  (.A(g21790), .Z(II29083) ) ;
INV     gate11425  (.A(II29083), .Z(g22533) ) ;
NAND2   gate11426  (.A(g20255), .B(g3722), .Z(g20728) ) ;
INV     gate11427  (.A(g20728), .Z(II29087) ) ;
INV     gate11428  (.A(II29087), .Z(g22537) ) ;
NAND2   gate11429  (.A(g20255), .B(g7085), .Z(g21772) ) ;
INV     gate11430  (.A(g21772), .Z(II29090) ) ;
INV     gate11431  (.A(II29090), .Z(g22540) ) ;
NAND2   gate11432  (.A(g20255), .B(g6838), .Z(g21791) ) ;
INV     gate11433  (.A(g21791), .Z(II29093) ) ;
INV     gate11434  (.A(II29093), .Z(g22543) ) ;
INV     gate11435  (.A(g21087), .Z(g22547) ) ;
NOR2    gate11436  (.A(g19601), .B(g17396), .Z(g20879) ) ;
INV     gate11437  (.A(g20879), .Z(II29098) ) ;
INV     gate11438  (.A(II29098), .Z(g22548) ) ;
NOR2    gate11439  (.A(g19602), .B(g17397), .Z(g20880) ) ;
INV     gate11440  (.A(g20880), .Z(II29101) ) ;
INV     gate11441  (.A(II29101), .Z(g22549) ) ;
NOR2    gate11442  (.A(g19603), .B(g17398), .Z(g20881) ) ;
INV     gate11443  (.A(g20881), .Z(II29104) ) ;
INV     gate11444  (.A(II29104), .Z(g22550) ) ;
NOR2    gate11445  (.A(g20503), .B(g16385), .Z(g21435) ) ;
INV     gate11446  (.A(g21435), .Z(II29107) ) ;
INV     gate11447  (.A(II29107), .Z(g22551) ) ;
NAND2   gate11448  (.A(g20198), .B(g3410), .Z(g20738) ) ;
INV     gate11449  (.A(g20738), .Z(II29110) ) ;
INV     gate11450  (.A(II29110), .Z(g22552) ) ;
NOR2    gate11451  (.A(g19614), .B(g17408), .Z(g20882) ) ;
INV     gate11452  (.A(g20882), .Z(II29116) ) ;
INV     gate11453  (.A(II29116), .Z(g22558) ) ;
NOR2    gate11454  (.A(g19615), .B(g17409), .Z(g20883) ) ;
INV     gate11455  (.A(g20883), .Z(II29119) ) ;
INV     gate11456  (.A(II29119), .Z(g22559) ) ;
NAND2   gate11457  (.A(g20228), .B(g3566), .Z(g20742) ) ;
INV     gate11458  (.A(g20742), .Z(II29122) ) ;
INV     gate11459  (.A(II29122), .Z(g22560) ) ;
NAND2   gate11460  (.A(g20228), .B(g6783), .Z(g21777) ) ;
INV     gate11461  (.A(g21777), .Z(II29125) ) ;
INV     gate11462  (.A(II29125), .Z(g22563) ) ;
NAND2   gate11463  (.A(g20255), .B(g3722), .Z(g20753) ) ;
INV     gate11464  (.A(g20753), .Z(II29129) ) ;
INV     gate11465  (.A(II29129), .Z(g22567) ) ;
NAND2   gate11466  (.A(g20255), .B(g7085), .Z(g21781) ) ;
INV     gate11467  (.A(g21781), .Z(II29132) ) ;
INV     gate11468  (.A(II29132), .Z(g22570) ) ;
NAND2   gate11469  (.A(g20255), .B(g6838), .Z(g21804) ) ;
INV     gate11470  (.A(g21804), .Z(II29135) ) ;
INV     gate11471  (.A(II29135), .Z(g22573) ) ;
NOR2    gate11472  (.A(g19160), .B(g10024), .Z(g20682) ) ;
INV     gate11473  (.A(g20682), .Z(II29142) ) ;
INV     gate11474  (.A(II29142), .Z(g22582) ) ;
NOR2    gate11475  (.A(g19626), .B(g17447), .Z(g20891) ) ;
INV     gate11476  (.A(g20891), .Z(II29145) ) ;
INV     gate11477  (.A(II29145), .Z(g22583) ) ;
NOR2    gate11478  (.A(g19627), .B(g17448), .Z(g20892) ) ;
INV     gate11479  (.A(g20892), .Z(II29148) ) ;
INV     gate11480  (.A(II29148), .Z(g22584) ) ;
NOR2    gate11481  (.A(g19628), .B(g17449), .Z(g20893) ) ;
INV     gate11482  (.A(g20893), .Z(II29151) ) ;
INV     gate11483  (.A(II29151), .Z(g22585) ) ;
NOR2    gate11484  (.A(g19629), .B(g17450), .Z(g20894) ) ;
INV     gate11485  (.A(g20894), .Z(II29154) ) ;
INV     gate11486  (.A(II29154), .Z(g22586) ) ;
INV     gate11487  (.A(g21099), .Z(g22588) ) ;
NOR2    gate11488  (.A(g19634), .B(g17462), .Z(g20896) ) ;
INV     gate11489  (.A(g20896), .Z(II29159) ) ;
INV     gate11490  (.A(II29159), .Z(g22589) ) ;
NOR2    gate11491  (.A(g19635), .B(g17463), .Z(g20897) ) ;
INV     gate11492  (.A(g20897), .Z(II29162) ) ;
INV     gate11493  (.A(II29162), .Z(g22590) ) ;
NOR2    gate11494  (.A(g19636), .B(g17464), .Z(g20898) ) ;
INV     gate11495  (.A(g20898), .Z(II29165) ) ;
INV     gate11496  (.A(II29165), .Z(g22591) ) ;
NAND2   gate11497  (.A(g20228), .B(g3566), .Z(g20775) ) ;
INV     gate11498  (.A(g20775), .Z(II29168) ) ;
INV     gate11499  (.A(II29168), .Z(g22592) ) ;
NOR2    gate11500  (.A(g19647), .B(g17474), .Z(g20899) ) ;
INV     gate11501  (.A(g20899), .Z(II29174) ) ;
INV     gate11502  (.A(II29174), .Z(g22598) ) ;
NOR2    gate11503  (.A(g19648), .B(g17475), .Z(g20900) ) ;
INV     gate11504  (.A(g20900), .Z(II29177) ) ;
INV     gate11505  (.A(II29177), .Z(g22599) ) ;
NAND2   gate11506  (.A(g20255), .B(g3722), .Z(g20779) ) ;
INV     gate11507  (.A(g20779), .Z(II29180) ) ;
INV     gate11508  (.A(II29180), .Z(g22600) ) ;
NAND2   gate11509  (.A(g20255), .B(g7085), .Z(g21792) ) ;
INV     gate11510  (.A(g21792), .Z(II29183) ) ;
INV     gate11511  (.A(II29183), .Z(g22603) ) ;
INV     gate11512  (.A(g21108), .Z(g22609) ) ;
NOR2    gate11513  (.A(g19660), .B(g17508), .Z(g20901) ) ;
INV     gate11514  (.A(g20901), .Z(II29191) ) ;
INV     gate11515  (.A(II29191), .Z(g22611) ) ;
NOR2    gate11516  (.A(g19661), .B(g17509), .Z(g20902) ) ;
INV     gate11517  (.A(g20902), .Z(II29194) ) ;
INV     gate11518  (.A(II29194), .Z(g22612) ) ;
NOR2    gate11519  (.A(g19662), .B(g17510), .Z(g20903) ) ;
INV     gate11520  (.A(g20903), .Z(II29197) ) ;
INV     gate11521  (.A(II29197), .Z(g22613) ) ;
NOR2    gate11522  (.A(g19165), .B(g10133), .Z(g20717) ) ;
INV     gate11523  (.A(g20717), .Z(II29203) ) ;
INV     gate11524  (.A(II29203), .Z(g22619) ) ;
NOR2    gate11525  (.A(g19666), .B(g17527), .Z(g20910) ) ;
INV     gate11526  (.A(g20910), .Z(II29206) ) ;
INV     gate11527  (.A(II29206), .Z(g22620) ) ;
NOR2    gate11528  (.A(g19667), .B(g17528), .Z(g20911) ) ;
INV     gate11529  (.A(g20911), .Z(II29209) ) ;
INV     gate11530  (.A(II29209), .Z(g22621) ) ;
NOR2    gate11531  (.A(g19668), .B(g17529), .Z(g20912) ) ;
INV     gate11532  (.A(g20912), .Z(II29212) ) ;
INV     gate11533  (.A(II29212), .Z(g22622) ) ;
NOR2    gate11534  (.A(g19669), .B(g17530), .Z(g20913) ) ;
INV     gate11535  (.A(g20913), .Z(II29215) ) ;
INV     gate11536  (.A(II29215), .Z(g22623) ) ;
INV     gate11537  (.A(g21113), .Z(g22625) ) ;
NOR2    gate11538  (.A(g19674), .B(g17542), .Z(g20915) ) ;
INV     gate11539  (.A(g20915), .Z(II29220) ) ;
INV     gate11540  (.A(II29220), .Z(g22626) ) ;
NOR2    gate11541  (.A(g19675), .B(g17543), .Z(g20916) ) ;
INV     gate11542  (.A(g20916), .Z(II29223) ) ;
INV     gate11543  (.A(II29223), .Z(g22627) ) ;
NOR2    gate11544  (.A(g19676), .B(g17544), .Z(g20917) ) ;
INV     gate11545  (.A(g20917), .Z(II29226) ) ;
INV     gate11546  (.A(II29226), .Z(g22628) ) ;
NAND2   gate11547  (.A(g20255), .B(g3722), .Z(g20805) ) ;
INV     gate11548  (.A(g20805), .Z(II29229) ) ;
INV     gate11549  (.A(II29229), .Z(g22629) ) ;
NOR2    gate11550  (.A(g19687), .B(g17554), .Z(g20918) ) ;
INV     gate11551  (.A(g20918), .Z(II29235) ) ;
INV     gate11552  (.A(II29235), .Z(g22635) ) ;
NOR2    gate11553  (.A(g19688), .B(g17555), .Z(g20919) ) ;
INV     gate11554  (.A(g20919), .Z(II29238) ) ;
INV     gate11555  (.A(II29238), .Z(g22636) ) ;
NOR2    gate11556  (.A(g19697), .B(g17576), .Z(g20921) ) ;
INV     gate11557  (.A(g20921), .Z(II29243) ) ;
INV     gate11558  (.A(II29243), .Z(g22639) ) ;
NOR2    gate11559  (.A(g19698), .B(g17577), .Z(g20922) ) ;
INV     gate11560  (.A(g20922), .Z(II29246) ) ;
INV     gate11561  (.A(II29246), .Z(g22640) ) ;
NOR2    gate11562  (.A(g19699), .B(g17578), .Z(g20923) ) ;
INV     gate11563  (.A(g20923), .Z(II29249) ) ;
INV     gate11564  (.A(II29249), .Z(g22641) ) ;
NOR2    gate11565  (.A(g19700), .B(g15257), .Z(g20924) ) ;
INV     gate11566  (.A(g20924), .Z(II29252) ) ;
INV     gate11567  (.A(II29252), .Z(g22642) ) ;
INV     gate11568  (.A(g21125), .Z(g22645) ) ;
NOR2    gate11569  (.A(g19708), .B(g17598), .Z(g20925) ) ;
INV     gate11570  (.A(g20925), .Z(II29259) ) ;
INV     gate11571  (.A(II29259), .Z(g22647) ) ;
NOR2    gate11572  (.A(g19709), .B(g17599), .Z(g20926) ) ;
INV     gate11573  (.A(g20926), .Z(II29262) ) ;
INV     gate11574  (.A(II29262), .Z(g22648) ) ;
NOR2    gate11575  (.A(g19710), .B(g17600), .Z(g20927) ) ;
INV     gate11576  (.A(g20927), .Z(II29265) ) ;
INV     gate11577  (.A(II29265), .Z(g22649) ) ;
NOR2    gate11578  (.A(g19171), .B(g10238), .Z(g20752) ) ;
INV     gate11579  (.A(g20752), .Z(II29271) ) ;
INV     gate11580  (.A(II29271), .Z(g22655) ) ;
NOR2    gate11581  (.A(g19714), .B(g17617), .Z(g20934) ) ;
INV     gate11582  (.A(g20934), .Z(II29274) ) ;
INV     gate11583  (.A(II29274), .Z(g22656) ) ;
NOR2    gate11584  (.A(g19715), .B(g17618), .Z(g20935) ) ;
INV     gate11585  (.A(g20935), .Z(II29277) ) ;
INV     gate11586  (.A(II29277), .Z(g22657) ) ;
NOR2    gate11587  (.A(g19716), .B(g17619), .Z(g20936) ) ;
INV     gate11588  (.A(g20936), .Z(II29280) ) ;
INV     gate11589  (.A(II29280), .Z(g22658) ) ;
NOR2    gate11590  (.A(g19717), .B(g17620), .Z(g20937) ) ;
INV     gate11591  (.A(g20937), .Z(II29283) ) ;
INV     gate11592  (.A(II29283), .Z(g22659) ) ;
INV     gate11593  (.A(g21130), .Z(g22661) ) ;
NOR2    gate11594  (.A(g19722), .B(g17632), .Z(g20939) ) ;
INV     gate11595  (.A(g20939), .Z(II29288) ) ;
INV     gate11596  (.A(II29288), .Z(g22662) ) ;
NOR2    gate11597  (.A(g19723), .B(g17633), .Z(g20940) ) ;
INV     gate11598  (.A(g20940), .Z(II29291) ) ;
INV     gate11599  (.A(II29291), .Z(g22663) ) ;
NOR2    gate11600  (.A(g19724), .B(g17634), .Z(g20941) ) ;
INV     gate11601  (.A(g20941), .Z(II29294) ) ;
INV     gate11602  (.A(II29294), .Z(g22664) ) ;
NOR2    gate11603  (.A(g19731), .B(g17652), .Z(g20944) ) ;
INV     gate11604  (.A(g20944), .Z(II29301) ) ;
INV     gate11605  (.A(II29301), .Z(g22669) ) ;
NOR2    gate11606  (.A(g19732), .B(g17653), .Z(g20945) ) ;
INV     gate11607  (.A(g20945), .Z(II29304) ) ;
INV     gate11608  (.A(II29304), .Z(g22670) ) ;
NOR2    gate11609  (.A(g19733), .B(g17654), .Z(g20946) ) ;
INV     gate11610  (.A(g20946), .Z(II29307) ) ;
INV     gate11611  (.A(II29307), .Z(g22671) ) ;
NOR2    gate11612  (.A(g19734), .B(g15335), .Z(g20947) ) ;
INV     gate11613  (.A(g20947), .Z(II29310) ) ;
INV     gate11614  (.A(II29310), .Z(g22672) ) ;
NOR2    gate11615  (.A(g19735), .B(g15336), .Z(g20948) ) ;
INV     gate11616  (.A(g20948), .Z(II29313) ) ;
INV     gate11617  (.A(II29313), .Z(g22673) ) ;
NOR2    gate11618  (.A(g19741), .B(g17673), .Z(g20949) ) ;
INV     gate11619  (.A(g20949), .Z(II29317) ) ;
INV     gate11620  (.A(II29317), .Z(g22675) ) ;
NOR2    gate11621  (.A(g19742), .B(g17674), .Z(g20950) ) ;
INV     gate11622  (.A(g20950), .Z(II29320) ) ;
INV     gate11623  (.A(II29320), .Z(g22676) ) ;
NOR2    gate11624  (.A(g19743), .B(g17675), .Z(g20951) ) ;
INV     gate11625  (.A(g20951), .Z(II29323) ) ;
INV     gate11626  (.A(II29323), .Z(g22677) ) ;
NOR2    gate11627  (.A(g19744), .B(g15349), .Z(g20952) ) ;
INV     gate11628  (.A(g20952), .Z(II29326) ) ;
INV     gate11629  (.A(II29326), .Z(g22678) ) ;
INV     gate11630  (.A(g21144), .Z(g22681) ) ;
NOR2    gate11631  (.A(g19752), .B(g17695), .Z(g20953) ) ;
INV     gate11632  (.A(g20953), .Z(II29333) ) ;
INV     gate11633  (.A(II29333), .Z(g22683) ) ;
NOR2    gate11634  (.A(g19753), .B(g17696), .Z(g20954) ) ;
INV     gate11635  (.A(g20954), .Z(II29336) ) ;
INV     gate11636  (.A(II29336), .Z(g22684) ) ;
NOR2    gate11637  (.A(g19754), .B(g17697), .Z(g20955) ) ;
INV     gate11638  (.A(g20955), .Z(II29339) ) ;
INV     gate11639  (.A(II29339), .Z(g22685) ) ;
NOR2    gate11640  (.A(g19177), .B(g10340), .Z(g20789) ) ;
INV     gate11641  (.A(g20789), .Z(II29345) ) ;
INV     gate11642  (.A(II29345), .Z(g22691) ) ;
NOR2    gate11643  (.A(g19758), .B(g17714), .Z(g20962) ) ;
INV     gate11644  (.A(g20962), .Z(II29348) ) ;
INV     gate11645  (.A(II29348), .Z(g22692) ) ;
NOR2    gate11646  (.A(g19759), .B(g17715), .Z(g20963) ) ;
INV     gate11647  (.A(g20963), .Z(II29351) ) ;
INV     gate11648  (.A(II29351), .Z(g22693) ) ;
NOR2    gate11649  (.A(g19760), .B(g17716), .Z(g20964) ) ;
INV     gate11650  (.A(g20964), .Z(II29354) ) ;
INV     gate11651  (.A(II29354), .Z(g22694) ) ;
NOR2    gate11652  (.A(g19761), .B(g17717), .Z(g20965) ) ;
INV     gate11653  (.A(g20965), .Z(II29357) ) ;
INV     gate11654  (.A(II29357), .Z(g22695) ) ;
NOR2    gate11655  (.A(g19830), .B(g13004), .Z(g21796) ) ;
INV     gate11656  (.A(g21796), .Z(II29360) ) ;
INV     gate11657  (.A(II29360), .Z(g22696) ) ;
NOR2    gate11658  (.A(g19765), .B(g17734), .Z(g20966) ) ;
INV     gate11659  (.A(g20966), .Z(II29366) ) ;
INV     gate11660  (.A(II29366), .Z(g22702) ) ;
NOR2    gate11661  (.A(g19766), .B(g17735), .Z(g20967) ) ;
INV     gate11662  (.A(g20967), .Z(II29369) ) ;
INV     gate11663  (.A(II29369), .Z(g22703) ) ;
NOR2    gate11664  (.A(g19767), .B(g17736), .Z(g20968) ) ;
INV     gate11665  (.A(g20968), .Z(II29372) ) ;
INV     gate11666  (.A(II29372), .Z(g22704) ) ;
NOR2    gate11667  (.A(g19768), .B(g15402), .Z(g20969) ) ;
INV     gate11668  (.A(g20969), .Z(II29375) ) ;
INV     gate11669  (.A(II29375), .Z(g22705) ) ;
NOR2    gate11670  (.A(g19769), .B(g15403), .Z(g20970) ) ;
INV     gate11671  (.A(g20970), .Z(II29378) ) ;
INV     gate11672  (.A(II29378), .Z(g22706) ) ;
NOR2    gate11673  (.A(g19774), .B(g17752), .Z(g20972) ) ;
INV     gate11674  (.A(g20972), .Z(II29383) ) ;
INV     gate11675  (.A(II29383), .Z(g22709) ) ;
NOR2    gate11676  (.A(g19775), .B(g17753), .Z(g20973) ) ;
INV     gate11677  (.A(g20973), .Z(II29386) ) ;
INV     gate11678  (.A(II29386), .Z(g22710) ) ;
NOR2    gate11679  (.A(g19776), .B(g17754), .Z(g20974) ) ;
INV     gate11680  (.A(g20974), .Z(II29389) ) ;
INV     gate11681  (.A(II29389), .Z(g22711) ) ;
NOR2    gate11682  (.A(g19777), .B(g15421), .Z(g20975) ) ;
INV     gate11683  (.A(g20975), .Z(II29392) ) ;
INV     gate11684  (.A(II29392), .Z(g22712) ) ;
NOR2    gate11685  (.A(g19778), .B(g15422), .Z(g20976) ) ;
INV     gate11686  (.A(g20976), .Z(II29395) ) ;
INV     gate11687  (.A(II29395), .Z(g22713) ) ;
NOR2    gate11688  (.A(g19784), .B(g17773), .Z(g20977) ) ;
INV     gate11689  (.A(g20977), .Z(II29399) ) ;
INV     gate11690  (.A(II29399), .Z(g22715) ) ;
NOR2    gate11691  (.A(g19785), .B(g17774), .Z(g20978) ) ;
INV     gate11692  (.A(g20978), .Z(II29402) ) ;
INV     gate11693  (.A(II29402), .Z(g22716) ) ;
NOR2    gate11694  (.A(g19786), .B(g17775), .Z(g20979) ) ;
INV     gate11695  (.A(g20979), .Z(II29405) ) ;
INV     gate11696  (.A(II29405), .Z(g22717) ) ;
NOR2    gate11697  (.A(g19787), .B(g15435), .Z(g20980) ) ;
INV     gate11698  (.A(g20980), .Z(II29408) ) ;
INV     gate11699  (.A(II29408), .Z(g22718) ) ;
INV     gate11700  (.A(g21164), .Z(g22721) ) ;
NOR2    gate11701  (.A(g19795), .B(g17795), .Z(g20981) ) ;
INV     gate11702  (.A(g20981), .Z(II29415) ) ;
INV     gate11703  (.A(II29415), .Z(g22723) ) ;
NOR2    gate11704  (.A(g19796), .B(g17796), .Z(g20982) ) ;
INV     gate11705  (.A(g20982), .Z(II29418) ) ;
INV     gate11706  (.A(II29418), .Z(g22724) ) ;
NOR2    gate11707  (.A(g19797), .B(g17797), .Z(g20983) ) ;
INV     gate11708  (.A(g20983), .Z(II29421) ) ;
INV     gate11709  (.A(II29421), .Z(g22725) ) ;
NOR2    gate11710  (.A(g19802), .B(g17812), .Z(g20989) ) ;
INV     gate11711  (.A(g20989), .Z(II29426) ) ;
INV     gate11712  (.A(II29426), .Z(g22728) ) ;
NOR2    gate11713  (.A(g19803), .B(g17813), .Z(g20990) ) ;
INV     gate11714  (.A(g20990), .Z(II29429) ) ;
INV     gate11715  (.A(II29429), .Z(g22729) ) ;
NOR2    gate11716  (.A(g19804), .B(g17814), .Z(g20991) ) ;
INV     gate11717  (.A(g20991), .Z(II29432) ) ;
INV     gate11718  (.A(II29432), .Z(g22730) ) ;
NOR2    gate11719  (.A(g19805), .B(g15470), .Z(g20992) ) ;
INV     gate11720  (.A(g20992), .Z(II29435) ) ;
INV     gate11721  (.A(II29435), .Z(g22731) ) ;
NOR2    gate11722  (.A(g19807), .B(g17835), .Z(g20993) ) ;
INV     gate11723  (.A(g20993), .Z(II29439) ) ;
INV     gate11724  (.A(II29439), .Z(g22733) ) ;
NOR2    gate11725  (.A(g19808), .B(g17836), .Z(g20994) ) ;
INV     gate11726  (.A(g20994), .Z(II29442) ) ;
INV     gate11727  (.A(II29442), .Z(g22734) ) ;
NOR2    gate11728  (.A(g19809), .B(g17837), .Z(g20995) ) ;
INV     gate11729  (.A(g20995), .Z(II29445) ) ;
INV     gate11730  (.A(II29445), .Z(g22735) ) ;
NOR2    gate11731  (.A(g19810), .B(g15486), .Z(g20996) ) ;
INV     gate11732  (.A(g20996), .Z(II29448) ) ;
INV     gate11733  (.A(II29448), .Z(g22736) ) ;
NOR2    gate11734  (.A(g19811), .B(g15487), .Z(g20997) ) ;
INV     gate11735  (.A(g20997), .Z(II29451) ) ;
INV     gate11736  (.A(II29451), .Z(g22737) ) ;
NOR2    gate11737  (.A(g19816), .B(g17853), .Z(g20999) ) ;
INV     gate11738  (.A(g20999), .Z(II29456) ) ;
INV     gate11739  (.A(II29456), .Z(g22740) ) ;
NOR2    gate11740  (.A(g19817), .B(g17854), .Z(g21000) ) ;
INV     gate11741  (.A(g21000), .Z(II29459) ) ;
INV     gate11742  (.A(II29459), .Z(g22741) ) ;
NOR2    gate11743  (.A(g19818), .B(g17855), .Z(g21001) ) ;
INV     gate11744  (.A(g21001), .Z(II29462) ) ;
INV     gate11745  (.A(II29462), .Z(g22742) ) ;
NOR2    gate11746  (.A(g19819), .B(g15505), .Z(g21002) ) ;
INV     gate11747  (.A(g21002), .Z(II29465) ) ;
INV     gate11748  (.A(II29465), .Z(g22743) ) ;
NOR2    gate11749  (.A(g19820), .B(g15506), .Z(g21003) ) ;
INV     gate11750  (.A(g21003), .Z(II29468) ) ;
INV     gate11751  (.A(II29468), .Z(g22744) ) ;
NOR2    gate11752  (.A(g19826), .B(g17874), .Z(g21004) ) ;
INV     gate11753  (.A(g21004), .Z(II29472) ) ;
INV     gate11754  (.A(II29472), .Z(g22746) ) ;
NOR2    gate11755  (.A(g19827), .B(g17875), .Z(g21005) ) ;
INV     gate11756  (.A(g21005), .Z(II29475) ) ;
INV     gate11757  (.A(II29475), .Z(g22747) ) ;
NOR2    gate11758  (.A(g19828), .B(g17876), .Z(g21006) ) ;
INV     gate11759  (.A(g21006), .Z(II29478) ) ;
INV     gate11760  (.A(II29478), .Z(g22748) ) ;
NOR2    gate11761  (.A(g19829), .B(g15519), .Z(g21007) ) ;
INV     gate11762  (.A(g21007), .Z(II29481) ) ;
INV     gate11763  (.A(II29481), .Z(g22749) ) ;
NAND2   gate11764  (.A(g20008), .B(g3013), .Z(g21903) ) ;
INV     gate11765  (.A(g21903), .Z(II29484) ) ;
INV     gate11766  (.A(II29484), .Z(g22750) ) ;
INV     gate11767  (.A(g21184), .Z(g22753) ) ;
NOR2    gate11768  (.A(g19839), .B(g17900), .Z(g21009) ) ;
INV     gate11769  (.A(g21009), .Z(II29490) ) ;
INV     gate11770  (.A(II29490), .Z(g22756) ) ;
NOR2    gate11771  (.A(g19840), .B(g17901), .Z(g21010) ) ;
INV     gate11772  (.A(g21010), .Z(II29493) ) ;
INV     gate11773  (.A(II29493), .Z(g22757) ) ;
NOR2    gate11774  (.A(g19841), .B(g17902), .Z(g21011) ) ;
INV     gate11775  (.A(g21011), .Z(II29496) ) ;
INV     gate11776  (.A(II29496), .Z(g22758) ) ;
NOR2    gate11777  (.A(g19846), .B(g17924), .Z(g21015) ) ;
INV     gate11778  (.A(g21015), .Z(II29500) ) ;
INV     gate11779  (.A(II29500), .Z(g22760) ) ;
NOR2    gate11780  (.A(g19847), .B(g17925), .Z(g21016) ) ;
INV     gate11781  (.A(g21016), .Z(II29503) ) ;
INV     gate11782  (.A(II29503), .Z(g22761) ) ;
NOR2    gate11783  (.A(g19848), .B(g17926), .Z(g21017) ) ;
INV     gate11784  (.A(g21017), .Z(II29506) ) ;
INV     gate11785  (.A(II29506), .Z(g22762) ) ;
NOR2    gate11786  (.A(g19849), .B(g15556), .Z(g21018) ) ;
INV     gate11787  (.A(g21018), .Z(II29509) ) ;
INV     gate11788  (.A(II29509), .Z(g22763) ) ;
NOR2    gate11789  (.A(g19851), .B(g17947), .Z(g21019) ) ;
INV     gate11790  (.A(g21019), .Z(II29513) ) ;
INV     gate11791  (.A(II29513), .Z(g22765) ) ;
NOR2    gate11792  (.A(g19852), .B(g17948), .Z(g21020) ) ;
INV     gate11793  (.A(g21020), .Z(II29516) ) ;
INV     gate11794  (.A(II29516), .Z(g22766) ) ;
NOR2    gate11795  (.A(g19853), .B(g17949), .Z(g21021) ) ;
INV     gate11796  (.A(g21021), .Z(II29519) ) ;
INV     gate11797  (.A(II29519), .Z(g22767) ) ;
NOR2    gate11798  (.A(g19854), .B(g15572), .Z(g21022) ) ;
INV     gate11799  (.A(g21022), .Z(II29522) ) ;
INV     gate11800  (.A(II29522), .Z(g22768) ) ;
NOR2    gate11801  (.A(g19855), .B(g15573), .Z(g21023) ) ;
INV     gate11802  (.A(g21023), .Z(II29525) ) ;
INV     gate11803  (.A(II29525), .Z(g22769) ) ;
NOR2    gate11804  (.A(g19860), .B(g17965), .Z(g21025) ) ;
INV     gate11805  (.A(g21025), .Z(II29530) ) ;
INV     gate11806  (.A(II29530), .Z(g22772) ) ;
NOR2    gate11807  (.A(g19861), .B(g17966), .Z(g21026) ) ;
INV     gate11808  (.A(g21026), .Z(II29533) ) ;
INV     gate11809  (.A(II29533), .Z(g22773) ) ;
NOR2    gate11810  (.A(g19862), .B(g17967), .Z(g21027) ) ;
INV     gate11811  (.A(g21027), .Z(II29536) ) ;
INV     gate11812  (.A(II29536), .Z(g22774) ) ;
NOR2    gate11813  (.A(g19863), .B(g15591), .Z(g21028) ) ;
INV     gate11814  (.A(g21028), .Z(II29539) ) ;
INV     gate11815  (.A(II29539), .Z(g22775) ) ;
NOR2    gate11816  (.A(g19864), .B(g15592), .Z(g21029) ) ;
INV     gate11817  (.A(g21029), .Z(II29542) ) ;
INV     gate11818  (.A(II29542), .Z(g22776) ) ;
INV     gate11819  (.A(g21796), .Z(g22777) ) ;
NOR2    gate11820  (.A(g19869), .B(g17989), .Z(g21031) ) ;
INV     gate11821  (.A(g21031), .Z(II29547) ) ;
INV     gate11822  (.A(II29547), .Z(g22785) ) ;
NOR2    gate11823  (.A(g19870), .B(g17990), .Z(g21032) ) ;
INV     gate11824  (.A(g21032), .Z(II29550) ) ;
INV     gate11825  (.A(II29550), .Z(g22786) ) ;
INV     gate11826  (.A(g21199), .Z(g22787) ) ;
NOR2    gate11827  (.A(g19872), .B(g18011), .Z(g21033) ) ;
INV     gate11828  (.A(g21033), .Z(II29556) ) ;
INV     gate11829  (.A(II29556), .Z(g22790) ) ;
NOR2    gate11830  (.A(g19873), .B(g18012), .Z(g21034) ) ;
INV     gate11831  (.A(g21034), .Z(II29559) ) ;
INV     gate11832  (.A(II29559), .Z(g22791) ) ;
NOR2    gate11833  (.A(g19874), .B(g18013), .Z(g21035) ) ;
INV     gate11834  (.A(g21035), .Z(II29562) ) ;
INV     gate11835  (.A(II29562), .Z(g22792) ) ;
NOR2    gate11836  (.A(g19879), .B(g18035), .Z(g21039) ) ;
INV     gate11837  (.A(g21039), .Z(II29566) ) ;
INV     gate11838  (.A(II29566), .Z(g22794) ) ;
NOR2    gate11839  (.A(g19880), .B(g18036), .Z(g21040) ) ;
INV     gate11840  (.A(g21040), .Z(II29569) ) ;
INV     gate11841  (.A(II29569), .Z(g22795) ) ;
NOR2    gate11842  (.A(g19881), .B(g18037), .Z(g21041) ) ;
INV     gate11843  (.A(g21041), .Z(II29572) ) ;
INV     gate11844  (.A(II29572), .Z(g22796) ) ;
NOR2    gate11845  (.A(g19882), .B(g15634), .Z(g21042) ) ;
INV     gate11846  (.A(g21042), .Z(II29575) ) ;
INV     gate11847  (.A(II29575), .Z(g22797) ) ;
NOR2    gate11848  (.A(g19884), .B(g18058), .Z(g21043) ) ;
INV     gate11849  (.A(g21043), .Z(II29579) ) ;
INV     gate11850  (.A(II29579), .Z(g22799) ) ;
NOR2    gate11851  (.A(g19885), .B(g18059), .Z(g21044) ) ;
INV     gate11852  (.A(g21044), .Z(II29582) ) ;
INV     gate11853  (.A(II29582), .Z(g22800) ) ;
NOR2    gate11854  (.A(g19886), .B(g18060), .Z(g21045) ) ;
INV     gate11855  (.A(g21045), .Z(II29585) ) ;
INV     gate11856  (.A(II29585), .Z(g22801) ) ;
NOR2    gate11857  (.A(g19887), .B(g15650), .Z(g21046) ) ;
INV     gate11858  (.A(g21046), .Z(II29588) ) ;
INV     gate11859  (.A(II29588), .Z(g22802) ) ;
NOR2    gate11860  (.A(g19888), .B(g15651), .Z(g21047) ) ;
INV     gate11861  (.A(g21047), .Z(II29591) ) ;
INV     gate11862  (.A(II29591), .Z(g22803) ) ;
NOR2    gate11863  (.A(g19317), .B(g19356), .Z(g21894) ) ;
INV     gate11864  (.A(g21894), .Z(g22805) ) ;
NOR2    gate11865  (.A(g16567), .B(g19957), .Z(g21615) ) ;
INV     gate11866  (.A(g21615), .Z(g22806) ) ;
NAND4   gate11867  (.A(g14256), .B(g15177), .C(g19871), .D(g19842), .Z(g21720) ) ;
INV     gate11868  (.A(g21720), .Z(II29600) ) ;
INV     gate11869  (.A(II29600), .Z(g22812) ) ;
NOR2    gate11870  (.A(g19895), .B(g18088), .Z(g21051) ) ;
INV     gate11871  (.A(g21051), .Z(II29603) ) ;
INV     gate11872  (.A(II29603), .Z(g22824) ) ;
NOR2    gate11873  (.A(g20486), .B(g13266), .Z(g21364) ) ;
INV     gate11874  (.A(g21364), .Z(II29606) ) ;
INV     gate11875  (.A(II29606), .Z(g22825) ) ;
NOR2    gate11876  (.A(g19900), .B(g18106), .Z(g21052) ) ;
INV     gate11877  (.A(g21052), .Z(II29610) ) ;
INV     gate11878  (.A(II29610), .Z(g22827) ) ;
NOR2    gate11879  (.A(g19901), .B(g18107), .Z(g21053) ) ;
INV     gate11880  (.A(g21053), .Z(II29613) ) ;
INV     gate11881  (.A(II29613), .Z(g22828) ) ;
INV     gate11882  (.A(g21214), .Z(g22829) ) ;
NOR2    gate11883  (.A(g19903), .B(g18128), .Z(g21054) ) ;
INV     gate11884  (.A(g21054), .Z(II29619) ) ;
INV     gate11885  (.A(II29619), .Z(g22832) ) ;
NOR2    gate11886  (.A(g19904), .B(g18129), .Z(g21055) ) ;
INV     gate11887  (.A(g21055), .Z(II29622) ) ;
INV     gate11888  (.A(II29622), .Z(g22833) ) ;
NOR2    gate11889  (.A(g19905), .B(g18130), .Z(g21056) ) ;
INV     gate11890  (.A(g21056), .Z(II29625) ) ;
INV     gate11891  (.A(II29625), .Z(g22834) ) ;
NOR2    gate11892  (.A(g19910), .B(g18152), .Z(g21060) ) ;
INV     gate11893  (.A(g21060), .Z(II29629) ) ;
INV     gate11894  (.A(II29629), .Z(g22836) ) ;
NOR2    gate11895  (.A(g19911), .B(g18153), .Z(g21061) ) ;
INV     gate11896  (.A(g21061), .Z(II29632) ) ;
INV     gate11897  (.A(II29632), .Z(g22837) ) ;
NOR2    gate11898  (.A(g19912), .B(g18154), .Z(g21062) ) ;
INV     gate11899  (.A(g21062), .Z(II29635) ) ;
INV     gate11900  (.A(II29635), .Z(g22838) ) ;
NOR2    gate11901  (.A(g19913), .B(g15710), .Z(g21063) ) ;
INV     gate11902  (.A(g21063), .Z(II29638) ) ;
INV     gate11903  (.A(II29638), .Z(g22839) ) ;
NAND2   gate11904  (.A(g19219), .B(g15959), .Z(g20825) ) ;
INV     gate11905  (.A(g20825), .Z(II29641) ) ;
INV     gate11906  (.A(II29641), .Z(g22840) ) ;
NOR2    gate11907  (.A(g19285), .B(g19316), .Z(g21889) ) ;
INV     gate11908  (.A(g21889), .Z(g22843) ) ;
NOR2    gate11909  (.A(g16591), .B(g19987), .Z(g21643) ) ;
INV     gate11910  (.A(g21643), .Z(g22847) ) ;
NAND4   gate11911  (.A(g14378), .B(g15263), .C(g19902), .D(g19875), .Z(g21746) ) ;
INV     gate11912  (.A(g21746), .Z(II29653) ) ;
INV     gate11913  (.A(II29653), .Z(g22852) ) ;
NOR2    gate11914  (.A(g19920), .B(g18204), .Z(g21070) ) ;
INV     gate11915  (.A(g21070), .Z(II29656) ) ;
INV     gate11916  (.A(II29656), .Z(g22864) ) ;
NOR2    gate11917  (.A(g19925), .B(g18222), .Z(g21071) ) ;
INV     gate11918  (.A(g21071), .Z(II29660) ) ;
INV     gate11919  (.A(II29660), .Z(g22866) ) ;
NOR2    gate11920  (.A(g19926), .B(g18223), .Z(g21072) ) ;
INV     gate11921  (.A(g21072), .Z(II29663) ) ;
INV     gate11922  (.A(II29663), .Z(g22867) ) ;
INV     gate11923  (.A(g21222), .Z(g22868) ) ;
NOR2    gate11924  (.A(g19928), .B(g18244), .Z(g21073) ) ;
INV     gate11925  (.A(g21073), .Z(II29669) ) ;
INV     gate11926  (.A(II29669), .Z(g22871) ) ;
NOR2    gate11927  (.A(g19929), .B(g18245), .Z(g21074) ) ;
INV     gate11928  (.A(g21074), .Z(II29672) ) ;
INV     gate11929  (.A(II29672), .Z(g22872) ) ;
NOR2    gate11930  (.A(g19930), .B(g18246), .Z(g21075) ) ;
INV     gate11931  (.A(g21075), .Z(II29675) ) ;
INV     gate11932  (.A(II29675), .Z(g22873) ) ;
NOR2    gate11933  (.A(g19260), .B(g19284), .Z(g21884) ) ;
INV     gate11934  (.A(g21884), .Z(g22875) ) ;
NOR2    gate11935  (.A(g16611), .B(g20025), .Z(g21674) ) ;
INV     gate11936  (.A(g21674), .Z(g22882) ) ;
NAND4   gate11937  (.A(g14490), .B(g15355), .C(g19927), .D(g19906), .Z(g21770) ) ;
INV     gate11938  (.A(g21770), .Z(II29687) ) ;
INV     gate11939  (.A(II29687), .Z(g22887) ) ;
NOR2    gate11940  (.A(g19935), .B(g18311), .Z(g21080) ) ;
INV     gate11941  (.A(g21080), .Z(II29690) ) ;
INV     gate11942  (.A(II29690), .Z(g22899) ) ;
NOR2    gate11943  (.A(g19940), .B(g18329), .Z(g21081) ) ;
INV     gate11944  (.A(g21081), .Z(II29694) ) ;
INV     gate11945  (.A(II29694), .Z(g22901) ) ;
NOR2    gate11946  (.A(g19941), .B(g18330), .Z(g21082) ) ;
INV     gate11947  (.A(g21082), .Z(II29697) ) ;
INV     gate11948  (.A(II29697), .Z(g22902) ) ;
NAND2   gate11949  (.A(g20153), .B(g2903), .Z(g20700) ) ;
INV     gate11950  (.A(g20700), .Z(II29700) ) ;
INV     gate11951  (.A(II29700), .Z(g22903) ) ;
NOR2    gate11952  (.A(g19830), .B(g15780), .Z(g21711) ) ;
INV     gate11953  (.A(g21711), .Z(g22907) ) ;
NOR2    gate11954  (.A(g16629), .B(g20067), .Z(g21703) ) ;
INV     gate11955  (.A(g21703), .Z(g22917) ) ;
NAND4   gate11956  (.A(g14577), .B(g15441), .C(g19942), .D(g19931), .Z(g21786) ) ;
INV     gate11957  (.A(g21786), .Z(II29712) ) ;
INV     gate11958  (.A(II29712), .Z(g22922) ) ;
NOR2    gate11959  (.A(g19952), .B(g18404), .Z(g21094) ) ;
INV     gate11960  (.A(g21094), .Z(II29715) ) ;
INV     gate11961  (.A(II29715), .Z(g22934) ) ;
INV     gate11962  (.A(g21851), .Z(II29724) ) ;
INV     gate11963  (.A(II29724), .Z(g22945) ) ;
NOR2    gate11964  (.A(g3919), .B(g19830), .Z(g20877) ) ;
INV     gate11965  (.A(g20877), .Z(II29727) ) ;
INV     gate11966  (.A(II29727), .Z(g22948) ) ;
NOR2    gate11967  (.A(g20507), .B(g18352), .Z(g21665) ) ;
INV     gate11968  (.A(g21665), .Z(g22949) ) ;
NOR2    gate11969  (.A(g20507), .B(g18430), .Z(g21739) ) ;
INV     gate11970  (.A(g21739), .Z(g22954) ) ;
NOR2    gate11971  (.A(g20526), .B(g18447), .Z(g21694) ) ;
INV     gate11972  (.A(g21694), .Z(g22958) ) ;
NOR2    gate11973  (.A(g20526), .B(g18503), .Z(g21763) ) ;
INV     gate11974  (.A(g21763), .Z(g22962) ) ;
NOR2    gate11975  (.A(g20545), .B(g18520), .Z(g21730) ) ;
INV     gate11976  (.A(g21730), .Z(g22966) ) ;
NOR2    gate11977  (.A(g5394), .B(g19830), .Z(g20884) ) ;
INV     gate11978  (.A(g20884), .Z(II29736) ) ;
INV     gate11979  (.A(II29736), .Z(g22970) ) ;
NOR2    gate11980  (.A(g20545), .B(g18567), .Z(g21779) ) ;
INV     gate11981  (.A(g21779), .Z(g22971) ) ;
NOR2    gate11982  (.A(g19070), .B(g18584), .Z(g21756) ) ;
INV     gate11983  (.A(g21756), .Z(g22975) ) ;
NOR2    gate11984  (.A(g20480), .B(g13247), .Z(g21346) ) ;
INV     gate11985  (.A(g21346), .Z(II29741) ) ;
INV     gate11986  (.A(II29741), .Z(g22979) ) ;
NOR2    gate11987  (.A(g19070), .B(g18617), .Z(g21794) ) ;
INV     gate11988  (.A(g21794), .Z(g22980) ) ;
INV     gate11989  (.A(g21382), .Z(g22986) ) ;
INV     gate11990  (.A(g21404), .Z(g22988) ) ;
INV     gate11991  (.A(g21415), .Z(g22989) ) ;
INV     gate11992  (.A(g21429), .Z(g22991) ) ;
INV     gate11993  (.A(g21441), .Z(g22995) ) ;
INV     gate11994  (.A(g21449), .Z(g22996) ) ;
INV     gate11995  (.A(g21458), .Z(g22998) ) ;
INV     gate11996  (.A(g21473), .Z(g23001) ) ;
INV     gate11997  (.A(g21477), .Z(g23002) ) ;
INV     gate11998  (.A(g21483), .Z(g23006) ) ;
INV     gate11999  (.A(g21491), .Z(g23007) ) ;
INV     gate12000  (.A(g21498), .Z(g23008) ) ;
INV     gate12001  (.A(g21505), .Z(g23012) ) ;
INV     gate12002  (.A(g21514), .Z(g23015) ) ;
INV     gate12003  (.A(g21518), .Z(g23016) ) ;
INV     gate12004  (.A(g21524), .Z(g23020) ) ;
INV     gate12005  (.A(g21530), .Z(g23021) ) ;
INV     gate12006  (.A(g21537), .Z(g23024) ) ;
INV     gate12007  (.A(g21541), .Z(g23028) ) ;
INV     gate12008  (.A(g21550), .Z(g23031) ) ;
INV     gate12009  (.A(g21554), .Z(g23032) ) ;
INV     gate12010  (.A(g21558), .Z(g23036) ) ;
INV     gate12011  (.A(g21561), .Z(g23037) ) ;
INV     gate12012  (.A(g21566), .Z(g23038) ) ;
INV     gate12013  (.A(g21573), .Z(g23041) ) ;
INV     gate12014  (.A(g21577), .Z(g23045) ) ;
INV     gate12015  (.A(g21586), .Z(g23048) ) ;
INV     gate12016  (.A(g21590), .Z(g23049) ) ;
INV     gate12017  (.A(g21432), .Z(II29797) ) ;
INV     gate12018  (.A(II29797), .Z(g23050) ) ;
INV     gate12019  (.A(g21435), .Z(II29802) ) ;
INV     gate12020  (.A(II29802), .Z(g23055) ) ;
INV     gate12021  (.A(g21594), .Z(g23056) ) ;
INV     gate12022  (.A(g21599), .Z(g23057) ) ;
INV     gate12023  (.A(g21606), .Z(g23060) ) ;
INV     gate12024  (.A(g21612), .Z(g23064) ) ;
INV     gate12025  (.A(g21467), .Z(II29812) ) ;
INV     gate12026  (.A(II29812), .Z(g23065) ) ;
INV     gate12027  (.A(g21470), .Z(II29817) ) ;
INV     gate12028  (.A(II29817), .Z(g23068) ) ;
INV     gate12029  (.A(g21619), .Z(g23069) ) ;
INV     gate12030  (.A(g21623), .Z(g23074) ) ;
INV     gate12031  (.A(g21628), .Z(g23075) ) ;
INV     gate12032  (.A(g21502), .Z(II29827) ) ;
INV     gate12033  (.A(II29827), .Z(g23078) ) ;
INV     gate12034  (.A(g21640), .Z(g23079) ) ;
INV     gate12035  (.A(g21647), .Z(g23082) ) ;
INV     gate12036  (.A(g21651), .Z(g23087) ) ;
INV     gate12037  (.A(g21655), .Z(g23088) ) ;
INV     gate12038  (.A(g21316), .Z(II29841) ) ;
INV     gate12039  (.A(II29841), .Z(g23094) ) ;
INV     gate12040  (.A(g21671), .Z(g23095) ) ;
INV     gate12041  (.A(g21678), .Z(g23098) ) ;
INV     gate12042  (.A(g21682), .Z(g23103) ) ;
INV     gate12043  (.A(g21331), .Z(II29852) ) ;
INV     gate12044  (.A(II29852), .Z(g23105) ) ;
INV     gate12045  (.A(g21700), .Z(g23112) ) ;
INV     gate12046  (.A(g21708), .Z(g23115) ) ;
INV     gate12047  (.A(g21346), .Z(II29863) ) ;
INV     gate12048  (.A(II29863), .Z(g23116) ) ;
INV     gate12049  (.A(g21364), .Z(II29872) ) ;
INV     gate12050  (.A(II29872), .Z(g23125) ) ;
INV     gate12051  (.A(g21385), .Z(II29881) ) ;
INV     gate12052  (.A(II29881), .Z(g23134) ) ;
INV     gate12053  (.A(g21825), .Z(g23140) ) ;
INV     gate12054  (.A(g21825), .Z(g23141) ) ;
INV     gate12055  (.A(g21825), .Z(g23142) ) ;
INV     gate12056  (.A(g21825), .Z(g23143) ) ;
INV     gate12057  (.A(g21825), .Z(g23144) ) ;
INV     gate12058  (.A(g21825), .Z(g23145) ) ;
INV     gate12059  (.A(g21825), .Z(g23146) ) ;
INV     gate12060  (.A(g21825), .Z(g23147) ) ;
INV     gate12061  (.A(g23116), .Z(II29897) ) ;
INV     gate12062  (.A(g23125), .Z(II29900) ) ;
INV     gate12063  (.A(g23134), .Z(II29903) ) ;
INV     gate12064  (.A(g21967), .Z(II29906) ) ;
INV     gate12065  (.A(g23050), .Z(II29909) ) ;
INV     gate12066  (.A(g23065), .Z(II29912) ) ;
INV     gate12067  (.A(g23055), .Z(II29915) ) ;
INV     gate12068  (.A(g23068), .Z(II29918) ) ;
INV     gate12069  (.A(g23078), .Z(II29921) ) ;
INV     gate12070  (.A(g23094), .Z(II29924) ) ;
INV     gate12071  (.A(g23105), .Z(II29927) ) ;
INV     gate12072  (.A(g22176), .Z(II29930) ) ;
INV     gate12073  (.A(g22082), .Z(II29933) ) ;
INV     gate12074  (.A(g22582), .Z(II29936) ) ;
INV     gate12075  (.A(g22518), .Z(II29939) ) ;
INV     gate12076  (.A(g22548), .Z(II29942) ) ;
INV     gate12077  (.A(g22583), .Z(II29945) ) ;
INV     gate12078  (.A(g22549), .Z(II29948) ) ;
INV     gate12079  (.A(g22584), .Z(II29951) ) ;
INV     gate12080  (.A(g22611), .Z(II29954) ) ;
INV     gate12081  (.A(g22585), .Z(II29957) ) ;
INV     gate12082  (.A(g22612), .Z(II29960) ) ;
INV     gate12083  (.A(g22639), .Z(II29963) ) ;
INV     gate12084  (.A(g22613), .Z(II29966) ) ;
INV     gate12085  (.A(g22640), .Z(II29969) ) ;
INV     gate12086  (.A(g22669), .Z(II29972) ) ;
INV     gate12087  (.A(g22641), .Z(II29975) ) ;
INV     gate12088  (.A(g22670), .Z(II29978) ) ;
INV     gate12089  (.A(g22702), .Z(II29981) ) ;
INV     gate12090  (.A(g22671), .Z(II29984) ) ;
INV     gate12091  (.A(g22703), .Z(II29987) ) ;
INV     gate12092  (.A(g22728), .Z(II29990) ) ;
INV     gate12093  (.A(g22704), .Z(II29993) ) ;
INV     gate12094  (.A(g22729), .Z(II29996) ) ;
INV     gate12095  (.A(g22756), .Z(II29999) ) ;
INV     gate12096  (.A(g22730), .Z(II30002) ) ;
INV     gate12097  (.A(g22757), .Z(II30005) ) ;
INV     gate12098  (.A(g22785), .Z(II30008) ) ;
INV     gate12099  (.A(g22758), .Z(II30011) ) ;
INV     gate12100  (.A(g22786), .Z(II30014) ) ;
INV     gate12101  (.A(g22824), .Z(II30017) ) ;
INV     gate12102  (.A(g22519), .Z(II30020) ) ;
INV     gate12103  (.A(g22550), .Z(II30023) ) ;
INV     gate12104  (.A(g22586), .Z(II30026) ) ;
INV     gate12105  (.A(g22642), .Z(II30029) ) ;
INV     gate12106  (.A(g22672), .Z(II30032) ) ;
INV     gate12107  (.A(g22705), .Z(II30035) ) ;
INV     gate12108  (.A(g22673), .Z(II30038) ) ;
INV     gate12109  (.A(g22706), .Z(II30041) ) ;
INV     gate12110  (.A(g22731), .Z(II30044) ) ;
INV     gate12111  (.A(g22107), .Z(II30047) ) ;
INV     gate12112  (.A(g22619), .Z(II30050) ) ;
INV     gate12113  (.A(g22558), .Z(II30053) ) ;
INV     gate12114  (.A(g22589), .Z(II30056) ) ;
INV     gate12115  (.A(g22620), .Z(II30059) ) ;
INV     gate12116  (.A(g22590), .Z(II30062) ) ;
INV     gate12117  (.A(g22621), .Z(II30065) ) ;
INV     gate12118  (.A(g22647), .Z(II30068) ) ;
INV     gate12119  (.A(g22622), .Z(II30071) ) ;
INV     gate12120  (.A(g22648), .Z(II30074) ) ;
INV     gate12121  (.A(g22675), .Z(II30077) ) ;
INV     gate12122  (.A(g22649), .Z(II30080) ) ;
INV     gate12123  (.A(g22676), .Z(II30083) ) ;
INV     gate12124  (.A(g22709), .Z(II30086) ) ;
INV     gate12125  (.A(g22677), .Z(II30089) ) ;
INV     gate12126  (.A(g22710), .Z(II30092) ) ;
INV     gate12127  (.A(g22733), .Z(II30095) ) ;
INV     gate12128  (.A(g22711), .Z(II30098) ) ;
INV     gate12129  (.A(g22734), .Z(II30101) ) ;
INV     gate12130  (.A(g22760), .Z(II30104) ) ;
INV     gate12131  (.A(g22735), .Z(II30107) ) ;
INV     gate12132  (.A(g22761), .Z(II30110) ) ;
INV     gate12133  (.A(g22790), .Z(II30113) ) ;
INV     gate12134  (.A(g22762), .Z(II30116) ) ;
INV     gate12135  (.A(g22791), .Z(II30119) ) ;
INV     gate12136  (.A(g22827), .Z(II30122) ) ;
INV     gate12137  (.A(g22792), .Z(II30125) ) ;
INV     gate12138  (.A(g22828), .Z(II30128) ) ;
INV     gate12139  (.A(g22864), .Z(II30131) ) ;
INV     gate12140  (.A(g22559), .Z(II30134) ) ;
INV     gate12141  (.A(g22591), .Z(II30137) ) ;
INV     gate12142  (.A(g22623), .Z(II30140) ) ;
INV     gate12143  (.A(g22678), .Z(II30143) ) ;
INV     gate12144  (.A(g22712), .Z(II30146) ) ;
INV     gate12145  (.A(g22736), .Z(II30149) ) ;
INV     gate12146  (.A(g22713), .Z(II30152) ) ;
INV     gate12147  (.A(g22737), .Z(II30155) ) ;
INV     gate12148  (.A(g22763), .Z(II30158) ) ;
INV     gate12149  (.A(g22133), .Z(II30161) ) ;
INV     gate12150  (.A(g22655), .Z(II30164) ) ;
INV     gate12151  (.A(g22598), .Z(II30167) ) ;
INV     gate12152  (.A(g22626), .Z(II30170) ) ;
INV     gate12153  (.A(g22656), .Z(II30173) ) ;
INV     gate12154  (.A(g22627), .Z(II30176) ) ;
INV     gate12155  (.A(g22657), .Z(II30179) ) ;
INV     gate12156  (.A(g22683), .Z(II30182) ) ;
INV     gate12157  (.A(g22658), .Z(II30185) ) ;
INV     gate12158  (.A(g22684), .Z(II30188) ) ;
INV     gate12159  (.A(g22715), .Z(II30191) ) ;
INV     gate12160  (.A(g22685), .Z(II30194) ) ;
INV     gate12161  (.A(g22716), .Z(II30197) ) ;
INV     gate12162  (.A(g22740), .Z(II30200) ) ;
INV     gate12163  (.A(g22717), .Z(II30203) ) ;
INV     gate12164  (.A(g22741), .Z(II30206) ) ;
INV     gate12165  (.A(g22765), .Z(II30209) ) ;
INV     gate12166  (.A(g22742), .Z(II30212) ) ;
INV     gate12167  (.A(g22766), .Z(II30215) ) ;
INV     gate12168  (.A(g22794), .Z(II30218) ) ;
INV     gate12169  (.A(g22767), .Z(II30221) ) ;
INV     gate12170  (.A(g22795), .Z(II30224) ) ;
INV     gate12171  (.A(g22832), .Z(II30227) ) ;
INV     gate12172  (.A(g22796), .Z(II30230) ) ;
INV     gate12173  (.A(g22833), .Z(II30233) ) ;
INV     gate12174  (.A(g22866), .Z(II30236) ) ;
INV     gate12175  (.A(g22834), .Z(II30239) ) ;
INV     gate12176  (.A(g22867), .Z(II30242) ) ;
INV     gate12177  (.A(g22899), .Z(II30245) ) ;
INV     gate12178  (.A(g22599), .Z(II30248) ) ;
INV     gate12179  (.A(g22628), .Z(II30251) ) ;
INV     gate12180  (.A(g22659), .Z(II30254) ) ;
INV     gate12181  (.A(g22718), .Z(II30257) ) ;
INV     gate12182  (.A(g22743), .Z(II30260) ) ;
INV     gate12183  (.A(g22768), .Z(II30263) ) ;
INV     gate12184  (.A(g22744), .Z(II30266) ) ;
INV     gate12185  (.A(g22769), .Z(II30269) ) ;
INV     gate12186  (.A(g22797), .Z(II30272) ) ;
INV     gate12187  (.A(g22156), .Z(II30275) ) ;
INV     gate12188  (.A(g22691), .Z(II30278) ) ;
INV     gate12189  (.A(g22635), .Z(II30281) ) ;
INV     gate12190  (.A(g22662), .Z(II30284) ) ;
INV     gate12191  (.A(g22692), .Z(II30287) ) ;
INV     gate12192  (.A(g22663), .Z(II30290) ) ;
INV     gate12193  (.A(g22693), .Z(II30293) ) ;
INV     gate12194  (.A(g22723), .Z(II30296) ) ;
INV     gate12195  (.A(g22694), .Z(II30299) ) ;
INV     gate12196  (.A(g22724), .Z(II30302) ) ;
INV     gate12197  (.A(g22746), .Z(II30305) ) ;
INV     gate12198  (.A(g22725), .Z(II30308) ) ;
INV     gate12199  (.A(g22747), .Z(II30311) ) ;
INV     gate12200  (.A(g22772), .Z(II30314) ) ;
INV     gate12201  (.A(g22748), .Z(II30317) ) ;
INV     gate12202  (.A(g22773), .Z(II30320) ) ;
INV     gate12203  (.A(g22799), .Z(II30323) ) ;
INV     gate12204  (.A(g22774), .Z(II30326) ) ;
INV     gate12205  (.A(g22800), .Z(II30329) ) ;
INV     gate12206  (.A(g22836), .Z(II30332) ) ;
INV     gate12207  (.A(g22801), .Z(II30335) ) ;
INV     gate12208  (.A(g22837), .Z(II30338) ) ;
INV     gate12209  (.A(g22871), .Z(II30341) ) ;
INV     gate12210  (.A(g22838), .Z(II30344) ) ;
INV     gate12211  (.A(g22872), .Z(II30347) ) ;
INV     gate12212  (.A(g22901), .Z(II30350) ) ;
INV     gate12213  (.A(g22873), .Z(II30353) ) ;
INV     gate12214  (.A(g22902), .Z(II30356) ) ;
INV     gate12215  (.A(g22934), .Z(II30359) ) ;
INV     gate12216  (.A(g22636), .Z(II30362) ) ;
INV     gate12217  (.A(g22664), .Z(II30365) ) ;
INV     gate12218  (.A(g22695), .Z(II30368) ) ;
INV     gate12219  (.A(g22749), .Z(II30371) ) ;
INV     gate12220  (.A(g22775), .Z(II30374) ) ;
INV     gate12221  (.A(g22802), .Z(II30377) ) ;
INV     gate12222  (.A(g22776), .Z(II30380) ) ;
INV     gate12223  (.A(g22803), .Z(II30383) ) ;
INV     gate12224  (.A(g22839), .Z(II30386) ) ;
INV     gate12225  (.A(g22225), .Z(II30389) ) ;
INV     gate12226  (.A(g22226), .Z(II30392) ) ;
INV     gate12227  (.A(g22253), .Z(II30395) ) ;
INV     gate12228  (.A(g22840), .Z(II30398) ) ;
INV     gate12229  (.A(g22444), .Z(II30401) ) ;
INV     gate12230  (.A(g22948), .Z(II30404) ) ;
INV     gate12231  (.A(g22970), .Z(II30407) ) ;
OR3     gate12232  (.A(g21800), .B(g21788), .C(g21844), .Z(g23052) ) ;
INV     gate12233  (.A(g23052), .Z(g23403) ) ;
OR3     gate12234  (.A(g21808), .B(g21802), .C(g21846), .Z(g23071) ) ;
INV     gate12235  (.A(g23071), .Z(g23410) ) ;
OR3     gate12236  (.A(g21815), .B(g21810), .C(g21849), .Z(g23084) ) ;
INV     gate12237  (.A(g23084), .Z(g23415) ) ;
OR2     gate12238  (.A(g21806), .B(g21799), .Z(g23089) ) ;
INV     gate12239  (.A(g23089), .Z(g23420) ) ;
OR3     gate12240  (.A(g21821), .B(g21817), .C(g21856), .Z(g23100) ) ;
INV     gate12241  (.A(g23100), .Z(g23424) ) ;
OR2     gate12242  (.A(g21813), .B(g21807), .Z(g23107) ) ;
INV     gate12243  (.A(g23107), .Z(g23429) ) ;
OR2     gate12244  (.A(g21819), .B(g21814), .Z(g23120) ) ;
INV     gate12245  (.A(g23120), .Z(g23435) ) ;
NOR2    gate12246  (.A(g16909), .B(g21067), .Z(g23000) ) ;
INV     gate12247  (.A(g23000), .Z(II30467) ) ;
INV     gate12248  (.A(II30467), .Z(g23438) ) ;
NOR2    gate12249  (.A(g17117), .B(g21188), .Z(g23117) ) ;
INV     gate12250  (.A(g23117), .Z(II30470) ) ;
INV     gate12251  (.A(II30470), .Z(g23439) ) ;
OR2     gate12252  (.A(g21823), .B(g21820), .Z(g23129) ) ;
INV     gate12253  (.A(g23129), .Z(g23441) ) ;
INV     gate12254  (.A(g22945), .Z(g23444) ) ;
NAND2   gate12255  (.A(g21238), .B(g83), .Z(g22876) ) ;
INV     gate12256  (.A(g22876), .Z(II30476) ) ;
INV     gate12257  (.A(II30476), .Z(g23448) ) ;
NOR2    gate12258  (.A(g16939), .B(g21077), .Z(g23014) ) ;
INV     gate12259  (.A(g23014), .Z(II30480) ) ;
INV     gate12260  (.A(II30480), .Z(g23452) ) ;
NOR2    gate12261  (.A(g17144), .B(g21203), .Z(g23126) ) ;
INV     gate12262  (.A(g23126), .Z(II30483) ) ;
INV     gate12263  (.A(II30483), .Z(g23453) ) ;
NOR2    gate12264  (.A(g16968), .B(g21086), .Z(g23022) ) ;
INV     gate12265  (.A(g23022), .Z(II30486) ) ;
INV     gate12266  (.A(II30486), .Z(g23454) ) ;
NAND2   gate12267  (.A(g21246), .B(g771), .Z(g22911) ) ;
INV     gate12268  (.A(g22911), .Z(II30489) ) ;
INV     gate12269  (.A(II30489), .Z(g23455) ) ;
NOR2    gate12270  (.A(g16970), .B(g21091), .Z(g23030) ) ;
INV     gate12271  (.A(g23030), .Z(II30493) ) ;
INV     gate12272  (.A(II30493), .Z(g23459) ) ;
NOR2    gate12273  (.A(g17167), .B(g21218), .Z(g23137) ) ;
INV     gate12274  (.A(g23137), .Z(II30496) ) ;
INV     gate12275  (.A(II30496), .Z(g23460) ) ;
NOR2    gate12276  (.A(g16989), .B(g21098), .Z(g23039) ) ;
INV     gate12277  (.A(g23039), .Z(II30501) ) ;
INV     gate12278  (.A(II30501), .Z(g23463) ) ;
NAND2   gate12279  (.A(g21255), .B(g1457), .Z(g22936) ) ;
INV     gate12280  (.A(g22936), .Z(II30504) ) ;
INV     gate12281  (.A(II30504), .Z(g23464) ) ;
NOR2    gate12282  (.A(g16991), .B(g21103), .Z(g23047) ) ;
INV     gate12283  (.A(g23047), .Z(II30508) ) ;
INV     gate12284  (.A(II30508), .Z(g23468) ) ;
NOR2    gate12285  (.A(g17182), .B(g21226), .Z(g21970) ) ;
INV     gate12286  (.A(g21970), .Z(II30511) ) ;
INV     gate12287  (.A(II30511), .Z(g23469) ) ;
NAND2   gate12288  (.A(II28727), .B(II28728), .Z(g22188) ) ;
INV     gate12289  (.A(g22188), .Z(g23470) ) ;
NOR2    gate12290  (.A(g16999), .B(g21112), .Z(g23058) ) ;
INV     gate12291  (.A(g23058), .Z(II30516) ) ;
INV     gate12292  (.A(II30516), .Z(g23472) ) ;
NAND2   gate12293  (.A(g21263), .B(g2151), .Z(g22942) ) ;
INV     gate12294  (.A(g22942), .Z(II30519) ) ;
INV     gate12295  (.A(II30519), .Z(g23473) ) ;
NOR2    gate12296  (.A(g17015), .B(g21122), .Z(g23067) ) ;
INV     gate12297  (.A(g23067), .Z(II30525) ) ;
INV     gate12298  (.A(II30525), .Z(g23481) ) ;
NAND2   gate12299  (.A(II28742), .B(II28743), .Z(g22197) ) ;
INV     gate12300  (.A(g22197), .Z(g23482) ) ;
NOR2    gate12301  (.A(g17023), .B(g21129), .Z(g23076) ) ;
INV     gate12302  (.A(g23076), .Z(II30531) ) ;
INV     gate12303  (.A(II30531), .Z(g23485) ) ;
NOR2    gate12304  (.A(g17045), .B(g21141), .Z(g23081) ) ;
INV     gate12305  (.A(g23081), .Z(II30536) ) ;
INV     gate12306  (.A(II30536), .Z(g23492) ) ;
NAND2   gate12307  (.A(II28754), .B(II28755), .Z(g22203) ) ;
INV     gate12308  (.A(g22203), .Z(g23493) ) ;
NOR2    gate12309  (.A(g17055), .B(g21154), .Z(g23092) ) ;
INV     gate12310  (.A(g23092), .Z(II30544) ) ;
INV     gate12311  (.A(II30544), .Z(g23500) ) ;
NOR2    gate12312  (.A(g17056), .B(g21155), .Z(g23093) ) ;
INV     gate12313  (.A(g23093), .Z(II30547) ) ;
INV     gate12314  (.A(II30547), .Z(g23501) ) ;
NOR2    gate12315  (.A(g17079), .B(g21161), .Z(g23097) ) ;
INV     gate12316  (.A(g23097), .Z(II30552) ) ;
INV     gate12317  (.A(II30552), .Z(g23508) ) ;
NAND2   gate12318  (.A(II28766), .B(II28767), .Z(g22209) ) ;
INV     gate12319  (.A(g22209), .Z(g23509) ) ;
NOR2    gate12320  (.A(g17090), .B(g21174), .Z(g23110) ) ;
INV     gate12321  (.A(g23110), .Z(II30560) ) ;
INV     gate12322  (.A(II30560), .Z(g23516) ) ;
NOR2    gate12323  (.A(g17091), .B(g21175), .Z(g23111) ) ;
INV     gate12324  (.A(g23111), .Z(II30563) ) ;
INV     gate12325  (.A(II30563), .Z(g23517) ) ;
NOR2    gate12326  (.A(g17114), .B(g21181), .Z(g23114) ) ;
INV     gate12327  (.A(g23114), .Z(II30568) ) ;
INV     gate12328  (.A(II30568), .Z(g23524) ) ;
NOR2    gate12329  (.A(g17128), .B(g21194), .Z(g23123) ) ;
INV     gate12330  (.A(g23123), .Z(II30575) ) ;
INV     gate12331  (.A(II30575), .Z(g23531) ) ;
NOR2    gate12332  (.A(g17129), .B(g21195), .Z(g23124) ) ;
INV     gate12333  (.A(g23124), .Z(II30578) ) ;
INV     gate12334  (.A(II30578), .Z(g23532) ) ;
NOR2    gate12335  (.A(g17155), .B(g21209), .Z(g23132) ) ;
INV     gate12336  (.A(g23132), .Z(II30586) ) ;
INV     gate12337  (.A(II30586), .Z(g23542) ) ;
NOR2    gate12338  (.A(g17156), .B(g21210), .Z(g23133) ) ;
INV     gate12339  (.A(g23133), .Z(II30589) ) ;
INV     gate12340  (.A(II30589), .Z(g23543) ) ;
NOR2    gate12341  (.A(g21284), .B(g19549), .Z(g22025) ) ;
INV     gate12342  (.A(g22025), .Z(II30594) ) ;
INV     gate12343  (.A(II30594), .Z(g23546) ) ;
NOR2    gate12344  (.A(g21290), .B(g19553), .Z(g22027) ) ;
INV     gate12345  (.A(g22027), .Z(II30598) ) ;
INV     gate12346  (.A(II30598), .Z(g23548) ) ;
NOR2    gate12347  (.A(g21291), .B(g19554), .Z(g22028) ) ;
INV     gate12348  (.A(g22028), .Z(II30601) ) ;
INV     gate12349  (.A(II30601), .Z(g23549) ) ;
NOR2    gate12350  (.A(g21292), .B(g19555), .Z(g22029) ) ;
INV     gate12351  (.A(g22029), .Z(II30607) ) ;
INV     gate12352  (.A(II30607), .Z(g23553) ) ;
NOR2    gate12353  (.A(g21298), .B(g19557), .Z(g22030) ) ;
INV     gate12354  (.A(g22030), .Z(II30611) ) ;
INV     gate12355  (.A(II30611), .Z(g23555) ) ;
NOR2    gate12356  (.A(g21299), .B(g19558), .Z(g22031) ) ;
INV     gate12357  (.A(g22031), .Z(II30614) ) ;
INV     gate12358  (.A(II30614), .Z(g23556) ) ;
NOR2    gate12359  (.A(g21300), .B(g19559), .Z(g22032) ) ;
INV     gate12360  (.A(g22032), .Z(II30617) ) ;
INV     gate12361  (.A(II30617), .Z(g23557) ) ;
NOR2    gate12362  (.A(g21301), .B(g19560), .Z(g22033) ) ;
INV     gate12363  (.A(g22033), .Z(II30623) ) ;
INV     gate12364  (.A(II30623), .Z(g23561) ) ;
NOR2    gate12365  (.A(g21302), .B(g19561), .Z(g22034) ) ;
INV     gate12366  (.A(g22034), .Z(II30626) ) ;
INV     gate12367  (.A(II30626), .Z(g23562) ) ;
NOR2    gate12368  (.A(g21303), .B(g19562), .Z(g22035) ) ;
INV     gate12369  (.A(g22035), .Z(II30632) ) ;
INV     gate12370  (.A(II30632), .Z(g23566) ) ;
NOR2    gate12371  (.A(g21304), .B(g19564), .Z(g22037) ) ;
INV     gate12372  (.A(g22037), .Z(II30636) ) ;
INV     gate12373  (.A(II30636), .Z(g23568) ) ;
NOR2    gate12374  (.A(g21305), .B(g19565), .Z(g22038) ) ;
INV     gate12375  (.A(g22038), .Z(II30639) ) ;
INV     gate12376  (.A(II30639), .Z(g23569) ) ;
NOR2    gate12377  (.A(g21306), .B(g19566), .Z(g22039) ) ;
INV     gate12378  (.A(g22039), .Z(II30642) ) ;
INV     gate12379  (.A(II30642), .Z(g23570) ) ;
NOR2    gate12380  (.A(g21307), .B(g19567), .Z(g22040) ) ;
INV     gate12381  (.A(g22040), .Z(II30648) ) ;
INV     gate12382  (.A(II30648), .Z(g23574) ) ;
NOR2    gate12383  (.A(g21308), .B(g19568), .Z(g22041) ) ;
INV     gate12384  (.A(g22041), .Z(II30651) ) ;
INV     gate12385  (.A(II30651), .Z(g23575) ) ;
NOR2    gate12386  (.A(g21309), .B(g19569), .Z(g22042) ) ;
INV     gate12387  (.A(g22042), .Z(II30654) ) ;
INV     gate12388  (.A(II30654), .Z(g23576) ) ;
NOR2    gate12389  (.A(g21310), .B(g19570), .Z(g22043) ) ;
INV     gate12390  (.A(g22043), .Z(II30660) ) ;
INV     gate12391  (.A(II30660), .Z(g23580) ) ;
NOR2    gate12392  (.A(g21311), .B(g19571), .Z(g22044) ) ;
INV     gate12393  (.A(g22044), .Z(II30663) ) ;
INV     gate12394  (.A(II30663), .Z(g23581) ) ;
NOR2    gate12395  (.A(g21312), .B(g19572), .Z(g22045) ) ;
INV     gate12396  (.A(g22045), .Z(II30669) ) ;
INV     gate12397  (.A(II30669), .Z(g23585) ) ;
NOR2    gate12398  (.A(g21313), .B(g19574), .Z(g22047) ) ;
INV     gate12399  (.A(g22047), .Z(II30673) ) ;
INV     gate12400  (.A(II30673), .Z(g23587) ) ;
NOR2    gate12401  (.A(g21314), .B(g19575), .Z(g22048) ) ;
INV     gate12402  (.A(g22048), .Z(II30676) ) ;
INV     gate12403  (.A(II30676), .Z(g23588) ) ;
NOR2    gate12404  (.A(g21315), .B(g19576), .Z(g22049) ) ;
INV     gate12405  (.A(g22049), .Z(II30679) ) ;
INV     gate12406  (.A(II30679), .Z(g23589) ) ;
NOR2    gate12407  (.A(g20878), .B(g10024), .Z(g23136) ) ;
INV     gate12408  (.A(g23136), .Z(II30686) ) ;
INV     gate12409  (.A(II30686), .Z(g23594) ) ;
NOR2    gate12410  (.A(g21319), .B(g19586), .Z(g22054) ) ;
INV     gate12411  (.A(g22054), .Z(II30689) ) ;
INV     gate12412  (.A(II30689), .Z(g23595) ) ;
NOR2    gate12413  (.A(g21320), .B(g19587), .Z(g22055) ) ;
INV     gate12414  (.A(g22055), .Z(II30692) ) ;
INV     gate12415  (.A(II30692), .Z(g23596) ) ;
NOR2    gate12416  (.A(g21321), .B(g19588), .Z(g22056) ) ;
INV     gate12417  (.A(g22056), .Z(II30695) ) ;
INV     gate12418  (.A(II30695), .Z(g23597) ) ;
NOR2    gate12419  (.A(g21322), .B(g19589), .Z(g22057) ) ;
INV     gate12420  (.A(g22057), .Z(II30701) ) ;
INV     gate12421  (.A(II30701), .Z(g23601) ) ;
NOR2    gate12422  (.A(g21323), .B(g19590), .Z(g22058) ) ;
INV     gate12423  (.A(g22058), .Z(II30704) ) ;
INV     gate12424  (.A(II30704), .Z(g23602) ) ;
NOR2    gate12425  (.A(g21324), .B(g19591), .Z(g22059) ) ;
INV     gate12426  (.A(g22059), .Z(II30707) ) ;
INV     gate12427  (.A(II30707), .Z(g23603) ) ;
NOR2    gate12428  (.A(g21325), .B(g19592), .Z(g22060) ) ;
INV     gate12429  (.A(g22060), .Z(II30713) ) ;
INV     gate12430  (.A(II30713), .Z(g23607) ) ;
NOR2    gate12431  (.A(g21326), .B(g19593), .Z(g22061) ) ;
INV     gate12432  (.A(g22061), .Z(II30716) ) ;
INV     gate12433  (.A(II30716), .Z(g23608) ) ;
NOR2    gate12434  (.A(g21328), .B(g19597), .Z(g22063) ) ;
INV     gate12435  (.A(g22063), .Z(II30722) ) ;
INV     gate12436  (.A(II30722), .Z(g23612) ) ;
NOR2    gate12437  (.A(g21329), .B(g19598), .Z(g22064) ) ;
INV     gate12438  (.A(g22064), .Z(II30725) ) ;
INV     gate12439  (.A(II30725), .Z(g23613) ) ;
NOR2    gate12440  (.A(g21330), .B(g19599), .Z(g22065) ) ;
INV     gate12441  (.A(g22065), .Z(II30728) ) ;
INV     gate12442  (.A(II30728), .Z(g23614) ) ;
NOR2    gate12443  (.A(g21334), .B(g19604), .Z(g22066) ) ;
INV     gate12444  (.A(g22066), .Z(II30735) ) ;
INV     gate12445  (.A(II30735), .Z(g23619) ) ;
NOR2    gate12446  (.A(g21335), .B(g19605), .Z(g22067) ) ;
INV     gate12447  (.A(g22067), .Z(II30738) ) ;
INV     gate12448  (.A(II30738), .Z(g23620) ) ;
NOR2    gate12449  (.A(g21336), .B(g19606), .Z(g22068) ) ;
INV     gate12450  (.A(g22068), .Z(II30741) ) ;
INV     gate12451  (.A(II30741), .Z(g23621) ) ;
NOR2    gate12452  (.A(g20895), .B(g10133), .Z(g21969) ) ;
INV     gate12453  (.A(g21969), .Z(II30748) ) ;
INV     gate12454  (.A(II30748), .Z(g23626) ) ;
NOR2    gate12455  (.A(g21337), .B(g19616), .Z(g22073) ) ;
INV     gate12456  (.A(g22073), .Z(II30751) ) ;
INV     gate12457  (.A(II30751), .Z(g23627) ) ;
NOR2    gate12458  (.A(g21338), .B(g19617), .Z(g22074) ) ;
INV     gate12459  (.A(g22074), .Z(II30754) ) ;
INV     gate12460  (.A(II30754), .Z(g23628) ) ;
NOR2    gate12461  (.A(g21339), .B(g19618), .Z(g22075) ) ;
INV     gate12462  (.A(g22075), .Z(II30757) ) ;
INV     gate12463  (.A(II30757), .Z(g23629) ) ;
NOR2    gate12464  (.A(g21340), .B(g19619), .Z(g22076) ) ;
INV     gate12465  (.A(g22076), .Z(II30763) ) ;
INV     gate12466  (.A(II30763), .Z(g23633) ) ;
NOR2    gate12467  (.A(g21341), .B(g19620), .Z(g22077) ) ;
INV     gate12468  (.A(g22077), .Z(II30766) ) ;
INV     gate12469  (.A(II30766), .Z(g23634) ) ;
NOR2    gate12470  (.A(g21342), .B(g19621), .Z(g22078) ) ;
INV     gate12471  (.A(g22078), .Z(II30769) ) ;
INV     gate12472  (.A(II30769), .Z(g23635) ) ;
NOR2    gate12473  (.A(g21343), .B(g19623), .Z(g22079) ) ;
INV     gate12474  (.A(g22079), .Z(II30776) ) ;
INV     gate12475  (.A(II30776), .Z(g23640) ) ;
NOR2    gate12476  (.A(g21344), .B(g19624), .Z(g22080) ) ;
INV     gate12477  (.A(g22080), .Z(II30779) ) ;
INV     gate12478  (.A(II30779), .Z(g23641) ) ;
NOR2    gate12479  (.A(g21345), .B(g19625), .Z(g22081) ) ;
INV     gate12480  (.A(g22081), .Z(II30782) ) ;
INV     gate12481  (.A(II30782), .Z(g23642) ) ;
NOR2    gate12482  (.A(g17012), .B(g21891), .Z(g22454) ) ;
INV     gate12483  (.A(g22454), .Z(II30786) ) ;
INV     gate12484  (.A(II30786), .Z(g23644) ) ;
NOR2    gate12485  (.A(g21349), .B(g19630), .Z(g22087) ) ;
INV     gate12486  (.A(g22087), .Z(II30797) ) ;
INV     gate12487  (.A(II30797), .Z(g23661) ) ;
NOR2    gate12488  (.A(g21350), .B(g19631), .Z(g22088) ) ;
INV     gate12489  (.A(g22088), .Z(II30800) ) ;
INV     gate12490  (.A(II30800), .Z(g23662) ) ;
NOR2    gate12491  (.A(g21351), .B(g19632), .Z(g22089) ) ;
INV     gate12492  (.A(g22089), .Z(II30803) ) ;
INV     gate12493  (.A(II30803), .Z(g23663) ) ;
NOR2    gate12494  (.A(g21352), .B(g19637), .Z(g22090) ) ;
INV     gate12495  (.A(g22090), .Z(II30810) ) ;
INV     gate12496  (.A(II30810), .Z(g23668) ) ;
NOR2    gate12497  (.A(g21353), .B(g19638), .Z(g22091) ) ;
INV     gate12498  (.A(g22091), .Z(II30813) ) ;
INV     gate12499  (.A(II30813), .Z(g23669) ) ;
NOR2    gate12500  (.A(g21354), .B(g19639), .Z(g22092) ) ;
INV     gate12501  (.A(g22092), .Z(II30816) ) ;
INV     gate12502  (.A(II30816), .Z(g23670) ) ;
NOR2    gate12503  (.A(g20914), .B(g10238), .Z(g21972) ) ;
INV     gate12504  (.A(g21972), .Z(II30823) ) ;
INV     gate12505  (.A(II30823), .Z(g23675) ) ;
NOR2    gate12506  (.A(g21355), .B(g19649), .Z(g22097) ) ;
INV     gate12507  (.A(g22097), .Z(II30826) ) ;
INV     gate12508  (.A(II30826), .Z(g23676) ) ;
NOR2    gate12509  (.A(g21356), .B(g19650), .Z(g22098) ) ;
INV     gate12510  (.A(g22098), .Z(II30829) ) ;
INV     gate12511  (.A(II30829), .Z(g23677) ) ;
NOR2    gate12512  (.A(g21357), .B(g19651), .Z(g22099) ) ;
INV     gate12513  (.A(g22099), .Z(II30832) ) ;
INV     gate12514  (.A(II30832), .Z(g23678) ) ;
NOR2    gate12515  (.A(g21360), .B(g19653), .Z(g22100) ) ;
INV     gate12516  (.A(g22100), .Z(II30838) ) ;
INV     gate12517  (.A(II30838), .Z(g23682) ) ;
NOR2    gate12518  (.A(g21361), .B(g19654), .Z(g22101) ) ;
INV     gate12519  (.A(g22101), .Z(II30841) ) ;
INV     gate12520  (.A(II30841), .Z(g23683) ) ;
NOR2    gate12521  (.A(g21362), .B(g19655), .Z(g22102) ) ;
INV     gate12522  (.A(g22102), .Z(II30844) ) ;
INV     gate12523  (.A(II30844), .Z(g23684) ) ;
NOR2    gate12524  (.A(g21363), .B(g19656), .Z(g22103) ) ;
INV     gate12525  (.A(g22103), .Z(II30847) ) ;
INV     gate12526  (.A(II30847), .Z(g23685) ) ;
NOR2    gate12527  (.A(g21367), .B(g19663), .Z(g22104) ) ;
INV     gate12528  (.A(g22104), .Z(II30854) ) ;
INV     gate12529  (.A(II30854), .Z(g23690) ) ;
NOR2    gate12530  (.A(g21368), .B(g19664), .Z(g22105) ) ;
INV     gate12531  (.A(g22105), .Z(II30857) ) ;
INV     gate12532  (.A(II30857), .Z(g23691) ) ;
NOR2    gate12533  (.A(g21369), .B(g19665), .Z(g22106) ) ;
INV     gate12534  (.A(g22106), .Z(II30860) ) ;
INV     gate12535  (.A(II30860), .Z(g23692) ) ;
NOR2    gate12536  (.A(g17042), .B(g21899), .Z(g22493) ) ;
INV     gate12537  (.A(g22493), .Z(II30864) ) ;
INV     gate12538  (.A(II30864), .Z(g23694) ) ;
NOR2    gate12539  (.A(g21370), .B(g19670), .Z(g22112) ) ;
INV     gate12540  (.A(g22112), .Z(II30875) ) ;
INV     gate12541  (.A(II30875), .Z(g23711) ) ;
NOR2    gate12542  (.A(g21371), .B(g19671), .Z(g22113) ) ;
INV     gate12543  (.A(g22113), .Z(II30878) ) ;
INV     gate12544  (.A(II30878), .Z(g23712) ) ;
NOR2    gate12545  (.A(g21372), .B(g19672), .Z(g22114) ) ;
INV     gate12546  (.A(g22114), .Z(II30881) ) ;
INV     gate12547  (.A(II30881), .Z(g23713) ) ;
NOR2    gate12548  (.A(g21373), .B(g19677), .Z(g22115) ) ;
INV     gate12549  (.A(g22115), .Z(II30888) ) ;
INV     gate12550  (.A(II30888), .Z(g23718) ) ;
NOR2    gate12551  (.A(g21374), .B(g19678), .Z(g22116) ) ;
INV     gate12552  (.A(g22116), .Z(II30891) ) ;
INV     gate12553  (.A(II30891), .Z(g23719) ) ;
NOR2    gate12554  (.A(g21375), .B(g19679), .Z(g22117) ) ;
INV     gate12555  (.A(g22117), .Z(II30894) ) ;
INV     gate12556  (.A(II30894), .Z(g23720) ) ;
NOR2    gate12557  (.A(g20938), .B(g10340), .Z(g21974) ) ;
INV     gate12558  (.A(g21974), .Z(II30901) ) ;
INV     gate12559  (.A(II30901), .Z(g23725) ) ;
NOR2    gate12560  (.A(g21378), .B(g19692), .Z(g22122) ) ;
INV     gate12561  (.A(g22122), .Z(II30905) ) ;
INV     gate12562  (.A(II30905), .Z(g23727) ) ;
NOR2    gate12563  (.A(g21379), .B(g19693), .Z(g22123) ) ;
INV     gate12564  (.A(g22123), .Z(II30908) ) ;
INV     gate12565  (.A(II30908), .Z(g23728) ) ;
NOR2    gate12566  (.A(g21380), .B(g19694), .Z(g22124) ) ;
INV     gate12567  (.A(g22124), .Z(II30911) ) ;
INV     gate12568  (.A(II30911), .Z(g23729) ) ;
NOR2    gate12569  (.A(g21381), .B(g19695), .Z(g22125) ) ;
INV     gate12570  (.A(g22125), .Z(II30914) ) ;
INV     gate12571  (.A(II30914), .Z(g23730) ) ;
INV     gate12572  (.A(g22806), .Z(II30917) ) ;
INV     gate12573  (.A(II30917), .Z(g23731) ) ;
NOR2    gate12574  (.A(g21389), .B(g19701), .Z(g22126) ) ;
INV     gate12575  (.A(g22126), .Z(II30922) ) ;
INV     gate12576  (.A(II30922), .Z(g23736) ) ;
NOR2    gate12577  (.A(g21390), .B(g19702), .Z(g22127) ) ;
INV     gate12578  (.A(g22127), .Z(II30925) ) ;
INV     gate12579  (.A(II30925), .Z(g23737) ) ;
NOR2    gate12580  (.A(g21391), .B(g19703), .Z(g22128) ) ;
INV     gate12581  (.A(g22128), .Z(II30928) ) ;
INV     gate12582  (.A(II30928), .Z(g23738) ) ;
NOR2    gate12583  (.A(g21392), .B(g19704), .Z(g22129) ) ;
INV     gate12584  (.A(g22129), .Z(II30931) ) ;
INV     gate12585  (.A(II30931), .Z(g23739) ) ;
NOR2    gate12586  (.A(g21393), .B(g19711), .Z(g22130) ) ;
INV     gate12587  (.A(g22130), .Z(II30938) ) ;
INV     gate12588  (.A(II30938), .Z(g23744) ) ;
NOR2    gate12589  (.A(g21394), .B(g19712), .Z(g22131) ) ;
INV     gate12590  (.A(g22131), .Z(II30941) ) ;
INV     gate12591  (.A(II30941), .Z(g23745) ) ;
NOR2    gate12592  (.A(g21395), .B(g19713), .Z(g22132) ) ;
INV     gate12593  (.A(g22132), .Z(II30944) ) ;
INV     gate12594  (.A(II30944), .Z(g23746) ) ;
NOR2    gate12595  (.A(g17076), .B(g21911), .Z(g22536) ) ;
INV     gate12596  (.A(g22536), .Z(II30948) ) ;
INV     gate12597  (.A(II30948), .Z(g23748) ) ;
NOR2    gate12598  (.A(g21396), .B(g19718), .Z(g22138) ) ;
INV     gate12599  (.A(g22138), .Z(II30959) ) ;
INV     gate12600  (.A(II30959), .Z(g23765) ) ;
NOR2    gate12601  (.A(g21397), .B(g19719), .Z(g22139) ) ;
INV     gate12602  (.A(g22139), .Z(II30962) ) ;
INV     gate12603  (.A(II30962), .Z(g23766) ) ;
NOR2    gate12604  (.A(g21398), .B(g19720), .Z(g22140) ) ;
INV     gate12605  (.A(g22140), .Z(II30965) ) ;
INV     gate12606  (.A(II30965), .Z(g23767) ) ;
NOR2    gate12607  (.A(g21401), .B(g19727), .Z(g22141) ) ;
INV     gate12608  (.A(g22141), .Z(II30973) ) ;
INV     gate12609  (.A(II30973), .Z(g23773) ) ;
NOR2    gate12610  (.A(g21402), .B(g19728), .Z(g22142) ) ;
INV     gate12611  (.A(g22142), .Z(II30976) ) ;
INV     gate12612  (.A(II30976), .Z(g23774) ) ;
NOR2    gate12613  (.A(g21403), .B(g19729), .Z(g22143) ) ;
INV     gate12614  (.A(g22143), .Z(II30979) ) ;
INV     gate12615  (.A(II30979), .Z(g23775) ) ;
NAND2   gate12616  (.A(g21636), .B(g672), .Z(g22992) ) ;
INV     gate12617  (.A(g22992), .Z(II30985) ) ;
INV     gate12618  (.A(II30985), .Z(g23779) ) ;
NOR2    gate12619  (.A(g21411), .B(g19736), .Z(g22145) ) ;
INV     gate12620  (.A(g22145), .Z(II30988) ) ;
INV     gate12621  (.A(II30988), .Z(g23782) ) ;
NOR2    gate12622  (.A(g21412), .B(g19737), .Z(g22146) ) ;
INV     gate12623  (.A(g22146), .Z(II30991) ) ;
INV     gate12624  (.A(II30991), .Z(g23783) ) ;
NOR2    gate12625  (.A(g21413), .B(g19738), .Z(g22147) ) ;
INV     gate12626  (.A(g22147), .Z(II30994) ) ;
INV     gate12627  (.A(II30994), .Z(g23784) ) ;
NOR2    gate12628  (.A(g21414), .B(g19739), .Z(g22148) ) ;
INV     gate12629  (.A(g22148), .Z(II30997) ) ;
INV     gate12630  (.A(II30997), .Z(g23785) ) ;
INV     gate12631  (.A(g22847), .Z(II31000) ) ;
INV     gate12632  (.A(II31000), .Z(g23786) ) ;
NOR2    gate12633  (.A(g21419), .B(g19745), .Z(g22149) ) ;
INV     gate12634  (.A(g22149), .Z(II31005) ) ;
INV     gate12635  (.A(II31005), .Z(g23791) ) ;
NOR2    gate12636  (.A(g21420), .B(g19746), .Z(g22150) ) ;
INV     gate12637  (.A(g22150), .Z(II31008) ) ;
INV     gate12638  (.A(II31008), .Z(g23792) ) ;
NOR2    gate12639  (.A(g21421), .B(g19747), .Z(g22151) ) ;
INV     gate12640  (.A(g22151), .Z(II31011) ) ;
INV     gate12641  (.A(II31011), .Z(g23793) ) ;
NOR2    gate12642  (.A(g21422), .B(g19748), .Z(g22152) ) ;
INV     gate12643  (.A(g22152), .Z(II31014) ) ;
INV     gate12644  (.A(II31014), .Z(g23794) ) ;
NOR2    gate12645  (.A(g21423), .B(g19755), .Z(g22153) ) ;
INV     gate12646  (.A(g22153), .Z(II31021) ) ;
INV     gate12647  (.A(II31021), .Z(g23799) ) ;
NOR2    gate12648  (.A(g21424), .B(g19756), .Z(g22154) ) ;
INV     gate12649  (.A(g22154), .Z(II31024) ) ;
INV     gate12650  (.A(II31024), .Z(g23800) ) ;
NOR2    gate12651  (.A(g21425), .B(g19757), .Z(g22155) ) ;
INV     gate12652  (.A(g22155), .Z(II31027) ) ;
INV     gate12653  (.A(II31027), .Z(g23801) ) ;
NOR2    gate12654  (.A(g17111), .B(g21925), .Z(g22576) ) ;
INV     gate12655  (.A(g22576), .Z(II31031) ) ;
INV     gate12656  (.A(II31031), .Z(g23803) ) ;
NOR2    gate12657  (.A(g21428), .B(g19764), .Z(g22161) ) ;
INV     gate12658  (.A(g22161), .Z(II31043) ) ;
INV     gate12659  (.A(II31043), .Z(g23821) ) ;
NOR2    gate12660  (.A(g21438), .B(g19770), .Z(g22162) ) ;
INV     gate12661  (.A(g22162), .Z(II31050) ) ;
INV     gate12662  (.A(II31050), .Z(g23826) ) ;
NOR2    gate12663  (.A(g21439), .B(g19771), .Z(g22163) ) ;
INV     gate12664  (.A(g22163), .Z(II31053) ) ;
INV     gate12665  (.A(II31053), .Z(g23827) ) ;
NOR2    gate12666  (.A(g21440), .B(g19772), .Z(g22164) ) ;
INV     gate12667  (.A(g22164), .Z(II31056) ) ;
INV     gate12668  (.A(II31056), .Z(g23828) ) ;
NAND2   gate12669  (.A(g21667), .B(g1358), .Z(g23003) ) ;
INV     gate12670  (.A(g23003), .Z(II31062) ) ;
INV     gate12671  (.A(II31062), .Z(g23832) ) ;
NOR2    gate12672  (.A(g21445), .B(g19779), .Z(g22166) ) ;
INV     gate12673  (.A(g22166), .Z(II31065) ) ;
INV     gate12674  (.A(II31065), .Z(g23835) ) ;
NOR2    gate12675  (.A(g21446), .B(g19780), .Z(g22167) ) ;
INV     gate12676  (.A(g22167), .Z(II31068) ) ;
INV     gate12677  (.A(II31068), .Z(g23836) ) ;
NOR2    gate12678  (.A(g21447), .B(g19781), .Z(g22168) ) ;
INV     gate12679  (.A(g22168), .Z(II31071) ) ;
INV     gate12680  (.A(II31071), .Z(g23837) ) ;
NOR2    gate12681  (.A(g21448), .B(g19782), .Z(g22169) ) ;
INV     gate12682  (.A(g22169), .Z(II31074) ) ;
INV     gate12683  (.A(II31074), .Z(g23838) ) ;
INV     gate12684  (.A(g22882), .Z(II31077) ) ;
INV     gate12685  (.A(II31077), .Z(g23839) ) ;
NOR2    gate12686  (.A(g21453), .B(g19788), .Z(g22170) ) ;
INV     gate12687  (.A(g22170), .Z(II31082) ) ;
INV     gate12688  (.A(II31082), .Z(g23844) ) ;
NOR2    gate12689  (.A(g21454), .B(g19789), .Z(g22171) ) ;
INV     gate12690  (.A(g22171), .Z(II31085) ) ;
INV     gate12691  (.A(II31085), .Z(g23845) ) ;
NOR2    gate12692  (.A(g21455), .B(g19790), .Z(g22172) ) ;
INV     gate12693  (.A(g22172), .Z(II31088) ) ;
INV     gate12694  (.A(II31088), .Z(g23846) ) ;
NOR2    gate12695  (.A(g21456), .B(g19791), .Z(g22173) ) ;
INV     gate12696  (.A(g22173), .Z(II31091) ) ;
INV     gate12697  (.A(II31091), .Z(g23847) ) ;
INV     gate12698  (.A(g22300), .Z(g23853) ) ;
NOR2    gate12699  (.A(g21476), .B(g19806), .Z(g22177) ) ;
INV     gate12700  (.A(g22177), .Z(II31102) ) ;
INV     gate12701  (.A(II31102), .Z(g23856) ) ;
NOR2    gate12702  (.A(g21480), .B(g19812), .Z(g22178) ) ;
INV     gate12703  (.A(g22178), .Z(II31109) ) ;
INV     gate12704  (.A(II31109), .Z(g23861) ) ;
NOR2    gate12705  (.A(g21481), .B(g19813), .Z(g22179) ) ;
INV     gate12706  (.A(g22179), .Z(II31112) ) ;
INV     gate12707  (.A(II31112), .Z(g23862) ) ;
NOR2    gate12708  (.A(g21482), .B(g19814), .Z(g22180) ) ;
INV     gate12709  (.A(g22180), .Z(II31115) ) ;
INV     gate12710  (.A(II31115), .Z(g23863) ) ;
NAND2   gate12711  (.A(g21696), .B(g2052), .Z(g23017) ) ;
INV     gate12712  (.A(g23017), .Z(II31121) ) ;
INV     gate12713  (.A(II31121), .Z(g23867) ) ;
NOR2    gate12714  (.A(g21487), .B(g19821), .Z(g22182) ) ;
INV     gate12715  (.A(g22182), .Z(II31124) ) ;
INV     gate12716  (.A(II31124), .Z(g23870) ) ;
NOR2    gate12717  (.A(g21488), .B(g19822), .Z(g22183) ) ;
INV     gate12718  (.A(g22183), .Z(II31127) ) ;
INV     gate12719  (.A(II31127), .Z(g23871) ) ;
NOR2    gate12720  (.A(g21489), .B(g19823), .Z(g22184) ) ;
INV     gate12721  (.A(g22184), .Z(II31130) ) ;
INV     gate12722  (.A(II31130), .Z(g23872) ) ;
NOR2    gate12723  (.A(g21490), .B(g19824), .Z(g22185) ) ;
INV     gate12724  (.A(g22185), .Z(II31133) ) ;
INV     gate12725  (.A(II31133), .Z(g23873) ) ;
INV     gate12726  (.A(g22917), .Z(II31136) ) ;
INV     gate12727  (.A(II31136), .Z(g23874) ) ;
INV     gate12728  (.A(g22777), .Z(II31141) ) ;
INV     gate12729  (.A(II31141), .Z(g23879) ) ;
NOR2    gate12730  (.A(g21903), .B(g7466), .Z(g22935) ) ;
INV     gate12731  (.A(g22935), .Z(II31144) ) ;
INV     gate12732  (.A(II31144), .Z(g23882) ) ;
AND4    gate12733  (.A(g21135), .B(g21118), .C(g21106), .D(II28609), .Z(g22062) ) ;
INV     gate12734  (.A(g22062), .Z(g23885) ) ;
INV     gate12735  (.A(g22328), .Z(g23887) ) ;
NOR2    gate12736  (.A(g21517), .B(g19850), .Z(g22191) ) ;
INV     gate12737  (.A(g22191), .Z(II31152) ) ;
INV     gate12738  (.A(II31152), .Z(g23890) ) ;
NOR2    gate12739  (.A(g21521), .B(g19856), .Z(g22192) ) ;
INV     gate12740  (.A(g22192), .Z(II31159) ) ;
INV     gate12741  (.A(II31159), .Z(g23895) ) ;
NOR2    gate12742  (.A(g21522), .B(g19857), .Z(g22193) ) ;
INV     gate12743  (.A(g22193), .Z(II31162) ) ;
INV     gate12744  (.A(II31162), .Z(g23896) ) ;
NOR2    gate12745  (.A(g21523), .B(g19858), .Z(g22194) ) ;
INV     gate12746  (.A(g22194), .Z(II31165) ) ;
INV     gate12747  (.A(II31165), .Z(g23897) ) ;
NAND2   gate12748  (.A(g21732), .B(g2746), .Z(g23033) ) ;
INV     gate12749  (.A(g23033), .Z(II31171) ) ;
INV     gate12750  (.A(II31171), .Z(g23901) ) ;
AND4    gate12751  (.A(g21117), .B(g21105), .C(g21096), .D(II28594), .Z(g22046) ) ;
INV     gate12752  (.A(g22046), .Z(g23905) ) ;
INV     gate12753  (.A(g22353), .Z(g23908) ) ;
NOR2    gate12754  (.A(g21553), .B(g19883), .Z(g22200) ) ;
INV     gate12755  (.A(g22200), .Z(II31181) ) ;
INV     gate12756  (.A(II31181), .Z(g23911) ) ;
NAND2   gate12757  (.A(g21048), .B(g18623), .Z(g21989) ) ;
INV     gate12758  (.A(g21989), .Z(II31188) ) ;
INV     gate12759  (.A(II31188), .Z(g23916) ) ;
AND4    gate12760  (.A(g21104), .B(g21095), .C(g21084), .D(II28582), .Z(g22036) ) ;
INV     gate12761  (.A(g22036), .Z(g23918) ) ;
NOR2    gate12762  (.A(g21892), .B(g18982), .Z(g22578) ) ;
INV     gate12763  (.A(g22578), .Z(II31195) ) ;
INV     gate12764  (.A(II31195), .Z(g23923) ) ;
INV     gate12765  (.A(g22376), .Z(g23940) ) ;
NAND2   gate12766  (.A(g21065), .B(g21711), .Z(g22002) ) ;
INV     gate12767  (.A(g22002), .Z(II31205) ) ;
INV     gate12768  (.A(II31205), .Z(g23943) ) ;
NOR2    gate12769  (.A(g21900), .B(g18990), .Z(g22615) ) ;
INV     gate12770  (.A(g22615), .Z(II31213) ) ;
INV     gate12771  (.A(II31213), .Z(g23955) ) ;
NOR2    gate12772  (.A(g21912), .B(g18997), .Z(g22651) ) ;
INV     gate12773  (.A(g22651), .Z(II31226) ) ;
INV     gate12774  (.A(II31226), .Z(g23984) ) ;
NOR2    gate12775  (.A(g21083), .B(g18407), .Z(g22026) ) ;
INV     gate12776  (.A(g22026), .Z(II31232) ) ;
INV     gate12777  (.A(II31232), .Z(g24000) ) ;
NOR2    gate12778  (.A(g21639), .B(g19949), .Z(g22218) ) ;
INV     gate12779  (.A(g22218), .Z(II31235) ) ;
INV     gate12780  (.A(II31235), .Z(g24001) ) ;
NOR2    gate12781  (.A(g21926), .B(g19010), .Z(g22687) ) ;
INV     gate12782  (.A(g22687), .Z(II31244) ) ;
INV     gate12783  (.A(II31244), .Z(g24014) ) ;
NOR2    gate12784  (.A(g20700), .B(g7595), .Z(g22953) ) ;
INV     gate12785  (.A(g22953), .Z(II31250) ) ;
INV     gate12786  (.A(II31250), .Z(g24030) ) ;
NOR2    gate12787  (.A(g21666), .B(g19971), .Z(g22231) ) ;
INV     gate12788  (.A(g22231), .Z(II31253) ) ;
INV     gate12789  (.A(II31253), .Z(g24033) ) ;
NOR2    gate12790  (.A(g21670), .B(g19976), .Z(g22234) ) ;
INV     gate12791  (.A(g22234), .Z(II31257) ) ;
INV     gate12792  (.A(II31257), .Z(g24035) ) ;
NOR3    gate12793  (.A(g14256), .B(g14175), .C(g21123), .Z(g23023) ) ;
INV     gate12794  (.A(g23023), .Z(g24047) ) ;
NOR2    gate12795  (.A(g21687), .B(g19983), .Z(g22242) ) ;
INV     gate12796  (.A(g22242), .Z(II31266) ) ;
INV     gate12797  (.A(II31266), .Z(g24051) ) ;
NOR2    gate12798  (.A(g21695), .B(g20001), .Z(g22247) ) ;
INV     gate12799  (.A(g22247), .Z(II31270) ) ;
INV     gate12800  (.A(II31270), .Z(g24053) ) ;
NOR2    gate12801  (.A(g21699), .B(g20006), .Z(g22249) ) ;
INV     gate12802  (.A(g22249), .Z(II31274) ) ;
INV     gate12803  (.A(II31274), .Z(g24055) ) ;
NOR3    gate12804  (.A(g14378), .B(g14290), .C(g21142), .Z(g23040) ) ;
INV     gate12805  (.A(g23040), .Z(g24060) ) ;
NOR2    gate12806  (.A(g21723), .B(g20021), .Z(g22263) ) ;
INV     gate12807  (.A(g22263), .Z(II31282) ) ;
INV     gate12808  (.A(II31282), .Z(g24064) ) ;
NOR2    gate12809  (.A(g21731), .B(g20039), .Z(g22267) ) ;
INV     gate12810  (.A(g22267), .Z(II31286) ) ;
INV     gate12811  (.A(II31286), .Z(g24066) ) ;
NOR2    gate12812  (.A(g21735), .B(g20044), .Z(g22269) ) ;
INV     gate12813  (.A(g22269), .Z(II31290) ) ;
INV     gate12814  (.A(II31290), .Z(g24068) ) ;
NOR3    gate12815  (.A(g14490), .B(g14412), .C(g21162), .Z(g23059) ) ;
INV     gate12816  (.A(g23059), .Z(g24073) ) ;
NOR2    gate12817  (.A(g21749), .B(g20063), .Z(g22280) ) ;
INV     gate12818  (.A(g22280), .Z(II31298) ) ;
INV     gate12819  (.A(II31298), .Z(g24077) ) ;
NOR2    gate12820  (.A(g21757), .B(g20081), .Z(g22284) ) ;
INV     gate12821  (.A(g22284), .Z(II31302) ) ;
INV     gate12822  (.A(II31302), .Z(g24079) ) ;
NOR3    gate12823  (.A(g14577), .B(g14524), .C(g21182), .Z(g23077) ) ;
INV     gate12824  (.A(g23077), .Z(g24084) ) ;
NOR2    gate12825  (.A(g21773), .B(g20104), .Z(g22299) ) ;
INV     gate12826  (.A(g22299), .Z(II31310) ) ;
INV     gate12827  (.A(II31310), .Z(g24088) ) ;
NAND3   gate12828  (.A(g14442), .B(g21149), .C(g10694), .Z(g22339) ) ;
INV     gate12829  (.A(g22339), .Z(g24094) ) ;
NAND3   gate12830  (.A(g14529), .B(g21169), .C(g10714), .Z(g22362) ) ;
INV     gate12831  (.A(g22362), .Z(g24095) ) ;
INV     gate12832  (.A(g22405), .Z(g24096) ) ;
NAND3   gate12833  (.A(g14584), .B(g21189), .C(g10735), .Z(g22382) ) ;
INV     gate12834  (.A(g22382), .Z(g24097) ) ;
INV     gate12835  (.A(g22409), .Z(g24098) ) ;
INV     gate12836  (.A(g22412), .Z(g24099) ) ;
INV     gate12837  (.A(g22415), .Z(g24101) ) ;
INV     gate12838  (.A(g22418), .Z(g24102) ) ;
NAND3   gate12839  (.A(g14618), .B(g21204), .C(g10754), .Z(g22397) ) ;
INV     gate12840  (.A(g22397), .Z(g24103) ) ;
INV     gate12841  (.A(g22422), .Z(g24104) ) ;
INV     gate12842  (.A(g22425), .Z(g24105) ) ;
INV     gate12843  (.A(g22428), .Z(g24106) ) ;
INV     gate12844  (.A(g22431), .Z(g24107) ) ;
INV     gate12845  (.A(g22434), .Z(g24108) ) ;
INV     gate12846  (.A(g22437), .Z(g24110) ) ;
INV     gate12847  (.A(g22440), .Z(g24111) ) ;
INV     gate12848  (.A(g22445), .Z(g24112) ) ;
INV     gate12849  (.A(g22448), .Z(g24113) ) ;
INV     gate12850  (.A(g22451), .Z(g24114) ) ;
NAND3   gate12851  (.A(g21211), .B(g14442), .C(g10694), .Z(g22381) ) ;
INV     gate12852  (.A(g22381), .Z(g24115) ) ;
INV     gate12853  (.A(g22455), .Z(g24121) ) ;
INV     gate12854  (.A(g22458), .Z(g24122) ) ;
INV     gate12855  (.A(g22461), .Z(g24123) ) ;
INV     gate12856  (.A(g22464), .Z(g24124) ) ;
INV     gate12857  (.A(g22467), .Z(g24125) ) ;
INV     gate12858  (.A(g22470), .Z(g24127) ) ;
INV     gate12859  (.A(g22473), .Z(g24128) ) ;
INV     gate12860  (.A(g22477), .Z(g24129) ) ;
INV     gate12861  (.A(g22480), .Z(g24130) ) ;
INV     gate12862  (.A(g22484), .Z(g24131) ) ;
INV     gate12863  (.A(g22487), .Z(g24132) ) ;
INV     gate12864  (.A(g22490), .Z(g24133) ) ;
NAND3   gate12865  (.A(g21219), .B(g14529), .C(g10714), .Z(g22396) ) ;
INV     gate12866  (.A(g22396), .Z(g24134) ) ;
INV     gate12867  (.A(g22494), .Z(g24140) ) ;
INV     gate12868  (.A(g22497), .Z(g24141) ) ;
INV     gate12869  (.A(g22500), .Z(g24142) ) ;
INV     gate12870  (.A(g22503), .Z(g24143) ) ;
INV     gate12871  (.A(g22506), .Z(g24144) ) ;
INV     gate12872  (.A(g22509), .Z(g24146) ) ;
INV     gate12873  (.A(g22512), .Z(g24147) ) ;
INV     gate12874  (.A(g22520), .Z(g24148) ) ;
INV     gate12875  (.A(g22523), .Z(g24149) ) ;
INV     gate12876  (.A(g22527), .Z(g24150) ) ;
INV     gate12877  (.A(g22530), .Z(g24151) ) ;
INV     gate12878  (.A(g22533), .Z(g24152) ) ;
NAND3   gate12879  (.A(g21230), .B(g14584), .C(g10735), .Z(g22399) ) ;
INV     gate12880  (.A(g22399), .Z(g24153) ) ;
INV     gate12881  (.A(g22537), .Z(g24159) ) ;
INV     gate12882  (.A(g22540), .Z(g24160) ) ;
INV     gate12883  (.A(g22543), .Z(g24161) ) ;
INV     gate12884  (.A(g22552), .Z(g24162) ) ;
INV     gate12885  (.A(g22560), .Z(g24163) ) ;
INV     gate12886  (.A(g22563), .Z(g24164) ) ;
INV     gate12887  (.A(g22567), .Z(g24165) ) ;
INV     gate12888  (.A(g22570), .Z(g24166) ) ;
INV     gate12889  (.A(g22573), .Z(g24167) ) ;
NAND3   gate12890  (.A(g21235), .B(g14618), .C(g10754), .Z(g22400) ) ;
INV     gate12891  (.A(g22400), .Z(g24168) ) ;
INV     gate12892  (.A(g22592), .Z(g24175) ) ;
INV     gate12893  (.A(g22600), .Z(g24176) ) ;
INV     gate12894  (.A(g22603), .Z(g24177) ) ;
INV     gate12895  (.A(g22629), .Z(g24180) ) ;
OR4     gate12896  (.A(g562), .B(g559), .C(g12451), .D(g21851), .Z(g22811) ) ;
INV     gate12897  (.A(g22811), .Z(II31387) ) ;
INV     gate12898  (.A(II31387), .Z(g24183) ) ;
INV     gate12899  (.A(g22696), .Z(g24210) ) ;
INV     gate12900  (.A(g22750), .Z(g24220) ) ;
INV     gate12901  (.A(g22578), .Z(II31417) ) ;
INV     gate12902  (.A(II31417), .Z(g24233) ) ;
INV     gate12903  (.A(g22615), .Z(II31426) ) ;
INV     gate12904  (.A(II31426), .Z(g24240) ) ;
INV     gate12905  (.A(g22651), .Z(II31436) ) ;
INV     gate12906  (.A(II31436), .Z(g24248) ) ;
INV     gate12907  (.A(g22903), .Z(g24251) ) ;
INV     gate12908  (.A(g22687), .Z(II31445) ) ;
INV     gate12909  (.A(II31445), .Z(g24255) ) ;
INV     gate12910  (.A(g23682), .Z(II31451) ) ;
INV     gate12911  (.A(g23727), .Z(II31454) ) ;
INV     gate12912  (.A(g23773), .Z(II31457) ) ;
INV     gate12913  (.A(g23728), .Z(II31460) ) ;
INV     gate12914  (.A(g23774), .Z(II31463) ) ;
INV     gate12915  (.A(g23821), .Z(II31466) ) ;
INV     gate12916  (.A(g23546), .Z(II31469) ) ;
INV     gate12917  (.A(g23548), .Z(II31472) ) ;
INV     gate12918  (.A(g23555), .Z(II31475) ) ;
INV     gate12919  (.A(g23549), .Z(II31478) ) ;
INV     gate12920  (.A(g23556), .Z(II31481) ) ;
INV     gate12921  (.A(g23568), .Z(II31484) ) ;
INV     gate12922  (.A(g23557), .Z(II31487) ) ;
INV     gate12923  (.A(g23569), .Z(II31490) ) ;
INV     gate12924  (.A(g23587), .Z(II31493) ) ;
INV     gate12925  (.A(g23570), .Z(II31496) ) ;
INV     gate12926  (.A(g23588), .Z(II31499) ) ;
INV     gate12927  (.A(g23612), .Z(II31502) ) ;
INV     gate12928  (.A(g23589), .Z(II31505) ) ;
INV     gate12929  (.A(g23613), .Z(II31508) ) ;
INV     gate12930  (.A(g23640), .Z(II31511) ) ;
INV     gate12931  (.A(g23614), .Z(II31514) ) ;
INV     gate12932  (.A(g23641), .Z(II31517) ) ;
INV     gate12933  (.A(g23683), .Z(II31520) ) ;
INV     gate12934  (.A(g23642), .Z(II31523) ) ;
INV     gate12935  (.A(g23684), .Z(II31526) ) ;
INV     gate12936  (.A(g23729), .Z(II31529) ) ;
INV     gate12937  (.A(g23685), .Z(II31532) ) ;
INV     gate12938  (.A(g23730), .Z(II31535) ) ;
INV     gate12939  (.A(g23775), .Z(II31538) ) ;
INV     gate12940  (.A(g23500), .Z(II31541) ) ;
INV     gate12941  (.A(g23438), .Z(II31544) ) ;
INV     gate12942  (.A(g23454), .Z(II31547) ) ;
INV     gate12943  (.A(g23481), .Z(II31550) ) ;
INV     gate12944  (.A(g23501), .Z(II31553) ) ;
INV     gate12945  (.A(g23439), .Z(II31556) ) ;
INV     gate12946  (.A(g24233), .Z(II31559) ) ;
INV     gate12947  (.A(g23594), .Z(II31562) ) ;
INV     gate12948  (.A(g24001), .Z(II31565) ) ;
INV     gate12949  (.A(g24033), .Z(II31568) ) ;
INV     gate12950  (.A(g24051), .Z(II31571) ) ;
INV     gate12951  (.A(g23736), .Z(II31574) ) ;
INV     gate12952  (.A(g23782), .Z(II31577) ) ;
INV     gate12953  (.A(g23826), .Z(II31580) ) ;
INV     gate12954  (.A(g23783), .Z(II31583) ) ;
INV     gate12955  (.A(g23827), .Z(II31586) ) ;
INV     gate12956  (.A(g23856), .Z(II31589) ) ;
INV     gate12957  (.A(g23553), .Z(II31592) ) ;
INV     gate12958  (.A(g23561), .Z(II31595) ) ;
INV     gate12959  (.A(g23574), .Z(II31598) ) ;
INV     gate12960  (.A(g23562), .Z(II31601) ) ;
INV     gate12961  (.A(g23575), .Z(II31604) ) ;
INV     gate12962  (.A(g23595), .Z(II31607) ) ;
INV     gate12963  (.A(g23576), .Z(II31610) ) ;
INV     gate12964  (.A(g23596), .Z(II31613) ) ;
INV     gate12965  (.A(g23619), .Z(II31616) ) ;
INV     gate12966  (.A(g23597), .Z(II31619) ) ;
INV     gate12967  (.A(g23620), .Z(II31622) ) ;
INV     gate12968  (.A(g23661), .Z(II31625) ) ;
INV     gate12969  (.A(g23621), .Z(II31628) ) ;
INV     gate12970  (.A(g23662), .Z(II31631) ) ;
INV     gate12971  (.A(g23690), .Z(II31634) ) ;
INV     gate12972  (.A(g23663), .Z(II31637) ) ;
INV     gate12973  (.A(g23691), .Z(II31640) ) ;
INV     gate12974  (.A(g23737), .Z(II31643) ) ;
INV     gate12975  (.A(g23692), .Z(II31646) ) ;
INV     gate12976  (.A(g23738), .Z(II31649) ) ;
INV     gate12977  (.A(g23784), .Z(II31652) ) ;
INV     gate12978  (.A(g23739), .Z(II31655) ) ;
INV     gate12979  (.A(g23785), .Z(II31658) ) ;
INV     gate12980  (.A(g23828), .Z(II31661) ) ;
INV     gate12981  (.A(g23516), .Z(II31664) ) ;
INV     gate12982  (.A(g23452), .Z(II31667) ) ;
INV     gate12983  (.A(g23463), .Z(II31670) ) ;
INV     gate12984  (.A(g23492), .Z(II31673) ) ;
INV     gate12985  (.A(g23517), .Z(II31676) ) ;
INV     gate12986  (.A(g23453), .Z(II31679) ) ;
INV     gate12987  (.A(g24240), .Z(II31682) ) ;
INV     gate12988  (.A(g23626), .Z(II31685) ) ;
INV     gate12989  (.A(g24035), .Z(II31688) ) ;
INV     gate12990  (.A(g24053), .Z(II31691) ) ;
INV     gate12991  (.A(g24064), .Z(II31694) ) ;
INV     gate12992  (.A(g23791), .Z(II31697) ) ;
INV     gate12993  (.A(g23835), .Z(II31700) ) ;
INV     gate12994  (.A(g23861), .Z(II31703) ) ;
INV     gate12995  (.A(g23836), .Z(II31706) ) ;
INV     gate12996  (.A(g23862), .Z(II31709) ) ;
INV     gate12997  (.A(g23890), .Z(II31712) ) ;
INV     gate12998  (.A(g23566), .Z(II31715) ) ;
INV     gate12999  (.A(g23580), .Z(II31718) ) ;
INV     gate13000  (.A(g23601), .Z(II31721) ) ;
INV     gate13001  (.A(g23581), .Z(II31724) ) ;
INV     gate13002  (.A(g23602), .Z(II31727) ) ;
INV     gate13003  (.A(g23627), .Z(II31730) ) ;
INV     gate13004  (.A(g23603), .Z(II31733) ) ;
INV     gate13005  (.A(g23628), .Z(II31736) ) ;
INV     gate13006  (.A(g23668), .Z(II31739) ) ;
INV     gate13007  (.A(g23629), .Z(II31742) ) ;
INV     gate13008  (.A(g23669), .Z(II31745) ) ;
INV     gate13009  (.A(g23711), .Z(II31748) ) ;
INV     gate13010  (.A(g23670), .Z(II31751) ) ;
INV     gate13011  (.A(g23712), .Z(II31754) ) ;
INV     gate13012  (.A(g23744), .Z(II31757) ) ;
INV     gate13013  (.A(g23713), .Z(II31760) ) ;
INV     gate13014  (.A(g23745), .Z(II31763) ) ;
INV     gate13015  (.A(g23792), .Z(II31766) ) ;
INV     gate13016  (.A(g23746), .Z(II31769) ) ;
INV     gate13017  (.A(g23793), .Z(II31772) ) ;
INV     gate13018  (.A(g23837), .Z(II31775) ) ;
INV     gate13019  (.A(g23794), .Z(II31778) ) ;
INV     gate13020  (.A(g23838), .Z(II31781) ) ;
INV     gate13021  (.A(g23863), .Z(II31784) ) ;
INV     gate13022  (.A(g23531), .Z(II31787) ) ;
INV     gate13023  (.A(g23459), .Z(II31790) ) ;
INV     gate13024  (.A(g23472), .Z(II31793) ) ;
INV     gate13025  (.A(g23508), .Z(II31796) ) ;
INV     gate13026  (.A(g23532), .Z(II31799) ) ;
INV     gate13027  (.A(g23460), .Z(II31802) ) ;
INV     gate13028  (.A(g24248), .Z(II31805) ) ;
INV     gate13029  (.A(g23675), .Z(II31808) ) ;
INV     gate13030  (.A(g24055), .Z(II31811) ) ;
INV     gate13031  (.A(g24066), .Z(II31814) ) ;
INV     gate13032  (.A(g24077), .Z(II31817) ) ;
INV     gate13033  (.A(g23844), .Z(II31820) ) ;
INV     gate13034  (.A(g23870), .Z(II31823) ) ;
INV     gate13035  (.A(g23895), .Z(II31826) ) ;
INV     gate13036  (.A(g23871), .Z(II31829) ) ;
INV     gate13037  (.A(g23896), .Z(II31832) ) ;
INV     gate13038  (.A(g23911), .Z(II31835) ) ;
INV     gate13039  (.A(g23585), .Z(II31838) ) ;
INV     gate13040  (.A(g23607), .Z(II31841) ) ;
INV     gate13041  (.A(g23633), .Z(II31844) ) ;
INV     gate13042  (.A(g23608), .Z(II31847) ) ;
INV     gate13043  (.A(g23634), .Z(II31850) ) ;
INV     gate13044  (.A(g23676), .Z(II31853) ) ;
INV     gate13045  (.A(g23635), .Z(II31856) ) ;
INV     gate13046  (.A(g23677), .Z(II31859) ) ;
INV     gate13047  (.A(g23718), .Z(II31862) ) ;
INV     gate13048  (.A(g23678), .Z(II31865) ) ;
INV     gate13049  (.A(g23719), .Z(II31868) ) ;
INV     gate13050  (.A(g23765), .Z(II31871) ) ;
INV     gate13051  (.A(g23720), .Z(II31874) ) ;
INV     gate13052  (.A(g23766), .Z(II31877) ) ;
INV     gate13053  (.A(g23799), .Z(II31880) ) ;
INV     gate13054  (.A(g23767), .Z(II31883) ) ;
INV     gate13055  (.A(g23800), .Z(II31886) ) ;
INV     gate13056  (.A(g23845), .Z(II31889) ) ;
INV     gate13057  (.A(g23801), .Z(II31892) ) ;
INV     gate13058  (.A(g23846), .Z(II31895) ) ;
INV     gate13059  (.A(g23872), .Z(II31898) ) ;
INV     gate13060  (.A(g23847), .Z(II31901) ) ;
INV     gate13061  (.A(g23873), .Z(II31904) ) ;
INV     gate13062  (.A(g23897), .Z(II31907) ) ;
INV     gate13063  (.A(g23542), .Z(II31910) ) ;
INV     gate13064  (.A(g23468), .Z(II31913) ) ;
INV     gate13065  (.A(g23485), .Z(II31916) ) ;
INV     gate13066  (.A(g23524), .Z(II31919) ) ;
INV     gate13067  (.A(g23543), .Z(II31922) ) ;
INV     gate13068  (.A(g23469), .Z(II31925) ) ;
INV     gate13069  (.A(g24255), .Z(II31928) ) ;
INV     gate13070  (.A(g23725), .Z(II31931) ) ;
INV     gate13071  (.A(g24068), .Z(II31934) ) ;
INV     gate13072  (.A(g24079), .Z(II31937) ) ;
INV     gate13073  (.A(g24088), .Z(II31940) ) ;
INV     gate13074  (.A(g24000), .Z(II31943) ) ;
INV     gate13075  (.A(g23916), .Z(II31946) ) ;
INV     gate13076  (.A(g23943), .Z(II31949) ) ;
INV     gate13077  (.A(g24183), .Z(g24482) ) ;
NOR2    gate13078  (.A(g17506), .B(g22581), .Z(g23399) ) ;
INV     gate13079  (.A(g23399), .Z(II32042) ) ;
INV     gate13080  (.A(II32042), .Z(g24518) ) ;
NOR2    gate13081  (.A(g17597), .B(g22618), .Z(g23406) ) ;
INV     gate13082  (.A(g23406), .Z(II32057) ) ;
INV     gate13083  (.A(II32057), .Z(g24531) ) ;
NOR2    gate13084  (.A(g16894), .B(g22206), .Z(g24174) ) ;
INV     gate13085  (.A(g24174), .Z(II32067) ) ;
INV     gate13086  (.A(II32067), .Z(g24539) ) ;
NOR2    gate13087  (.A(g17694), .B(g22654), .Z(g23413) ) ;
INV     gate13088  (.A(g23413), .Z(II32074) ) ;
INV     gate13089  (.A(II32074), .Z(g24544) ) ;
NOR2    gate13090  (.A(g16908), .B(g22211), .Z(g24178) ) ;
INV     gate13091  (.A(g24178), .Z(II32081) ) ;
INV     gate13092  (.A(II32081), .Z(g24549) ) ;
NOR2    gate13093  (.A(g16923), .B(g22214), .Z(g24179) ) ;
INV     gate13094  (.A(g24179), .Z(II32085) ) ;
INV     gate13095  (.A(II32085), .Z(g24551) ) ;
NOR2    gate13096  (.A(g17794), .B(g22690), .Z(g23418) ) ;
INV     gate13097  (.A(g23418), .Z(II32092) ) ;
INV     gate13098  (.A(II32092), .Z(g24556) ) ;
NOR2    gate13099  (.A(g16938), .B(g22220), .Z(g24181) ) ;
INV     gate13100  (.A(g24181), .Z(II32098) ) ;
INV     gate13101  (.A(II32098), .Z(g24560) ) ;
NOR2    gate13102  (.A(g16953), .B(g22223), .Z(g24182) ) ;
INV     gate13103  (.A(g24182), .Z(II32102) ) ;
INV     gate13104  (.A(II32102), .Z(g24562) ) ;
NOR2    gate13105  (.A(g16966), .B(g22228), .Z(g24206) ) ;
INV     gate13106  (.A(g24206), .Z(II32109) ) ;
INV     gate13107  (.A(II32109), .Z(g24567) ) ;
NOR2    gate13108  (.A(g16967), .B(g22229), .Z(g24207) ) ;
INV     gate13109  (.A(g24207), .Z(II32112) ) ;
INV     gate13110  (.A(II32112), .Z(g24568) ) ;
NOR2    gate13111  (.A(g16969), .B(g22235), .Z(g24208) ) ;
INV     gate13112  (.A(g24208), .Z(II32116) ) ;
INV     gate13113  (.A(II32116), .Z(g24570) ) ;
NOR2    gate13114  (.A(g16984), .B(g22238), .Z(g24209) ) ;
INV     gate13115  (.A(g24209), .Z(II32120) ) ;
INV     gate13116  (.A(II32120), .Z(g24572) ) ;
NOR2    gate13117  (.A(g16987), .B(g22244), .Z(g24212) ) ;
INV     gate13118  (.A(g24212), .Z(II32126) ) ;
INV     gate13119  (.A(II32126), .Z(g24576) ) ;
NOR2    gate13120  (.A(g16988), .B(g22245), .Z(g24213) ) ;
INV     gate13121  (.A(g24213), .Z(II32129) ) ;
INV     gate13122  (.A(II32129), .Z(g24577) ) ;
NOR2    gate13123  (.A(g16990), .B(g22250), .Z(g24214) ) ;
INV     gate13124  (.A(g24214), .Z(II32133) ) ;
INV     gate13125  (.A(II32133), .Z(g24579) ) ;
NOR2    gate13126  (.A(g16993), .B(g22254), .Z(g24215) ) ;
INV     gate13127  (.A(g24215), .Z(II32137) ) ;
INV     gate13128  (.A(II32137), .Z(g24581) ) ;
NOR2    gate13129  (.A(g16994), .B(g22255), .Z(g24216) ) ;
INV     gate13130  (.A(g24216), .Z(II32140) ) ;
INV     gate13131  (.A(II32140), .Z(g24582) ) ;
NOR2    gate13132  (.A(g16997), .B(g22264), .Z(g24218) ) ;
INV     gate13133  (.A(g24218), .Z(II32143) ) ;
INV     gate13134  (.A(II32143), .Z(g24583) ) ;
NOR2    gate13135  (.A(g16998), .B(g22265), .Z(g24219) ) ;
INV     gate13136  (.A(g24219), .Z(II32146) ) ;
INV     gate13137  (.A(II32146), .Z(g24584) ) ;
NOR2    gate13138  (.A(g17017), .B(g22272), .Z(g24222) ) ;
INV     gate13139  (.A(g24222), .Z(II32150) ) ;
INV     gate13140  (.A(II32150), .Z(g24586) ) ;
NOR2    gate13141  (.A(g17018), .B(g22273), .Z(g24223) ) ;
INV     gate13142  (.A(g24223), .Z(II32153) ) ;
INV     gate13143  (.A(II32153), .Z(g24587) ) ;
NOR2    gate13144  (.A(g17021), .B(g22281), .Z(g24225) ) ;
INV     gate13145  (.A(g24225), .Z(II32156) ) ;
INV     gate13146  (.A(II32156), .Z(g24588) ) ;
NOR2    gate13147  (.A(g17022), .B(g22282), .Z(g24226) ) ;
INV     gate13148  (.A(g24226), .Z(II32159) ) ;
INV     gate13149  (.A(II32159), .Z(g24589) ) ;
NOR2    gate13150  (.A(g17028), .B(g22285), .Z(g24228) ) ;
INV     gate13151  (.A(g24228), .Z(II32164) ) ;
INV     gate13152  (.A(II32164), .Z(g24592) ) ;
NOR2    gate13153  (.A(g17047), .B(g22291), .Z(g24230) ) ;
INV     gate13154  (.A(g24230), .Z(II32167) ) ;
INV     gate13155  (.A(II32167), .Z(g24593) ) ;
NOR2    gate13156  (.A(g17048), .B(g22292), .Z(g24231) ) ;
INV     gate13157  (.A(g24231), .Z(II32170) ) ;
INV     gate13158  (.A(II32170), .Z(g24594) ) ;
NOR2    gate13159  (.A(g17062), .B(g22305), .Z(g24235) ) ;
INV     gate13160  (.A(g24235), .Z(II32175) ) ;
INV     gate13161  (.A(II32175), .Z(g24597) ) ;
NOR2    gate13162  (.A(g17081), .B(g22311), .Z(g24237) ) ;
INV     gate13163  (.A(g24237), .Z(II32178) ) ;
INV     gate13164  (.A(II32178), .Z(g24598) ) ;
NOR2    gate13165  (.A(g17082), .B(g22312), .Z(g24238) ) ;
INV     gate13166  (.A(g24238), .Z(II32181) ) ;
INV     gate13167  (.A(II32181), .Z(g24599) ) ;
NOR2    gate13168  (.A(g22876), .B(g5606), .Z(g23497) ) ;
INV     gate13169  (.A(g23497), .Z(II32184) ) ;
INV     gate13170  (.A(II32184), .Z(g24600) ) ;
NOR2    gate13171  (.A(g17097), .B(g22333), .Z(g24243) ) ;
INV     gate13172  (.A(g24243), .Z(II32189) ) ;
INV     gate13173  (.A(II32189), .Z(g24605) ) ;
NOR2    gate13174  (.A(g22911), .B(g5631), .Z(g23513) ) ;
INV     gate13175  (.A(g23513), .Z(II32193) ) ;
INV     gate13176  (.A(II32193), .Z(g24607) ) ;
NOR2    gate13177  (.A(g17135), .B(g22358), .Z(g24250) ) ;
INV     gate13178  (.A(g24250), .Z(II32198) ) ;
INV     gate13179  (.A(II32198), .Z(g24612) ) ;
NOR2    gate13180  (.A(g22936), .B(g5659), .Z(g23528) ) ;
INV     gate13181  (.A(g23528), .Z(II32203) ) ;
INV     gate13182  (.A(II32203), .Z(g24619) ) ;
NOR2    gate13183  (.A(g22942), .B(g5697), .Z(g23539) ) ;
INV     gate13184  (.A(g23539), .Z(II32210) ) ;
INV     gate13185  (.A(II32210), .Z(g24630) ) ;
INV     gate13186  (.A(g23470), .Z(g24648) ) ;
INV     gate13187  (.A(g23482), .Z(g24668) ) ;
INV     gate13188  (.A(g23493), .Z(g24687) ) ;
INV     gate13189  (.A(g23509), .Z(g24704) ) ;
OR2     gate13190  (.A(g22666), .B(g23140), .Z(g23919) ) ;
INV     gate13191  (.A(g23919), .Z(II32248) ) ;
INV     gate13192  (.A(g23919), .Z(II32251) ) ;
INV     gate13193  (.A(II32251), .Z(g24735) ) ;
NOR2    gate13194  (.A(g22992), .B(g6707), .Z(g23950) ) ;
INV     gate13195  (.A(g23950), .Z(II32281) ) ;
INV     gate13196  (.A(II32281), .Z(g24763) ) ;
NOR2    gate13197  (.A(g23003), .B(g7009), .Z(g23979) ) ;
INV     gate13198  (.A(g23979), .Z(II32320) ) ;
INV     gate13199  (.A(II32320), .Z(g24784) ) ;
NOR2    gate13200  (.A(g23017), .B(g7259), .Z(g24009) ) ;
INV     gate13201  (.A(g24009), .Z(II32365) ) ;
INV     gate13202  (.A(II32365), .Z(g24805) ) ;
INV     gate13203  (.A(g23448), .Z(g24815) ) ;
NOR2    gate13204  (.A(g17393), .B(g22517), .Z(g23385) ) ;
INV     gate13205  (.A(g23385), .Z(II32388) ) ;
INV     gate13206  (.A(II32388), .Z(g24816) ) ;
NOR2    gate13207  (.A(g23033), .B(g7455), .Z(g24043) ) ;
INV     gate13208  (.A(g24043), .Z(II32419) ) ;
INV     gate13209  (.A(II32419), .Z(g24827) ) ;
INV     gate13210  (.A(g23455), .Z(g24834) ) ;
NOR2    gate13211  (.A(g17460), .B(g22557), .Z(g23392) ) ;
INV     gate13212  (.A(g23392), .Z(II32439) ) ;
INV     gate13213  (.A(II32439), .Z(g24835) ) ;
INV     gate13214  (.A(g23464), .Z(g24850) ) ;
NOR2    gate13215  (.A(g17540), .B(g22597), .Z(g23400) ) ;
INV     gate13216  (.A(g23400), .Z(II32487) ) ;
INV     gate13217  (.A(II32487), .Z(g24851) ) ;
NOR2    gate13218  (.A(g22144), .B(g10024), .Z(g23324) ) ;
INV     gate13219  (.A(g23324), .Z(II32506) ) ;
INV     gate13220  (.A(II32506), .Z(g24856) ) ;
INV     gate13221  (.A(g23473), .Z(g24864) ) ;
NOR2    gate13222  (.A(g17630), .B(g22634), .Z(g23407) ) ;
INV     gate13223  (.A(g23407), .Z(II32535) ) ;
INV     gate13224  (.A(II32535), .Z(g24865) ) ;
NOR2    gate13225  (.A(g22165), .B(g10133), .Z(g23329) ) ;
INV     gate13226  (.A(g23329), .Z(II32556) ) ;
INV     gate13227  (.A(II32556), .Z(g24872) ) ;
NOR2    gate13228  (.A(g22186), .B(g22777), .Z(g23330) ) ;
INV     gate13229  (.A(g23330), .Z(II32583) ) ;
INV     gate13230  (.A(II32583), .Z(g24879) ) ;
NOR2    gate13231  (.A(g22181), .B(g10238), .Z(g23339) ) ;
INV     gate13232  (.A(g23339), .Z(II32604) ) ;
INV     gate13233  (.A(II32604), .Z(g24886) ) ;
NAND3   gate13234  (.A(g22844), .B(g14442), .C(g10694), .Z(g23486) ) ;
INV     gate13235  (.A(g23486), .Z(g24893) ) ;
NOR2    gate13236  (.A(g22195), .B(g10340), .Z(g23348) ) ;
INV     gate13237  (.A(g23348), .Z(II32642) ) ;
INV     gate13238  (.A(II32642), .Z(g24903) ) ;
NAND3   gate13239  (.A(g10694), .B(g14442), .C(g22316), .Z(g23495) ) ;
INV     gate13240  (.A(g23495), .Z(g24912) ) ;
NAND3   gate13241  (.A(g22879), .B(g14529), .C(g10714), .Z(g23502) ) ;
INV     gate13242  (.A(g23502), .Z(g24916) ) ;
NAND3   gate13243  (.A(g10714), .B(g14529), .C(g22341), .Z(g23511) ) ;
INV     gate13244  (.A(g23511), .Z(g24929) ) ;
NAND3   gate13245  (.A(g22914), .B(g14584), .C(g10735), .Z(g23518) ) ;
INV     gate13246  (.A(g23518), .Z(g24933) ) ;
NAND2   gate13247  (.A(II30791), .B(II30792), .Z(g23660) ) ;
INV     gate13248  (.A(g23660), .Z(g24939) ) ;
NAND3   gate13249  (.A(g10735), .B(g14584), .C(g22364), .Z(g23526) ) ;
INV     gate13250  (.A(g23526), .Z(g24941) ) ;
NAND3   gate13251  (.A(g22939), .B(g14618), .C(g10754), .Z(g23533) ) ;
INV     gate13252  (.A(g23533), .Z(g24945) ) ;
NOR2    gate13253  (.A(g22210), .B(g20127), .Z(g23357) ) ;
INV     gate13254  (.A(g23357), .Z(II32704) ) ;
INV     gate13255  (.A(II32704), .Z(g24949) ) ;
NAND2   gate13256  (.A(II30869), .B(II30870), .Z(g23710) ) ;
INV     gate13257  (.A(g23710), .Z(g24950) ) ;
NAND3   gate13258  (.A(g10754), .B(g14618), .C(g22384), .Z(g23537) ) ;
INV     gate13259  (.A(g23537), .Z(g24952) ) ;
NOR2    gate13260  (.A(g22227), .B(g18407), .Z(g23358) ) ;
INV     gate13261  (.A(g23358), .Z(II32716) ) ;
INV     gate13262  (.A(II32716), .Z(g24956) ) ;
NOR2    gate13263  (.A(g22216), .B(g22907), .Z(g23359) ) ;
INV     gate13264  (.A(g23359), .Z(II32719) ) ;
INV     gate13265  (.A(II32719), .Z(g24957) ) ;
NAND3   gate13266  (.A(g22809), .B(g14442), .C(g10694), .Z(g23478) ) ;
INV     gate13267  (.A(g23478), .Z(g24958) ) ;
NAND2   gate13268  (.A(II30953), .B(II30954), .Z(g23764) ) ;
INV     gate13269  (.A(g23764), .Z(g24962) ) ;
NAND3   gate13270  (.A(g22850), .B(g14529), .C(g10714), .Z(g23489) ) ;
INV     gate13271  (.A(g23489), .Z(g24969) ) ;
NAND2   gate13272  (.A(II31036), .B(II31037), .Z(g23819) ) ;
INV     gate13273  (.A(g23819), .Z(g24973) ) ;
NAND3   gate13274  (.A(g22885), .B(g14584), .C(g10735), .Z(g23505) ) ;
INV     gate13275  (.A(g23505), .Z(g24982) ) ;
NAND3   gate13276  (.A(g22920), .B(g14618), .C(g10754), .Z(g23521) ) ;
INV     gate13277  (.A(g23521), .Z(g24993) ) ;
INV     gate13278  (.A(g23731), .Z(g25087) ) ;
INV     gate13279  (.A(g23779), .Z(g25094) ) ;
INV     gate13280  (.A(g23786), .Z(g25095) ) ;
NOR2    gate13281  (.A(g21990), .B(g20809), .Z(g24059) ) ;
INV     gate13282  (.A(g24059), .Z(II32829) ) ;
INV     gate13283  (.A(II32829), .Z(g25103) ) ;
INV     gate13284  (.A(g23832), .Z(g25104) ) ;
INV     gate13285  (.A(g23839), .Z(g25105) ) ;
NOR2    gate13286  (.A(g22004), .B(g20826), .Z(g24072) ) ;
INV     gate13287  (.A(g24072), .Z(II32835) ) ;
INV     gate13288  (.A(II32835), .Z(g25109) ) ;
INV     gate13289  (.A(g23867), .Z(g25110) ) ;
INV     gate13290  (.A(g23874), .Z(g25111) ) ;
INV     gate13291  (.A(g23879), .Z(g25115) ) ;
INV     gate13292  (.A(g23882), .Z(g25116) ) ;
INV     gate13293  (.A(g23644), .Z(II32844) ) ;
INV     gate13294  (.A(II32844), .Z(g25118) ) ;
NOR2    gate13295  (.A(g22015), .B(g20836), .Z(g24083) ) ;
INV     gate13296  (.A(g24083), .Z(II32847) ) ;
INV     gate13297  (.A(II32847), .Z(g25119) ) ;
INV     gate13298  (.A(g23901), .Z(g25120) ) ;
INV     gate13299  (.A(g23694), .Z(II32851) ) ;
INV     gate13300  (.A(II32851), .Z(g25121) ) ;
NOR2    gate13301  (.A(g22020), .B(g20840), .Z(g24092) ) ;
INV     gate13302  (.A(g24092), .Z(II32854) ) ;
INV     gate13303  (.A(II32854), .Z(g25122) ) ;
INV     gate13304  (.A(g23748), .Z(II32857) ) ;
INV     gate13305  (.A(II32857), .Z(g25123) ) ;
INV     gate13306  (.A(g23803), .Z(II32860) ) ;
INV     gate13307  (.A(II32860), .Z(g25124) ) ;
INV     gate13308  (.A(g24030), .Z(g25126) ) ;
INV     gate13309  (.A(g25118), .Z(II32868) ) ;
INV     gate13310  (.A(g24518), .Z(II32871) ) ;
INV     gate13311  (.A(g24539), .Z(II32874) ) ;
INV     gate13312  (.A(g24567), .Z(II32877) ) ;
INV     gate13313  (.A(g24581), .Z(II32880) ) ;
INV     gate13314  (.A(g24592), .Z(II32883) ) ;
INV     gate13315  (.A(g24549), .Z(II32886) ) ;
INV     gate13316  (.A(g24568), .Z(II32889) ) ;
INV     gate13317  (.A(g24582), .Z(II32892) ) ;
INV     gate13318  (.A(g24816), .Z(II32895) ) ;
INV     gate13319  (.A(g24856), .Z(II32898) ) ;
INV     gate13320  (.A(g25121), .Z(II32901) ) ;
INV     gate13321  (.A(g24531), .Z(II32904) ) ;
INV     gate13322  (.A(g24551), .Z(II32907) ) ;
INV     gate13323  (.A(g24576), .Z(II32910) ) ;
INV     gate13324  (.A(g24586), .Z(II32913) ) ;
INV     gate13325  (.A(g24597), .Z(II32916) ) ;
INV     gate13326  (.A(g24560), .Z(II32919) ) ;
INV     gate13327  (.A(g24577), .Z(II32922) ) ;
INV     gate13328  (.A(g24587), .Z(II32925) ) ;
INV     gate13329  (.A(g24835), .Z(II32928) ) ;
INV     gate13330  (.A(g24872), .Z(II32931) ) ;
INV     gate13331  (.A(g25123), .Z(II32934) ) ;
INV     gate13332  (.A(g24544), .Z(II32937) ) ;
INV     gate13333  (.A(g24562), .Z(II32940) ) ;
INV     gate13334  (.A(g24583), .Z(II32943) ) ;
INV     gate13335  (.A(g24593), .Z(II32946) ) ;
INV     gate13336  (.A(g24605), .Z(II32949) ) ;
INV     gate13337  (.A(g24570), .Z(II32952) ) ;
INV     gate13338  (.A(g24584), .Z(II32955) ) ;
INV     gate13339  (.A(g24594), .Z(II32958) ) ;
INV     gate13340  (.A(g24851), .Z(II32961) ) ;
INV     gate13341  (.A(g24886), .Z(II32964) ) ;
INV     gate13342  (.A(g25124), .Z(II32967) ) ;
INV     gate13343  (.A(g24556), .Z(II32970) ) ;
INV     gate13344  (.A(g24572), .Z(II32973) ) ;
INV     gate13345  (.A(g24588), .Z(II32976) ) ;
INV     gate13346  (.A(g24598), .Z(II32979) ) ;
INV     gate13347  (.A(g24612), .Z(II32982) ) ;
INV     gate13348  (.A(g24579), .Z(II32985) ) ;
INV     gate13349  (.A(g24589), .Z(II32988) ) ;
INV     gate13350  (.A(g24599), .Z(II32991) ) ;
INV     gate13351  (.A(g24865), .Z(II32994) ) ;
INV     gate13352  (.A(g24903), .Z(II32997) ) ;
INV     gate13353  (.A(g24949), .Z(II33000) ) ;
INV     gate13354  (.A(g24956), .Z(II33003) ) ;
INV     gate13355  (.A(g24957), .Z(II33006) ) ;
INV     gate13356  (.A(g24879), .Z(II33009) ) ;
INV     gate13357  (.A(g25119), .Z(II33013) ) ;
INV     gate13358  (.A(II33013), .Z(g25179) ) ;
INV     gate13359  (.A(g25122), .Z(II33016) ) ;
INV     gate13360  (.A(II33016), .Z(g25180) ) ;
INV     gate13361  (.A(g24912), .Z(g25274) ) ;
INV     gate13362  (.A(g24929), .Z(g25283) ) ;
INV     gate13363  (.A(g24941), .Z(g25291) ) ;
NAND2   gate13364  (.A(g23497), .B(g74), .Z(g24975) ) ;
INV     gate13365  (.A(g24975), .Z(II33128) ) ;
INV     gate13366  (.A(II33128), .Z(g25296) ) ;
INV     gate13367  (.A(g24952), .Z(g25301) ) ;
NAND2   gate13368  (.A(II32587), .B(II32588), .Z(g24880) ) ;
INV     gate13369  (.A(g24880), .Z(g25305) ) ;
NAND2   gate13370  (.A(g23513), .B(g762), .Z(g24986) ) ;
INV     gate13371  (.A(g24986), .Z(II33136) ) ;
INV     gate13372  (.A(II33136), .Z(g25306) ) ;
NAND2   gate13373  (.A(II32547), .B(II32548), .Z(g24868) ) ;
INV     gate13374  (.A(g24868), .Z(g25313) ) ;
NAND2   gate13375  (.A(II32625), .B(II32626), .Z(g24897) ) ;
INV     gate13376  (.A(g24897), .Z(g25314) ) ;
NAND2   gate13377  (.A(g23528), .B(g1448), .Z(g24997) ) ;
INV     gate13378  (.A(g24997), .Z(II33145) ) ;
INV     gate13379  (.A(II33145), .Z(g25315) ) ;
NAND2   gate13380  (.A(II32510), .B(II32511), .Z(g24857) ) ;
INV     gate13381  (.A(g24857), .Z(g25319) ) ;
NAND2   gate13382  (.A(II32596), .B(II32597), .Z(g24883) ) ;
INV     gate13383  (.A(g24883), .Z(g25322) ) ;
NAND2   gate13384  (.A(II32660), .B(II32661), .Z(g24920) ) ;
INV     gate13385  (.A(g24920), .Z(g25323) ) ;
NAND2   gate13386  (.A(g23539), .B(g2142), .Z(g25005) ) ;
INV     gate13387  (.A(g25005), .Z(II33154) ) ;
INV     gate13388  (.A(II33154), .Z(g25324) ) ;
NOR2    gate13389  (.A(g24227), .B(g17001), .Z(g25027) ) ;
INV     gate13390  (.A(g25027), .Z(II33157) ) ;
INV     gate13391  (.A(II33157), .Z(g25327) ) ;
NAND2   gate13392  (.A(II32469), .B(II32470), .Z(g24844) ) ;
INV     gate13393  (.A(g24844), .Z(g25329) ) ;
NAND2   gate13394  (.A(II32560), .B(II32561), .Z(g24873) ) ;
INV     gate13395  (.A(g24873), .Z(g25330) ) ;
NAND2   gate13396  (.A(II32634), .B(II32635), .Z(g24900) ) ;
INV     gate13397  (.A(g24900), .Z(g25332) ) ;
NAND2   gate13398  (.A(II32687), .B(II32688), .Z(g24937) ) ;
INV     gate13399  (.A(g24937), .Z(g25333) ) ;
NAND2   gate13400  (.A(II32431), .B(II32432), .Z(g24832) ) ;
INV     gate13401  (.A(g24832), .Z(g25335) ) ;
NOR2    gate13402  (.A(g24234), .B(g17031), .Z(g25042) ) ;
INV     gate13403  (.A(g25042), .Z(II33168) ) ;
INV     gate13404  (.A(II33168), .Z(g25336) ) ;
NAND2   gate13405  (.A(II32519), .B(II32520), .Z(g24860) ) ;
INV     gate13406  (.A(g24860), .Z(g25338) ) ;
NAND2   gate13407  (.A(II32608), .B(II32609), .Z(g24887) ) ;
INV     gate13408  (.A(g24887), .Z(g25339) ) ;
NAND2   gate13409  (.A(II32669), .B(II32670), .Z(g24923) ) ;
INV     gate13410  (.A(g24923), .Z(g25341) ) ;
NAND2   gate13411  (.A(II32392), .B(II32393), .Z(g24817) ) ;
INV     gate13412  (.A(g24817), .Z(g25347) ) ;
NAND2   gate13413  (.A(II32479), .B(II32480), .Z(g24848) ) ;
INV     gate13414  (.A(g24848), .Z(g25349) ) ;
NOR2    gate13415  (.A(g24242), .B(g17065), .Z(g25056) ) ;
INV     gate13416  (.A(g25056), .Z(II33182) ) ;
INV     gate13417  (.A(II33182), .Z(g25350) ) ;
NAND2   gate13418  (.A(II32568), .B(II32569), .Z(g24875) ) ;
INV     gate13419  (.A(g24875), .Z(g25352) ) ;
NAND2   gate13420  (.A(II32646), .B(II32647), .Z(g24904) ) ;
INV     gate13421  (.A(g24904), .Z(g25353) ) ;
NAND2   gate13422  (.A(g24239), .B(g24244), .Z(g24814) ) ;
INV     gate13423  (.A(g24814), .Z(II33188) ) ;
INV     gate13424  (.A(II33188), .Z(g25354) ) ;
NAND2   gate13425  (.A(II32346), .B(II32347), .Z(g24797) ) ;
INV     gate13426  (.A(g24797), .Z(g25355) ) ;
NAND2   gate13427  (.A(II32444), .B(II32445), .Z(g24837) ) ;
INV     gate13428  (.A(g24837), .Z(g25361) ) ;
NAND2   gate13429  (.A(II32527), .B(II32528), .Z(g24862) ) ;
INV     gate13430  (.A(g24862), .Z(g25363) ) ;
NOR2    gate13431  (.A(g24249), .B(g17100), .Z(g25067) ) ;
INV     gate13432  (.A(g25067), .Z(II33198) ) ;
INV     gate13433  (.A(II33198), .Z(g25364) ) ;
NAND2   gate13434  (.A(II32616), .B(II32617), .Z(g24889) ) ;
INV     gate13435  (.A(g24889), .Z(g25366) ) ;
AND2    gate13436  (.A(g13568), .B(g24115), .Z(g24676) ) ;
INV     gate13437  (.A(g24676), .Z(g25367) ) ;
NAND2   gate13438  (.A(II32309), .B(II32310), .Z(g24778) ) ;
INV     gate13439  (.A(g24778), .Z(g25368) ) ;
NAND2   gate13440  (.A(g24245), .B(g24252), .Z(g24833) ) ;
INV     gate13441  (.A(g24833), .Z(II33205) ) ;
INV     gate13442  (.A(II33205), .Z(g25369) ) ;
NAND2   gate13443  (.A(II32401), .B(II32402), .Z(g24820) ) ;
INV     gate13444  (.A(g24820), .Z(g25370) ) ;
NAND2   gate13445  (.A(II32491), .B(II32492), .Z(g24852) ) ;
INV     gate13446  (.A(g24852), .Z(g25376) ) ;
NAND2   gate13447  (.A(II32576), .B(II32577), .Z(g24877) ) ;
INV     gate13448  (.A(g24877), .Z(g25378) ) ;
INV     gate13449  (.A(g24893), .Z(g25379) ) ;
NAND2   gate13450  (.A(II32285), .B(II32286), .Z(g24766) ) ;
INV     gate13451  (.A(g24766), .Z(g25383) ) ;
AND2    gate13452  (.A(g13576), .B(g24134), .Z(g24695) ) ;
INV     gate13453  (.A(g24695), .Z(g25384) ) ;
NAND2   gate13454  (.A(II32356), .B(II32357), .Z(g24801) ) ;
INV     gate13455  (.A(g24801), .Z(g25385) ) ;
NAND2   gate13456  (.A(g24254), .B(g24257), .Z(g24849) ) ;
INV     gate13457  (.A(g24849), .Z(II33219) ) ;
INV     gate13458  (.A(II33219), .Z(g25386) ) ;
NAND2   gate13459  (.A(II32452), .B(II32453), .Z(g24839) ) ;
INV     gate13460  (.A(g24839), .Z(g25387) ) ;
NAND2   gate13461  (.A(II32539), .B(II32540), .Z(g24866) ) ;
INV     gate13462  (.A(g24866), .Z(g25393) ) ;
NAND2   gate13463  (.A(II32266), .B(II32267), .Z(g24753) ) ;
INV     gate13464  (.A(g24753), .Z(g25394) ) ;
INV     gate13465  (.A(g24916), .Z(g25395) ) ;
NAND2   gate13466  (.A(II32324), .B(II32325), .Z(g24787) ) ;
INV     gate13467  (.A(g24787), .Z(g25399) ) ;
AND2    gate13468  (.A(g13585), .B(g24153), .Z(g24712) ) ;
INV     gate13469  (.A(g24712), .Z(g25400) ) ;
NAND2   gate13470  (.A(II32410), .B(II32411), .Z(g24823) ) ;
INV     gate13471  (.A(g24823), .Z(g25401) ) ;
NAND2   gate13472  (.A(g24258), .B(g23319), .Z(g24863) ) ;
INV     gate13473  (.A(g24863), .Z(II33232) ) ;
INV     gate13474  (.A(II33232), .Z(g25402) ) ;
NAND2   gate13475  (.A(II32499), .B(II32500), .Z(g24854) ) ;
INV     gate13476  (.A(g24854), .Z(g25403) ) ;
NAND2   gate13477  (.A(II32296), .B(II32297), .Z(g24771) ) ;
INV     gate13478  (.A(g24771), .Z(g25404) ) ;
INV     gate13479  (.A(g24933), .Z(g25405) ) ;
NAND2   gate13480  (.A(II32369), .B(II32370), .Z(g24808) ) ;
INV     gate13481  (.A(g24808), .Z(g25409) ) ;
AND2    gate13482  (.A(g13605), .B(g24168), .Z(g24723) ) ;
INV     gate13483  (.A(g24723), .Z(g25410) ) ;
NAND2   gate13484  (.A(II32461), .B(II32462), .Z(g24842) ) ;
INV     gate13485  (.A(g24842), .Z(g25411) ) ;
NAND2   gate13486  (.A(II32334), .B(II32335), .Z(g24791) ) ;
INV     gate13487  (.A(g24791), .Z(g25412) ) ;
INV     gate13488  (.A(g24945), .Z(g25413) ) ;
NAND2   gate13489  (.A(II32423), .B(II32424), .Z(g24830) ) ;
INV     gate13490  (.A(g24830), .Z(g25417) ) ;
NAND2   gate13491  (.A(II32379), .B(II32380), .Z(g24812) ) ;
INV     gate13492  (.A(g24812), .Z(g25419) ) ;
OR2     gate13493  (.A(g23639), .B(g23144), .Z(g24890) ) ;
INV     gate13494  (.A(g24890), .Z(II33246) ) ;
INV     gate13495  (.A(g24890), .Z(II33249) ) ;
INV     gate13496  (.A(II33249), .Z(g25421) ) ;
INV     gate13497  (.A(g24958), .Z(g25422) ) ;
NAND2   gate13498  (.A(g499), .B(g23376), .Z(g24616) ) ;
INV     gate13499  (.A(g24616), .Z(g25430) ) ;
INV     gate13500  (.A(g24969), .Z(g25431) ) ;
OR2     gate13501  (.A(g23726), .B(g23142), .Z(g24909) ) ;
INV     gate13502  (.A(g24909), .Z(II33257) ) ;
INV     gate13503  (.A(g24909), .Z(II33260) ) ;
INV     gate13504  (.A(II33260), .Z(g25436) ) ;
NAND2   gate13505  (.A(g1186), .B(g23387), .Z(g24627) ) ;
INV     gate13506  (.A(g24627), .Z(g25437) ) ;
INV     gate13507  (.A(g24982), .Z(g25438) ) ;
OR2     gate13508  (.A(g23772), .B(g23141), .Z(g24925) ) ;
INV     gate13509  (.A(g24925), .Z(II33265) ) ;
INV     gate13510  (.A(g24925), .Z(II33268) ) ;
INV     gate13511  (.A(II33268), .Z(g25443) ) ;
NAND2   gate13512  (.A(g1880), .B(g23394), .Z(g24641) ) ;
INV     gate13513  (.A(g24641), .Z(g25444) ) ;
INV     gate13514  (.A(g24993), .Z(g25445) ) ;
NAND2   gate13515  (.A(g2574), .B(g23402), .Z(g24660) ) ;
INV     gate13516  (.A(g24660), .Z(g25449) ) ;
NAND2   gate13517  (.A(g23950), .B(g679), .Z(g25088) ) ;
INV     gate13518  (.A(g25088), .Z(II33278) ) ;
INV     gate13519  (.A(II33278), .Z(g25454) ) ;
NAND2   gate13520  (.A(g23979), .B(g1365), .Z(g25096) ) ;
INV     gate13521  (.A(g25096), .Z(II33282) ) ;
INV     gate13522  (.A(II33282), .Z(g25458) ) ;
NOR2    gate13523  (.A(g23386), .B(g10024), .Z(g24426) ) ;
INV     gate13524  (.A(g24426), .Z(II33286) ) ;
INV     gate13525  (.A(II33286), .Z(g25462) ) ;
NAND2   gate13526  (.A(g24009), .B(g2059), .Z(g25106) ) ;
INV     gate13527  (.A(g25106), .Z(II33289) ) ;
INV     gate13528  (.A(II33289), .Z(g25463) ) ;
NAND2   gate13529  (.A(g23644), .B(g5438), .Z(g25008) ) ;
INV     gate13530  (.A(g25008), .Z(II33293) ) ;
INV     gate13531  (.A(II33293), .Z(g25467) ) ;
NOR2    gate13532  (.A(g23393), .B(g10133), .Z(g24430) ) ;
INV     gate13533  (.A(g24430), .Z(II33297) ) ;
INV     gate13534  (.A(II33297), .Z(g25471) ) ;
NAND2   gate13535  (.A(g24043), .B(g2753), .Z(g25112) ) ;
INV     gate13536  (.A(g25112), .Z(II33300) ) ;
INV     gate13537  (.A(II33300), .Z(g25472) ) ;
NAND2   gate13538  (.A(g23644), .B(g6448), .Z(g25004) ) ;
INV     gate13539  (.A(g25004), .Z(II33304) ) ;
INV     gate13540  (.A(II33304), .Z(g25476) ) ;
NAND2   gate13541  (.A(g23644), .B(g5438), .Z(g25011) ) ;
INV     gate13542  (.A(g25011), .Z(II33307) ) ;
INV     gate13543  (.A(II33307), .Z(g25479) ) ;
NAND2   gate13544  (.A(g23694), .B(g5473), .Z(g25014) ) ;
INV     gate13545  (.A(g25014), .Z(II33312) ) ;
INV     gate13546  (.A(II33312), .Z(g25484) ) ;
NOR2    gate13547  (.A(g23401), .B(g10238), .Z(g24434) ) ;
INV     gate13548  (.A(g24434), .Z(II33316) ) ;
INV     gate13549  (.A(II33316), .Z(g25488) ) ;
NAND2   gate13550  (.A(g23644), .B(g3306), .Z(g24442) ) ;
INV     gate13551  (.A(g24442), .Z(II33321) ) ;
INV     gate13552  (.A(II33321), .Z(g25493) ) ;
NAND2   gate13553  (.A(g23644), .B(g6448), .Z(g25009) ) ;
INV     gate13554  (.A(g25009), .Z(II33324) ) ;
INV     gate13555  (.A(II33324), .Z(g25496) ) ;
NAND2   gate13556  (.A(g23644), .B(g5438), .Z(g25017) ) ;
INV     gate13557  (.A(g25017), .Z(II33327) ) ;
INV     gate13558  (.A(II33327), .Z(g25499) ) ;
NAND2   gate13559  (.A(g23923), .B(g6486), .Z(g25019) ) ;
INV     gate13560  (.A(g25019), .Z(II33330) ) ;
INV     gate13561  (.A(II33330), .Z(g25502) ) ;
NAND2   gate13562  (.A(g23694), .B(g6713), .Z(g25010) ) ;
INV     gate13563  (.A(g25010), .Z(II33335) ) ;
INV     gate13564  (.A(II33335), .Z(g25507) ) ;
NAND2   gate13565  (.A(g23694), .B(g5473), .Z(g25021) ) ;
INV     gate13566  (.A(g25021), .Z(II33338) ) ;
INV     gate13567  (.A(II33338), .Z(g25510) ) ;
NAND2   gate13568  (.A(g23748), .B(g5512), .Z(g25024) ) ;
INV     gate13569  (.A(g25024), .Z(II33343) ) ;
INV     gate13570  (.A(II33343), .Z(g25515) ) ;
NOR2    gate13571  (.A(g23408), .B(g10340), .Z(g24438) ) ;
INV     gate13572  (.A(g24438), .Z(II33347) ) ;
INV     gate13573  (.A(II33347), .Z(g25519) ) ;
NAND2   gate13574  (.A(g23644), .B(g3306), .Z(g24443) ) ;
INV     gate13575  (.A(g24443), .Z(II33352) ) ;
INV     gate13576  (.A(II33352), .Z(g25524) ) ;
NAND2   gate13577  (.A(g23644), .B(g6448), .Z(g25012) ) ;
INV     gate13578  (.A(g25012), .Z(II33355) ) ;
INV     gate13579  (.A(II33355), .Z(g25527) ) ;
NAND2   gate13580  (.A(g23644), .B(g5438), .Z(g25028) ) ;
INV     gate13581  (.A(g25028), .Z(II33358) ) ;
INV     gate13582  (.A(II33358), .Z(g25530) ) ;
NAND2   gate13583  (.A(g23923), .B(g6643), .Z(g25013) ) ;
INV     gate13584  (.A(g25013), .Z(II33361) ) ;
INV     gate13585  (.A(II33361), .Z(g25533) ) ;
NAND2   gate13586  (.A(g23923), .B(g6486), .Z(g25029) ) ;
INV     gate13587  (.A(g25029), .Z(II33364) ) ;
INV     gate13588  (.A(II33364), .Z(g25536) ) ;
NAND2   gate13589  (.A(g23694), .B(g3462), .Z(g24444) ) ;
INV     gate13590  (.A(g24444), .Z(II33368) ) ;
INV     gate13591  (.A(II33368), .Z(g25540) ) ;
NAND2   gate13592  (.A(g23694), .B(g6713), .Z(g25015) ) ;
INV     gate13593  (.A(g25015), .Z(II33371) ) ;
INV     gate13594  (.A(II33371), .Z(g25543) ) ;
NAND2   gate13595  (.A(g23694), .B(g5473), .Z(g25031) ) ;
INV     gate13596  (.A(g25031), .Z(II33374) ) ;
INV     gate13597  (.A(II33374), .Z(g25546) ) ;
NAND2   gate13598  (.A(g23955), .B(g6751), .Z(g25033) ) ;
INV     gate13599  (.A(g25033), .Z(II33377) ) ;
INV     gate13600  (.A(II33377), .Z(g25549) ) ;
NAND2   gate13601  (.A(g23748), .B(g7015), .Z(g25016) ) ;
INV     gate13602  (.A(g25016), .Z(II33382) ) ;
INV     gate13603  (.A(II33382), .Z(g25554) ) ;
NAND2   gate13604  (.A(g23748), .B(g5512), .Z(g25035) ) ;
INV     gate13605  (.A(g25035), .Z(II33385) ) ;
INV     gate13606  (.A(II33385), .Z(g25557) ) ;
NAND2   gate13607  (.A(g23803), .B(g5556), .Z(g25038) ) ;
INV     gate13608  (.A(g25038), .Z(II33390) ) ;
INV     gate13609  (.A(II33390), .Z(g25562) ) ;
NAND2   gate13610  (.A(g23644), .B(g3306), .Z(g24447) ) ;
INV     gate13611  (.A(g24447), .Z(II33396) ) ;
INV     gate13612  (.A(II33396), .Z(g25573) ) ;
NAND2   gate13613  (.A(g23644), .B(g6448), .Z(g25018) ) ;
INV     gate13614  (.A(g25018), .Z(II33399) ) ;
INV     gate13615  (.A(II33399), .Z(g25576) ) ;
NAND2   gate13616  (.A(g23923), .B(g3338), .Z(g24448) ) ;
INV     gate13617  (.A(g24448), .Z(II33402) ) ;
INV     gate13618  (.A(II33402), .Z(g25579) ) ;
NAND2   gate13619  (.A(g23923), .B(g6643), .Z(g25020) ) ;
INV     gate13620  (.A(g25020), .Z(II33405) ) ;
INV     gate13621  (.A(II33405), .Z(g25582) ) ;
NAND2   gate13622  (.A(g23923), .B(g6486), .Z(g25040) ) ;
INV     gate13623  (.A(g25040), .Z(II33408) ) ;
INV     gate13624  (.A(II33408), .Z(g25585) ) ;
NOR2    gate13625  (.A(g15247), .B(g23735), .Z(g24491) ) ;
INV     gate13626  (.A(g24491), .Z(II33411) ) ;
INV     gate13627  (.A(II33411), .Z(g25588) ) ;
NAND2   gate13628  (.A(g23694), .B(g3462), .Z(g24449) ) ;
INV     gate13629  (.A(g24449), .Z(II33415) ) ;
INV     gate13630  (.A(II33415), .Z(g25590) ) ;
NAND2   gate13631  (.A(g23694), .B(g6713), .Z(g25022) ) ;
INV     gate13632  (.A(g25022), .Z(II33418) ) ;
INV     gate13633  (.A(II33418), .Z(g25593) ) ;
NAND2   gate13634  (.A(g23694), .B(g5473), .Z(g25043) ) ;
INV     gate13635  (.A(g25043), .Z(II33421) ) ;
INV     gate13636  (.A(II33421), .Z(g25596) ) ;
NAND2   gate13637  (.A(g23955), .B(g6945), .Z(g25023) ) ;
INV     gate13638  (.A(g25023), .Z(II33424) ) ;
INV     gate13639  (.A(II33424), .Z(g25599) ) ;
NAND2   gate13640  (.A(g23955), .B(g6751), .Z(g25044) ) ;
INV     gate13641  (.A(g25044), .Z(II33427) ) ;
INV     gate13642  (.A(II33427), .Z(g25602) ) ;
NAND2   gate13643  (.A(g23748), .B(g3618), .Z(g24450) ) ;
INV     gate13644  (.A(g24450), .Z(II33431) ) ;
INV     gate13645  (.A(II33431), .Z(g25606) ) ;
NAND2   gate13646  (.A(g23748), .B(g7015), .Z(g25025) ) ;
INV     gate13647  (.A(g25025), .Z(II33434) ) ;
INV     gate13648  (.A(II33434), .Z(g25609) ) ;
NAND2   gate13649  (.A(g23748), .B(g5512), .Z(g25046) ) ;
INV     gate13650  (.A(g25046), .Z(II33437) ) ;
INV     gate13651  (.A(II33437), .Z(g25612) ) ;
NAND2   gate13652  (.A(g23984), .B(g7053), .Z(g25048) ) ;
INV     gate13653  (.A(g25048), .Z(II33440) ) ;
INV     gate13654  (.A(II33440), .Z(g25615) ) ;
NAND2   gate13655  (.A(g23803), .B(g7265), .Z(g25026) ) ;
INV     gate13656  (.A(g25026), .Z(II33445) ) ;
INV     gate13657  (.A(II33445), .Z(g25620) ) ;
NAND2   gate13658  (.A(g23803), .B(g5556), .Z(g25050) ) ;
INV     gate13659  (.A(g25050), .Z(II33448) ) ;
INV     gate13660  (.A(II33448), .Z(g25623) ) ;
AND3    gate13661  (.A(g23545), .B(g21119), .C(g21227), .Z(g24478) ) ;
INV     gate13662  (.A(g24478), .Z(g25630) ) ;
NAND2   gate13663  (.A(g23644), .B(g3306), .Z(g24451) ) ;
INV     gate13664  (.A(g24451), .Z(II33457) ) ;
INV     gate13665  (.A(II33457), .Z(g25634) ) ;
NAND2   gate13666  (.A(g23923), .B(g3338), .Z(g24452) ) ;
INV     gate13667  (.A(g24452), .Z(II33460) ) ;
INV     gate13668  (.A(II33460), .Z(g25637) ) ;
NAND2   gate13669  (.A(g23923), .B(g6643), .Z(g25030) ) ;
INV     gate13670  (.A(g25030), .Z(II33463) ) ;
INV     gate13671  (.A(II33463), .Z(g25640) ) ;
NAND2   gate13672  (.A(g23923), .B(g6486), .Z(g25053) ) ;
INV     gate13673  (.A(g25053), .Z(II33466) ) ;
INV     gate13674  (.A(II33466), .Z(g25643) ) ;
NOR2    gate13675  (.A(g15324), .B(g23777), .Z(g24498) ) ;
INV     gate13676  (.A(g24498), .Z(II33469) ) ;
INV     gate13677  (.A(II33469), .Z(g25646) ) ;
NOR2    gate13678  (.A(g15325), .B(g23778), .Z(g24499) ) ;
INV     gate13679  (.A(g24499), .Z(II33472) ) ;
INV     gate13680  (.A(II33472), .Z(g25647) ) ;
NAND2   gate13681  (.A(g23694), .B(g3462), .Z(g24453) ) ;
INV     gate13682  (.A(g24453), .Z(II33476) ) ;
INV     gate13683  (.A(II33476), .Z(g25652) ) ;
NAND2   gate13684  (.A(g23694), .B(g6713), .Z(g25032) ) ;
INV     gate13685  (.A(g25032), .Z(II33479) ) ;
INV     gate13686  (.A(II33479), .Z(g25655) ) ;
NAND2   gate13687  (.A(g23955), .B(g3494), .Z(g24454) ) ;
INV     gate13688  (.A(g24454), .Z(II33482) ) ;
INV     gate13689  (.A(II33482), .Z(g25658) ) ;
NAND2   gate13690  (.A(g23955), .B(g6945), .Z(g25034) ) ;
INV     gate13691  (.A(g25034), .Z(II33485) ) ;
INV     gate13692  (.A(II33485), .Z(g25661) ) ;
NAND2   gate13693  (.A(g23955), .B(g6751), .Z(g25054) ) ;
INV     gate13694  (.A(g25054), .Z(II33488) ) ;
INV     gate13695  (.A(II33488), .Z(g25664) ) ;
NOR2    gate13696  (.A(g15339), .B(g23790), .Z(g24501) ) ;
INV     gate13697  (.A(g24501), .Z(II33491) ) ;
INV     gate13698  (.A(II33491), .Z(g25667) ) ;
NAND2   gate13699  (.A(g23748), .B(g3618), .Z(g24455) ) ;
INV     gate13700  (.A(g24455), .Z(II33495) ) ;
INV     gate13701  (.A(II33495), .Z(g25669) ) ;
NAND2   gate13702  (.A(g23748), .B(g7015), .Z(g25036) ) ;
INV     gate13703  (.A(g25036), .Z(II33498) ) ;
INV     gate13704  (.A(II33498), .Z(g25672) ) ;
NAND2   gate13705  (.A(g23748), .B(g5512), .Z(g25057) ) ;
INV     gate13706  (.A(g25057), .Z(II33501) ) ;
INV     gate13707  (.A(II33501), .Z(g25675) ) ;
NAND2   gate13708  (.A(g23984), .B(g7195), .Z(g25037) ) ;
INV     gate13709  (.A(g25037), .Z(II33504) ) ;
INV     gate13710  (.A(II33504), .Z(g25678) ) ;
NAND2   gate13711  (.A(g23984), .B(g7053), .Z(g25058) ) ;
INV     gate13712  (.A(g25058), .Z(II33507) ) ;
INV     gate13713  (.A(II33507), .Z(g25681) ) ;
NAND2   gate13714  (.A(g23803), .B(g3774), .Z(g24456) ) ;
INV     gate13715  (.A(g24456), .Z(II33511) ) ;
INV     gate13716  (.A(II33511), .Z(g25685) ) ;
NAND2   gate13717  (.A(g23803), .B(g7265), .Z(g25039) ) ;
INV     gate13718  (.A(g25039), .Z(II33514) ) ;
INV     gate13719  (.A(II33514), .Z(g25688) ) ;
NAND2   gate13720  (.A(g23803), .B(g5556), .Z(g25060) ) ;
INV     gate13721  (.A(g25060), .Z(II33517) ) ;
INV     gate13722  (.A(II33517), .Z(g25691) ) ;
NAND2   gate13723  (.A(g24014), .B(g7303), .Z(g25062) ) ;
INV     gate13724  (.A(g25062), .Z(II33520) ) ;
INV     gate13725  (.A(II33520), .Z(g25694) ) ;
INV     gate13726  (.A(g24600), .Z(g25698) ) ;
NAND2   gate13727  (.A(g23923), .B(g3338), .Z(g24457) ) ;
INV     gate13728  (.A(g24457), .Z(II33526) ) ;
INV     gate13729  (.A(II33526), .Z(g25700) ) ;
NAND2   gate13730  (.A(g23923), .B(g6643), .Z(g25041) ) ;
INV     gate13731  (.A(g25041), .Z(II33529) ) ;
INV     gate13732  (.A(II33529), .Z(g25703) ) ;
NOR2    gate13733  (.A(g15391), .B(g23824), .Z(g24507) ) ;
INV     gate13734  (.A(g24507), .Z(II33532) ) ;
INV     gate13735  (.A(II33532), .Z(g25706) ) ;
NOR2    gate13736  (.A(g15392), .B(g23825), .Z(g24508) ) ;
INV     gate13737  (.A(g24508), .Z(II33535) ) ;
INV     gate13738  (.A(II33535), .Z(g25707) ) ;
NAND2   gate13739  (.A(g23694), .B(g3462), .Z(g24458) ) ;
INV     gate13740  (.A(g24458), .Z(II33539) ) ;
INV     gate13741  (.A(II33539), .Z(g25711) ) ;
NAND2   gate13742  (.A(g23955), .B(g3494), .Z(g24459) ) ;
INV     gate13743  (.A(g24459), .Z(II33542) ) ;
INV     gate13744  (.A(II33542), .Z(g25714) ) ;
NAND2   gate13745  (.A(g23955), .B(g6945), .Z(g25045) ) ;
INV     gate13746  (.A(g25045), .Z(II33545) ) ;
INV     gate13747  (.A(II33545), .Z(g25717) ) ;
NAND2   gate13748  (.A(g23955), .B(g6751), .Z(g25064) ) ;
INV     gate13749  (.A(g25064), .Z(II33548) ) ;
INV     gate13750  (.A(II33548), .Z(g25720) ) ;
NOR2    gate13751  (.A(g15410), .B(g23830), .Z(g24510) ) ;
INV     gate13752  (.A(g24510), .Z(II33551) ) ;
INV     gate13753  (.A(II33551), .Z(g25723) ) ;
NOR2    gate13754  (.A(g15411), .B(g23831), .Z(g24511) ) ;
INV     gate13755  (.A(g24511), .Z(II33554) ) ;
INV     gate13756  (.A(II33554), .Z(g25724) ) ;
NAND2   gate13757  (.A(g23748), .B(g3618), .Z(g24460) ) ;
INV     gate13758  (.A(g24460), .Z(II33558) ) ;
INV     gate13759  (.A(II33558), .Z(g25729) ) ;
NAND2   gate13760  (.A(g23748), .B(g7015), .Z(g25047) ) ;
INV     gate13761  (.A(g25047), .Z(II33561) ) ;
INV     gate13762  (.A(II33561), .Z(g25732) ) ;
NAND2   gate13763  (.A(g23984), .B(g3650), .Z(g24461) ) ;
INV     gate13764  (.A(g24461), .Z(II33564) ) ;
INV     gate13765  (.A(II33564), .Z(g25735) ) ;
NAND2   gate13766  (.A(g23984), .B(g7195), .Z(g25049) ) ;
INV     gate13767  (.A(g25049), .Z(II33567) ) ;
INV     gate13768  (.A(II33567), .Z(g25738) ) ;
NAND2   gate13769  (.A(g23984), .B(g7053), .Z(g25065) ) ;
INV     gate13770  (.A(g25065), .Z(II33570) ) ;
INV     gate13771  (.A(II33570), .Z(g25741) ) ;
NOR2    gate13772  (.A(g15425), .B(g23843), .Z(g24513) ) ;
INV     gate13773  (.A(g24513), .Z(II33573) ) ;
INV     gate13774  (.A(II33573), .Z(g25744) ) ;
NAND2   gate13775  (.A(g23803), .B(g3774), .Z(g24462) ) ;
INV     gate13776  (.A(g24462), .Z(II33577) ) ;
INV     gate13777  (.A(II33577), .Z(g25746) ) ;
NAND2   gate13778  (.A(g23803), .B(g7265), .Z(g25051) ) ;
INV     gate13779  (.A(g25051), .Z(II33580) ) ;
INV     gate13780  (.A(II33580), .Z(g25749) ) ;
NAND2   gate13781  (.A(g23803), .B(g5556), .Z(g25068) ) ;
INV     gate13782  (.A(g25068), .Z(II33583) ) ;
INV     gate13783  (.A(II33583), .Z(g25752) ) ;
NAND2   gate13784  (.A(g24014), .B(g7391), .Z(g25052) ) ;
INV     gate13785  (.A(g25052), .Z(II33586) ) ;
INV     gate13786  (.A(II33586), .Z(g25755) ) ;
NAND2   gate13787  (.A(g24014), .B(g7303), .Z(g25069) ) ;
INV     gate13788  (.A(g25069), .Z(II33589) ) ;
INV     gate13789  (.A(II33589), .Z(g25758) ) ;
NOR2    gate13790  (.A(g23427), .B(g22777), .Z(g24445) ) ;
INV     gate13791  (.A(g24445), .Z(II33593) ) ;
INV     gate13792  (.A(II33593), .Z(g25762) ) ;
NOR2    gate13793  (.A(g23433), .B(g22907), .Z(g24446) ) ;
INV     gate13794  (.A(g24446), .Z(II33596) ) ;
INV     gate13795  (.A(II33596), .Z(g25763) ) ;
NAND2   gate13796  (.A(g23923), .B(g3338), .Z(g24463) ) ;
INV     gate13797  (.A(g24463), .Z(II33600) ) ;
INV     gate13798  (.A(II33600), .Z(g25767) ) ;
NOR2    gate13799  (.A(g15459), .B(g23855), .Z(g24519) ) ;
INV     gate13800  (.A(g24519), .Z(II33603) ) ;
INV     gate13801  (.A(II33603), .Z(g25770) ) ;
INV     gate13802  (.A(g24607), .Z(g25771) ) ;
NAND2   gate13803  (.A(g23955), .B(g3494), .Z(g24464) ) ;
INV     gate13804  (.A(g24464), .Z(II33608) ) ;
INV     gate13805  (.A(II33608), .Z(g25773) ) ;
NAND2   gate13806  (.A(g23955), .B(g6945), .Z(g25055) ) ;
INV     gate13807  (.A(g25055), .Z(II33611) ) ;
INV     gate13808  (.A(II33611), .Z(g25776) ) ;
NOR2    gate13809  (.A(g15475), .B(g23859), .Z(g24521) ) ;
INV     gate13810  (.A(g24521), .Z(II33614) ) ;
INV     gate13811  (.A(II33614), .Z(g25779) ) ;
NOR2    gate13812  (.A(g15476), .B(g23860), .Z(g24522) ) ;
INV     gate13813  (.A(g24522), .Z(II33617) ) ;
INV     gate13814  (.A(II33617), .Z(g25780) ) ;
NAND2   gate13815  (.A(g23748), .B(g3618), .Z(g24465) ) ;
INV     gate13816  (.A(g24465), .Z(II33621) ) ;
INV     gate13817  (.A(II33621), .Z(g25784) ) ;
NAND2   gate13818  (.A(g23984), .B(g3650), .Z(g24466) ) ;
INV     gate13819  (.A(g24466), .Z(II33624) ) ;
INV     gate13820  (.A(II33624), .Z(g25787) ) ;
NAND2   gate13821  (.A(g23984), .B(g7195), .Z(g25059) ) ;
INV     gate13822  (.A(g25059), .Z(II33627) ) ;
INV     gate13823  (.A(II33627), .Z(g25790) ) ;
NAND2   gate13824  (.A(g23984), .B(g7053), .Z(g25071) ) ;
INV     gate13825  (.A(g25071), .Z(II33630) ) ;
INV     gate13826  (.A(II33630), .Z(g25793) ) ;
NOR2    gate13827  (.A(g15494), .B(g23865), .Z(g24524) ) ;
INV     gate13828  (.A(g24524), .Z(II33633) ) ;
INV     gate13829  (.A(II33633), .Z(g25796) ) ;
NOR2    gate13830  (.A(g15495), .B(g23866), .Z(g24525) ) ;
INV     gate13831  (.A(g24525), .Z(II33636) ) ;
INV     gate13832  (.A(II33636), .Z(g25797) ) ;
NAND2   gate13833  (.A(g23803), .B(g3774), .Z(g24467) ) ;
INV     gate13834  (.A(g24467), .Z(II33640) ) ;
INV     gate13835  (.A(II33640), .Z(g25802) ) ;
NAND2   gate13836  (.A(g23803), .B(g7265), .Z(g25061) ) ;
INV     gate13837  (.A(g25061), .Z(II33643) ) ;
INV     gate13838  (.A(II33643), .Z(g25805) ) ;
NAND2   gate13839  (.A(g24014), .B(g3806), .Z(g24468) ) ;
INV     gate13840  (.A(g24468), .Z(II33646) ) ;
INV     gate13841  (.A(II33646), .Z(g25808) ) ;
NAND2   gate13842  (.A(g24014), .B(g7391), .Z(g25063) ) ;
INV     gate13843  (.A(g25063), .Z(II33649) ) ;
INV     gate13844  (.A(II33649), .Z(g25811) ) ;
NAND2   gate13845  (.A(g24014), .B(g7303), .Z(g25072) ) ;
INV     gate13846  (.A(g25072), .Z(II33652) ) ;
INV     gate13847  (.A(II33652), .Z(g25814) ) ;
NOR2    gate13848  (.A(g15509), .B(g23878), .Z(g24527) ) ;
INV     gate13849  (.A(g24527), .Z(II33655) ) ;
INV     gate13850  (.A(II33655), .Z(g25817) ) ;
NAND2   gate13851  (.A(g23955), .B(g3494), .Z(g24469) ) ;
INV     gate13852  (.A(g24469), .Z(II33659) ) ;
INV     gate13853  (.A(II33659), .Z(g25821) ) ;
NOR2    gate13854  (.A(g15545), .B(g23889), .Z(g24532) ) ;
INV     gate13855  (.A(g24532), .Z(II33662) ) ;
INV     gate13856  (.A(II33662), .Z(g25824) ) ;
INV     gate13857  (.A(g24619), .Z(g25825) ) ;
NAND2   gate13858  (.A(g23984), .B(g3650), .Z(g24470) ) ;
INV     gate13859  (.A(g24470), .Z(II33667) ) ;
INV     gate13860  (.A(II33667), .Z(g25827) ) ;
NAND2   gate13861  (.A(g23984), .B(g7195), .Z(g25066) ) ;
INV     gate13862  (.A(g25066), .Z(II33670) ) ;
INV     gate13863  (.A(II33670), .Z(g25830) ) ;
NOR2    gate13864  (.A(g15561), .B(g23893), .Z(g24534) ) ;
INV     gate13865  (.A(g24534), .Z(II33673) ) ;
INV     gate13866  (.A(II33673), .Z(g25833) ) ;
NOR2    gate13867  (.A(g15562), .B(g23894), .Z(g24535) ) ;
INV     gate13868  (.A(g24535), .Z(II33676) ) ;
INV     gate13869  (.A(II33676), .Z(g25834) ) ;
NAND2   gate13870  (.A(g23803), .B(g3774), .Z(g24471) ) ;
INV     gate13871  (.A(g24471), .Z(II33680) ) ;
INV     gate13872  (.A(II33680), .Z(g25838) ) ;
NAND2   gate13873  (.A(g24014), .B(g3806), .Z(g24472) ) ;
INV     gate13874  (.A(g24472), .Z(II33683) ) ;
INV     gate13875  (.A(II33683), .Z(g25841) ) ;
NAND2   gate13876  (.A(g24014), .B(g7391), .Z(g25070) ) ;
INV     gate13877  (.A(g25070), .Z(II33686) ) ;
INV     gate13878  (.A(II33686), .Z(g25844) ) ;
NAND2   gate13879  (.A(g24014), .B(g7303), .Z(g25074) ) ;
INV     gate13880  (.A(g25074), .Z(II33689) ) ;
INV     gate13881  (.A(II33689), .Z(g25847) ) ;
NOR2    gate13882  (.A(g15580), .B(g23899), .Z(g24537) ) ;
INV     gate13883  (.A(g24537), .Z(II33692) ) ;
INV     gate13884  (.A(II33692), .Z(g25850) ) ;
NOR2    gate13885  (.A(g15581), .B(g23900), .Z(g24538) ) ;
INV     gate13886  (.A(g24538), .Z(II33695) ) ;
INV     gate13887  (.A(II33695), .Z(g25851) ) ;
NAND2   gate13888  (.A(g23984), .B(g3650), .Z(g24474) ) ;
INV     gate13889  (.A(g24474), .Z(II33700) ) ;
INV     gate13890  (.A(II33700), .Z(g25856) ) ;
NOR2    gate13891  (.A(g15623), .B(g23910), .Z(g24545) ) ;
INV     gate13892  (.A(g24545), .Z(II33703) ) ;
INV     gate13893  (.A(II33703), .Z(g25859) ) ;
INV     gate13894  (.A(g24630), .Z(g25860) ) ;
NAND2   gate13895  (.A(g24014), .B(g3806), .Z(g24475) ) ;
INV     gate13896  (.A(g24475), .Z(II33708) ) ;
INV     gate13897  (.A(II33708), .Z(g25862) ) ;
NAND2   gate13898  (.A(g24014), .B(g7391), .Z(g25073) ) ;
INV     gate13899  (.A(g25073), .Z(II33711) ) ;
INV     gate13900  (.A(II33711), .Z(g25865) ) ;
NOR2    gate13901  (.A(g15639), .B(g23914), .Z(g24547) ) ;
INV     gate13902  (.A(g24547), .Z(II33714) ) ;
INV     gate13903  (.A(II33714), .Z(g25868) ) ;
NOR2    gate13904  (.A(g15640), .B(g23915), .Z(g24548) ) ;
INV     gate13905  (.A(g24548), .Z(II33717) ) ;
INV     gate13906  (.A(II33717), .Z(g25869) ) ;
NAND2   gate13907  (.A(g24014), .B(g3806), .Z(g24477) ) ;
INV     gate13908  (.A(g24477), .Z(II33723) ) ;
INV     gate13909  (.A(II33723), .Z(g25877) ) ;
NOR2    gate13910  (.A(g15699), .B(g23942), .Z(g24557) ) ;
INV     gate13911  (.A(g24557), .Z(II33726) ) ;
INV     gate13912  (.A(II33726), .Z(g25880) ) ;
NOR2    gate13913  (.A(g23461), .B(g18407), .Z(g24473) ) ;
INV     gate13914  (.A(g24473), .Z(II33732) ) ;
INV     gate13915  (.A(II33732), .Z(g25886) ) ;
NOR2    gate13916  (.A(g23477), .B(g20127), .Z(g24476) ) ;
INV     gate13917  (.A(g24476), .Z(II33737) ) ;
INV     gate13918  (.A(II33737), .Z(g25891) ) ;
INV     gate13919  (.A(g24939), .Z(g25895) ) ;
NAND2   gate13920  (.A(II32678), .B(II32679), .Z(g24928) ) ;
INV     gate13921  (.A(g24928), .Z(g25899) ) ;
INV     gate13922  (.A(g24950), .Z(g25903) ) ;
NAND2   gate13923  (.A(II32696), .B(II32697), .Z(g24940) ) ;
INV     gate13924  (.A(g24940), .Z(g25907) ) ;
INV     gate13925  (.A(g24962), .Z(g25911) ) ;
NAND2   gate13926  (.A(II32709), .B(II32710), .Z(g24951) ) ;
INV     gate13927  (.A(g24951), .Z(g25915) ) ;
INV     gate13928  (.A(g24973), .Z(g25919) ) ;
NAND2   gate13929  (.A(II32725), .B(II32726), .Z(g24963) ) ;
INV     gate13930  (.A(g24963), .Z(g25923) ) ;
INV     gate13931  (.A(g24763), .Z(g25937) ) ;
INV     gate13932  (.A(g24784), .Z(g25939) ) ;
INV     gate13933  (.A(g24805), .Z(g25942) ) ;
INV     gate13934  (.A(g24827), .Z(g25945) ) ;
INV     gate13935  (.A(g24735), .Z(g25952) ) ;
INV     gate13936  (.A(g25103), .Z(II33790) ) ;
INV     gate13937  (.A(II33790), .Z(g25976) ) ;
INV     gate13938  (.A(g25109), .Z(II33798) ) ;
INV     gate13939  (.A(II33798), .Z(g25982) ) ;
INV     gate13940  (.A(g25327), .Z(II33801) ) ;
INV     gate13941  (.A(g25976), .Z(II33804) ) ;
INV     gate13942  (.A(g25588), .Z(II33807) ) ;
INV     gate13943  (.A(g25646), .Z(II33810) ) ;
INV     gate13944  (.A(g25706), .Z(II33813) ) ;
INV     gate13945  (.A(g25647), .Z(II33816) ) ;
INV     gate13946  (.A(g25707), .Z(II33819) ) ;
INV     gate13947  (.A(g25770), .Z(II33822) ) ;
INV     gate13948  (.A(g25462), .Z(II33825) ) ;
INV     gate13949  (.A(g25336), .Z(II33828) ) ;
INV     gate13950  (.A(g25982), .Z(II33831) ) ;
INV     gate13951  (.A(g25667), .Z(II33834) ) ;
INV     gate13952  (.A(g25723), .Z(II33837) ) ;
INV     gate13953  (.A(g25779), .Z(II33840) ) ;
INV     gate13954  (.A(g25724), .Z(II33843) ) ;
INV     gate13955  (.A(g25780), .Z(II33846) ) ;
INV     gate13956  (.A(g25824), .Z(II33849) ) ;
INV     gate13957  (.A(g25471), .Z(II33852) ) ;
INV     gate13958  (.A(g25350), .Z(II33855) ) ;
INV     gate13959  (.A(g25179), .Z(II33858) ) ;
INV     gate13960  (.A(g25744), .Z(II33861) ) ;
INV     gate13961  (.A(g25796), .Z(II33864) ) ;
INV     gate13962  (.A(g25833), .Z(II33867) ) ;
INV     gate13963  (.A(g25797), .Z(II33870) ) ;
INV     gate13964  (.A(g25834), .Z(II33873) ) ;
INV     gate13965  (.A(g25859), .Z(II33876) ) ;
INV     gate13966  (.A(g25488), .Z(II33879) ) ;
INV     gate13967  (.A(g25364), .Z(II33882) ) ;
INV     gate13968  (.A(g25180), .Z(II33885) ) ;
INV     gate13969  (.A(g25817), .Z(II33888) ) ;
INV     gate13970  (.A(g25850), .Z(II33891) ) ;
INV     gate13971  (.A(g25868), .Z(II33894) ) ;
INV     gate13972  (.A(g25851), .Z(II33897) ) ;
INV     gate13973  (.A(g25869), .Z(II33900) ) ;
INV     gate13974  (.A(g25880), .Z(II33903) ) ;
INV     gate13975  (.A(g25519), .Z(II33906) ) ;
INV     gate13976  (.A(g25886), .Z(II33909) ) ;
INV     gate13977  (.A(g25891), .Z(II33912) ) ;
INV     gate13978  (.A(g25762), .Z(II33915) ) ;
INV     gate13979  (.A(g25763), .Z(II33918) ) ;
NOR2    gate13980  (.A(g24975), .B(g5623), .Z(g25343) ) ;
INV     gate13981  (.A(g25343), .Z(II33954) ) ;
INV     gate13982  (.A(II33954), .Z(g26056) ) ;
NOR2    gate13983  (.A(g24986), .B(g5651), .Z(g25357) ) ;
INV     gate13984  (.A(g25357), .Z(II33961) ) ;
INV     gate13985  (.A(II33961), .Z(g26063) ) ;
NOR2    gate13986  (.A(g24997), .B(g5689), .Z(g25372) ) ;
INV     gate13987  (.A(g25372), .Z(II33968) ) ;
INV     gate13988  (.A(II33968), .Z(g26070) ) ;
NOR2    gate13989  (.A(g25005), .B(g5741), .Z(g25389) ) ;
INV     gate13990  (.A(g25389), .Z(II33974) ) ;
INV     gate13991  (.A(II33974), .Z(g26076) ) ;
NOR2    gate13992  (.A(g25125), .B(g17001), .Z(g25932) ) ;
INV     gate13993  (.A(g25932), .Z(II33984) ) ;
INV     gate13994  (.A(II33984), .Z(g26086) ) ;
NOR4    gate13995  (.A(g4456), .B(g25078), .C(g18429), .D(g16075), .Z(g25870) ) ;
INV     gate13996  (.A(g25870), .Z(II33990) ) ;
INV     gate13997  (.A(II33990), .Z(g26092) ) ;
NOR2    gate13998  (.A(g25127), .B(g17031), .Z(g25935) ) ;
INV     gate13999  (.A(g25935), .Z(II33995) ) ;
INV     gate14000  (.A(II33995), .Z(g26102) ) ;
OR2     gate14001  (.A(g24759), .B(g23146), .Z(g25490) ) ;
INV     gate14002  (.A(g25490), .Z(II33999) ) ;
INV     gate14003  (.A(g25490), .Z(II34002) ) ;
INV     gate14004  (.A(II34002), .Z(g26105) ) ;
NOR4    gate14005  (.A(g4632), .B(g25082), .C(g18502), .D(g16113), .Z(g25882) ) ;
INV     gate14006  (.A(g25882), .Z(II34009) ) ;
INV     gate14007  (.A(II34009), .Z(g26114) ) ;
NOR2    gate14008  (.A(g25129), .B(g17065), .Z(g25938) ) ;
INV     gate14009  (.A(g25938), .Z(II34012) ) ;
INV     gate14010  (.A(II34012), .Z(g26118) ) ;
NOR4    gate14011  (.A(g4809), .B(g25091), .C(g18566), .D(g16164), .Z(g25887) ) ;
INV     gate14012  (.A(g25887), .Z(II34017) ) ;
INV     gate14013  (.A(II34017), .Z(g26121) ) ;
NOR2    gate14014  (.A(g24428), .B(g17100), .Z(g25940) ) ;
INV     gate14015  (.A(g25940), .Z(II34020) ) ;
INV     gate14016  (.A(II34020), .Z(g26125) ) ;
NOR4    gate14017  (.A(g4985), .B(g25099), .C(g18616), .D(g16223), .Z(g25892) ) ;
INV     gate14018  (.A(g25892), .Z(II34026) ) ;
INV     gate14019  (.A(II34026), .Z(g26131) ) ;
OR2     gate14020  (.A(g24813), .B(g23145), .Z(g25520) ) ;
INV     gate14021  (.A(g25520), .Z(II34029) ) ;
INV     gate14022  (.A(g25520), .Z(II34032) ) ;
INV     gate14023  (.A(II34032), .Z(g26136) ) ;
OR2     gate14024  (.A(g24843), .B(g23143), .Z(g25566) ) ;
INV     gate14025  (.A(g25566), .Z(II34041) ) ;
INV     gate14026  (.A(g25566), .Z(II34044) ) ;
INV     gate14027  (.A(II34044), .Z(g26150) ) ;
NOR2    gate14028  (.A(g24745), .B(g23547), .Z(g25204) ) ;
INV     gate14029  (.A(g25204), .Z(II34051) ) ;
INV     gate14030  (.A(II34051), .Z(g26159) ) ;
NOR2    gate14031  (.A(g24746), .B(g23550), .Z(g25206) ) ;
INV     gate14032  (.A(g25206), .Z(II34056) ) ;
INV     gate14033  (.A(II34056), .Z(g26164) ) ;
NOR2    gate14034  (.A(g24747), .B(g23551), .Z(g25207) ) ;
INV     gate14035  (.A(g25207), .Z(II34059) ) ;
INV     gate14036  (.A(II34059), .Z(g26165) ) ;
NOR2    gate14037  (.A(g24749), .B(g23554), .Z(g25209) ) ;
INV     gate14038  (.A(g25209), .Z(II34063) ) ;
INV     gate14039  (.A(II34063), .Z(g26167) ) ;
NOR2    gate14040  (.A(g24750), .B(g23558), .Z(g25211) ) ;
INV     gate14041  (.A(g25211), .Z(II34068) ) ;
INV     gate14042  (.A(II34068), .Z(g26172) ) ;
NOR2    gate14043  (.A(g24751), .B(g23559), .Z(g25212) ) ;
INV     gate14044  (.A(g25212), .Z(II34071) ) ;
INV     gate14045  (.A(II34071), .Z(g26173) ) ;
NOR2    gate14046  (.A(g24752), .B(g23560), .Z(g25213) ) ;
INV     gate14047  (.A(g25213), .Z(II34074) ) ;
INV     gate14048  (.A(II34074), .Z(g26174) ) ;
NAND2   gate14049  (.A(g22806), .B(g24517), .Z(g25954) ) ;
INV     gate14050  (.A(g25954), .Z(II34077) ) ;
INV     gate14051  (.A(II34077), .Z(g26175) ) ;
NOR2    gate14052  (.A(g25088), .B(g6157), .Z(g25539) ) ;
INV     gate14053  (.A(g25539), .Z(II34080) ) ;
INV     gate14054  (.A(II34080), .Z(g26178) ) ;
NOR2    gate14055  (.A(g24754), .B(g23563), .Z(g25214) ) ;
INV     gate14056  (.A(g25214), .Z(II34083) ) ;
INV     gate14057  (.A(II34083), .Z(g26181) ) ;
NOR2    gate14058  (.A(g24755), .B(g23564), .Z(g25215) ) ;
INV     gate14059  (.A(g25215), .Z(II34086) ) ;
INV     gate14060  (.A(II34086), .Z(g26182) ) ;
NOR2    gate14061  (.A(g24758), .B(g23567), .Z(g25217) ) ;
INV     gate14062  (.A(g25217), .Z(II34091) ) ;
INV     gate14063  (.A(II34091), .Z(g26187) ) ;
INV     gate14064  (.A(g25952), .Z(g26189) ) ;
NOR2    gate14065  (.A(g24760), .B(g23571), .Z(g25218) ) ;
INV     gate14066  (.A(g25218), .Z(II34096) ) ;
INV     gate14067  (.A(II34096), .Z(g26190) ) ;
NOR2    gate14068  (.A(g24761), .B(g23572), .Z(g25219) ) ;
INV     gate14069  (.A(g25219), .Z(II34099) ) ;
INV     gate14070  (.A(II34099), .Z(g26191) ) ;
NOR2    gate14071  (.A(g24762), .B(g23573), .Z(g25220) ) ;
INV     gate14072  (.A(g25220), .Z(II34102) ) ;
INV     gate14073  (.A(II34102), .Z(g26192) ) ;
NOR2    gate14074  (.A(g24767), .B(g23577), .Z(g25221) ) ;
INV     gate14075  (.A(g25221), .Z(II34105) ) ;
INV     gate14076  (.A(II34105), .Z(g26193) ) ;
NOR2    gate14077  (.A(g24768), .B(g23578), .Z(g25222) ) ;
INV     gate14078  (.A(g25222), .Z(II34108) ) ;
INV     gate14079  (.A(II34108), .Z(g26194) ) ;
NOR2    gate14080  (.A(g24769), .B(g23579), .Z(g25223) ) ;
INV     gate14081  (.A(g25223), .Z(II34111) ) ;
INV     gate14082  (.A(II34111), .Z(g26195) ) ;
NAND2   gate14083  (.A(g22847), .B(g24530), .Z(g25958) ) ;
INV     gate14084  (.A(g25958), .Z(II34114) ) ;
INV     gate14085  (.A(II34114), .Z(g26196) ) ;
NOR2    gate14086  (.A(g25096), .B(g6184), .Z(g25605) ) ;
INV     gate14087  (.A(g25605), .Z(II34118) ) ;
INV     gate14088  (.A(II34118), .Z(g26202) ) ;
NOR2    gate14089  (.A(g24772), .B(g23582), .Z(g25224) ) ;
INV     gate14090  (.A(g25224), .Z(II34121) ) ;
INV     gate14091  (.A(II34121), .Z(g26205) ) ;
NOR2    gate14092  (.A(g24773), .B(g23583), .Z(g25225) ) ;
INV     gate14093  (.A(g25225), .Z(II34124) ) ;
INV     gate14094  (.A(II34124), .Z(g26206) ) ;
NOR2    gate14095  (.A(g24775), .B(g23586), .Z(g25227) ) ;
INV     gate14096  (.A(g25227), .Z(II34128) ) ;
INV     gate14097  (.A(II34128), .Z(g26208) ) ;
INV     gate14098  (.A(g25296), .Z(g26209) ) ;
NOR2    gate14099  (.A(g24776), .B(g23590), .Z(g25228) ) ;
INV     gate14100  (.A(g25228), .Z(II34132) ) ;
INV     gate14101  (.A(II34132), .Z(g26210) ) ;
NOR2    gate14102  (.A(g24777), .B(g23591), .Z(g25229) ) ;
INV     gate14103  (.A(g25229), .Z(II34135) ) ;
INV     gate14104  (.A(II34135), .Z(g26211) ) ;
NOR2    gate14105  (.A(g24779), .B(g23598), .Z(g25230) ) ;
INV     gate14106  (.A(g25230), .Z(II34140) ) ;
INV     gate14107  (.A(II34140), .Z(g26214) ) ;
NOR2    gate14108  (.A(g24780), .B(g23599), .Z(g25231) ) ;
INV     gate14109  (.A(g25231), .Z(II34143) ) ;
INV     gate14110  (.A(II34143), .Z(g26215) ) ;
NOR2    gate14111  (.A(g24781), .B(g23600), .Z(g25232) ) ;
INV     gate14112  (.A(g25232), .Z(II34146) ) ;
INV     gate14113  (.A(II34146), .Z(g26216) ) ;
NOR2    gate14114  (.A(g24788), .B(g23604), .Z(g25233) ) ;
INV     gate14115  (.A(g25233), .Z(II34150) ) ;
INV     gate14116  (.A(II34150), .Z(g26220) ) ;
NOR2    gate14117  (.A(g24789), .B(g23605), .Z(g25234) ) ;
INV     gate14118  (.A(g25234), .Z(II34153) ) ;
INV     gate14119  (.A(II34153), .Z(g26221) ) ;
NOR2    gate14120  (.A(g24790), .B(g23606), .Z(g25235) ) ;
INV     gate14121  (.A(g25235), .Z(II34156) ) ;
INV     gate14122  (.A(II34156), .Z(g26222) ) ;
NAND2   gate14123  (.A(g22882), .B(g24543), .Z(g25964) ) ;
INV     gate14124  (.A(g25964), .Z(II34159) ) ;
INV     gate14125  (.A(II34159), .Z(g26223) ) ;
NOR2    gate14126  (.A(g25106), .B(g6216), .Z(g25684) ) ;
INV     gate14127  (.A(g25684), .Z(II34162) ) ;
INV     gate14128  (.A(II34162), .Z(g26226) ) ;
NOR2    gate14129  (.A(g24792), .B(g23609), .Z(g25236) ) ;
INV     gate14130  (.A(g25236), .Z(II34165) ) ;
INV     gate14131  (.A(II34165), .Z(g26229) ) ;
NOR2    gate14132  (.A(g24793), .B(g23610), .Z(g25237) ) ;
INV     gate14133  (.A(g25237), .Z(II34168) ) ;
INV     gate14134  (.A(II34168), .Z(g26230) ) ;
NOR2    gate14135  (.A(g24796), .B(g23615), .Z(g25239) ) ;
INV     gate14136  (.A(g25239), .Z(II34172) ) ;
INV     gate14137  (.A(II34172), .Z(g26232) ) ;
INV     gate14138  (.A(g25306), .Z(g26237) ) ;
NOR2    gate14139  (.A(g24798), .B(g23622), .Z(g25240) ) ;
INV     gate14140  (.A(g25240), .Z(II34180) ) ;
INV     gate14141  (.A(II34180), .Z(g26238) ) ;
NOR2    gate14142  (.A(g24799), .B(g23623), .Z(g25241) ) ;
INV     gate14143  (.A(g25241), .Z(II34183) ) ;
INV     gate14144  (.A(II34183), .Z(g26239) ) ;
NOR2    gate14145  (.A(g24802), .B(g23630), .Z(g25242) ) ;
INV     gate14146  (.A(g25242), .Z(II34189) ) ;
INV     gate14147  (.A(II34189), .Z(g26245) ) ;
NOR2    gate14148  (.A(g24803), .B(g23631), .Z(g25243) ) ;
INV     gate14149  (.A(g25243), .Z(II34192) ) ;
INV     gate14150  (.A(II34192), .Z(g26246) ) ;
NOR2    gate14151  (.A(g24804), .B(g23632), .Z(g25244) ) ;
INV     gate14152  (.A(g25244), .Z(II34195) ) ;
INV     gate14153  (.A(II34195), .Z(g26247) ) ;
NOR2    gate14154  (.A(g24809), .B(g23636), .Z(g25245) ) ;
INV     gate14155  (.A(g25245), .Z(II34198) ) ;
INV     gate14156  (.A(II34198), .Z(g26248) ) ;
NOR2    gate14157  (.A(g24810), .B(g23637), .Z(g25246) ) ;
INV     gate14158  (.A(g25246), .Z(II34201) ) ;
INV     gate14159  (.A(II34201), .Z(g26249) ) ;
NOR2    gate14160  (.A(g24811), .B(g23638), .Z(g25247) ) ;
INV     gate14161  (.A(g25247), .Z(II34204) ) ;
INV     gate14162  (.A(II34204), .Z(g26250) ) ;
NAND2   gate14163  (.A(g22917), .B(g24555), .Z(g25969) ) ;
INV     gate14164  (.A(g25969), .Z(II34207) ) ;
INV     gate14165  (.A(II34207), .Z(g26251) ) ;
NOR2    gate14166  (.A(g25112), .B(g6305), .Z(g25761) ) ;
INV     gate14167  (.A(g25761), .Z(II34210) ) ;
INV     gate14168  (.A(II34210), .Z(g26254) ) ;
NOR2    gate14169  (.A(g24818), .B(g23664), .Z(g25248) ) ;
INV     gate14170  (.A(g25248), .Z(II34220) ) ;
INV     gate14171  (.A(II34220), .Z(g26264) ) ;
INV     gate14172  (.A(g25315), .Z(g26275) ) ;
NOR2    gate14173  (.A(g24821), .B(g23671), .Z(g25249) ) ;
INV     gate14174  (.A(g25249), .Z(II34230) ) ;
INV     gate14175  (.A(II34230), .Z(g26276) ) ;
NOR2    gate14176  (.A(g24822), .B(g23672), .Z(g25250) ) ;
INV     gate14177  (.A(g25250), .Z(II34233) ) ;
INV     gate14178  (.A(II34233), .Z(g26277) ) ;
NOR2    gate14179  (.A(g24824), .B(g23679), .Z(g25251) ) ;
INV     gate14180  (.A(g25251), .Z(II34238) ) ;
INV     gate14181  (.A(II34238), .Z(g26280) ) ;
NOR2    gate14182  (.A(g24825), .B(g23680), .Z(g25252) ) ;
INV     gate14183  (.A(g25252), .Z(II34241) ) ;
INV     gate14184  (.A(II34241), .Z(g26281) ) ;
NOR2    gate14185  (.A(g24826), .B(g23681), .Z(g25253) ) ;
INV     gate14186  (.A(g25253), .Z(II34244) ) ;
INV     gate14187  (.A(II34244), .Z(g26282) ) ;
NOR2    gate14188  (.A(g24492), .B(g10024), .Z(g25185) ) ;
INV     gate14189  (.A(g25185), .Z(II34254) ) ;
INV     gate14190  (.A(II34254), .Z(g26294) ) ;
NOR2    gate14191  (.A(g24838), .B(g23714), .Z(g25255) ) ;
INV     gate14192  (.A(g25255), .Z(II34266) ) ;
INV     gate14193  (.A(II34266), .Z(g26308) ) ;
INV     gate14194  (.A(g25324), .Z(g26313) ) ;
NOR2    gate14195  (.A(g24840), .B(g23721), .Z(g25256) ) ;
INV     gate14196  (.A(g25256), .Z(II34274) ) ;
INV     gate14197  (.A(II34274), .Z(g26314) ) ;
NOR2    gate14198  (.A(g24841), .B(g23722), .Z(g25257) ) ;
INV     gate14199  (.A(g25257), .Z(II34277) ) ;
INV     gate14200  (.A(II34277), .Z(g26315) ) ;
NOR2    gate14201  (.A(g24502), .B(g10133), .Z(g25189) ) ;
INV     gate14202  (.A(g25189), .Z(II34296) ) ;
INV     gate14203  (.A(II34296), .Z(g26341) ) ;
NOR2    gate14204  (.A(g24853), .B(g23768), .Z(g25259) ) ;
INV     gate14205  (.A(g25259), .Z(II34306) ) ;
INV     gate14206  (.A(II34306), .Z(g26349) ) ;
NOR2    gate14207  (.A(g24878), .B(g23852), .Z(g25265) ) ;
INV     gate14208  (.A(g25265), .Z(II34313) ) ;
INV     gate14209  (.A(II34313), .Z(g26354) ) ;
NOR2    gate14210  (.A(g24516), .B(g22777), .Z(g25191) ) ;
INV     gate14211  (.A(g25191), .Z(II34316) ) ;
INV     gate14212  (.A(II34316), .Z(g26355) ) ;
NAND2   gate14213  (.A(g24965), .B(g5438), .Z(g25928) ) ;
INV     gate14214  (.A(g25928), .Z(II34321) ) ;
INV     gate14215  (.A(II34321), .Z(g26358) ) ;
NOR2    gate14216  (.A(g24858), .B(g17737), .Z(g25260) ) ;
INV     gate14217  (.A(g25260), .Z(II34327) ) ;
INV     gate14218  (.A(II34327), .Z(g26364) ) ;
NOR2    gate14219  (.A(g24514), .B(g10238), .Z(g25194) ) ;
INV     gate14220  (.A(g25194), .Z(II34343) ) ;
INV     gate14221  (.A(II34343), .Z(g26385) ) ;
NAND2   gate14222  (.A(g24965), .B(g6448), .Z(g25927) ) ;
INV     gate14223  (.A(g25927), .Z(II34353) ) ;
INV     gate14224  (.A(II34353), .Z(g26393) ) ;
NOR2    gate14225  (.A(g24869), .B(g17824), .Z(g25262) ) ;
INV     gate14226  (.A(g25262), .Z(II34358) ) ;
INV     gate14227  (.A(II34358), .Z(g26398) ) ;
NAND2   gate14228  (.A(g24978), .B(g5473), .Z(g25930) ) ;
INV     gate14229  (.A(g25930), .Z(II34363) ) ;
INV     gate14230  (.A(II34363), .Z(g26401) ) ;
NOR2    gate14231  (.A(g24874), .B(g17838), .Z(g25263) ) ;
INV     gate14232  (.A(g25263), .Z(II34369) ) ;
INV     gate14233  (.A(II34369), .Z(g26407) ) ;
NOR2    gate14234  (.A(g24528), .B(g10340), .Z(g25197) ) ;
INV     gate14235  (.A(g25197), .Z(II34385) ) ;
INV     gate14236  (.A(II34385), .Z(g26428) ) ;
NAND2   gate14237  (.A(g24965), .B(g3306), .Z(g25200) ) ;
INV     gate14238  (.A(g25200), .Z(II34388) ) ;
INV     gate14239  (.A(II34388), .Z(g26429) ) ;
NOR2    gate14240  (.A(g24881), .B(g17912), .Z(g25266) ) ;
INV     gate14241  (.A(g25266), .Z(II34392) ) ;
INV     gate14242  (.A(II34392), .Z(g26433) ) ;
NAND2   gate14243  (.A(g24978), .B(g6713), .Z(g25929) ) ;
INV     gate14244  (.A(g25929), .Z(II34395) ) ;
INV     gate14245  (.A(II34395), .Z(g26434) ) ;
NOR2    gate14246  (.A(g24884), .B(g17936), .Z(g25267) ) ;
INV     gate14247  (.A(g25267), .Z(II34400) ) ;
INV     gate14248  (.A(II34400), .Z(g26439) ) ;
NAND2   gate14249  (.A(g24989), .B(g5512), .Z(g25933) ) ;
INV     gate14250  (.A(g25933), .Z(II34405) ) ;
INV     gate14251  (.A(II34405), .Z(g26442) ) ;
NOR2    gate14252  (.A(g24888), .B(g17950), .Z(g25268) ) ;
INV     gate14253  (.A(g25268), .Z(II34411) ) ;
INV     gate14254  (.A(II34411), .Z(g26448) ) ;
NAND2   gate14255  (.A(g24978), .B(g3462), .Z(g25203) ) ;
INV     gate14256  (.A(g25203), .Z(II34421) ) ;
INV     gate14257  (.A(II34421), .Z(g26461) ) ;
NOR2    gate14258  (.A(g24898), .B(g18023), .Z(g25270) ) ;
INV     gate14259  (.A(g25270), .Z(II34425) ) ;
INV     gate14260  (.A(II34425), .Z(g26465) ) ;
NAND2   gate14261  (.A(g24989), .B(g7015), .Z(g25931) ) ;
INV     gate14262  (.A(g25931), .Z(II34428) ) ;
INV     gate14263  (.A(II34428), .Z(g26466) ) ;
NOR2    gate14264  (.A(g24901), .B(g18047), .Z(g25271) ) ;
INV     gate14265  (.A(g25271), .Z(II34433) ) ;
INV     gate14266  (.A(II34433), .Z(g26471) ) ;
NAND2   gate14267  (.A(g25000), .B(g5556), .Z(g25936) ) ;
INV     gate14268  (.A(g25936), .Z(II34438) ) ;
INV     gate14269  (.A(II34438), .Z(g26474) ) ;
NOR2    gate14270  (.A(g24905), .B(g18061), .Z(g25272) ) ;
INV     gate14271  (.A(g25272), .Z(II34444) ) ;
INV     gate14272  (.A(II34444), .Z(g26480) ) ;
NOR2    gate14273  (.A(g25076), .B(g21615), .Z(g25764) ) ;
INV     gate14274  (.A(g25764), .Z(g26481) ) ;
NAND2   gate14275  (.A(g24989), .B(g3618), .Z(g25205) ) ;
INV     gate14276  (.A(g25205), .Z(II34449) ) ;
INV     gate14277  (.A(II34449), .Z(g26485) ) ;
NOR2    gate14278  (.A(g24921), .B(g18140), .Z(g25279) ) ;
INV     gate14279  (.A(g25279), .Z(II34453) ) ;
INV     gate14280  (.A(II34453), .Z(g26489) ) ;
NAND2   gate14281  (.A(g25000), .B(g7265), .Z(g25934) ) ;
INV     gate14282  (.A(g25934), .Z(II34456) ) ;
INV     gate14283  (.A(II34456), .Z(g26490) ) ;
NOR2    gate14284  (.A(g24924), .B(g18164), .Z(g25280) ) ;
INV     gate14285  (.A(g25280), .Z(II34461) ) ;
INV     gate14286  (.A(II34461), .Z(g26495) ) ;
NOR2    gate14287  (.A(g24558), .B(g20127), .Z(g25199) ) ;
INV     gate14288  (.A(g25199), .Z(II34464) ) ;
INV     gate14289  (.A(II34464), .Z(g26496) ) ;
NOR2    gate14290  (.A(g25077), .B(g21643), .Z(g25818) ) ;
INV     gate14291  (.A(g25818), .Z(g26497) ) ;
NAND2   gate14292  (.A(g25000), .B(g3774), .Z(g25210) ) ;
INV     gate14293  (.A(g25210), .Z(II34469) ) ;
INV     gate14294  (.A(II34469), .Z(g26501) ) ;
NOR2    gate14295  (.A(g24938), .B(g18256), .Z(g25288) ) ;
INV     gate14296  (.A(g25288), .Z(II34473) ) ;
INV     gate14297  (.A(II34473), .Z(g26505) ) ;
NOR2    gate14298  (.A(g24575), .B(g18407), .Z(g25201) ) ;
INV     gate14299  (.A(g25201), .Z(II34476) ) ;
INV     gate14300  (.A(II34476), .Z(g26506) ) ;
NOR2    gate14301  (.A(g24566), .B(g22907), .Z(g25202) ) ;
INV     gate14302  (.A(g25202), .Z(II34479) ) ;
INV     gate14303  (.A(II34479), .Z(g26507) ) ;
NAND4   gate14304  (.A(g21211), .B(g14442), .C(g10694), .D(g24590), .Z(g25312) ) ;
INV     gate14305  (.A(g25312), .Z(g26508) ) ;
NOR2    gate14306  (.A(g25081), .B(g21674), .Z(g25853) ) ;
INV     gate14307  (.A(g25853), .Z(g26512) ) ;
NAND4   gate14308  (.A(g21219), .B(g14529), .C(g10714), .D(g24595), .Z(g25320) ) ;
INV     gate14309  (.A(g25320), .Z(g26516) ) ;
NOR2    gate14310  (.A(g25085), .B(g21703), .Z(g25874) ) ;
INV     gate14311  (.A(g25874), .Z(g26520) ) ;
NAND4   gate14312  (.A(g21230), .B(g14584), .C(g10735), .D(g24603), .Z(g25331) ) ;
INV     gate14313  (.A(g25331), .Z(g26521) ) ;
NAND4   gate14314  (.A(g21235), .B(g14618), .C(g10754), .D(g24610), .Z(g25340) ) ;
INV     gate14315  (.A(g25340), .Z(g26525) ) ;
INV     gate14316  (.A(g25454), .Z(g26533) ) ;
INV     gate14317  (.A(g25458), .Z(g26538) ) ;
INV     gate14318  (.A(g25463), .Z(g26539) ) ;
INV     gate14319  (.A(g25467), .Z(g26540) ) ;
INV     gate14320  (.A(g25472), .Z(g26542) ) ;
INV     gate14321  (.A(g25476), .Z(g26543) ) ;
INV     gate14322  (.A(g25479), .Z(g26544) ) ;
INV     gate14323  (.A(g25484), .Z(g26546) ) ;
NOR2    gate14324  (.A(g16018), .B(g25086), .Z(g25450) ) ;
INV     gate14325  (.A(g25450), .Z(II34505) ) ;
INV     gate14326  (.A(II34505), .Z(g26548) ) ;
INV     gate14327  (.A(g25421), .Z(g26549) ) ;
INV     gate14328  (.A(g25493), .Z(g26550) ) ;
INV     gate14329  (.A(g25496), .Z(g26551) ) ;
INV     gate14330  (.A(g25499), .Z(g26552) ) ;
INV     gate14331  (.A(g25502), .Z(g26554) ) ;
INV     gate14332  (.A(g25507), .Z(g26555) ) ;
INV     gate14333  (.A(g25510), .Z(g26556) ) ;
INV     gate14334  (.A(g25515), .Z(g26558) ) ;
INV     gate14335  (.A(g25524), .Z(g26561) ) ;
INV     gate14336  (.A(g25527), .Z(g26562) ) ;
INV     gate14337  (.A(g25530), .Z(g26563) ) ;
INV     gate14338  (.A(g25533), .Z(g26564) ) ;
INV     gate14339  (.A(g25536), .Z(g26565) ) ;
INV     gate14340  (.A(g25540), .Z(g26566) ) ;
INV     gate14341  (.A(g25543), .Z(g26567) ) ;
INV     gate14342  (.A(g25546), .Z(g26568) ) ;
INV     gate14343  (.A(g25549), .Z(g26570) ) ;
INV     gate14344  (.A(g25554), .Z(g26571) ) ;
INV     gate14345  (.A(g25557), .Z(g26572) ) ;
INV     gate14346  (.A(g25562), .Z(g26574) ) ;
NOR2    gate14347  (.A(g16048), .B(g25102), .Z(g25451) ) ;
INV     gate14348  (.A(g25451), .Z(II34535) ) ;
INV     gate14349  (.A(II34535), .Z(g26576) ) ;
INV     gate14350  (.A(g25436), .Z(g26577) ) ;
INV     gate14351  (.A(g25573), .Z(g26578) ) ;
INV     gate14352  (.A(g25576), .Z(g26579) ) ;
INV     gate14353  (.A(g25579), .Z(g26580) ) ;
INV     gate14354  (.A(g25582), .Z(g26581) ) ;
INV     gate14355  (.A(g25585), .Z(g26582) ) ;
INV     gate14356  (.A(g25590), .Z(g26584) ) ;
INV     gate14357  (.A(g25593), .Z(g26585) ) ;
INV     gate14358  (.A(g25596), .Z(g26586) ) ;
INV     gate14359  (.A(g25599), .Z(g26587) ) ;
INV     gate14360  (.A(g25602), .Z(g26588) ) ;
INV     gate14361  (.A(g25606), .Z(g26589) ) ;
INV     gate14362  (.A(g25609), .Z(g26590) ) ;
INV     gate14363  (.A(g25612), .Z(g26591) ) ;
INV     gate14364  (.A(g25615), .Z(g26593) ) ;
INV     gate14365  (.A(g25620), .Z(g26594) ) ;
INV     gate14366  (.A(g25623), .Z(g26595) ) ;
INV     gate14367  (.A(g25443), .Z(g26597) ) ;
INV     gate14368  (.A(g25634), .Z(g26598) ) ;
INV     gate14369  (.A(g25637), .Z(g26599) ) ;
INV     gate14370  (.A(g25640), .Z(g26600) ) ;
INV     gate14371  (.A(g25643), .Z(g26601) ) ;
INV     gate14372  (.A(g25652), .Z(g26602) ) ;
INV     gate14373  (.A(g25655), .Z(g26603) ) ;
INV     gate14374  (.A(g25658), .Z(g26604) ) ;
INV     gate14375  (.A(g25661), .Z(g26605) ) ;
INV     gate14376  (.A(g25664), .Z(g26606) ) ;
INV     gate14377  (.A(g25669), .Z(g26608) ) ;
INV     gate14378  (.A(g25672), .Z(g26609) ) ;
INV     gate14379  (.A(g25675), .Z(g26610) ) ;
INV     gate14380  (.A(g25678), .Z(g26611) ) ;
INV     gate14381  (.A(g25681), .Z(g26612) ) ;
INV     gate14382  (.A(g25685), .Z(g26613) ) ;
INV     gate14383  (.A(g25688), .Z(g26614) ) ;
INV     gate14384  (.A(g25691), .Z(g26615) ) ;
INV     gate14385  (.A(g25694), .Z(g26617) ) ;
NOR2    gate14386  (.A(g16101), .B(g25117), .Z(g25452) ) ;
INV     gate14387  (.A(g25452), .Z(II34579) ) ;
INV     gate14388  (.A(II34579), .Z(g26618) ) ;
INV     gate14389  (.A(g25700), .Z(g26619) ) ;
INV     gate14390  (.A(g25703), .Z(g26620) ) ;
INV     gate14391  (.A(g25711), .Z(g26621) ) ;
INV     gate14392  (.A(g25714), .Z(g26622) ) ;
INV     gate14393  (.A(g25717), .Z(g26623) ) ;
INV     gate14394  (.A(g25720), .Z(g26624) ) ;
INV     gate14395  (.A(g25729), .Z(g26625) ) ;
INV     gate14396  (.A(g25732), .Z(g26626) ) ;
INV     gate14397  (.A(g25735), .Z(g26627) ) ;
INV     gate14398  (.A(g25738), .Z(g26628) ) ;
INV     gate14399  (.A(g25741), .Z(g26629) ) ;
INV     gate14400  (.A(g25746), .Z(g26631) ) ;
INV     gate14401  (.A(g25749), .Z(g26632) ) ;
INV     gate14402  (.A(g25752), .Z(g26633) ) ;
INV     gate14403  (.A(g25755), .Z(g26634) ) ;
INV     gate14404  (.A(g25758), .Z(g26635) ) ;
INV     gate14405  (.A(g25767), .Z(g26636) ) ;
INV     gate14406  (.A(g25773), .Z(g26637) ) ;
INV     gate14407  (.A(g25776), .Z(g26638) ) ;
INV     gate14408  (.A(g25784), .Z(g26639) ) ;
INV     gate14409  (.A(g25787), .Z(g26640) ) ;
INV     gate14410  (.A(g25790), .Z(g26641) ) ;
INV     gate14411  (.A(g25793), .Z(g26642) ) ;
INV     gate14412  (.A(g25802), .Z(g26643) ) ;
INV     gate14413  (.A(g25805), .Z(g26644) ) ;
INV     gate14414  (.A(g25808), .Z(g26645) ) ;
INV     gate14415  (.A(g25811), .Z(g26646) ) ;
INV     gate14416  (.A(g25814), .Z(g26647) ) ;
INV     gate14417  (.A(g25821), .Z(g26648) ) ;
INV     gate14418  (.A(g25827), .Z(g26649) ) ;
INV     gate14419  (.A(g25830), .Z(g26650) ) ;
INV     gate14420  (.A(g25838), .Z(g26651) ) ;
INV     gate14421  (.A(g25841), .Z(g26652) ) ;
INV     gate14422  (.A(g25844), .Z(g26653) ) ;
INV     gate14423  (.A(g25847), .Z(g26654) ) ;
INV     gate14424  (.A(g25856), .Z(g26656) ) ;
INV     gate14425  (.A(g25862), .Z(g26657) ) ;
INV     gate14426  (.A(g25865), .Z(g26658) ) ;
INV     gate14427  (.A(g25877), .Z(g26662) ) ;
INV     gate14428  (.A(g26086), .Z(II34641) ) ;
INV     gate14429  (.A(g26159), .Z(II34644) ) ;
INV     gate14430  (.A(g26164), .Z(II34647) ) ;
INV     gate14431  (.A(g26172), .Z(II34650) ) ;
INV     gate14432  (.A(g26165), .Z(II34653) ) ;
INV     gate14433  (.A(g26173), .Z(II34656) ) ;
INV     gate14434  (.A(g26190), .Z(II34659) ) ;
INV     gate14435  (.A(g26174), .Z(II34662) ) ;
INV     gate14436  (.A(g26191), .Z(II34665) ) ;
INV     gate14437  (.A(g26210), .Z(II34668) ) ;
INV     gate14438  (.A(g26192), .Z(II34671) ) ;
INV     gate14439  (.A(g26211), .Z(II34674) ) ;
INV     gate14440  (.A(g26232), .Z(II34677) ) ;
INV     gate14441  (.A(g26294), .Z(II34680) ) ;
INV     gate14442  (.A(g26364), .Z(II34683) ) ;
INV     gate14443  (.A(g26398), .Z(II34686) ) ;
INV     gate14444  (.A(g26433), .Z(II34689) ) ;
INV     gate14445  (.A(g26102), .Z(II34692) ) ;
INV     gate14446  (.A(g26167), .Z(II34695) ) ;
INV     gate14447  (.A(g26181), .Z(II34698) ) ;
INV     gate14448  (.A(g26193), .Z(II34701) ) ;
INV     gate14449  (.A(g26182), .Z(II34704) ) ;
INV     gate14450  (.A(g26194), .Z(II34707) ) ;
INV     gate14451  (.A(g26214), .Z(II34710) ) ;
INV     gate14452  (.A(g26195), .Z(II34713) ) ;
INV     gate14453  (.A(g26215), .Z(II34716) ) ;
INV     gate14454  (.A(g26238), .Z(II34719) ) ;
INV     gate14455  (.A(g26216), .Z(II34722) ) ;
INV     gate14456  (.A(g26239), .Z(II34725) ) ;
INV     gate14457  (.A(g26264), .Z(II34728) ) ;
INV     gate14458  (.A(g26341), .Z(II34731) ) ;
INV     gate14459  (.A(g26407), .Z(II34734) ) ;
INV     gate14460  (.A(g26439), .Z(II34737) ) ;
INV     gate14461  (.A(g26465), .Z(II34740) ) ;
INV     gate14462  (.A(g26118), .Z(II34743) ) ;
INV     gate14463  (.A(g26187), .Z(II34746) ) ;
INV     gate14464  (.A(g26205), .Z(II34749) ) ;
INV     gate14465  (.A(g26220), .Z(II34752) ) ;
INV     gate14466  (.A(g26206), .Z(II34755) ) ;
INV     gate14467  (.A(g26221), .Z(II34758) ) ;
INV     gate14468  (.A(g26245), .Z(II34761) ) ;
INV     gate14469  (.A(g26222), .Z(II34764) ) ;
INV     gate14470  (.A(g26246), .Z(II34767) ) ;
INV     gate14471  (.A(g26276), .Z(II34770) ) ;
INV     gate14472  (.A(g26247), .Z(II34773) ) ;
INV     gate14473  (.A(g26277), .Z(II34776) ) ;
INV     gate14474  (.A(g26308), .Z(II34779) ) ;
INV     gate14475  (.A(g26385), .Z(II34782) ) ;
INV     gate14476  (.A(g26448), .Z(II34785) ) ;
INV     gate14477  (.A(g26471), .Z(II34788) ) ;
INV     gate14478  (.A(g26489), .Z(II34791) ) ;
INV     gate14479  (.A(g26125), .Z(II34794) ) ;
INV     gate14480  (.A(g26208), .Z(II34797) ) ;
INV     gate14481  (.A(g26229), .Z(II34800) ) ;
INV     gate14482  (.A(g26248), .Z(II34803) ) ;
INV     gate14483  (.A(g26230), .Z(II34806) ) ;
INV     gate14484  (.A(g26249), .Z(II34809) ) ;
INV     gate14485  (.A(g26280), .Z(II34812) ) ;
INV     gate14486  (.A(g26250), .Z(II34815) ) ;
INV     gate14487  (.A(g26281), .Z(II34818) ) ;
INV     gate14488  (.A(g26314), .Z(II34821) ) ;
INV     gate14489  (.A(g26282), .Z(II34824) ) ;
INV     gate14490  (.A(g26315), .Z(II34827) ) ;
INV     gate14491  (.A(g26349), .Z(II34830) ) ;
INV     gate14492  (.A(g26428), .Z(II34833) ) ;
INV     gate14493  (.A(g26480), .Z(II34836) ) ;
INV     gate14494  (.A(g26495), .Z(II34839) ) ;
INV     gate14495  (.A(g26505), .Z(II34842) ) ;
INV     gate14496  (.A(g26496), .Z(II34845) ) ;
INV     gate14497  (.A(g26506), .Z(II34848) ) ;
INV     gate14498  (.A(g26354), .Z(II34851) ) ;
INV     gate14499  (.A(g26507), .Z(II34854) ) ;
INV     gate14500  (.A(g26355), .Z(II34857) ) ;
INV     gate14501  (.A(g26548), .Z(II34860) ) ;
INV     gate14502  (.A(g26576), .Z(II34863) ) ;
INV     gate14503  (.A(g26618), .Z(II34866) ) ;
NOR2    gate14504  (.A(g25963), .B(g13320), .Z(g26217) ) ;
INV     gate14505  (.A(g26217), .Z(II34872) ) ;
INV     gate14506  (.A(II34872), .Z(g26757) ) ;
NOR2    gate14507  (.A(g25968), .B(g13340), .Z(g26240) ) ;
INV     gate14508  (.A(g26240), .Z(II34879) ) ;
INV     gate14509  (.A(II34879), .Z(g26762) ) ;
NOR2    gate14510  (.A(g25977), .B(g13385), .Z(g26295) ) ;
INV     gate14511  (.A(g26295), .Z(II34901) ) ;
INV     gate14512  (.A(II34901), .Z(g26782) ) ;
NOR2    gate14513  (.A(g25972), .B(g13360), .Z(g26265) ) ;
INV     gate14514  (.A(g26265), .Z(II34909) ) ;
INV     gate14515  (.A(II34909), .Z(g26788) ) ;
INV     gate14516  (.A(g26240), .Z(II34916) ) ;
INV     gate14517  (.A(II34916), .Z(g26793) ) ;
INV     gate14518  (.A(g26217), .Z(II34921) ) ;
INV     gate14519  (.A(II34921), .Z(g26796) ) ;
NOR2    gate14520  (.A(g25321), .B(g8869), .Z(g26534) ) ;
INV     gate14521  (.A(g26534), .Z(II34946) ) ;
INV     gate14522  (.A(II34946), .Z(g26819) ) ;
NOR2    gate14523  (.A(g13755), .B(g25269), .Z(g26541) ) ;
INV     gate14524  (.A(g26541), .Z(II34957) ) ;
INV     gate14525  (.A(II34957), .Z(g26828) ) ;
NOR2    gate14526  (.A(g13790), .B(g25277), .Z(g26545) ) ;
INV     gate14527  (.A(g26545), .Z(II34961) ) ;
INV     gate14528  (.A(II34961), .Z(g26830) ) ;
NOR2    gate14529  (.A(g13796), .B(g25278), .Z(g26547) ) ;
INV     gate14530  (.A(g26547), .Z(II34964) ) ;
INV     gate14531  (.A(II34964), .Z(g26831) ) ;
NOR2    gate14532  (.A(g13816), .B(g25282), .Z(g26553) ) ;
INV     gate14533  (.A(g26553), .Z(II34967) ) ;
INV     gate14534  (.A(II34967), .Z(g26832) ) ;
NOR2    gate14535  (.A(g13818), .B(g25286), .Z(g26557) ) ;
INV     gate14536  (.A(g26557), .Z(II34971) ) ;
INV     gate14537  (.A(II34971), .Z(g26834) ) ;
NOR2    gate14538  (.A(g25953), .B(g16212), .Z(g26168) ) ;
INV     gate14539  (.A(g26168), .Z(II34974) ) ;
INV     gate14540  (.A(II34974), .Z(g26835) ) ;
NOR2    gate14541  (.A(g13824), .B(g25287), .Z(g26559) ) ;
INV     gate14542  (.A(g26559), .Z(II34977) ) ;
INV     gate14543  (.A(II34977), .Z(g26836) ) ;
NAND2   gate14544  (.A(g25343), .B(g65), .Z(g26458) ) ;
INV     gate14545  (.A(g26458), .Z(II34980) ) ;
INV     gate14546  (.A(II34980), .Z(g26837) ) ;
NOR2    gate14547  (.A(g13837), .B(g25290), .Z(g26569) ) ;
INV     gate14548  (.A(g26569), .Z(II34983) ) ;
INV     gate14549  (.A(II34983), .Z(g26840) ) ;
NOR2    gate14550  (.A(g25951), .B(g16162), .Z(g26160) ) ;
INV     gate14551  (.A(g26160), .Z(II34986) ) ;
INV     gate14552  (.A(II34986), .Z(g26841) ) ;
NOR2    gate14553  (.A(g13839), .B(g25294), .Z(g26573) ) ;
INV     gate14554  (.A(g26573), .Z(II34990) ) ;
INV     gate14555  (.A(II34990), .Z(g26843) ) ;
NOR2    gate14556  (.A(g13845), .B(g25295), .Z(g26575) ) ;
INV     gate14557  (.A(g26575), .Z(II34993) ) ;
INV     gate14558  (.A(II34993), .Z(g26844) ) ;
NAND2   gate14559  (.A(g25357), .B(g753), .Z(g26482) ) ;
INV     gate14560  (.A(g26482), .Z(II34997) ) ;
INV     gate14561  (.A(II34997), .Z(g26846) ) ;
NOR2    gate14562  (.A(g25981), .B(g13481), .Z(g26336) ) ;
INV     gate14563  (.A(g26336), .Z(II35000) ) ;
INV     gate14564  (.A(II35000), .Z(g26849) ) ;
NOR2    gate14565  (.A(g13851), .B(g25300), .Z(g26592) ) ;
INV     gate14566  (.A(g26592), .Z(II35003) ) ;
INV     gate14567  (.A(II35003), .Z(g26850) ) ;
NOR2    gate14568  (.A(g13853), .B(g25304), .Z(g26596) ) ;
INV     gate14569  (.A(g26596), .Z(II35007) ) ;
INV     gate14570  (.A(II35007), .Z(g26852) ) ;
NOR2    gate14571  (.A(g25978), .B(g16451), .Z(g26304) ) ;
INV     gate14572  (.A(g26304), .Z(II35011) ) ;
INV     gate14573  (.A(II35011), .Z(g26854) ) ;
NAND2   gate14574  (.A(g25372), .B(g1439), .Z(g26498) ) ;
INV     gate14575  (.A(g26498), .Z(II35014) ) ;
INV     gate14576  (.A(II35014), .Z(g26855) ) ;
NOR2    gate14577  (.A(g13860), .B(g25310), .Z(g26616) ) ;
INV     gate14578  (.A(g26616), .Z(II35017) ) ;
INV     gate14579  (.A(II35017), .Z(g26858) ) ;
NAND2   gate14580  (.A(g25389), .B(g2133), .Z(g26513) ) ;
INV     gate14581  (.A(g26513), .Z(II35028) ) ;
INV     gate14582  (.A(II35028), .Z(g26861) ) ;
NOR2    gate14583  (.A(g25962), .B(g17001), .Z(g26529) ) ;
INV     gate14584  (.A(g26529), .Z(II35031) ) ;
INV     gate14585  (.A(II35031), .Z(g26864) ) ;
NOR2    gate14586  (.A(g25967), .B(g17031), .Z(g26530) ) ;
INV     gate14587  (.A(g26530), .Z(II35049) ) ;
INV     gate14588  (.A(II35049), .Z(g26868) ) ;
NOR2    gate14589  (.A(g25328), .B(g17084), .Z(g26655) ) ;
INV     gate14590  (.A(g26655), .Z(II35053) ) ;
INV     gate14591  (.A(II35053), .Z(g26872) ) ;
NOR2    gate14592  (.A(g25974), .B(g17065), .Z(g26531) ) ;
INV     gate14593  (.A(g26531), .Z(II35064) ) ;
INV     gate14594  (.A(II35064), .Z(g26875) ) ;
NOR2    gate14595  (.A(g25334), .B(g17116), .Z(g26659) ) ;
INV     gate14596  (.A(g26659), .Z(II35067) ) ;
INV     gate14597  (.A(II35067), .Z(g26876) ) ;
NOR2    gate14598  (.A(g25337), .B(g17122), .Z(g26661) ) ;
INV     gate14599  (.A(g26661), .Z(II35072) ) ;
INV     gate14600  (.A(II35072), .Z(g26881) ) ;
NOR2    gate14601  (.A(g25979), .B(g17100), .Z(g26532) ) ;
INV     gate14602  (.A(g26532), .Z(II35076) ) ;
INV     gate14603  (.A(II35076), .Z(g26883) ) ;
NOR2    gate14604  (.A(g25346), .B(g17138), .Z(g26664) ) ;
INV     gate14605  (.A(g26664), .Z(II35079) ) ;
INV     gate14606  (.A(II35079), .Z(g26884) ) ;
NOR2    gate14607  (.A(g25348), .B(g17143), .Z(g26665) ) ;
INV     gate14608  (.A(g26665), .Z(II35083) ) ;
INV     gate14609  (.A(II35083), .Z(g26886) ) ;
NOR2    gate14610  (.A(g25351), .B(g17149), .Z(g26667) ) ;
INV     gate14611  (.A(g26667), .Z(II35087) ) ;
INV     gate14612  (.A(II35087), .Z(g26890) ) ;
NOR2    gate14613  (.A(g25360), .B(g17161), .Z(g26669) ) ;
INV     gate14614  (.A(g26669), .Z(II35092) ) ;
INV     gate14615  (.A(II35092), .Z(g26895) ) ;
NOR2    gate14616  (.A(g25362), .B(g17166), .Z(g26670) ) ;
INV     gate14617  (.A(g26670), .Z(II35095) ) ;
INV     gate14618  (.A(II35095), .Z(g26896) ) ;
NOR2    gate14619  (.A(g25365), .B(g17172), .Z(g26672) ) ;
INV     gate14620  (.A(g26672), .Z(II35099) ) ;
INV     gate14621  (.A(II35099), .Z(g26900) ) ;
NOR2    gate14622  (.A(g25375), .B(g17176), .Z(g26675) ) ;
INV     gate14623  (.A(g26675), .Z(II35106) ) ;
INV     gate14624  (.A(II35106), .Z(g26909) ) ;
NOR2    gate14625  (.A(g25377), .B(g17181), .Z(g26676) ) ;
INV     gate14626  (.A(g26676), .Z(II35109) ) ;
INV     gate14627  (.A(II35109), .Z(g26910) ) ;
NOR2    gate14628  (.A(g25392), .B(g17193), .Z(g26025) ) ;
INV     gate14629  (.A(g26025), .Z(II35116) ) ;
INV     gate14630  (.A(II35116), .Z(g26921) ) ;
NOR2    gate14631  (.A(g25954), .B(g24486), .Z(g26283) ) ;
INV     gate14632  (.A(g26283), .Z(g26922) ) ;
NOR2    gate14633  (.A(g25958), .B(g24493), .Z(g26327) ) ;
INV     gate14634  (.A(g26327), .Z(g26935) ) ;
NOR2    gate14635  (.A(g25964), .B(g24503), .Z(g26374) ) ;
INV     gate14636  (.A(g26374), .Z(g26944) ) ;
NOR2    gate14637  (.A(g25969), .B(g24515), .Z(g26417) ) ;
INV     gate14638  (.A(g26417), .Z(g26950) ) ;
NOR2    gate14639  (.A(g25208), .B(g10024), .Z(g26660) ) ;
INV     gate14640  (.A(g26660), .Z(II35136) ) ;
INV     gate14641  (.A(II35136), .Z(g26953) ) ;
INV     gate14642  (.A(g26549), .Z(g26954) ) ;
NOR2    gate14643  (.A(g25216), .B(g10133), .Z(g26666) ) ;
INV     gate14644  (.A(g26666), .Z(II35141) ) ;
INV     gate14645  (.A(II35141), .Z(g26956) ) ;
INV     gate14646  (.A(g26577), .Z(g26957) ) ;
NOR2    gate14647  (.A(g25226), .B(g10238), .Z(g26671) ) ;
INV     gate14648  (.A(g26671), .Z(II35146) ) ;
INV     gate14649  (.A(II35146), .Z(g26959) ) ;
INV     gate14650  (.A(g26597), .Z(g26960) ) ;
NOR2    gate14651  (.A(g25238), .B(g10340), .Z(g26677) ) ;
INV     gate14652  (.A(g26677), .Z(II35153) ) ;
INV     gate14653  (.A(II35153), .Z(g26964) ) ;
NOR2    gate14654  (.A(g25973), .B(g16423), .Z(g26272) ) ;
INV     gate14655  (.A(g26272), .Z(II35172) ) ;
INV     gate14656  (.A(II35172), .Z(g26983) ) ;
INV     gate14657  (.A(g26056), .Z(g26987) ) ;
INV     gate14658  (.A(g26063), .Z(g27010) ) ;
INV     gate14659  (.A(g26070), .Z(g27036) ) ;
INV     gate14660  (.A(g26076), .Z(g27064) ) ;
NOR2    gate14661  (.A(g25628), .B(g24906), .Z(g26048) ) ;
INV     gate14662  (.A(g26048), .Z(II35254) ) ;
INV     gate14663  (.A(II35254), .Z(g27075) ) ;
NOR2    gate14664  (.A(g25273), .B(g22777), .Z(g26031) ) ;
INV     gate14665  (.A(g26031), .Z(II35283) ) ;
INV     gate14666  (.A(II35283), .Z(g27102) ) ;
NOR2    gate14667  (.A(g25961), .B(g13291), .Z(g26199) ) ;
INV     gate14668  (.A(g26199), .Z(II35297) ) ;
INV     gate14669  (.A(II35297), .Z(g27114) ) ;
NOR2    gate14670  (.A(g25311), .B(g18407), .Z(g26037) ) ;
INV     gate14671  (.A(g26037), .Z(II35301) ) ;
INV     gate14672  (.A(II35301), .Z(g27116) ) ;
INV     gate14673  (.A(g26534), .Z(II35313) ) ;
INV     gate14674  (.A(II35313), .Z(g27126) ) ;
NOR2    gate14675  (.A(g25957), .B(g13270), .Z(g26183) ) ;
INV     gate14676  (.A(g26183), .Z(II35319) ) ;
INV     gate14677  (.A(II35319), .Z(g27132) ) ;
INV     gate14678  (.A(g26105), .Z(g27133) ) ;
INV     gate14679  (.A(g26175), .Z(g27134) ) ;
INV     gate14680  (.A(g26178), .Z(g27135) ) ;
INV     gate14681  (.A(g26196), .Z(g27136) ) ;
INV     gate14682  (.A(g26202), .Z(g27137) ) ;
INV     gate14683  (.A(g26223), .Z(g27138) ) ;
INV     gate14684  (.A(g26226), .Z(g27139) ) ;
INV     gate14685  (.A(g26136), .Z(g27140) ) ;
INV     gate14686  (.A(g26251), .Z(g27141) ) ;
INV     gate14687  (.A(g26254), .Z(g27142) ) ;
INV     gate14688  (.A(g26150), .Z(g27143) ) ;
NAND2   gate14689  (.A(g23644), .B(g25354), .Z(g26106) ) ;
INV     gate14690  (.A(g26106), .Z(II35334) ) ;
INV     gate14691  (.A(II35334), .Z(g27145) ) ;
INV     gate14692  (.A(g26358), .Z(g27146) ) ;
INV     gate14693  (.A(g26393), .Z(g27148) ) ;
NAND2   gate14694  (.A(g23694), .B(g25369), .Z(g26120) ) ;
INV     gate14695  (.A(g26120), .Z(II35341) ) ;
INV     gate14696  (.A(II35341), .Z(g27150) ) ;
INV     gate14697  (.A(g26401), .Z(g27151) ) ;
INV     gate14698  (.A(g26429), .Z(g27153) ) ;
INV     gate14699  (.A(g26265), .Z(II35347) ) ;
INV     gate14700  (.A(II35347), .Z(g27154) ) ;
INV     gate14701  (.A(g26434), .Z(g27155) ) ;
INV     gate14702  (.A(g26272), .Z(II35351) ) ;
INV     gate14703  (.A(II35351), .Z(g27156) ) ;
NAND2   gate14704  (.A(g23748), .B(g25386), .Z(g26130) ) ;
INV     gate14705  (.A(g26130), .Z(II35355) ) ;
INV     gate14706  (.A(II35355), .Z(g27158) ) ;
INV     gate14707  (.A(g26442), .Z(g27159) ) ;
INV     gate14708  (.A(g26295), .Z(II35360) ) ;
INV     gate14709  (.A(II35360), .Z(g27161) ) ;
INV     gate14710  (.A(g26461), .Z(g27162) ) ;
INV     gate14711  (.A(g26304), .Z(II35364) ) ;
INV     gate14712  (.A(II35364), .Z(g27163) ) ;
INV     gate14713  (.A(g26466), .Z(g27164) ) ;
NAND2   gate14714  (.A(g23803), .B(g25402), .Z(g26144) ) ;
INV     gate14715  (.A(g26144), .Z(II35369) ) ;
INV     gate14716  (.A(II35369), .Z(g27166) ) ;
INV     gate14717  (.A(g26474), .Z(g27167) ) ;
INV     gate14718  (.A(g26189), .Z(II35373) ) ;
INV     gate14719  (.A(II35373), .Z(g27168) ) ;
INV     gate14720  (.A(g26336), .Z(II35376) ) ;
INV     gate14721  (.A(II35376), .Z(g27171) ) ;
INV     gate14722  (.A(g26485), .Z(g27172) ) ;
INV     gate14723  (.A(g26490), .Z(g27173) ) ;
INV     gate14724  (.A(g26160), .Z(II35383) ) ;
INV     gate14725  (.A(II35383), .Z(g27176) ) ;
INV     gate14726  (.A(g26501), .Z(g27177) ) ;
INV     gate14727  (.A(g26168), .Z(II35389) ) ;
INV     gate14728  (.A(II35389), .Z(g27180) ) ;
INV     gate14729  (.A(g26183), .Z(II35394) ) ;
INV     gate14730  (.A(II35394), .Z(g27183) ) ;
INV     gate14731  (.A(g26199), .Z(II35399) ) ;
INV     gate14732  (.A(II35399), .Z(g27186) ) ;
INV     gate14733  (.A(g26864), .Z(II35404) ) ;
INV     gate14734  (.A(g27145), .Z(II35407) ) ;
INV     gate14735  (.A(g26872), .Z(II35410) ) ;
INV     gate14736  (.A(g26876), .Z(II35413) ) ;
INV     gate14737  (.A(g26884), .Z(II35416) ) ;
INV     gate14738  (.A(g26828), .Z(II35419) ) ;
INV     gate14739  (.A(g26830), .Z(II35422) ) ;
INV     gate14740  (.A(g26832), .Z(II35425) ) ;
INV     gate14741  (.A(g26953), .Z(II35428) ) ;
INV     gate14742  (.A(g26868), .Z(II35431) ) ;
INV     gate14743  (.A(g27150), .Z(II35434) ) ;
INV     gate14744  (.A(g27183), .Z(II35437) ) ;
INV     gate14745  (.A(g27186), .Z(II35440) ) ;
INV     gate14746  (.A(g26757), .Z(II35443) ) ;
INV     gate14747  (.A(g26762), .Z(II35446) ) ;
INV     gate14748  (.A(g27154), .Z(II35449) ) ;
INV     gate14749  (.A(g27161), .Z(II35452) ) ;
INV     gate14750  (.A(g26881), .Z(II35455) ) ;
INV     gate14751  (.A(g26886), .Z(II35458) ) ;
INV     gate14752  (.A(g26895), .Z(II35461) ) ;
INV     gate14753  (.A(g26831), .Z(II35464) ) ;
INV     gate14754  (.A(g26834), .Z(II35467) ) ;
INV     gate14755  (.A(g26840), .Z(II35470) ) ;
INV     gate14756  (.A(g27156), .Z(II35473) ) ;
INV     gate14757  (.A(g27163), .Z(II35476) ) ;
INV     gate14758  (.A(g27171), .Z(II35479) ) ;
INV     gate14759  (.A(g27176), .Z(II35482) ) ;
INV     gate14760  (.A(g27180), .Z(II35485) ) ;
INV     gate14761  (.A(g26819), .Z(II35488) ) ;
INV     gate14762  (.A(g26956), .Z(II35491) ) ;
INV     gate14763  (.A(g26875), .Z(II35494) ) ;
INV     gate14764  (.A(g27158), .Z(II35497) ) ;
INV     gate14765  (.A(g26890), .Z(II35500) ) ;
INV     gate14766  (.A(g26896), .Z(II35503) ) ;
INV     gate14767  (.A(g26909), .Z(II35506) ) ;
INV     gate14768  (.A(g26836), .Z(II35509) ) ;
INV     gate14769  (.A(g26843), .Z(II35512) ) ;
INV     gate14770  (.A(g26850), .Z(II35515) ) ;
INV     gate14771  (.A(g26959), .Z(II35518) ) ;
INV     gate14772  (.A(g26883), .Z(II35521) ) ;
INV     gate14773  (.A(g27166), .Z(II35524) ) ;
INV     gate14774  (.A(g26900), .Z(II35527) ) ;
INV     gate14775  (.A(g26910), .Z(II35530) ) ;
INV     gate14776  (.A(g26921), .Z(II35533) ) ;
INV     gate14777  (.A(g26844), .Z(II35536) ) ;
INV     gate14778  (.A(g26852), .Z(II35539) ) ;
INV     gate14779  (.A(g26858), .Z(II35542) ) ;
INV     gate14780  (.A(g26964), .Z(II35545) ) ;
INV     gate14781  (.A(g27116), .Z(II35548) ) ;
INV     gate14782  (.A(g27075), .Z(II35551) ) ;
INV     gate14783  (.A(g27102), .Z(II35554) ) ;
INV     gate14784  (.A(g27126), .Z(g27349) ) ;
NOR2    gate14785  (.A(g26560), .B(g17001), .Z(g27120) ) ;
INV     gate14786  (.A(g27120), .Z(II35667) ) ;
INV     gate14787  (.A(II35667), .Z(g27353) ) ;
NOR2    gate14788  (.A(g26583), .B(g17031), .Z(g27123) ) ;
INV     gate14789  (.A(g27123), .Z(II35673) ) ;
INV     gate14790  (.A(II35673), .Z(g27357) ) ;
NOR2    gate14791  (.A(g26607), .B(g17065), .Z(g27129) ) ;
INV     gate14792  (.A(g27129), .Z(II35678) ) ;
INV     gate14793  (.A(II35678), .Z(g27360) ) ;
NOR2    gate14794  (.A(g26458), .B(g5642), .Z(g26869) ) ;
INV     gate14795  (.A(g26869), .Z(II35681) ) ;
INV     gate14796  (.A(II35681), .Z(g27361) ) ;
NOR2    gate14797  (.A(g26630), .B(g17100), .Z(g27131) ) ;
INV     gate14798  (.A(g27131), .Z(II35686) ) ;
INV     gate14799  (.A(II35686), .Z(g27366) ) ;
NOR2    gate14800  (.A(g26482), .B(g5680), .Z(g26878) ) ;
INV     gate14801  (.A(g26878), .Z(II35689) ) ;
INV     gate14802  (.A(II35689), .Z(g27367) ) ;
NOR2    gate14803  (.A(g26498), .B(g5732), .Z(g26887) ) ;
INV     gate14804  (.A(g26887), .Z(II35695) ) ;
INV     gate14805  (.A(II35695), .Z(g27373) ) ;
NOR2    gate14806  (.A(g26513), .B(g5790), .Z(g26897) ) ;
INV     gate14807  (.A(g26897), .Z(II35698) ) ;
INV     gate14808  (.A(II35698), .Z(g27376) ) ;
OR2     gate14809  (.A(g26157), .B(g23147), .Z(g26974) ) ;
INV     gate14810  (.A(g26974), .Z(II35708) ) ;
INV     gate14811  (.A(g26974), .Z(II35711) ) ;
INV     gate14812  (.A(II35711), .Z(g27381) ) ;
INV     gate14813  (.A(g27133), .Z(g27383) ) ;
INV     gate14814  (.A(g27140), .Z(g27384) ) ;
INV     gate14815  (.A(g27168), .Z(II35723) ) ;
INV     gate14816  (.A(II35723), .Z(g27385) ) ;
INV     gate14817  (.A(g27143), .Z(g27386) ) ;
NAND3   gate14818  (.A(g25631), .B(g26283), .C(g25569), .Z(g26902) ) ;
INV     gate14819  (.A(g26902), .Z(II35727) ) ;
INV     gate14820  (.A(II35727), .Z(g27387) ) ;
NAND4   gate14821  (.A(g25699), .B(g26283), .C(g25569), .D(g25631), .Z(g26892) ) ;
INV     gate14822  (.A(g26892), .Z(II35731) ) ;
INV     gate14823  (.A(II35731), .Z(g27391) ) ;
NAND3   gate14824  (.A(g25708), .B(g26327), .C(g25648), .Z(g26915) ) ;
INV     gate14825  (.A(g26915), .Z(II35737) ) ;
INV     gate14826  (.A(II35737), .Z(g27397) ) ;
NAND2   gate14827  (.A(g26320), .B(g5438), .Z(g27118) ) ;
INV     gate14828  (.A(g27118), .Z(II35741) ) ;
INV     gate14829  (.A(II35741), .Z(g27401) ) ;
NAND4   gate14830  (.A(g25772), .B(g26327), .C(g25648), .D(g25708), .Z(g26906) ) ;
INV     gate14831  (.A(g26906), .Z(II35744) ) ;
INV     gate14832  (.A(II35744), .Z(g27404) ) ;
NAND3   gate14833  (.A(g25781), .B(g26374), .C(g25725), .Z(g26928) ) ;
INV     gate14834  (.A(g26928), .Z(II35750) ) ;
INV     gate14835  (.A(II35750), .Z(g27410) ) ;
NAND2   gate14836  (.A(g26320), .B(g6448), .Z(g27117) ) ;
INV     gate14837  (.A(g27117), .Z(II35756) ) ;
INV     gate14838  (.A(II35756), .Z(g27416) ) ;
NAND2   gate14839  (.A(g26367), .B(g5473), .Z(g27121) ) ;
INV     gate14840  (.A(g27121), .Z(II35759) ) ;
INV     gate14841  (.A(II35759), .Z(g27419) ) ;
NAND4   gate14842  (.A(g25826), .B(g26374), .C(g25725), .D(g25781), .Z(g26918) ) ;
INV     gate14843  (.A(g26918), .Z(II35762) ) ;
INV     gate14844  (.A(II35762), .Z(g27422) ) ;
NAND3   gate14845  (.A(g25835), .B(g26417), .C(g25798), .Z(g26941) ) ;
INV     gate14846  (.A(g26941), .Z(II35768) ) ;
INV     gate14847  (.A(II35768), .Z(g27428) ) ;
NAND2   gate14848  (.A(g26320), .B(g3306), .Z(g26772) ) ;
INV     gate14849  (.A(g26772), .Z(II35772) ) ;
INV     gate14850  (.A(II35772), .Z(g27432) ) ;
NAND2   gate14851  (.A(g26367), .B(g6713), .Z(g27119) ) ;
INV     gate14852  (.A(g27119), .Z(II35777) ) ;
INV     gate14853  (.A(II35777), .Z(g27437) ) ;
NAND2   gate14854  (.A(g26410), .B(g5512), .Z(g27124) ) ;
INV     gate14855  (.A(g27124), .Z(II35780) ) ;
INV     gate14856  (.A(II35780), .Z(g27440) ) ;
NAND4   gate14857  (.A(g25861), .B(g26417), .C(g25798), .D(g25835), .Z(g26931) ) ;
INV     gate14858  (.A(g26931), .Z(II35783) ) ;
INV     gate14859  (.A(II35783), .Z(g27443) ) ;
INV     gate14860  (.A(g26837), .Z(g27449) ) ;
NAND2   gate14861  (.A(g26367), .B(g3462), .Z(g26779) ) ;
INV     gate14862  (.A(g26779), .Z(II35791) ) ;
INV     gate14863  (.A(II35791), .Z(g27451) ) ;
NAND2   gate14864  (.A(g26410), .B(g7015), .Z(g27122) ) ;
INV     gate14865  (.A(g27122), .Z(II35796) ) ;
INV     gate14866  (.A(II35796), .Z(g27456) ) ;
NAND2   gate14867  (.A(g26451), .B(g5556), .Z(g27130) ) ;
INV     gate14868  (.A(g27130), .Z(II35799) ) ;
INV     gate14869  (.A(II35799), .Z(g27459) ) ;
NOR2    gate14870  (.A(g15105), .B(g26213), .Z(g26803) ) ;
INV     gate14871  (.A(g26803), .Z(II35803) ) ;
INV     gate14872  (.A(II35803), .Z(g27463) ) ;
INV     gate14873  (.A(g26846), .Z(g27465) ) ;
NAND2   gate14874  (.A(g26410), .B(g3618), .Z(g26785) ) ;
INV     gate14875  (.A(g26785), .Z(II35809) ) ;
INV     gate14876  (.A(II35809), .Z(g27467) ) ;
NAND2   gate14877  (.A(g26451), .B(g7265), .Z(g27125) ) ;
INV     gate14878  (.A(g27125), .Z(II35814) ) ;
INV     gate14879  (.A(II35814), .Z(g27472) ) ;
INV     gate14880  (.A(g26922), .Z(II35817) ) ;
INV     gate14881  (.A(II35817), .Z(g27475) ) ;
NOR2    gate14882  (.A(g15172), .B(g26235), .Z(g26804) ) ;
INV     gate14883  (.A(g26804), .Z(II35821) ) ;
INV     gate14884  (.A(II35821), .Z(g27479) ) ;
NOR2    gate14885  (.A(g15173), .B(g26236), .Z(g26805) ) ;
INV     gate14886  (.A(g26805), .Z(II35824) ) ;
INV     gate14887  (.A(II35824), .Z(g27480) ) ;
NOR2    gate14888  (.A(g15197), .B(g26244), .Z(g26806) ) ;
INV     gate14889  (.A(g26806), .Z(II35829) ) ;
INV     gate14890  (.A(II35829), .Z(g27483) ) ;
INV     gate14891  (.A(g26855), .Z(g27484) ) ;
NAND2   gate14892  (.A(g26451), .B(g3774), .Z(g26792) ) ;
INV     gate14893  (.A(g26792), .Z(II35834) ) ;
INV     gate14894  (.A(II35834), .Z(g27486) ) ;
NAND2   gate14895  (.A(g25569), .B(g26283), .Z(g26911) ) ;
INV     gate14896  (.A(g26911), .Z(II35837) ) ;
INV     gate14897  (.A(II35837), .Z(g27489) ) ;
NOR2    gate14898  (.A(g15245), .B(g26261), .Z(g26807) ) ;
INV     gate14899  (.A(g26807), .Z(II35841) ) ;
INV     gate14900  (.A(II35841), .Z(g27493) ) ;
NOR2    gate14901  (.A(g15246), .B(g26262), .Z(g26808) ) ;
INV     gate14902  (.A(g26808), .Z(II35844) ) ;
INV     gate14903  (.A(II35844), .Z(g27494) ) ;
NOR2    gate14904  (.A(g26042), .B(g10024), .Z(g26776) ) ;
INV     gate14905  (.A(g26776), .Z(II35849) ) ;
INV     gate14906  (.A(II35849), .Z(g27497) ) ;
INV     gate14907  (.A(g26935), .Z(II35852) ) ;
INV     gate14908  (.A(II35852), .Z(g27498) ) ;
NOR2    gate14909  (.A(g15258), .B(g26270), .Z(g26809) ) ;
INV     gate14910  (.A(g26809), .Z(II35856) ) ;
INV     gate14911  (.A(II35856), .Z(g27502) ) ;
NOR2    gate14912  (.A(g15259), .B(g26271), .Z(g26810) ) ;
INV     gate14913  (.A(g26810), .Z(II35859) ) ;
INV     gate14914  (.A(II35859), .Z(g27503) ) ;
NOR2    gate14915  (.A(g15283), .B(g26279), .Z(g26811) ) ;
INV     gate14916  (.A(g26811), .Z(II35863) ) ;
INV     gate14917  (.A(II35863), .Z(g27505) ) ;
INV     gate14918  (.A(g26861), .Z(g27506) ) ;
NOR2    gate14919  (.A(g15321), .B(g26291), .Z(g26812) ) ;
INV     gate14920  (.A(g26812), .Z(II35868) ) ;
INV     gate14921  (.A(II35868), .Z(g27508) ) ;
NAND2   gate14922  (.A(g25648), .B(g26327), .Z(g26925) ) ;
INV     gate14923  (.A(g26925), .Z(II35872) ) ;
INV     gate14924  (.A(II35872), .Z(g27510) ) ;
NOR2    gate14925  (.A(g15337), .B(g26302), .Z(g26813) ) ;
INV     gate14926  (.A(g26813), .Z(II35876) ) ;
INV     gate14927  (.A(II35876), .Z(g27514) ) ;
NOR2    gate14928  (.A(g15338), .B(g26303), .Z(g26814) ) ;
INV     gate14929  (.A(g26814), .Z(II35879) ) ;
INV     gate14930  (.A(II35879), .Z(g27515) ) ;
NOR2    gate14931  (.A(g26044), .B(g10133), .Z(g26781) ) ;
INV     gate14932  (.A(g26781), .Z(II35883) ) ;
INV     gate14933  (.A(II35883), .Z(g27517) ) ;
INV     gate14934  (.A(g26944), .Z(II35886) ) ;
INV     gate14935  (.A(II35886), .Z(g27518) ) ;
NOR2    gate14936  (.A(g15350), .B(g26311), .Z(g26815) ) ;
INV     gate14937  (.A(g26815), .Z(II35890) ) ;
INV     gate14938  (.A(II35890), .Z(g27522) ) ;
NOR2    gate14939  (.A(g15351), .B(g26312), .Z(g26816) ) ;
INV     gate14940  (.A(g26816), .Z(II35893) ) ;
INV     gate14941  (.A(II35893), .Z(g27523) ) ;
NOR2    gate14942  (.A(g15375), .B(g26317), .Z(g26817) ) ;
INV     gate14943  (.A(g26817), .Z(II35897) ) ;
INV     gate14944  (.A(II35897), .Z(g27525) ) ;
NOR2    gate14945  (.A(g26049), .B(g22777), .Z(g26786) ) ;
INV     gate14946  (.A(g26786), .Z(II35900) ) ;
INV     gate14947  (.A(II35900), .Z(g27526) ) ;
NOR2    gate14948  (.A(g15407), .B(g26335), .Z(g26818) ) ;
INV     gate14949  (.A(g26818), .Z(II35915) ) ;
INV     gate14950  (.A(II35915), .Z(g27533) ) ;
NAND2   gate14951  (.A(g25725), .B(g26374), .Z(g26938) ) ;
INV     gate14952  (.A(g26938), .Z(II35919) ) ;
INV     gate14953  (.A(II35919), .Z(g27535) ) ;
NOR2    gate14954  (.A(g15423), .B(g26346), .Z(g26820) ) ;
INV     gate14955  (.A(g26820), .Z(II35923) ) ;
INV     gate14956  (.A(II35923), .Z(g27539) ) ;
NOR2    gate14957  (.A(g15424), .B(g26347), .Z(g26821) ) ;
INV     gate14958  (.A(g26821), .Z(II35926) ) ;
INV     gate14959  (.A(II35926), .Z(g27540) ) ;
NOR2    gate14960  (.A(g26046), .B(g10238), .Z(g26789) ) ;
INV     gate14961  (.A(g26789), .Z(II35930) ) ;
INV     gate14962  (.A(II35930), .Z(g27542) ) ;
INV     gate14963  (.A(g26950), .Z(II35933) ) ;
INV     gate14964  (.A(II35933), .Z(g27543) ) ;
NOR2    gate14965  (.A(g15436), .B(g26352), .Z(g26822) ) ;
INV     gate14966  (.A(g26822), .Z(II35937) ) ;
INV     gate14967  (.A(II35937), .Z(g27547) ) ;
NOR2    gate14968  (.A(g15437), .B(g26353), .Z(g26823) ) ;
INV     gate14969  (.A(g26823), .Z(II35940) ) ;
INV     gate14970  (.A(II35940), .Z(g27548) ) ;
NOR2    gate14971  (.A(g15491), .B(g26382), .Z(g26824) ) ;
INV     gate14972  (.A(g26824), .Z(II35953) ) ;
INV     gate14973  (.A(II35953), .Z(g27553) ) ;
NAND2   gate14974  (.A(g25798), .B(g26417), .Z(g26947) ) ;
INV     gate14975  (.A(g26947), .Z(II35957) ) ;
INV     gate14976  (.A(II35957), .Z(g27555) ) ;
NOR2    gate14977  (.A(g15507), .B(g26390), .Z(g26825) ) ;
INV     gate14978  (.A(g26825), .Z(II35961) ) ;
INV     gate14979  (.A(II35961), .Z(g27559) ) ;
NOR2    gate14980  (.A(g15508), .B(g26391), .Z(g26826) ) ;
INV     gate14981  (.A(g26826), .Z(II35964) ) ;
INV     gate14982  (.A(II35964), .Z(g27560) ) ;
NOR2    gate14983  (.A(g26050), .B(g10340), .Z(g26795) ) ;
INV     gate14984  (.A(g26795), .Z(II35968) ) ;
INV     gate14985  (.A(II35968), .Z(g27562) ) ;
NOR2    gate14986  (.A(g15577), .B(g26425), .Z(g26827) ) ;
INV     gate14987  (.A(g26827), .Z(II35983) ) ;
INV     gate14988  (.A(II35983), .Z(g27569) ) ;
NOR2    gate14989  (.A(g26055), .B(g18407), .Z(g26798) ) ;
INV     gate14990  (.A(g26798), .Z(II36008) ) ;
INV     gate14991  (.A(II36008), .Z(g27586) ) ;
INV     gate14992  (.A(g27168), .Z(g27589) ) ;
NOR2    gate14993  (.A(g23451), .B(g26052), .Z(g27144) ) ;
INV     gate14994  (.A(g27144), .Z(g27590) ) ;
NOR2    gate14995  (.A(g23462), .B(g26060), .Z(g27149) ) ;
INV     gate14996  (.A(g27149), .Z(g27595) ) ;
NOR2    gate14997  (.A(g23458), .B(g26054), .Z(g27147) ) ;
INV     gate14998  (.A(g27147), .Z(g27599) ) ;
NOR2    gate14999  (.A(g23471), .B(g26067), .Z(g27157) ) ;
INV     gate15000  (.A(g27157), .Z(g27604) ) ;
NOR2    gate15001  (.A(g23467), .B(g26062), .Z(g27152) ) ;
INV     gate15002  (.A(g27152), .Z(g27608) ) ;
NOR2    gate15003  (.A(g23484), .B(g26074), .Z(g27165) ) ;
INV     gate15004  (.A(g27165), .Z(g27613) ) ;
NOR2    gate15005  (.A(g23476), .B(g26069), .Z(g27160) ) ;
INV     gate15006  (.A(g27160), .Z(g27617) ) ;
NOR2    gate15007  (.A(g23494), .B(g26080), .Z(g27174) ) ;
INV     gate15008  (.A(g27174), .Z(g27622) ) ;
OR3     gate15009  (.A(g1248), .B(g1245), .C(g26534), .Z(g27113) ) ;
INV     gate15010  (.A(g27113), .Z(II36032) ) ;
INV     gate15011  (.A(II36032), .Z(g27632) ) ;
INV     gate15012  (.A(g26960), .Z(II36042) ) ;
INV     gate15013  (.A(II36042), .Z(g27662) ) ;
INV     gate15014  (.A(g26957), .Z(II36046) ) ;
INV     gate15015  (.A(II36046), .Z(g27667) ) ;
INV     gate15016  (.A(g26954), .Z(II36052) ) ;
INV     gate15017  (.A(II36052), .Z(g27674) ) ;
INV     gate15018  (.A(g27353), .Z(II36060) ) ;
INV     gate15019  (.A(g27463), .Z(II36063) ) ;
INV     gate15020  (.A(g27479), .Z(II36066) ) ;
INV     gate15021  (.A(g27493), .Z(II36069) ) ;
INV     gate15022  (.A(g27480), .Z(II36072) ) ;
INV     gate15023  (.A(g27494), .Z(II36075) ) ;
INV     gate15024  (.A(g27508), .Z(II36078) ) ;
INV     gate15025  (.A(g27497), .Z(II36081) ) ;
INV     gate15026  (.A(g27357), .Z(II36084) ) ;
INV     gate15027  (.A(g27483), .Z(II36087) ) ;
INV     gate15028  (.A(g27502), .Z(II36090) ) ;
INV     gate15029  (.A(g27514), .Z(II36093) ) ;
INV     gate15030  (.A(g27503), .Z(II36096) ) ;
INV     gate15031  (.A(g27515), .Z(II36099) ) ;
INV     gate15032  (.A(g27533), .Z(II36102) ) ;
INV     gate15033  (.A(g27517), .Z(II36105) ) ;
INV     gate15034  (.A(g27360), .Z(II36108) ) ;
INV     gate15035  (.A(g27505), .Z(II36111) ) ;
INV     gate15036  (.A(g27522), .Z(II36114) ) ;
INV     gate15037  (.A(g27539), .Z(II36117) ) ;
INV     gate15038  (.A(g27523), .Z(II36120) ) ;
INV     gate15039  (.A(g27540), .Z(II36123) ) ;
INV     gate15040  (.A(g27553), .Z(II36126) ) ;
INV     gate15041  (.A(g27542), .Z(II36129) ) ;
INV     gate15042  (.A(g27366), .Z(II36132) ) ;
INV     gate15043  (.A(g27525), .Z(II36135) ) ;
INV     gate15044  (.A(g27547), .Z(II36138) ) ;
INV     gate15045  (.A(g27559), .Z(II36141) ) ;
INV     gate15046  (.A(g27548), .Z(II36144) ) ;
INV     gate15047  (.A(g27560), .Z(II36147) ) ;
INV     gate15048  (.A(g27569), .Z(II36150) ) ;
INV     gate15049  (.A(g27562), .Z(II36153) ) ;
INV     gate15050  (.A(g27586), .Z(II36156) ) ;
INV     gate15051  (.A(g27526), .Z(II36159) ) ;
INV     gate15052  (.A(g27385), .Z(II36162) ) ;
INV     gate15053  (.A(g27632), .Z(g27748) ) ;
NAND2   gate15054  (.A(g26869), .B(g56), .Z(g27571) ) ;
INV     gate15055  (.A(g27571), .Z(II36213) ) ;
INV     gate15056  (.A(II36213), .Z(g27776) ) ;
NAND2   gate15057  (.A(g26878), .B(g744), .Z(g27580) ) ;
INV     gate15058  (.A(g27580), .Z(II36217) ) ;
INV     gate15059  (.A(II36217), .Z(g27780) ) ;
INV     gate15060  (.A(g27662), .Z(II36221) ) ;
INV     gate15061  (.A(II36221), .Z(g27784) ) ;
INV     gate15062  (.A(g27589), .Z(II36224) ) ;
INV     gate15063  (.A(II36224), .Z(g27785) ) ;
NOR2    gate15064  (.A(g27175), .B(g17001), .Z(g27594) ) ;
INV     gate15065  (.A(g27594), .Z(II36227) ) ;
INV     gate15066  (.A(II36227), .Z(g27786) ) ;
NAND2   gate15067  (.A(g26887), .B(g1430), .Z(g27583) ) ;
INV     gate15068  (.A(g27583), .Z(II36230) ) ;
INV     gate15069  (.A(II36230), .Z(g27787) ) ;
INV     gate15070  (.A(g27667), .Z(II36234) ) ;
INV     gate15071  (.A(II36234), .Z(g27791) ) ;
INV     gate15072  (.A(g27662), .Z(II36237) ) ;
INV     gate15073  (.A(II36237), .Z(g27792) ) ;
NOR2    gate15074  (.A(g27179), .B(g17031), .Z(g27603) ) ;
INV     gate15075  (.A(g27603), .Z(II36240) ) ;
INV     gate15076  (.A(II36240), .Z(g27793) ) ;
NAND2   gate15077  (.A(g26897), .B(g2124), .Z(g27587) ) ;
INV     gate15078  (.A(g27587), .Z(II36243) ) ;
INV     gate15079  (.A(II36243), .Z(g27794) ) ;
INV     gate15080  (.A(g27674), .Z(II36246) ) ;
INV     gate15081  (.A(II36246), .Z(g27797) ) ;
NOR2    gate15082  (.A(g27184), .B(g17065), .Z(g27612) ) ;
INV     gate15083  (.A(g27612), .Z(II36250) ) ;
INV     gate15084  (.A(II36250), .Z(g27799) ) ;
INV     gate15085  (.A(g27674), .Z(II36253) ) ;
INV     gate15086  (.A(II36253), .Z(g27800) ) ;
NOR2    gate15087  (.A(g27188), .B(g17100), .Z(g27621) ) ;
INV     gate15088  (.A(g27621), .Z(II36264) ) ;
INV     gate15089  (.A(II36264), .Z(g27805) ) ;
NAND2   gate15090  (.A(g26989), .B(g5438), .Z(g27395) ) ;
INV     gate15091  (.A(g27395), .Z(II36267) ) ;
INV     gate15092  (.A(II36267), .Z(g27806) ) ;
NAND2   gate15093  (.A(g26989), .B(g6448), .Z(g27390) ) ;
INV     gate15094  (.A(g27390), .Z(II36280) ) ;
INV     gate15095  (.A(II36280), .Z(g27817) ) ;
NAND2   gate15096  (.A(g27012), .B(g5473), .Z(g27408) ) ;
INV     gate15097  (.A(g27408), .Z(II36283) ) ;
INV     gate15098  (.A(II36283), .Z(g27820) ) ;
NAND2   gate15099  (.A(g26989), .B(g3306), .Z(g27626) ) ;
INV     gate15100  (.A(g27626), .Z(II36296) ) ;
INV     gate15101  (.A(II36296), .Z(g27831) ) ;
NAND2   gate15102  (.A(g27012), .B(g6713), .Z(g27400) ) ;
INV     gate15103  (.A(g27400), .Z(II36307) ) ;
INV     gate15104  (.A(II36307), .Z(g27839) ) ;
NAND2   gate15105  (.A(g27038), .B(g5512), .Z(g27426) ) ;
INV     gate15106  (.A(g27426), .Z(II36311) ) ;
INV     gate15107  (.A(II36311), .Z(g27843) ) ;
NAND2   gate15108  (.A(g27012), .B(g3462), .Z(g27627) ) ;
INV     gate15109  (.A(g27627), .Z(II36321) ) ;
INV     gate15110  (.A(II36321), .Z(g27847) ) ;
NAND2   gate15111  (.A(g27038), .B(g7015), .Z(g27413) ) ;
INV     gate15112  (.A(g27413), .Z(II36327) ) ;
INV     gate15113  (.A(II36327), .Z(g27858) ) ;
NAND2   gate15114  (.A(g27066), .B(g5556), .Z(g27447) ) ;
INV     gate15115  (.A(g27447), .Z(II36330) ) ;
INV     gate15116  (.A(II36330), .Z(g27861) ) ;
NAND2   gate15117  (.A(g27038), .B(g3618), .Z(g27628) ) ;
INV     gate15118  (.A(g27628), .Z(II36337) ) ;
INV     gate15119  (.A(II36337), .Z(g27872) ) ;
NAND2   gate15120  (.A(g27066), .B(g7265), .Z(g27431) ) ;
INV     gate15121  (.A(g27431), .Z(II36341) ) ;
INV     gate15122  (.A(II36341), .Z(g27879) ) ;
NAND2   gate15123  (.A(g27066), .B(g3774), .Z(g27630) ) ;
INV     gate15124  (.A(g27630), .Z(II36347) ) ;
INV     gate15125  (.A(II36347), .Z(g27889) ) ;
INV     gate15126  (.A(g27662), .Z(II36354) ) ;
INV     gate15127  (.A(II36354), .Z(g27903) ) ;
NOR2    gate15128  (.A(g26799), .B(g10024), .Z(g27672) ) ;
INV     gate15129  (.A(g27672), .Z(II36358) ) ;
INV     gate15130  (.A(II36358), .Z(g27905) ) ;
INV     gate15131  (.A(g27667), .Z(II36362) ) ;
INV     gate15132  (.A(II36362), .Z(g27907) ) ;
NOR2    gate15133  (.A(g26800), .B(g10133), .Z(g27678) ) ;
INV     gate15134  (.A(g27678), .Z(II36367) ) ;
INV     gate15135  (.A(II36367), .Z(g27910) ) ;
INV     gate15136  (.A(g27674), .Z(II36371) ) ;
INV     gate15137  (.A(II36371), .Z(g27912) ) ;
NOR2    gate15138  (.A(g26801), .B(g10238), .Z(g27682) ) ;
INV     gate15139  (.A(g27682), .Z(II36379) ) ;
INV     gate15140  (.A(II36379), .Z(g27918) ) ;
NOR2    gate15141  (.A(g26922), .B(g24708), .Z(g27563) ) ;
INV     gate15142  (.A(g27563), .Z(II36382) ) ;
INV     gate15143  (.A(II36382), .Z(g27919) ) ;
NOR2    gate15144  (.A(g26802), .B(g10340), .Z(g27243) ) ;
INV     gate15145  (.A(g27243), .Z(II36390) ) ;
INV     gate15146  (.A(II36390), .Z(g27927) ) ;
NOR2    gate15147  (.A(g26911), .B(g24717), .Z(g27572) ) ;
INV     gate15148  (.A(g27572), .Z(II36393) ) ;
INV     gate15149  (.A(II36393), .Z(g27928) ) ;
NOR2    gate15150  (.A(g26935), .B(g24720), .Z(g27574) ) ;
INV     gate15151  (.A(g27574), .Z(II36397) ) ;
INV     gate15152  (.A(II36397), .Z(g27932) ) ;
NOR2    gate15153  (.A(g26902), .B(g24613), .Z(g27450) ) ;
INV     gate15154  (.A(g27450), .Z(II36404) ) ;
INV     gate15155  (.A(II36404), .Z(g27939) ) ;
NOR2    gate15156  (.A(g26925), .B(g24728), .Z(g27581) ) ;
INV     gate15157  (.A(g27581), .Z(II36407) ) ;
INV     gate15158  (.A(II36407), .Z(g27942) ) ;
NOR2    gate15159  (.A(g26944), .B(g24731), .Z(g27582) ) ;
INV     gate15160  (.A(g27582), .Z(II36411) ) ;
INV     gate15161  (.A(II36411), .Z(g27946) ) ;
NOR2    gate15162  (.A(g26892), .B(g24622), .Z(g27462) ) ;
INV     gate15163  (.A(g27462), .Z(II36417) ) ;
INV     gate15164  (.A(II36417), .Z(g27952) ) ;
NOR2    gate15165  (.A(g26965), .B(g26212), .Z(g27253) ) ;
INV     gate15166  (.A(g27253), .Z(II36420) ) ;
INV     gate15167  (.A(II36420), .Z(g27955) ) ;
NOR2    gate15168  (.A(g26915), .B(g24624), .Z(g27466) ) ;
INV     gate15169  (.A(g27466), .Z(II36423) ) ;
INV     gate15170  (.A(II36423), .Z(g27956) ) ;
NOR2    gate15171  (.A(g26938), .B(g24736), .Z(g27584) ) ;
INV     gate15172  (.A(g27584), .Z(II36426) ) ;
INV     gate15173  (.A(II36426), .Z(g27959) ) ;
NOR2    gate15174  (.A(g26950), .B(g24739), .Z(g27585) ) ;
INV     gate15175  (.A(g27585), .Z(II36432) ) ;
INV     gate15176  (.A(II36432), .Z(g27965) ) ;
INV     gate15177  (.A(g27361), .Z(g27969) ) ;
NOR2    gate15178  (.A(g26969), .B(g26233), .Z(g27255) ) ;
INV     gate15179  (.A(g27255), .Z(II36438) ) ;
INV     gate15180  (.A(II36438), .Z(g27971) ) ;
NOR2    gate15181  (.A(g26970), .B(g26234), .Z(g27256) ) ;
INV     gate15182  (.A(g27256), .Z(II36441) ) ;
INV     gate15183  (.A(II36441), .Z(g27972) ) ;
NOR2    gate15184  (.A(g26906), .B(g24637), .Z(g27482) ) ;
INV     gate15185  (.A(g27482), .Z(II36444) ) ;
INV     gate15186  (.A(II36444), .Z(g27973) ) ;
NOR2    gate15187  (.A(g26971), .B(g26243), .Z(g27257) ) ;
INV     gate15188  (.A(g27257), .Z(II36447) ) ;
INV     gate15189  (.A(II36447), .Z(g27976) ) ;
NOR2    gate15190  (.A(g26928), .B(g24638), .Z(g27485) ) ;
INV     gate15191  (.A(g27485), .Z(II36450) ) ;
INV     gate15192  (.A(II36450), .Z(g27977) ) ;
NOR2    gate15193  (.A(g26947), .B(g24742), .Z(g27588) ) ;
INV     gate15194  (.A(g27588), .Z(II36454) ) ;
INV     gate15195  (.A(II36454), .Z(g27981) ) ;
NOR2    gate15196  (.A(g26977), .B(g26257), .Z(g27258) ) ;
INV     gate15197  (.A(g27258), .Z(II36459) ) ;
INV     gate15198  (.A(II36459), .Z(g27986) ) ;
NOR2    gate15199  (.A(g26978), .B(g26258), .Z(g27259) ) ;
INV     gate15200  (.A(g27259), .Z(II36462) ) ;
INV     gate15201  (.A(II36462), .Z(g27987) ) ;
NOR2    gate15202  (.A(g26979), .B(g26259), .Z(g27260) ) ;
INV     gate15203  (.A(g27260), .Z(II36465) ) ;
INV     gate15204  (.A(II36465), .Z(g27988) ) ;
NOR2    gate15205  (.A(g26980), .B(g26263), .Z(g27261) ) ;
INV     gate15206  (.A(g27261), .Z(II36468) ) ;
INV     gate15207  (.A(II36468), .Z(g27989) ) ;
INV     gate15208  (.A(g27367), .Z(g27990) ) ;
NOR2    gate15209  (.A(g26981), .B(g26268), .Z(g27262) ) ;
INV     gate15210  (.A(g27262), .Z(II36473) ) ;
INV     gate15211  (.A(II36473), .Z(g27992) ) ;
NOR2    gate15212  (.A(g26982), .B(g26269), .Z(g27263) ) ;
INV     gate15213  (.A(g27263), .Z(II36476) ) ;
INV     gate15214  (.A(II36476), .Z(g27993) ) ;
NOR2    gate15215  (.A(g26918), .B(g24656), .Z(g27504) ) ;
INV     gate15216  (.A(g27504), .Z(II36479) ) ;
INV     gate15217  (.A(II36479), .Z(g27994) ) ;
NOR2    gate15218  (.A(g26984), .B(g26278), .Z(g27264) ) ;
INV     gate15219  (.A(g27264), .Z(II36483) ) ;
INV     gate15220  (.A(II36483), .Z(g27998) ) ;
NOR2    gate15221  (.A(g26941), .B(g24657), .Z(g27507) ) ;
INV     gate15222  (.A(g27507), .Z(II36486) ) ;
INV     gate15223  (.A(II36486), .Z(g27999) ) ;
NOR2    gate15224  (.A(g26993), .B(g26288), .Z(g27265) ) ;
INV     gate15225  (.A(g27265), .Z(II36490) ) ;
INV     gate15226  (.A(II36490), .Z(g28003) ) ;
NOR2    gate15227  (.A(g26994), .B(g26289), .Z(g27266) ) ;
INV     gate15228  (.A(g27266), .Z(II36493) ) ;
INV     gate15229  (.A(II36493), .Z(g28004) ) ;
NOR2    gate15230  (.A(g26995), .B(g26290), .Z(g27267) ) ;
INV     gate15231  (.A(g27267), .Z(II36496) ) ;
INV     gate15232  (.A(II36496), .Z(g28005) ) ;
NOR2    gate15233  (.A(g26996), .B(g26292), .Z(g27268) ) ;
INV     gate15234  (.A(g27268), .Z(II36499) ) ;
INV     gate15235  (.A(II36499), .Z(g28006) ) ;
NOR2    gate15236  (.A(g26997), .B(g26293), .Z(g27269) ) ;
INV     gate15237  (.A(g27269), .Z(II36502) ) ;
INV     gate15238  (.A(II36502), .Z(g28007) ) ;
NOR2    gate15239  (.A(g26998), .B(g26298), .Z(g27270) ) ;
INV     gate15240  (.A(g27270), .Z(II36507) ) ;
INV     gate15241  (.A(II36507), .Z(g28010) ) ;
NOR2    gate15242  (.A(g26999), .B(g26299), .Z(g27271) ) ;
INV     gate15243  (.A(g27271), .Z(II36510) ) ;
INV     gate15244  (.A(II36510), .Z(g28011) ) ;
NOR2    gate15245  (.A(g27000), .B(g26300), .Z(g27272) ) ;
INV     gate15246  (.A(g27272), .Z(II36513) ) ;
INV     gate15247  (.A(II36513), .Z(g28012) ) ;
NOR2    gate15248  (.A(g27001), .B(g26307), .Z(g27273) ) ;
INV     gate15249  (.A(g27273), .Z(II36516) ) ;
INV     gate15250  (.A(II36516), .Z(g28013) ) ;
INV     gate15251  (.A(g27373), .Z(g28014) ) ;
NOR2    gate15252  (.A(g27002), .B(g26309), .Z(g27274) ) ;
INV     gate15253  (.A(g27274), .Z(II36521) ) ;
INV     gate15254  (.A(II36521), .Z(g28016) ) ;
NOR2    gate15255  (.A(g27003), .B(g26310), .Z(g27275) ) ;
INV     gate15256  (.A(g27275), .Z(II36524) ) ;
INV     gate15257  (.A(II36524), .Z(g28017) ) ;
NOR2    gate15258  (.A(g26931), .B(g24675), .Z(g27524) ) ;
INV     gate15259  (.A(g27524), .Z(II36527) ) ;
INV     gate15260  (.A(II36527), .Z(g28018) ) ;
NOR2    gate15261  (.A(g27004), .B(g26316), .Z(g27276) ) ;
INV     gate15262  (.A(g27276), .Z(II36530) ) ;
INV     gate15263  (.A(II36530), .Z(g28021) ) ;
NOR2    gate15264  (.A(g27005), .B(g26318), .Z(g27277) ) ;
INV     gate15265  (.A(g27277), .Z(II36533) ) ;
INV     gate15266  (.A(II36533), .Z(g28022) ) ;
NOR2    gate15267  (.A(g27006), .B(g26319), .Z(g27278) ) ;
INV     gate15268  (.A(g27278), .Z(II36536) ) ;
INV     gate15269  (.A(II36536), .Z(g28023) ) ;
NOR2    gate15270  (.A(g27007), .B(g26324), .Z(g27279) ) ;
INV     gate15271  (.A(g27279), .Z(II36539) ) ;
INV     gate15272  (.A(II36539), .Z(g28024) ) ;
NOR2    gate15273  (.A(g27008), .B(g26325), .Z(g27280) ) ;
INV     gate15274  (.A(g27280), .Z(II36542) ) ;
INV     gate15275  (.A(II36542), .Z(g28025) ) ;
NOR2    gate15276  (.A(g27009), .B(g26326), .Z(g27281) ) ;
INV     gate15277  (.A(g27281), .Z(II36545) ) ;
INV     gate15278  (.A(II36545), .Z(g28026) ) ;
NOR2    gate15279  (.A(g27016), .B(g26332), .Z(g27282) ) ;
INV     gate15280  (.A(g27282), .Z(II36551) ) ;
INV     gate15281  (.A(II36551), .Z(g28030) ) ;
NOR2    gate15282  (.A(g27017), .B(g26333), .Z(g27283) ) ;
INV     gate15283  (.A(g27283), .Z(II36554) ) ;
INV     gate15284  (.A(II36554), .Z(g28031) ) ;
NOR2    gate15285  (.A(g27018), .B(g26334), .Z(g27284) ) ;
INV     gate15286  (.A(g27284), .Z(II36557) ) ;
INV     gate15287  (.A(II36557), .Z(g28032) ) ;
NOR2    gate15288  (.A(g27019), .B(g26339), .Z(g27285) ) ;
INV     gate15289  (.A(g27285), .Z(II36560) ) ;
INV     gate15290  (.A(II36560), .Z(g28033) ) ;
NOR2    gate15291  (.A(g27020), .B(g26340), .Z(g27286) ) ;
INV     gate15292  (.A(g27286), .Z(II36563) ) ;
INV     gate15293  (.A(II36563), .Z(g28034) ) ;
NOR2    gate15294  (.A(g27021), .B(g26342), .Z(g27287) ) ;
INV     gate15295  (.A(g27287), .Z(II36568) ) ;
INV     gate15296  (.A(II36568), .Z(g28037) ) ;
NOR2    gate15297  (.A(g27022), .B(g26343), .Z(g27288) ) ;
INV     gate15298  (.A(g27288), .Z(II36571) ) ;
INV     gate15299  (.A(II36571), .Z(g28038) ) ;
NOR2    gate15300  (.A(g27023), .B(g26344), .Z(g27289) ) ;
INV     gate15301  (.A(g27289), .Z(II36574) ) ;
INV     gate15302  (.A(II36574), .Z(g28039) ) ;
NOR2    gate15303  (.A(g27024), .B(g26348), .Z(g27290) ) ;
INV     gate15304  (.A(g27290), .Z(II36577) ) ;
INV     gate15305  (.A(II36577), .Z(g28040) ) ;
INV     gate15306  (.A(g27376), .Z(g28041) ) ;
NOR2    gate15307  (.A(g27025), .B(g26350), .Z(g27291) ) ;
INV     gate15308  (.A(g27291), .Z(II36582) ) ;
INV     gate15309  (.A(II36582), .Z(g28043) ) ;
NOR2    gate15310  (.A(g27026), .B(g26351), .Z(g27292) ) ;
INV     gate15311  (.A(g27292), .Z(II36585) ) ;
INV     gate15312  (.A(II36585), .Z(g28044) ) ;
NOR2    gate15313  (.A(g27027), .B(g26357), .Z(g27293) ) ;
INV     gate15314  (.A(g27293), .Z(II36588) ) ;
INV     gate15315  (.A(II36588), .Z(g28045) ) ;
NOR2    gate15316  (.A(g27028), .B(g26361), .Z(g27294) ) ;
INV     gate15317  (.A(g27294), .Z(II36598) ) ;
INV     gate15318  (.A(II36598), .Z(g28047) ) ;
NOR2    gate15319  (.A(g27029), .B(g26362), .Z(g27295) ) ;
INV     gate15320  (.A(g27295), .Z(II36601) ) ;
INV     gate15321  (.A(II36601), .Z(g28048) ) ;
NOR2    gate15322  (.A(g27030), .B(g26363), .Z(g27296) ) ;
INV     gate15323  (.A(g27296), .Z(II36604) ) ;
INV     gate15324  (.A(II36604), .Z(g28049) ) ;
NOR2    gate15325  (.A(g27031), .B(g26365), .Z(g27297) ) ;
INV     gate15326  (.A(g27297), .Z(II36609) ) ;
INV     gate15327  (.A(II36609), .Z(g28052) ) ;
NOR2    gate15328  (.A(g27032), .B(g26366), .Z(g27298) ) ;
INV     gate15329  (.A(g27298), .Z(II36612) ) ;
INV     gate15330  (.A(II36612), .Z(g28053) ) ;
NOR2    gate15331  (.A(g27033), .B(g26371), .Z(g27299) ) ;
INV     gate15332  (.A(g27299), .Z(II36615) ) ;
INV     gate15333  (.A(II36615), .Z(g28054) ) ;
NOR2    gate15334  (.A(g27034), .B(g26372), .Z(g27300) ) ;
INV     gate15335  (.A(g27300), .Z(II36618) ) ;
INV     gate15336  (.A(II36618), .Z(g28055) ) ;
NOR2    gate15337  (.A(g27035), .B(g26373), .Z(g27301) ) ;
INV     gate15338  (.A(g27301), .Z(II36621) ) ;
INV     gate15339  (.A(II36621), .Z(g28056) ) ;
NOR2    gate15340  (.A(g27042), .B(g26379), .Z(g27302) ) ;
INV     gate15341  (.A(g27302), .Z(II36627) ) ;
INV     gate15342  (.A(II36627), .Z(g28060) ) ;
NOR2    gate15343  (.A(g27043), .B(g26380), .Z(g27303) ) ;
INV     gate15344  (.A(g27303), .Z(II36630) ) ;
INV     gate15345  (.A(II36630), .Z(g28061) ) ;
NOR2    gate15346  (.A(g27044), .B(g26381), .Z(g27304) ) ;
INV     gate15347  (.A(g27304), .Z(II36633) ) ;
INV     gate15348  (.A(II36633), .Z(g28062) ) ;
NOR2    gate15349  (.A(g27045), .B(g26383), .Z(g27305) ) ;
INV     gate15350  (.A(g27305), .Z(II36636) ) ;
INV     gate15351  (.A(II36636), .Z(g28063) ) ;
NOR2    gate15352  (.A(g27046), .B(g26384), .Z(g27306) ) ;
INV     gate15353  (.A(g27306), .Z(II36639) ) ;
INV     gate15354  (.A(II36639), .Z(g28064) ) ;
NOR2    gate15355  (.A(g27047), .B(g26386), .Z(g27307) ) ;
INV     gate15356  (.A(g27307), .Z(II36644) ) ;
INV     gate15357  (.A(II36644), .Z(g28067) ) ;
NOR2    gate15358  (.A(g27048), .B(g26387), .Z(g27308) ) ;
INV     gate15359  (.A(g27308), .Z(II36647) ) ;
INV     gate15360  (.A(II36647), .Z(g28068) ) ;
NOR2    gate15361  (.A(g27049), .B(g26388), .Z(g27309) ) ;
INV     gate15362  (.A(g27309), .Z(II36650) ) ;
INV     gate15363  (.A(II36650), .Z(g28069) ) ;
NOR2    gate15364  (.A(g27050), .B(g26392), .Z(g27310) ) ;
INV     gate15365  (.A(g27310), .Z(II36653) ) ;
INV     gate15366  (.A(II36653), .Z(g28070) ) ;
NOR2    gate15367  (.A(g27053), .B(g26396), .Z(g27311) ) ;
INV     gate15368  (.A(g27311), .Z(II36656) ) ;
INV     gate15369  (.A(II36656), .Z(g28071) ) ;
NOR2    gate15370  (.A(g27054), .B(g26397), .Z(g27312) ) ;
INV     gate15371  (.A(g27312), .Z(II36659) ) ;
INV     gate15372  (.A(II36659), .Z(g28072) ) ;
NOR2    gate15373  (.A(g27055), .B(g26400), .Z(g27313) ) ;
INV     gate15374  (.A(g27313), .Z(II36663) ) ;
INV     gate15375  (.A(II36663), .Z(g28074) ) ;
NOR2    gate15376  (.A(g27056), .B(g26404), .Z(g27314) ) ;
INV     gate15377  (.A(g27314), .Z(II36673) ) ;
INV     gate15378  (.A(II36673), .Z(g28076) ) ;
NOR2    gate15379  (.A(g27057), .B(g26405), .Z(g27315) ) ;
INV     gate15380  (.A(g27315), .Z(II36676) ) ;
INV     gate15381  (.A(II36676), .Z(g28077) ) ;
NOR2    gate15382  (.A(g27058), .B(g26406), .Z(g27316) ) ;
INV     gate15383  (.A(g27316), .Z(II36679) ) ;
INV     gate15384  (.A(II36679), .Z(g28078) ) ;
NOR2    gate15385  (.A(g27059), .B(g26408), .Z(g27317) ) ;
INV     gate15386  (.A(g27317), .Z(II36684) ) ;
INV     gate15387  (.A(II36684), .Z(g28081) ) ;
NOR2    gate15388  (.A(g27060), .B(g26409), .Z(g27318) ) ;
INV     gate15389  (.A(g27318), .Z(II36687) ) ;
INV     gate15390  (.A(II36687), .Z(g28082) ) ;
NOR2    gate15391  (.A(g27061), .B(g26414), .Z(g27319) ) ;
INV     gate15392  (.A(g27319), .Z(II36690) ) ;
INV     gate15393  (.A(II36690), .Z(g28083) ) ;
NOR2    gate15394  (.A(g27062), .B(g26415), .Z(g27320) ) ;
INV     gate15395  (.A(g27320), .Z(II36693) ) ;
INV     gate15396  (.A(II36693), .Z(g28084) ) ;
NOR2    gate15397  (.A(g27063), .B(g26416), .Z(g27321) ) ;
INV     gate15398  (.A(g27321), .Z(II36696) ) ;
INV     gate15399  (.A(II36696), .Z(g28085) ) ;
NOR2    gate15400  (.A(g27070), .B(g26422), .Z(g27322) ) ;
INV     gate15401  (.A(g27322), .Z(II36702) ) ;
INV     gate15402  (.A(II36702), .Z(g28089) ) ;
NOR2    gate15403  (.A(g27071), .B(g26423), .Z(g27323) ) ;
INV     gate15404  (.A(g27323), .Z(II36705) ) ;
INV     gate15405  (.A(II36705), .Z(g28090) ) ;
NOR2    gate15406  (.A(g27072), .B(g26424), .Z(g27324) ) ;
INV     gate15407  (.A(g27324), .Z(II36708) ) ;
INV     gate15408  (.A(II36708), .Z(g28091) ) ;
NOR2    gate15409  (.A(g27073), .B(g26426), .Z(g27325) ) ;
INV     gate15410  (.A(g27325), .Z(II36711) ) ;
INV     gate15411  (.A(II36711), .Z(g28092) ) ;
NOR2    gate15412  (.A(g27074), .B(g26427), .Z(g27326) ) ;
INV     gate15413  (.A(g27326), .Z(II36714) ) ;
INV     gate15414  (.A(II36714), .Z(g28093) ) ;
NOR2    gate15415  (.A(g27077), .B(g26432), .Z(g27327) ) ;
INV     gate15416  (.A(g27327), .Z(II36718) ) ;
INV     gate15417  (.A(II36718), .Z(g28095) ) ;
NOR2    gate15418  (.A(g27080), .B(g26437), .Z(g27328) ) ;
INV     gate15419  (.A(g27328), .Z(II36721) ) ;
INV     gate15420  (.A(II36721), .Z(g28096) ) ;
NOR2    gate15421  (.A(g27081), .B(g26438), .Z(g27329) ) ;
INV     gate15422  (.A(g27329), .Z(II36724) ) ;
INV     gate15423  (.A(II36724), .Z(g28097) ) ;
NOR2    gate15424  (.A(g27082), .B(g26441), .Z(g27330) ) ;
INV     gate15425  (.A(g27330), .Z(II36728) ) ;
INV     gate15426  (.A(II36728), .Z(g28099) ) ;
NOR2    gate15427  (.A(g27083), .B(g26445), .Z(g27331) ) ;
INV     gate15428  (.A(g27331), .Z(II36738) ) ;
INV     gate15429  (.A(II36738), .Z(g28101) ) ;
NOR2    gate15430  (.A(g27084), .B(g26446), .Z(g27332) ) ;
INV     gate15431  (.A(g27332), .Z(II36741) ) ;
INV     gate15432  (.A(II36741), .Z(g28102) ) ;
NOR2    gate15433  (.A(g27085), .B(g26447), .Z(g27333) ) ;
INV     gate15434  (.A(g27333), .Z(II36744) ) ;
INV     gate15435  (.A(II36744), .Z(g28103) ) ;
NOR2    gate15436  (.A(g27086), .B(g26449), .Z(g27334) ) ;
INV     gate15437  (.A(g27334), .Z(II36749) ) ;
INV     gate15438  (.A(II36749), .Z(g28106) ) ;
NOR2    gate15439  (.A(g27087), .B(g26450), .Z(g27335) ) ;
INV     gate15440  (.A(g27335), .Z(II36752) ) ;
INV     gate15441  (.A(II36752), .Z(g28107) ) ;
NOR2    gate15442  (.A(g27088), .B(g26455), .Z(g27336) ) ;
INV     gate15443  (.A(g27336), .Z(II36755) ) ;
INV     gate15444  (.A(II36755), .Z(g28108) ) ;
NOR2    gate15445  (.A(g27089), .B(g26456), .Z(g27337) ) ;
INV     gate15446  (.A(g27337), .Z(II36758) ) ;
INV     gate15447  (.A(II36758), .Z(g28109) ) ;
NOR2    gate15448  (.A(g27090), .B(g26457), .Z(g27338) ) ;
INV     gate15449  (.A(g27338), .Z(II36761) ) ;
INV     gate15450  (.A(II36761), .Z(g28110) ) ;
NOR2    gate15451  (.A(g27093), .B(g26464), .Z(g27339) ) ;
INV     gate15452  (.A(g27339), .Z(II36766) ) ;
INV     gate15453  (.A(II36766), .Z(g28113) ) ;
NOR2    gate15454  (.A(g27096), .B(g26469), .Z(g27340) ) ;
INV     gate15455  (.A(g27340), .Z(II36769) ) ;
INV     gate15456  (.A(II36769), .Z(g28114) ) ;
NOR2    gate15457  (.A(g27097), .B(g26470), .Z(g27341) ) ;
INV     gate15458  (.A(g27341), .Z(II36772) ) ;
INV     gate15459  (.A(II36772), .Z(g28115) ) ;
NOR2    gate15460  (.A(g27098), .B(g26473), .Z(g27342) ) ;
INV     gate15461  (.A(g27342), .Z(II36776) ) ;
INV     gate15462  (.A(II36776), .Z(g28117) ) ;
NOR2    gate15463  (.A(g27099), .B(g26477), .Z(g27343) ) ;
INV     gate15464  (.A(g27343), .Z(II36786) ) ;
INV     gate15465  (.A(II36786), .Z(g28119) ) ;
NOR2    gate15466  (.A(g27100), .B(g26478), .Z(g27344) ) ;
INV     gate15467  (.A(g27344), .Z(II36789) ) ;
INV     gate15468  (.A(II36789), .Z(g28120) ) ;
NOR2    gate15469  (.A(g27101), .B(g26479), .Z(g27345) ) ;
INV     gate15470  (.A(g27345), .Z(II36792) ) ;
INV     gate15471  (.A(II36792), .Z(g28121) ) ;
NOR2    gate15472  (.A(g27105), .B(g26488), .Z(g27346) ) ;
INV     gate15473  (.A(g27346), .Z(II36797) ) ;
INV     gate15474  (.A(II36797), .Z(g28124) ) ;
NOR2    gate15475  (.A(g27108), .B(g26493), .Z(g27347) ) ;
INV     gate15476  (.A(g27347), .Z(II36800) ) ;
INV     gate15477  (.A(II36800), .Z(g28125) ) ;
NOR2    gate15478  (.A(g27109), .B(g26494), .Z(g27348) ) ;
INV     gate15479  (.A(g27348), .Z(II36803) ) ;
INV     gate15480  (.A(II36803), .Z(g28126) ) ;
NAND2   gate15481  (.A(II35905), .B(II35906), .Z(g27528) ) ;
INV     gate15482  (.A(g27528), .Z(g28128) ) ;
NOR2    gate15483  (.A(g27112), .B(g26504), .Z(g27354) ) ;
INV     gate15484  (.A(g27354), .Z(II36808) ) ;
INV     gate15485  (.A(II36808), .Z(g28132) ) ;
NAND2   gate15486  (.A(II35945), .B(II35946), .Z(g27550) ) ;
INV     gate15487  (.A(g27550), .Z(g28133) ) ;
NAND2   gate15488  (.A(II35975), .B(II35976), .Z(g27566) ) ;
INV     gate15489  (.A(g27566), .Z(g28137) ) ;
NAND2   gate15490  (.A(II35993), .B(II35994), .Z(g27576) ) ;
INV     gate15491  (.A(g27576), .Z(g28141) ) ;
INV     gate15492  (.A(g27667), .Z(g28149) ) ;
INV     gate15493  (.A(g27387), .Z(g28150) ) ;
INV     gate15494  (.A(g27381), .Z(g28151) ) ;
INV     gate15495  (.A(g27391), .Z(g28152) ) ;
INV     gate15496  (.A(g27397), .Z(g28153) ) ;
INV     gate15497  (.A(g27401), .Z(g28154) ) ;
INV     gate15498  (.A(g27404), .Z(g28155) ) ;
INV     gate15499  (.A(g27410), .Z(g28156) ) ;
INV     gate15500  (.A(g27416), .Z(g28158) ) ;
INV     gate15501  (.A(g27419), .Z(g28159) ) ;
INV     gate15502  (.A(g27422), .Z(g28160) ) ;
INV     gate15503  (.A(g27428), .Z(g28161) ) ;
INV     gate15504  (.A(g27432), .Z(g28162) ) ;
INV     gate15505  (.A(g27437), .Z(g28163) ) ;
INV     gate15506  (.A(g27440), .Z(g28164) ) ;
INV     gate15507  (.A(g27443), .Z(g28165) ) ;
INV     gate15508  (.A(g27451), .Z(g28166) ) ;
INV     gate15509  (.A(g27456), .Z(g28167) ) ;
INV     gate15510  (.A(g27459), .Z(g28168) ) ;
INV     gate15511  (.A(g27467), .Z(g28169) ) ;
INV     gate15512  (.A(g27472), .Z(g28170) ) ;
INV     gate15513  (.A(g27475), .Z(g28172) ) ;
INV     gate15514  (.A(g27486), .Z(g28173) ) ;
INV     gate15515  (.A(g27489), .Z(g28174) ) ;
INV     gate15516  (.A(g27498), .Z(g28175) ) ;
INV     gate15517  (.A(g27510), .Z(g28177) ) ;
INV     gate15518  (.A(g27518), .Z(g28178) ) ;
INV     gate15519  (.A(g27383), .Z(II36848) ) ;
INV     gate15520  (.A(II36848), .Z(g28179) ) ;
INV     gate15521  (.A(g27535), .Z(g28186) ) ;
INV     gate15522  (.A(g27543), .Z(g28187) ) ;
INV     gate15523  (.A(g27555), .Z(g28190) ) ;
INV     gate15524  (.A(g27386), .Z(II36860) ) ;
INV     gate15525  (.A(II36860), .Z(g28194) ) ;
INV     gate15526  (.A(g27384), .Z(II36864) ) ;
INV     gate15527  (.A(II36864), .Z(g28200) ) ;
INV     gate15528  (.A(g27786), .Z(II36867) ) ;
INV     gate15529  (.A(g27955), .Z(II36870) ) ;
INV     gate15530  (.A(g27971), .Z(II36873) ) ;
INV     gate15531  (.A(g27986), .Z(II36876) ) ;
INV     gate15532  (.A(g27972), .Z(II36879) ) ;
INV     gate15533  (.A(g27987), .Z(II36882) ) ;
INV     gate15534  (.A(g28003), .Z(II36885) ) ;
INV     gate15535  (.A(g27988), .Z(II36888) ) ;
INV     gate15536  (.A(g28004), .Z(II36891) ) ;
INV     gate15537  (.A(g28022), .Z(II36894) ) ;
INV     gate15538  (.A(g28005), .Z(II36897) ) ;
INV     gate15539  (.A(g28023), .Z(II36900) ) ;
INV     gate15540  (.A(g28045), .Z(II36903) ) ;
INV     gate15541  (.A(g27989), .Z(II36906) ) ;
INV     gate15542  (.A(g28006), .Z(II36909) ) ;
INV     gate15543  (.A(g28024), .Z(II36912) ) ;
INV     gate15544  (.A(g28007), .Z(II36915) ) ;
INV     gate15545  (.A(g28025), .Z(II36918) ) ;
INV     gate15546  (.A(g28047), .Z(II36921) ) ;
INV     gate15547  (.A(g28026), .Z(II36924) ) ;
INV     gate15548  (.A(g28048), .Z(II36927) ) ;
INV     gate15549  (.A(g28071), .Z(II36930) ) ;
INV     gate15550  (.A(g28049), .Z(II36933) ) ;
INV     gate15551  (.A(g28072), .Z(II36936) ) ;
INV     gate15552  (.A(g28095), .Z(II36939) ) ;
INV     gate15553  (.A(g27905), .Z(II36942) ) ;
INV     gate15554  (.A(g27793), .Z(II36945) ) ;
INV     gate15555  (.A(g27976), .Z(II36948) ) ;
INV     gate15556  (.A(g27992), .Z(II36951) ) ;
INV     gate15557  (.A(g28010), .Z(II36954) ) ;
INV     gate15558  (.A(g27993), .Z(II36957) ) ;
INV     gate15559  (.A(g28011), .Z(II36960) ) ;
INV     gate15560  (.A(g28030), .Z(II36963) ) ;
INV     gate15561  (.A(g28012), .Z(II36966) ) ;
INV     gate15562  (.A(g28031), .Z(II36969) ) ;
INV     gate15563  (.A(g28052), .Z(II36972) ) ;
INV     gate15564  (.A(g28032), .Z(II36975) ) ;
INV     gate15565  (.A(g28053), .Z(II36978) ) ;
INV     gate15566  (.A(g28074), .Z(II36981) ) ;
INV     gate15567  (.A(g28013), .Z(II36984) ) ;
INV     gate15568  (.A(g28033), .Z(II36987) ) ;
INV     gate15569  (.A(g28054), .Z(II36990) ) ;
INV     gate15570  (.A(g28034), .Z(II36993) ) ;
INV     gate15571  (.A(g28055), .Z(II36996) ) ;
INV     gate15572  (.A(g28076), .Z(II36999) ) ;
INV     gate15573  (.A(g28056), .Z(II37002) ) ;
INV     gate15574  (.A(g28077), .Z(II37005) ) ;
INV     gate15575  (.A(g28096), .Z(II37008) ) ;
INV     gate15576  (.A(g28078), .Z(II37011) ) ;
INV     gate15577  (.A(g28097), .Z(II37014) ) ;
INV     gate15578  (.A(g28113), .Z(II37017) ) ;
INV     gate15579  (.A(g27910), .Z(II37020) ) ;
INV     gate15580  (.A(g27799), .Z(II37023) ) ;
INV     gate15581  (.A(g27998), .Z(II37026) ) ;
INV     gate15582  (.A(g28016), .Z(II37029) ) ;
INV     gate15583  (.A(g28037), .Z(II37032) ) ;
INV     gate15584  (.A(g28017), .Z(II37035) ) ;
INV     gate15585  (.A(g28038), .Z(II37038) ) ;
INV     gate15586  (.A(g28060), .Z(II37041) ) ;
INV     gate15587  (.A(g28039), .Z(II37044) ) ;
INV     gate15588  (.A(g28061), .Z(II37047) ) ;
INV     gate15589  (.A(g28081), .Z(II37050) ) ;
INV     gate15590  (.A(g28062), .Z(II37053) ) ;
INV     gate15591  (.A(g28082), .Z(II37056) ) ;
INV     gate15592  (.A(g28099), .Z(II37059) ) ;
INV     gate15593  (.A(g28040), .Z(II37062) ) ;
INV     gate15594  (.A(g28063), .Z(II37065) ) ;
INV     gate15595  (.A(g28083), .Z(II37068) ) ;
INV     gate15596  (.A(g28064), .Z(II37071) ) ;
INV     gate15597  (.A(g28084), .Z(II37074) ) ;
INV     gate15598  (.A(g28101), .Z(II37077) ) ;
INV     gate15599  (.A(g28085), .Z(II37080) ) ;
INV     gate15600  (.A(g28102), .Z(II37083) ) ;
INV     gate15601  (.A(g28114), .Z(II37086) ) ;
INV     gate15602  (.A(g28103), .Z(II37089) ) ;
INV     gate15603  (.A(g28115), .Z(II37092) ) ;
INV     gate15604  (.A(g28124), .Z(II37095) ) ;
INV     gate15605  (.A(g27918), .Z(II37098) ) ;
INV     gate15606  (.A(g27805), .Z(II37101) ) ;
INV     gate15607  (.A(g28021), .Z(II37104) ) ;
INV     gate15608  (.A(g28043), .Z(II37107) ) ;
INV     gate15609  (.A(g28067), .Z(II37110) ) ;
INV     gate15610  (.A(g28044), .Z(II37113) ) ;
INV     gate15611  (.A(g28068), .Z(II37116) ) ;
INV     gate15612  (.A(g28089), .Z(II37119) ) ;
INV     gate15613  (.A(g28069), .Z(II37122) ) ;
INV     gate15614  (.A(g28090), .Z(II37125) ) ;
INV     gate15615  (.A(g28106), .Z(II37128) ) ;
INV     gate15616  (.A(g28091), .Z(II37131) ) ;
INV     gate15617  (.A(g28107), .Z(II37134) ) ;
INV     gate15618  (.A(g28117), .Z(II37137) ) ;
INV     gate15619  (.A(g28070), .Z(II37140) ) ;
INV     gate15620  (.A(g28092), .Z(II37143) ) ;
INV     gate15621  (.A(g28108), .Z(II37146) ) ;
INV     gate15622  (.A(g28093), .Z(II37149) ) ;
INV     gate15623  (.A(g28109), .Z(II37152) ) ;
INV     gate15624  (.A(g28119), .Z(II37155) ) ;
INV     gate15625  (.A(g28110), .Z(II37158) ) ;
INV     gate15626  (.A(g28120), .Z(II37161) ) ;
INV     gate15627  (.A(g28125), .Z(II37164) ) ;
INV     gate15628  (.A(g28121), .Z(II37167) ) ;
INV     gate15629  (.A(g28126), .Z(II37170) ) ;
INV     gate15630  (.A(g28132), .Z(II37173) ) ;
INV     gate15631  (.A(g27927), .Z(II37176) ) ;
INV     gate15632  (.A(g27784), .Z(II37179) ) ;
INV     gate15633  (.A(g27791), .Z(II37182) ) ;
INV     gate15634  (.A(g27797), .Z(II37185) ) ;
INV     gate15635  (.A(g27785), .Z(II37188) ) ;
INV     gate15636  (.A(g27792), .Z(II37191) ) ;
INV     gate15637  (.A(g27800), .Z(II37194) ) ;
INV     gate15638  (.A(g27903), .Z(II37197) ) ;
INV     gate15639  (.A(g27907), .Z(II37200) ) ;
INV     gate15640  (.A(g27912), .Z(II37203) ) ;
INV     gate15641  (.A(g28194), .Z(II37228) ) ;
INV     gate15642  (.A(II37228), .Z(g28341) ) ;
INV     gate15643  (.A(g28200), .Z(II37232) ) ;
INV     gate15644  (.A(II37232), .Z(g28343) ) ;
INV     gate15645  (.A(g28179), .Z(II37238) ) ;
INV     gate15646  (.A(II37238), .Z(g28347) ) ;
INV     gate15647  (.A(g28200), .Z(II37252) ) ;
INV     gate15648  (.A(II37252), .Z(g28359) ) ;
INV     gate15649  (.A(g28179), .Z(II37260) ) ;
INV     gate15650  (.A(II37260), .Z(g28365) ) ;
INV     gate15651  (.A(g28200), .Z(II37266) ) ;
INV     gate15652  (.A(II37266), .Z(g28369) ) ;
NOR2    gate15653  (.A(g27629), .B(g17001), .Z(g28145) ) ;
INV     gate15654  (.A(g28145), .Z(II37269) ) ;
INV     gate15655  (.A(II37269), .Z(g28370) ) ;
INV     gate15656  (.A(g28179), .Z(II37273) ) ;
INV     gate15657  (.A(II37273), .Z(g28372) ) ;
NOR2    gate15658  (.A(g27631), .B(g17031), .Z(g28146) ) ;
INV     gate15659  (.A(g28146), .Z(II37277) ) ;
INV     gate15660  (.A(II37277), .Z(g28374) ) ;
INV     gate15661  (.A(g28179), .Z(II37280) ) ;
INV     gate15662  (.A(II37280), .Z(g28375) ) ;
NOR2    gate15663  (.A(g27655), .B(g17065), .Z(g28147) ) ;
INV     gate15664  (.A(g28147), .Z(II37284) ) ;
INV     gate15665  (.A(II37284), .Z(g28377) ) ;
NOR2    gate15666  (.A(g27658), .B(g17100), .Z(g28148) ) ;
INV     gate15667  (.A(g28148), .Z(II37291) ) ;
INV     gate15668  (.A(II37291), .Z(g28382) ) ;
INV     gate15669  (.A(g28149), .Z(II37319) ) ;
INV     gate15670  (.A(II37319), .Z(g28390) ) ;
INV     gate15671  (.A(g28194), .Z(II37330) ) ;
INV     gate15672  (.A(II37330), .Z(g28393) ) ;
INV     gate15673  (.A(g28194), .Z(II37334) ) ;
INV     gate15674  (.A(II37334), .Z(g28395) ) ;
INV     gate15675  (.A(g28151), .Z(g28419) ) ;
NOR2    gate15676  (.A(g27250), .B(g10024), .Z(g28199) ) ;
INV     gate15677  (.A(g28199), .Z(II37379) ) ;
INV     gate15678  (.A(II37379), .Z(g28432) ) ;
INV     gate15679  (.A(g28194), .Z(II37386) ) ;
INV     gate15680  (.A(II37386), .Z(g28437) ) ;
NOR2    gate15681  (.A(g27251), .B(g10133), .Z(g27718) ) ;
INV     gate15682  (.A(g27718), .Z(II37394) ) ;
INV     gate15683  (.A(II37394), .Z(g28443) ) ;
INV     gate15684  (.A(g28200), .Z(II37400) ) ;
INV     gate15685  (.A(II37400), .Z(g28447) ) ;
NOR2    gate15686  (.A(g27252), .B(g10238), .Z(g27722) ) ;
INV     gate15687  (.A(g27722), .Z(II37410) ) ;
INV     gate15688  (.A(II37410), .Z(g28455) ) ;
INV     gate15689  (.A(g28179), .Z(II37415) ) ;
INV     gate15690  (.A(II37415), .Z(g28458) ) ;
NOR2    gate15691  (.A(g27254), .B(g10340), .Z(g27724) ) ;
INV     gate15692  (.A(g27724), .Z(II37426) ) ;
INV     gate15693  (.A(II37426), .Z(g28467) ) ;
INV     gate15694  (.A(g27776), .Z(g28483) ) ;
INV     gate15695  (.A(g27780), .Z(g28491) ) ;
INV     gate15696  (.A(g27787), .Z(g28496) ) ;
NOR2    gate15697  (.A(g27495), .B(g27052), .Z(g27759) ) ;
INV     gate15698  (.A(g27759), .Z(II37459) ) ;
INV     gate15699  (.A(II37459), .Z(g28498) ) ;
INV     gate15700  (.A(g27794), .Z(g28500) ) ;
NOR2    gate15701  (.A(g27509), .B(g27076), .Z(g27760) ) ;
INV     gate15702  (.A(g27760), .Z(II37467) ) ;
INV     gate15703  (.A(II37467), .Z(g28524) ) ;
NOR2    gate15704  (.A(g27516), .B(g27079), .Z(g27761) ) ;
INV     gate15705  (.A(g27761), .Z(II37471) ) ;
INV     gate15706  (.A(II37471), .Z(g28526) ) ;
NOR2    gate15707  (.A(g27530), .B(g27091), .Z(g27762) ) ;
INV     gate15708  (.A(g27762), .Z(II37474) ) ;
INV     gate15709  (.A(II37474), .Z(g28527) ) ;
NOR2    gate15710  (.A(g27534), .B(g27092), .Z(g27763) ) ;
INV     gate15711  (.A(g27763), .Z(II37481) ) ;
INV     gate15712  (.A(II37481), .Z(g28552) ) ;
NOR2    gate15713  (.A(g27541), .B(g27095), .Z(g27764) ) ;
INV     gate15714  (.A(g27764), .Z(II37484) ) ;
INV     gate15715  (.A(II37484), .Z(g28553) ) ;
INV     gate15716  (.A(g27806), .Z(g28554) ) ;
NOR2    gate15717  (.A(g27552), .B(g27103), .Z(g27765) ) ;
INV     gate15718  (.A(g27765), .Z(II37488) ) ;
INV     gate15719  (.A(II37488), .Z(g28555) ) ;
NOR2    gate15720  (.A(g27554), .B(g27104), .Z(g27766) ) ;
INV     gate15721  (.A(g27766), .Z(II37494) ) ;
INV     gate15722  (.A(II37494), .Z(g28579) ) ;
NOR2    gate15723  (.A(g27561), .B(g27107), .Z(g27767) ) ;
INV     gate15724  (.A(g27767), .Z(II37497) ) ;
INV     gate15725  (.A(II37497), .Z(g28580) ) ;
INV     gate15726  (.A(g27817), .Z(g28581) ) ;
INV     gate15727  (.A(g27820), .Z(g28582) ) ;
NOR2    gate15728  (.A(g27568), .B(g27110), .Z(g27768) ) ;
INV     gate15729  (.A(g27768), .Z(II37502) ) ;
INV     gate15730  (.A(II37502), .Z(g28583) ) ;
NOR2    gate15731  (.A(g27570), .B(g27111), .Z(g27769) ) ;
INV     gate15732  (.A(g27769), .Z(II37508) ) ;
INV     gate15733  (.A(II37508), .Z(g28607) ) ;
INV     gate15734  (.A(g27831), .Z(g28608) ) ;
INV     gate15735  (.A(g27839), .Z(g28609) ) ;
INV     gate15736  (.A(g27843), .Z(g28610) ) ;
NOR2    gate15737  (.A(g27578), .B(g27115), .Z(g27771) ) ;
INV     gate15738  (.A(g27771), .Z(II37514) ) ;
INV     gate15739  (.A(II37514), .Z(g28611) ) ;
NAND2   gate15740  (.A(II36592), .B(II36593), .Z(g28046) ) ;
INV     gate15741  (.A(g28046), .Z(g28612) ) ;
INV     gate15742  (.A(g27847), .Z(g28616) ) ;
INV     gate15743  (.A(g27858), .Z(g28617) ) ;
INV     gate15744  (.A(g27861), .Z(g28618) ) ;
NAND2   gate15745  (.A(II36667), .B(II36668), .Z(g28075) ) ;
INV     gate15746  (.A(g28075), .Z(g28619) ) ;
INV     gate15747  (.A(g27872), .Z(g28623) ) ;
INV     gate15748  (.A(g27879), .Z(g28624) ) ;
NAND2   gate15749  (.A(II36732), .B(II36733), .Z(g28100) ) ;
INV     gate15750  (.A(g28100), .Z(g28625) ) ;
INV     gate15751  (.A(g27889), .Z(g28629) ) ;
NAND2   gate15752  (.A(II36780), .B(II36781), .Z(g28118) ) ;
INV     gate15753  (.A(g28118), .Z(g28630) ) ;
INV     gate15754  (.A(g28200), .Z(g28638) ) ;
INV     gate15755  (.A(g27919), .Z(g28639) ) ;
INV     gate15756  (.A(g27928), .Z(g28640) ) ;
INV     gate15757  (.A(g27932), .Z(g28641) ) ;
INV     gate15758  (.A(g27939), .Z(g28642) ) ;
INV     gate15759  (.A(g27942), .Z(g28643) ) ;
INV     gate15760  (.A(g27946), .Z(g28644) ) ;
INV     gate15761  (.A(g27952), .Z(g28645) ) ;
INV     gate15762  (.A(g27956), .Z(g28646) ) ;
INV     gate15763  (.A(g27959), .Z(g28647) ) ;
INV     gate15764  (.A(g27965), .Z(g28648) ) ;
INV     gate15765  (.A(g27973), .Z(g28649) ) ;
INV     gate15766  (.A(g27977), .Z(g28650) ) ;
INV     gate15767  (.A(g27981), .Z(g28651) ) ;
INV     gate15768  (.A(g27994), .Z(g28652) ) ;
INV     gate15769  (.A(g27999), .Z(g28653) ) ;
INV     gate15770  (.A(g28018), .Z(g28655) ) ;
INV     gate15771  (.A(g28370), .Z(II37566) ) ;
INV     gate15772  (.A(g28498), .Z(II37569) ) ;
INV     gate15773  (.A(g28524), .Z(II37572) ) ;
INV     gate15774  (.A(g28527), .Z(II37575) ) ;
INV     gate15775  (.A(g28432), .Z(II37578) ) ;
INV     gate15776  (.A(g28374), .Z(II37581) ) ;
INV     gate15777  (.A(g28526), .Z(II37584) ) ;
INV     gate15778  (.A(g28552), .Z(II37587) ) ;
INV     gate15779  (.A(g28555), .Z(II37590) ) ;
INV     gate15780  (.A(g28443), .Z(II37593) ) ;
INV     gate15781  (.A(g28377), .Z(II37596) ) ;
INV     gate15782  (.A(g28553), .Z(II37599) ) ;
INV     gate15783  (.A(g28579), .Z(II37602) ) ;
INV     gate15784  (.A(g28583), .Z(II37605) ) ;
INV     gate15785  (.A(g28455), .Z(II37608) ) ;
INV     gate15786  (.A(g28382), .Z(II37611) ) ;
INV     gate15787  (.A(g28580), .Z(II37614) ) ;
INV     gate15788  (.A(g28607), .Z(II37617) ) ;
INV     gate15789  (.A(g28611), .Z(II37620) ) ;
INV     gate15790  (.A(g28467), .Z(II37623) ) ;
INV     gate15791  (.A(g28393), .Z(II37626) ) ;
INV     gate15792  (.A(g28369), .Z(II37629) ) ;
INV     gate15793  (.A(g28372), .Z(II37632) ) ;
INV     gate15794  (.A(g28390), .Z(II37635) ) ;
INV     gate15795  (.A(g28395), .Z(II37638) ) ;
INV     gate15796  (.A(g28375), .Z(II37641) ) ;
INV     gate15797  (.A(g28341), .Z(II37644) ) ;
INV     gate15798  (.A(g28343), .Z(II37647) ) ;
INV     gate15799  (.A(g28347), .Z(II37650) ) ;
INV     gate15800  (.A(g28359), .Z(II37653) ) ;
INV     gate15801  (.A(g28365), .Z(II37656) ) ;
INV     gate15802  (.A(g28437), .Z(II37659) ) ;
INV     gate15803  (.A(g28447), .Z(II37662) ) ;
INV     gate15804  (.A(g28458), .Z(II37665) ) ;
NOR2    gate15805  (.A(g27244), .B(g27723), .Z(g28495) ) ;
INV     gate15806  (.A(g28495), .Z(g28720) ) ;
NOR2    gate15807  (.A(g27240), .B(g27721), .Z(g28490) ) ;
INV     gate15808  (.A(g28490), .Z(g28721) ) ;
NOR2    gate15809  (.A(g26030), .B(g27728), .Z(g28528) ) ;
INV     gate15810  (.A(g28528), .Z(g28723) ) ;
NOR2    gate15811  (.A(g26027), .B(g27725), .Z(g28499) ) ;
INV     gate15812  (.A(g28499), .Z(g28725) ) ;
NOR2    gate15813  (.A(g26756), .B(g27720), .Z(g28489) ) ;
INV     gate15814  (.A(g28489), .Z(g28727) ) ;
NOR2    gate15815  (.A(g27671), .B(g28193), .Z(g28470) ) ;
INV     gate15816  (.A(g28470), .Z(g28730) ) ;
NOR2    gate15817  (.A(g27245), .B(g27726), .Z(g28525) ) ;
INV     gate15818  (.A(g28525), .Z(g28734) ) ;
NOR2    gate15819  (.A(g26755), .B(g27719), .Z(g28488) ) ;
INV     gate15820  (.A(g28488), .Z(g28740) ) ;
OR2     gate15821  (.A(g26481), .B(g27738), .Z(g28512) ) ;
INV     gate15822  (.A(g28512), .Z(II37702) ) ;
INV     gate15823  (.A(II37702), .Z(g28741) ) ;
INV     gate15824  (.A(g28512), .Z(II37712) ) ;
INV     gate15825  (.A(II37712), .Z(g28751) ) ;
OR2     gate15826  (.A(g26497), .B(g27743), .Z(g28540) ) ;
INV     gate15827  (.A(g28540), .Z(II37716) ) ;
INV     gate15828  (.A(II37716), .Z(g28755) ) ;
INV     gate15829  (.A(g28540), .Z(II37725) ) ;
INV     gate15830  (.A(II37725), .Z(g28764) ) ;
OR2     gate15831  (.A(g26512), .B(g27751), .Z(g28567) ) ;
INV     gate15832  (.A(g28567), .Z(II37729) ) ;
INV     gate15833  (.A(II37729), .Z(g28768) ) ;
INV     gate15834  (.A(g28567), .Z(II37736) ) ;
INV     gate15835  (.A(II37736), .Z(g28775) ) ;
OR2     gate15836  (.A(g26520), .B(g27756), .Z(g28595) ) ;
INV     gate15837  (.A(g28595), .Z(II37740) ) ;
INV     gate15838  (.A(II37740), .Z(g28779) ) ;
INV     gate15839  (.A(g28595), .Z(II37746) ) ;
INV     gate15840  (.A(II37746), .Z(g28785) ) ;
INV     gate15841  (.A(g28512), .Z(II37752) ) ;
INV     gate15842  (.A(II37752), .Z(g28791) ) ;
INV     gate15843  (.A(g28512), .Z(II37757) ) ;
INV     gate15844  (.A(II37757), .Z(g28796) ) ;
INV     gate15845  (.A(g28540), .Z(II37760) ) ;
INV     gate15846  (.A(II37760), .Z(g28799) ) ;
INV     gate15847  (.A(g28512), .Z(II37765) ) ;
INV     gate15848  (.A(II37765), .Z(g28804) ) ;
INV     gate15849  (.A(g28540), .Z(II37768) ) ;
INV     gate15850  (.A(II37768), .Z(g28807) ) ;
INV     gate15851  (.A(g28567), .Z(II37771) ) ;
INV     gate15852  (.A(II37771), .Z(g28810) ) ;
INV     gate15853  (.A(g28540), .Z(II37775) ) ;
INV     gate15854  (.A(II37775), .Z(g28814) ) ;
INV     gate15855  (.A(g28567), .Z(II37778) ) ;
INV     gate15856  (.A(II37778), .Z(g28817) ) ;
INV     gate15857  (.A(g28595), .Z(II37781) ) ;
INV     gate15858  (.A(II37781), .Z(g28820) ) ;
INV     gate15859  (.A(g28567), .Z(II37784) ) ;
INV     gate15860  (.A(II37784), .Z(g28823) ) ;
INV     gate15861  (.A(g28595), .Z(II37787) ) ;
INV     gate15862  (.A(II37787), .Z(g28826) ) ;
INV     gate15863  (.A(g28595), .Z(II37790) ) ;
INV     gate15864  (.A(II37790), .Z(g28829) ) ;
INV     gate15865  (.A(g28638), .Z(II37793) ) ;
INV     gate15866  (.A(II37793), .Z(g28832) ) ;
NOR2    gate15867  (.A(g28185), .B(g17001), .Z(g28634) ) ;
INV     gate15868  (.A(g28634), .Z(II37796) ) ;
INV     gate15869  (.A(II37796), .Z(g28833) ) ;
NOR2    gate15870  (.A(g28189), .B(g17031), .Z(g28635) ) ;
INV     gate15871  (.A(g28635), .Z(II37800) ) ;
INV     gate15872  (.A(II37800), .Z(g28835) ) ;
NOR2    gate15873  (.A(g28191), .B(g17065), .Z(g28636) ) ;
INV     gate15874  (.A(g28636), .Z(II37804) ) ;
INV     gate15875  (.A(II37804), .Z(g28837) ) ;
NOR2    gate15876  (.A(g28192), .B(g17100), .Z(g28637) ) ;
INV     gate15877  (.A(g28637), .Z(II37808) ) ;
INV     gate15878  (.A(II37808), .Z(g28839) ) ;
NOR2    gate15879  (.A(g24676), .B(g27801), .Z(g28409) ) ;
INV     gate15880  (.A(g28409), .Z(g28855) ) ;
NOR2    gate15881  (.A(g24695), .B(g27809), .Z(g28413) ) ;
INV     gate15882  (.A(g28413), .Z(g28859) ) ;
NOR2    gate15883  (.A(g24712), .B(g27830), .Z(g28417) ) ;
INV     gate15884  (.A(g28417), .Z(g28863) ) ;
NOR2    gate15885  (.A(g24723), .B(g27846), .Z(g28418) ) ;
INV     gate15886  (.A(g28418), .Z(g28867) ) ;
OR2     gate15887  (.A(g27738), .B(g25764), .Z(g28501) ) ;
INV     gate15888  (.A(g28501), .Z(II37842) ) ;
INV     gate15889  (.A(II37842), .Z(g28871) ) ;
INV     gate15890  (.A(g28501), .Z(II37846) ) ;
INV     gate15891  (.A(II37846), .Z(g28877) ) ;
NOR2    gate15892  (.A(g27736), .B(g10024), .Z(g28668) ) ;
INV     gate15893  (.A(g28668), .Z(II37851) ) ;
INV     gate15894  (.A(II37851), .Z(g28882) ) ;
OR2     gate15895  (.A(g27743), .B(g25818), .Z(g28529) ) ;
INV     gate15896  (.A(g28529), .Z(II37854) ) ;
INV     gate15897  (.A(II37854), .Z(g28883) ) ;
INV     gate15898  (.A(g28501), .Z(II37858) ) ;
INV     gate15899  (.A(II37858), .Z(g28889) ) ;
INV     gate15900  (.A(g28529), .Z(II37863) ) ;
INV     gate15901  (.A(II37863), .Z(g28894) ) ;
NOR2    gate15902  (.A(g27742), .B(g10133), .Z(g28321) ) ;
INV     gate15903  (.A(g28321), .Z(II37868) ) ;
INV     gate15904  (.A(II37868), .Z(g28899) ) ;
OR2     gate15905  (.A(g27751), .B(g25853), .Z(g28556) ) ;
INV     gate15906  (.A(g28556), .Z(II37871) ) ;
INV     gate15907  (.A(II37871), .Z(g28900) ) ;
INV     gate15908  (.A(g28501), .Z(II37875) ) ;
INV     gate15909  (.A(II37875), .Z(g28906) ) ;
INV     gate15910  (.A(g28529), .Z(II37880) ) ;
INV     gate15911  (.A(II37880), .Z(g28911) ) ;
INV     gate15912  (.A(g28556), .Z(II37885) ) ;
INV     gate15913  (.A(II37885), .Z(g28916) ) ;
NOR2    gate15914  (.A(g27747), .B(g10238), .Z(g28325) ) ;
INV     gate15915  (.A(g28325), .Z(II37891) ) ;
INV     gate15916  (.A(II37891), .Z(g28924) ) ;
OR2     gate15917  (.A(g27756), .B(g25874), .Z(g28584) ) ;
INV     gate15918  (.A(g28584), .Z(II37894) ) ;
INV     gate15919  (.A(II37894), .Z(g28925) ) ;
INV     gate15920  (.A(g28501), .Z(II37897) ) ;
INV     gate15921  (.A(II37897), .Z(g28928) ) ;
INV     gate15922  (.A(g28529), .Z(II37901) ) ;
INV     gate15923  (.A(II37901), .Z(g28932) ) ;
INV     gate15924  (.A(g28556), .Z(II37906) ) ;
INV     gate15925  (.A(II37906), .Z(g28937) ) ;
INV     gate15926  (.A(g28584), .Z(II37912) ) ;
INV     gate15927  (.A(II37912), .Z(g28945) ) ;
NOR2    gate15928  (.A(g27755), .B(g10340), .Z(g28328) ) ;
INV     gate15929  (.A(g28328), .Z(II37917) ) ;
INV     gate15930  (.A(II37917), .Z(g28950) ) ;
INV     gate15931  (.A(g28501), .Z(II37920) ) ;
INV     gate15932  (.A(II37920), .Z(g28951) ) ;
INV     gate15933  (.A(g28529), .Z(II37924) ) ;
INV     gate15934  (.A(II37924), .Z(g28955) ) ;
INV     gate15935  (.A(g28556), .Z(II37928) ) ;
INV     gate15936  (.A(II37928), .Z(g28959) ) ;
INV     gate15937  (.A(g28584), .Z(II37934) ) ;
INV     gate15938  (.A(II37934), .Z(g28967) ) ;
INV     gate15939  (.A(g28501), .Z(II37939) ) ;
INV     gate15940  (.A(II37939), .Z(g28972) ) ;
INV     gate15941  (.A(g28501), .Z(II37942) ) ;
INV     gate15942  (.A(II37942), .Z(g28975) ) ;
INV     gate15943  (.A(g28529), .Z(II37946) ) ;
INV     gate15944  (.A(II37946), .Z(g28979) ) ;
INV     gate15945  (.A(g28556), .Z(II37950) ) ;
INV     gate15946  (.A(II37950), .Z(g28983) ) ;
INV     gate15947  (.A(g28584), .Z(II37956) ) ;
INV     gate15948  (.A(II37956), .Z(g28993) ) ;
INV     gate15949  (.A(g28501), .Z(II37961) ) ;
INV     gate15950  (.A(II37961), .Z(g28998) ) ;
INV     gate15951  (.A(g28529), .Z(II37965) ) ;
INV     gate15952  (.A(II37965), .Z(g29002) ) ;
INV     gate15953  (.A(g28529), .Z(II37968) ) ;
INV     gate15954  (.A(II37968), .Z(g29005) ) ;
INV     gate15955  (.A(g28556), .Z(II37973) ) ;
INV     gate15956  (.A(II37973), .Z(g29010) ) ;
INV     gate15957  (.A(g28584), .Z(II37978) ) ;
INV     gate15958  (.A(II37978), .Z(g29019) ) ;
INV     gate15959  (.A(g28501), .Z(II37982) ) ;
INV     gate15960  (.A(II37982), .Z(g29023) ) ;
INV     gate15961  (.A(g28529), .Z(II37986) ) ;
INV     gate15962  (.A(II37986), .Z(g29027) ) ;
INV     gate15963  (.A(g28556), .Z(II37991) ) ;
INV     gate15964  (.A(II37991), .Z(g29032) ) ;
INV     gate15965  (.A(g28556), .Z(II37994) ) ;
INV     gate15966  (.A(II37994), .Z(g29035) ) ;
INV     gate15967  (.A(g28584), .Z(II37999) ) ;
INV     gate15968  (.A(II37999), .Z(g29042) ) ;
INV     gate15969  (.A(g28529), .Z(II38003) ) ;
INV     gate15970  (.A(II38003), .Z(g29046) ) ;
INV     gate15971  (.A(g28556), .Z(II38007) ) ;
INV     gate15972  (.A(II38007), .Z(g29050) ) ;
INV     gate15973  (.A(g28584), .Z(II38011) ) ;
INV     gate15974  (.A(II38011), .Z(g29054) ) ;
INV     gate15975  (.A(g28584), .Z(II38014) ) ;
INV     gate15976  (.A(II38014), .Z(g29057) ) ;
NOR2    gate15977  (.A(g15460), .B(g28008), .Z(g28342) ) ;
INV     gate15978  (.A(g28342), .Z(II38018) ) ;
INV     gate15979  (.A(II38018), .Z(g29061) ) ;
INV     gate15980  (.A(g28556), .Z(II38024) ) ;
INV     gate15981  (.A(II38024), .Z(g29065) ) ;
INV     gate15982  (.A(g28584), .Z(II38028) ) ;
INV     gate15983  (.A(II38028), .Z(g29069) ) ;
NOR2    gate15984  (.A(g15526), .B(g28027), .Z(g28344) ) ;
INV     gate15985  (.A(g28344), .Z(II38032) ) ;
INV     gate15986  (.A(II38032), .Z(g29073) ) ;
NOR2    gate15987  (.A(g15527), .B(g28028), .Z(g28345) ) ;
INV     gate15988  (.A(g28345), .Z(II38035) ) ;
INV     gate15989  (.A(II38035), .Z(g29074) ) ;
NOR2    gate15990  (.A(g15546), .B(g28035), .Z(g28346) ) ;
INV     gate15991  (.A(g28346), .Z(II38038) ) ;
INV     gate15992  (.A(II38038), .Z(g29075) ) ;
INV     gate15993  (.A(g28584), .Z(II38042) ) ;
INV     gate15994  (.A(II38042), .Z(g29077) ) ;
NOR2    gate15995  (.A(g15594), .B(g28050), .Z(g28348) ) ;
INV     gate15996  (.A(g28348), .Z(II38046) ) ;
INV     gate15997  (.A(II38046), .Z(g29081) ) ;
NOR2    gate15998  (.A(g15595), .B(g28051), .Z(g28349) ) ;
INV     gate15999  (.A(g28349), .Z(II38049) ) ;
INV     gate16000  (.A(II38049), .Z(g29082) ) ;
NOR2    gate16001  (.A(g15604), .B(g28057), .Z(g28350) ) ;
INV     gate16002  (.A(g28350), .Z(II38053) ) ;
INV     gate16003  (.A(II38053), .Z(g29084) ) ;
NOR2    gate16004  (.A(g15605), .B(g28058), .Z(g28351) ) ;
INV     gate16005  (.A(g28351), .Z(II38056) ) ;
INV     gate16006  (.A(II38056), .Z(g29085) ) ;
NOR2    gate16007  (.A(g15624), .B(g28065), .Z(g28352) ) ;
INV     gate16008  (.A(g28352), .Z(II38059) ) ;
INV     gate16009  (.A(II38059), .Z(g29086) ) ;
NOR2    gate16010  (.A(g15666), .B(g28073), .Z(g28353) ) ;
INV     gate16011  (.A(g28353), .Z(II38064) ) ;
INV     gate16012  (.A(II38064), .Z(g29089) ) ;
NOR2    gate16013  (.A(g15670), .B(g28079), .Z(g28354) ) ;
INV     gate16014  (.A(g28354), .Z(II38068) ) ;
INV     gate16015  (.A(II38068), .Z(g29091) ) ;
NOR2    gate16016  (.A(g15671), .B(g28080), .Z(g28355) ) ;
INV     gate16017  (.A(g28355), .Z(II38071) ) ;
INV     gate16018  (.A(II38071), .Z(g29092) ) ;
NOR2    gate16019  (.A(g15680), .B(g28086), .Z(g28356) ) ;
INV     gate16020  (.A(g28356), .Z(II38074) ) ;
INV     gate16021  (.A(II38074), .Z(g29093) ) ;
NOR2    gate16022  (.A(g15681), .B(g28087), .Z(g28357) ) ;
INV     gate16023  (.A(g28357), .Z(II38077) ) ;
INV     gate16024  (.A(II38077), .Z(g29094) ) ;
NOR2    gate16025  (.A(g15700), .B(g28094), .Z(g28358) ) ;
INV     gate16026  (.A(g28358), .Z(II38080) ) ;
INV     gate16027  (.A(II38080), .Z(g29095) ) ;
NOR2    gate16028  (.A(g15725), .B(g28098), .Z(g28360) ) ;
INV     gate16029  (.A(g28360), .Z(II38085) ) ;
INV     gate16030  (.A(II38085), .Z(g29098) ) ;
NOR2    gate16031  (.A(g15729), .B(g28104), .Z(g28361) ) ;
INV     gate16032  (.A(g28361), .Z(II38088) ) ;
INV     gate16033  (.A(II38088), .Z(g29099) ) ;
NOR2    gate16034  (.A(g15730), .B(g28105), .Z(g28362) ) ;
INV     gate16035  (.A(g28362), .Z(II38091) ) ;
INV     gate16036  (.A(II38091), .Z(g29100) ) ;
NOR2    gate16037  (.A(g15739), .B(g28111), .Z(g28363) ) ;
INV     gate16038  (.A(g28363), .Z(II38094) ) ;
INV     gate16039  (.A(II38094), .Z(g29101) ) ;
NOR2    gate16040  (.A(g15740), .B(g28112), .Z(g28364) ) ;
INV     gate16041  (.A(g28364), .Z(II38097) ) ;
INV     gate16042  (.A(II38097), .Z(g29102) ) ;
NOR2    gate16043  (.A(g15765), .B(g28116), .Z(g28366) ) ;
INV     gate16044  (.A(g28366), .Z(II38101) ) ;
INV     gate16045  (.A(II38101), .Z(g29104) ) ;
NOR2    gate16046  (.A(g15769), .B(g28122), .Z(g28367) ) ;
INV     gate16047  (.A(g28367), .Z(II38104) ) ;
INV     gate16048  (.A(II38104), .Z(g29105) ) ;
NOR2    gate16049  (.A(g15770), .B(g28123), .Z(g28368) ) ;
INV     gate16050  (.A(g28368), .Z(II38107) ) ;
INV     gate16051  (.A(II38107), .Z(g29106) ) ;
NOR2    gate16052  (.A(g15793), .B(g28127), .Z(g28371) ) ;
INV     gate16053  (.A(g28371), .Z(II38111) ) ;
INV     gate16054  (.A(II38111), .Z(g29108) ) ;
NOR2    gate16055  (.A(g16031), .B(g28171), .Z(g28420) ) ;
INV     gate16056  (.A(g28420), .Z(II38119) ) ;
INV     gate16057  (.A(II38119), .Z(g29117) ) ;
NOR2    gate16058  (.A(g16068), .B(g28176), .Z(g28421) ) ;
INV     gate16059  (.A(g28421), .Z(II38122) ) ;
INV     gate16060  (.A(II38122), .Z(g29118) ) ;
NOR2    gate16061  (.A(g16133), .B(g28188), .Z(g28425) ) ;
INV     gate16062  (.A(g28425), .Z(II38125) ) ;
INV     gate16063  (.A(II38125), .Z(g29119) ) ;
INV     gate16064  (.A(g28419), .Z(II38128) ) ;
INV     gate16065  (.A(II38128), .Z(g29120) ) ;
INV     gate16066  (.A(g28833), .Z(II38136) ) ;
INV     gate16067  (.A(g29061), .Z(II38139) ) ;
INV     gate16068  (.A(g29073), .Z(II38142) ) ;
INV     gate16069  (.A(g29081), .Z(II38145) ) ;
INV     gate16070  (.A(g29074), .Z(II38148) ) ;
INV     gate16071  (.A(g29082), .Z(II38151) ) ;
INV     gate16072  (.A(g29089), .Z(II38154) ) ;
INV     gate16073  (.A(g28882), .Z(II38157) ) ;
INV     gate16074  (.A(g28835), .Z(II38160) ) ;
INV     gate16075  (.A(g29075), .Z(II38163) ) ;
INV     gate16076  (.A(g29084), .Z(II38166) ) ;
INV     gate16077  (.A(g29091), .Z(II38169) ) ;
INV     gate16078  (.A(g29085), .Z(II38172) ) ;
INV     gate16079  (.A(g29092), .Z(II38175) ) ;
INV     gate16080  (.A(g29098), .Z(II38178) ) ;
INV     gate16081  (.A(g28899), .Z(II38181) ) ;
INV     gate16082  (.A(g28837), .Z(II38184) ) ;
INV     gate16083  (.A(g29086), .Z(II38187) ) ;
INV     gate16084  (.A(g29093), .Z(II38190) ) ;
INV     gate16085  (.A(g29099), .Z(II38193) ) ;
INV     gate16086  (.A(g29094), .Z(II38196) ) ;
INV     gate16087  (.A(g29100), .Z(II38199) ) ;
INV     gate16088  (.A(g29104), .Z(II38202) ) ;
INV     gate16089  (.A(g28924), .Z(II38205) ) ;
INV     gate16090  (.A(g28839), .Z(II38208) ) ;
INV     gate16091  (.A(g29095), .Z(II38211) ) ;
INV     gate16092  (.A(g29101), .Z(II38214) ) ;
INV     gate16093  (.A(g29105), .Z(II38217) ) ;
INV     gate16094  (.A(g29102), .Z(II38220) ) ;
INV     gate16095  (.A(g29106), .Z(II38223) ) ;
INV     gate16096  (.A(g29108), .Z(II38226) ) ;
INV     gate16097  (.A(g28950), .Z(II38229) ) ;
INV     gate16098  (.A(g29117), .Z(II38232) ) ;
INV     gate16099  (.A(g29118), .Z(II38235) ) ;
INV     gate16100  (.A(g29119), .Z(II38238) ) ;
INV     gate16101  (.A(g28832), .Z(II38241) ) ;
NOR2    gate16102  (.A(g28662), .B(g13322), .Z(g28920) ) ;
INV     gate16103  (.A(g28920), .Z(II38245) ) ;
INV     gate16104  (.A(II38245), .Z(g29168) ) ;
NOR2    gate16105  (.A(g28663), .B(g13343), .Z(g28941) ) ;
INV     gate16106  (.A(g28941), .Z(II38250) ) ;
INV     gate16107  (.A(II38250), .Z(g29171) ) ;
NOR2    gate16108  (.A(g28664), .B(g13365), .Z(g28963) ) ;
INV     gate16109  (.A(g28963), .Z(II38258) ) ;
INV     gate16110  (.A(II38258), .Z(g29177) ) ;
NOR2    gate16111  (.A(g28671), .B(g11607), .Z(g29013) ) ;
INV     gate16112  (.A(g29013), .Z(II38272) ) ;
INV     gate16113  (.A(II38272), .Z(g29189) ) ;
NOR2    gate16114  (.A(g28666), .B(g13390), .Z(g28987) ) ;
INV     gate16115  (.A(g28987), .Z(II38275) ) ;
INV     gate16116  (.A(II38275), .Z(g29190) ) ;
INV     gate16117  (.A(g28963), .Z(II38278) ) ;
INV     gate16118  (.A(II38278), .Z(g29191) ) ;
NOR3    gate16119  (.A(g26673), .B(g27241), .C(g28323), .Z(g28954) ) ;
INV     gate16120  (.A(g28954), .Z(g29192) ) ;
INV     gate16121  (.A(g28941), .Z(II38282) ) ;
INV     gate16122  (.A(II38282), .Z(g29193) ) ;
NOR2    gate16123  (.A(g28381), .B(g8907), .Z(g29113) ) ;
INV     gate16124  (.A(g29113), .Z(II38321) ) ;
INV     gate16125  (.A(II38321), .Z(g29230) ) ;
INV     gate16126  (.A(g29120), .Z(II38330) ) ;
INV     gate16127  (.A(II38330), .Z(g29237) ) ;
INV     gate16128  (.A(g29120), .Z(II38339) ) ;
INV     gate16129  (.A(II38339), .Z(g29244) ) ;
NOR2    gate16130  (.A(g28659), .B(g16277), .Z(g28886) ) ;
INV     gate16131  (.A(g28886), .Z(II38342) ) ;
INV     gate16132  (.A(II38342), .Z(g29245) ) ;
NOR2    gate16133  (.A(g28654), .B(g17001), .Z(g29109) ) ;
INV     gate16134  (.A(g29109), .Z(II38345) ) ;
INV     gate16135  (.A(II38345), .Z(g29246) ) ;
NOR2    gate16136  (.A(g28657), .B(g16221), .Z(g28874) ) ;
INV     gate16137  (.A(g28874), .Z(II38348) ) ;
INV     gate16138  (.A(II38348), .Z(g29247) ) ;
NOR2    gate16139  (.A(g28656), .B(g17031), .Z(g29110) ) ;
INV     gate16140  (.A(g29110), .Z(II38352) ) ;
INV     gate16141  (.A(II38352), .Z(g29249) ) ;
NOR2    gate16142  (.A(g28322), .B(g13500), .Z(g29039) ) ;
INV     gate16143  (.A(g29039), .Z(II38355) ) ;
INV     gate16144  (.A(II38355), .Z(g29250) ) ;
NOR2    gate16145  (.A(g28658), .B(g17065), .Z(g29111) ) ;
INV     gate16146  (.A(g29111), .Z(II38360) ) ;
INV     gate16147  (.A(II38360), .Z(g29253) ) ;
NOR2    gate16148  (.A(g28672), .B(g13487), .Z(g29016) ) ;
INV     gate16149  (.A(g29016), .Z(II38363) ) ;
INV     gate16150  (.A(II38363), .Z(g29254) ) ;
NOR2    gate16151  (.A(g28661), .B(g17100), .Z(g29112) ) ;
INV     gate16152  (.A(g29112), .Z(II38369) ) ;
INV     gate16153  (.A(II38369), .Z(g29258) ) ;
INV     gate16154  (.A(g28741), .Z(g29266) ) ;
INV     gate16155  (.A(g28734), .Z(II38386) ) ;
INV     gate16156  (.A(II38386), .Z(g29267) ) ;
INV     gate16157  (.A(g28751), .Z(g29268) ) ;
INV     gate16158  (.A(g28755), .Z(g29269) ) ;
INV     gate16159  (.A(g28730), .Z(II38391) ) ;
INV     gate16160  (.A(II38391), .Z(g29270) ) ;
INV     gate16161  (.A(g28764), .Z(g29271) ) ;
INV     gate16162  (.A(g28768), .Z(g29272) ) ;
INV     gate16163  (.A(g28727), .Z(II38396) ) ;
INV     gate16164  (.A(II38396), .Z(g29273) ) ;
INV     gate16165  (.A(g28775), .Z(g29274) ) ;
INV     gate16166  (.A(g28779), .Z(g29275) ) ;
INV     gate16167  (.A(g28725), .Z(II38401) ) ;
INV     gate16168  (.A(II38401), .Z(g29276) ) ;
INV     gate16169  (.A(g28785), .Z(g29277) ) ;
INV     gate16170  (.A(g28723), .Z(II38405) ) ;
INV     gate16171  (.A(II38405), .Z(g29278) ) ;
INV     gate16172  (.A(g28721), .Z(II38408) ) ;
INV     gate16173  (.A(II38408), .Z(g29279) ) ;
INV     gate16174  (.A(g28791), .Z(g29280) ) ;
INV     gate16175  (.A(g28720), .Z(II38412) ) ;
INV     gate16176  (.A(II38412), .Z(g29281) ) ;
INV     gate16177  (.A(g28796), .Z(g29282) ) ;
INV     gate16178  (.A(g28799), .Z(g29283) ) ;
INV     gate16179  (.A(g28804), .Z(g29285) ) ;
INV     gate16180  (.A(g28807), .Z(g29286) ) ;
INV     gate16181  (.A(g28810), .Z(g29287) ) ;
INV     gate16182  (.A(g28740), .Z(II38421) ) ;
INV     gate16183  (.A(II38421), .Z(g29288) ) ;
INV     gate16184  (.A(g28814), .Z(g29290) ) ;
INV     gate16185  (.A(g28817), .Z(g29291) ) ;
INV     gate16186  (.A(g28820), .Z(g29292) ) ;
NOR2    gate16187  (.A(g14894), .B(g28426), .Z(g28732) ) ;
INV     gate16188  (.A(g28732), .Z(II38428) ) ;
INV     gate16189  (.A(II38428), .Z(g29293) ) ;
INV     gate16190  (.A(g28823), .Z(g29295) ) ;
INV     gate16191  (.A(g28826), .Z(g29296) ) ;
NOR2    gate16192  (.A(g14957), .B(g28430), .Z(g28735) ) ;
INV     gate16193  (.A(g28735), .Z(II38434) ) ;
INV     gate16194  (.A(II38434), .Z(g29297) ) ;
NOR2    gate16195  (.A(g28427), .B(g27913), .Z(g28736) ) ;
INV     gate16196  (.A(g28736), .Z(II38437) ) ;
INV     gate16197  (.A(II38437), .Z(g29298) ) ;
NOR2    gate16198  (.A(g14975), .B(g28433), .Z(g28738) ) ;
INV     gate16199  (.A(g28738), .Z(II38440) ) ;
INV     gate16200  (.A(II38440), .Z(g29299) ) ;
INV     gate16201  (.A(g28829), .Z(g29301) ) ;
NOR2    gate16202  (.A(g15030), .B(g28439), .Z(g28744) ) ;
INV     gate16203  (.A(g28744), .Z(II38447) ) ;
INV     gate16204  (.A(II38447), .Z(g29304) ) ;
NOR2    gate16205  (.A(g28431), .B(g27922), .Z(g28745) ) ;
INV     gate16206  (.A(g28745), .Z(II38450) ) ;
INV     gate16207  (.A(II38450), .Z(g29305) ) ;
NOR2    gate16208  (.A(g15046), .B(g28441), .Z(g28746) ) ;
INV     gate16209  (.A(g28746), .Z(II38453) ) ;
INV     gate16210  (.A(II38453), .Z(g29306) ) ;
NOR2    gate16211  (.A(g28434), .B(g27923), .Z(g28747) ) ;
INV     gate16212  (.A(g28747), .Z(II38456) ) ;
INV     gate16213  (.A(II38456), .Z(g29307) ) ;
NOR2    gate16214  (.A(g15064), .B(g28444), .Z(g28749) ) ;
INV     gate16215  (.A(g28749), .Z(II38459) ) ;
INV     gate16216  (.A(II38459), .Z(g29308) ) ;
INV     gate16217  (.A(g29120), .Z(II38462) ) ;
INV     gate16218  (.A(II38462), .Z(g29309) ) ;
NOR2    gate16219  (.A(g28440), .B(g27931), .Z(g28754) ) ;
INV     gate16220  (.A(g28754), .Z(II38466) ) ;
INV     gate16221  (.A(II38466), .Z(g29311) ) ;
NOR2    gate16222  (.A(g15126), .B(g28451), .Z(g28758) ) ;
INV     gate16223  (.A(g28758), .Z(II38471) ) ;
INV     gate16224  (.A(II38471), .Z(g29314) ) ;
NOR2    gate16225  (.A(g28442), .B(g27935), .Z(g28759) ) ;
INV     gate16226  (.A(g28759), .Z(II38474) ) ;
INV     gate16227  (.A(II38474), .Z(g29315) ) ;
NOR2    gate16228  (.A(g15142), .B(g28453), .Z(g28760) ) ;
INV     gate16229  (.A(g28760), .Z(II38477) ) ;
INV     gate16230  (.A(II38477), .Z(g29316) ) ;
NOR2    gate16231  (.A(g28445), .B(g27936), .Z(g28761) ) ;
INV     gate16232  (.A(g28761), .Z(II38480) ) ;
INV     gate16233  (.A(II38480), .Z(g29317) ) ;
NOR2    gate16234  (.A(g28667), .B(g16457), .Z(g28990) ) ;
INV     gate16235  (.A(g28990), .Z(II38483) ) ;
INV     gate16236  (.A(II38483), .Z(g29318) ) ;
NOR2    gate16237  (.A(g15160), .B(g28456), .Z(g28763) ) ;
INV     gate16238  (.A(g28763), .Z(II38486) ) ;
INV     gate16239  (.A(II38486), .Z(g29319) ) ;
NOR2    gate16240  (.A(g28452), .B(g27945), .Z(g28767) ) ;
INV     gate16241  (.A(g28767), .Z(II38491) ) ;
INV     gate16242  (.A(II38491), .Z(g29322) ) ;
NOR2    gate16243  (.A(g15218), .B(g28463), .Z(g28771) ) ;
INV     gate16244  (.A(g28771), .Z(II38496) ) ;
INV     gate16245  (.A(II38496), .Z(g29325) ) ;
NOR2    gate16246  (.A(g28454), .B(g27949), .Z(g28772) ) ;
INV     gate16247  (.A(g28772), .Z(II38499) ) ;
INV     gate16248  (.A(II38499), .Z(g29326) ) ;
NOR2    gate16249  (.A(g15234), .B(g28465), .Z(g28773) ) ;
INV     gate16250  (.A(g28773), .Z(II38502) ) ;
INV     gate16251  (.A(II38502), .Z(g29327) ) ;
NOR2    gate16252  (.A(g28457), .B(g27951), .Z(g28774) ) ;
INV     gate16253  (.A(g28774), .Z(II38505) ) ;
INV     gate16254  (.A(II38505), .Z(g29328) ) ;
NOR2    gate16255  (.A(g28464), .B(g27963), .Z(g28778) ) ;
INV     gate16256  (.A(g28778), .Z(II38510) ) ;
INV     gate16257  (.A(II38510), .Z(g29331) ) ;
NOR2    gate16258  (.A(g15304), .B(g28475), .Z(g28782) ) ;
INV     gate16259  (.A(g28782), .Z(II38515) ) ;
INV     gate16260  (.A(II38515), .Z(g29334) ) ;
NOR2    gate16261  (.A(g28466), .B(g27968), .Z(g28783) ) ;
INV     gate16262  (.A(g28783), .Z(II38518) ) ;
INV     gate16263  (.A(II38518), .Z(g29335) ) ;
NOR2    gate16264  (.A(g28476), .B(g27984), .Z(g28788) ) ;
INV     gate16265  (.A(g28788), .Z(II38524) ) ;
INV     gate16266  (.A(II38524), .Z(g29339) ) ;
INV     gate16267  (.A(g28920), .Z(II38536) ) ;
INV     gate16268  (.A(II38536), .Z(g29349) ) ;
INV     gate16269  (.A(g29113), .Z(II38539) ) ;
INV     gate16270  (.A(II38539), .Z(g29350) ) ;
INV     gate16271  (.A(g29120), .Z(g29356) ) ;
INV     gate16272  (.A(g29120), .Z(g29358) ) ;
NOR2    gate16273  (.A(g28660), .B(g13295), .Z(g28903) ) ;
INV     gate16274  (.A(g28903), .Z(II38548) ) ;
INV     gate16275  (.A(II38548), .Z(g29359) ) ;
INV     gate16276  (.A(g28871), .Z(g29360) ) ;
INV     gate16277  (.A(g28877), .Z(g29361) ) ;
INV     gate16278  (.A(g28883), .Z(g29362) ) ;
INV     gate16279  (.A(g28889), .Z(g29363) ) ;
INV     gate16280  (.A(g28894), .Z(g29364) ) ;
INV     gate16281  (.A(g28900), .Z(g29365) ) ;
INV     gate16282  (.A(g28906), .Z(g29366) ) ;
INV     gate16283  (.A(g28911), .Z(g29367) ) ;
INV     gate16284  (.A(g28916), .Z(g29368) ) ;
INV     gate16285  (.A(g28925), .Z(g29369) ) ;
INV     gate16286  (.A(g28928), .Z(g29370) ) ;
INV     gate16287  (.A(g28932), .Z(g29371) ) ;
INV     gate16288  (.A(g28937), .Z(g29372) ) ;
INV     gate16289  (.A(g28945), .Z(g29373) ) ;
INV     gate16290  (.A(g28951), .Z(g29374) ) ;
INV     gate16291  (.A(g28955), .Z(g29375) ) ;
INV     gate16292  (.A(g28959), .Z(g29376) ) ;
INV     gate16293  (.A(g28967), .Z(g29377) ) ;
INV     gate16294  (.A(g28972), .Z(g29378) ) ;
INV     gate16295  (.A(g28975), .Z(g29379) ) ;
INV     gate16296  (.A(g28979), .Z(g29380) ) ;
INV     gate16297  (.A(g28983), .Z(g29381) ) ;
INV     gate16298  (.A(g28993), .Z(g29382) ) ;
INV     gate16299  (.A(g28998), .Z(g29383) ) ;
INV     gate16300  (.A(g29002), .Z(g29384) ) ;
INV     gate16301  (.A(g29005), .Z(g29385) ) ;
INV     gate16302  (.A(g29010), .Z(g29386) ) ;
INV     gate16303  (.A(g29019), .Z(g29387) ) ;
INV     gate16304  (.A(g29023), .Z(g29388) ) ;
INV     gate16305  (.A(g29027), .Z(g29389) ) ;
INV     gate16306  (.A(g29032), .Z(g29390) ) ;
INV     gate16307  (.A(g29035), .Z(g29391) ) ;
INV     gate16308  (.A(g29042), .Z(g29392) ) ;
INV     gate16309  (.A(g29046), .Z(g29393) ) ;
INV     gate16310  (.A(g29050), .Z(g29394) ) ;
INV     gate16311  (.A(g29054), .Z(g29395) ) ;
INV     gate16312  (.A(g29057), .Z(g29396) ) ;
INV     gate16313  (.A(g29065), .Z(g29397) ) ;
INV     gate16314  (.A(g29069), .Z(g29398) ) ;
INV     gate16315  (.A(g28987), .Z(II38591) ) ;
INV     gate16316  (.A(II38591), .Z(g29400) ) ;
INV     gate16317  (.A(g28990), .Z(II38594) ) ;
INV     gate16318  (.A(II38594), .Z(g29401) ) ;
INV     gate16319  (.A(g29077), .Z(g29402) ) ;
INV     gate16320  (.A(g29013), .Z(II38599) ) ;
INV     gate16321  (.A(II38599), .Z(g29404) ) ;
INV     gate16322  (.A(g29016), .Z(II38602) ) ;
INV     gate16323  (.A(II38602), .Z(g29405) ) ;
INV     gate16324  (.A(g29039), .Z(II38606) ) ;
INV     gate16325  (.A(II38606), .Z(g29407) ) ;
INV     gate16326  (.A(g28874), .Z(II38609) ) ;
INV     gate16327  (.A(II38609), .Z(g29408) ) ;
INV     gate16328  (.A(g28886), .Z(II38613) ) ;
INV     gate16329  (.A(II38613), .Z(g29410) ) ;
INV     gate16330  (.A(g28903), .Z(II38617) ) ;
INV     gate16331  (.A(II38617), .Z(g29412) ) ;
INV     gate16332  (.A(g29246), .Z(II38620) ) ;
INV     gate16333  (.A(g29293), .Z(II38623) ) ;
INV     gate16334  (.A(g29297), .Z(II38626) ) ;
INV     gate16335  (.A(g29304), .Z(II38629) ) ;
INV     gate16336  (.A(g29298), .Z(II38632) ) ;
INV     gate16337  (.A(g29305), .Z(II38635) ) ;
INV     gate16338  (.A(g29311), .Z(II38638) ) ;
INV     gate16339  (.A(g29249), .Z(II38641) ) ;
INV     gate16340  (.A(g29299), .Z(II38644) ) ;
INV     gate16341  (.A(g29306), .Z(II38647) ) ;
INV     gate16342  (.A(g29314), .Z(II38650) ) ;
INV     gate16343  (.A(g29307), .Z(II38653) ) ;
INV     gate16344  (.A(g29315), .Z(II38656) ) ;
INV     gate16345  (.A(g29322), .Z(II38659) ) ;
INV     gate16346  (.A(g29253), .Z(II38662) ) ;
INV     gate16347  (.A(g29412), .Z(II38665) ) ;
INV     gate16348  (.A(g29168), .Z(II38668) ) ;
INV     gate16349  (.A(g29171), .Z(II38671) ) ;
INV     gate16350  (.A(g29177), .Z(II38674) ) ;
INV     gate16351  (.A(g29400), .Z(II38677) ) ;
INV     gate16352  (.A(g29404), .Z(II38680) ) ;
INV     gate16353  (.A(g29308), .Z(II38683) ) ;
INV     gate16354  (.A(g29316), .Z(II38686) ) ;
INV     gate16355  (.A(g29325), .Z(II38689) ) ;
INV     gate16356  (.A(g29317), .Z(II38692) ) ;
INV     gate16357  (.A(g29326), .Z(II38695) ) ;
INV     gate16358  (.A(g29331), .Z(II38698) ) ;
INV     gate16359  (.A(g29401), .Z(II38701) ) ;
INV     gate16360  (.A(g29405), .Z(II38704) ) ;
INV     gate16361  (.A(g29407), .Z(II38707) ) ;
INV     gate16362  (.A(g29408), .Z(II38710) ) ;
INV     gate16363  (.A(g29410), .Z(II38713) ) ;
INV     gate16364  (.A(g29230), .Z(II38716) ) ;
INV     gate16365  (.A(g29258), .Z(II38719) ) ;
INV     gate16366  (.A(g29319), .Z(II38722) ) ;
INV     gate16367  (.A(g29327), .Z(II38725) ) ;
INV     gate16368  (.A(g29334), .Z(II38728) ) ;
INV     gate16369  (.A(g29328), .Z(II38731) ) ;
INV     gate16370  (.A(g29335), .Z(II38734) ) ;
INV     gate16371  (.A(g29339), .Z(II38737) ) ;
INV     gate16372  (.A(g29288), .Z(II38740) ) ;
INV     gate16373  (.A(g29267), .Z(II38743) ) ;
INV     gate16374  (.A(g29270), .Z(II38746) ) ;
INV     gate16375  (.A(g29273), .Z(II38749) ) ;
INV     gate16376  (.A(g29276), .Z(II38752) ) ;
INV     gate16377  (.A(g29278), .Z(II38755) ) ;
INV     gate16378  (.A(g29279), .Z(II38758) ) ;
INV     gate16379  (.A(g29281), .Z(II38761) ) ;
INV     gate16380  (.A(g29237), .Z(II38764) ) ;
INV     gate16381  (.A(g29244), .Z(II38767) ) ;
INV     gate16382  (.A(g29309), .Z(II38770) ) ;
INV     gate16383  (.A(g29350), .Z(g29491) ) ;
INV     gate16384  (.A(g29358), .Z(II38801) ) ;
INV     gate16385  (.A(II38801), .Z(g29495) ) ;
NOR2    gate16386  (.A(g29126), .B(g17001), .Z(g29353) ) ;
INV     gate16387  (.A(g29353), .Z(II38804) ) ;
INV     gate16388  (.A(II38804), .Z(g29496) ) ;
INV     gate16389  (.A(g29356), .Z(II38807) ) ;
INV     gate16390  (.A(II38807), .Z(g29497) ) ;
NOR2    gate16391  (.A(g29127), .B(g17031), .Z(g29354) ) ;
INV     gate16392  (.A(g29354), .Z(II38817) ) ;
INV     gate16393  (.A(II38817), .Z(g29499) ) ;
NOR2    gate16394  (.A(g29128), .B(g17065), .Z(g29355) ) ;
INV     gate16395  (.A(g29355), .Z(II38827) ) ;
INV     gate16396  (.A(II38827), .Z(g29501) ) ;
NOR2    gate16397  (.A(g29129), .B(g17100), .Z(g29357) ) ;
INV     gate16398  (.A(g29357), .Z(II38838) ) ;
INV     gate16399  (.A(II38838), .Z(g29504) ) ;
NOR2    gate16400  (.A(g28841), .B(g28396), .Z(g29167) ) ;
INV     gate16401  (.A(g29167), .Z(II38848) ) ;
INV     gate16402  (.A(II38848), .Z(g29506) ) ;
NOR2    gate16403  (.A(g28843), .B(g28398), .Z(g29169) ) ;
INV     gate16404  (.A(g29169), .Z(II38851) ) ;
INV     gate16405  (.A(II38851), .Z(g29507) ) ;
NOR2    gate16406  (.A(g28844), .B(g28399), .Z(g29170) ) ;
INV     gate16407  (.A(g29170), .Z(II38854) ) ;
INV     gate16408  (.A(II38854), .Z(g29508) ) ;
NOR2    gate16409  (.A(g28846), .B(g28401), .Z(g29172) ) ;
INV     gate16410  (.A(g29172), .Z(II38857) ) ;
INV     gate16411  (.A(II38857), .Z(g29509) ) ;
NOR2    gate16412  (.A(g28847), .B(g28402), .Z(g29173) ) ;
INV     gate16413  (.A(g29173), .Z(II38860) ) ;
INV     gate16414  (.A(II38860), .Z(g29510) ) ;
NOR2    gate16415  (.A(g28848), .B(g28404), .Z(g29178) ) ;
INV     gate16416  (.A(g29178), .Z(II38863) ) ;
INV     gate16417  (.A(II38863), .Z(g29511) ) ;
NOR2    gate16418  (.A(g28849), .B(g28405), .Z(g29179) ) ;
INV     gate16419  (.A(g29179), .Z(II38866) ) ;
INV     gate16420  (.A(II38866), .Z(g29512) ) ;
NOR2    gate16421  (.A(g28850), .B(g28407), .Z(g29181) ) ;
INV     gate16422  (.A(g29181), .Z(II38869) ) ;
INV     gate16423  (.A(II38869), .Z(g29513) ) ;
NOR2    gate16424  (.A(g28851), .B(g28408), .Z(g29182) ) ;
INV     gate16425  (.A(g29182), .Z(II38872) ) ;
INV     gate16426  (.A(II38872), .Z(g29514) ) ;
NOR2    gate16427  (.A(g28852), .B(g28411), .Z(g29184) ) ;
INV     gate16428  (.A(g29184), .Z(II38875) ) ;
INV     gate16429  (.A(II38875), .Z(g29515) ) ;
NOR2    gate16430  (.A(g28853), .B(g28412), .Z(g29185) ) ;
INV     gate16431  (.A(g29185), .Z(II38878) ) ;
INV     gate16432  (.A(II38878), .Z(g29516) ) ;
NOR2    gate16433  (.A(g28854), .B(g28416), .Z(g29187) ) ;
INV     gate16434  (.A(g29187), .Z(II38881) ) ;
INV     gate16435  (.A(II38881), .Z(g29517) ) ;
INV     gate16436  (.A(g29192), .Z(II38885) ) ;
INV     gate16437  (.A(II38885), .Z(g29519) ) ;
NOR2    gate16438  (.A(g14958), .B(g28881), .Z(g29194) ) ;
INV     gate16439  (.A(g29194), .Z(II38898) ) ;
INV     gate16440  (.A(II38898), .Z(g29530) ) ;
NOR2    gate16441  (.A(g15031), .B(g28893), .Z(g29197) ) ;
INV     gate16442  (.A(g29197), .Z(II38905) ) ;
INV     gate16443  (.A(II38905), .Z(g29535) ) ;
NOR2    gate16444  (.A(g15047), .B(g28898), .Z(g29198) ) ;
INV     gate16445  (.A(g29198), .Z(II38909) ) ;
INV     gate16446  (.A(II38909), .Z(g29537) ) ;
NOR2    gate16447  (.A(g15104), .B(g28910), .Z(g29201) ) ;
INV     gate16448  (.A(g29201), .Z(II38916) ) ;
INV     gate16449  (.A(II38916), .Z(g29542) ) ;
NOR2    gate16450  (.A(g15127), .B(g28915), .Z(g29204) ) ;
INV     gate16451  (.A(g29204), .Z(II38920) ) ;
INV     gate16452  (.A(II38920), .Z(g29544) ) ;
NOR2    gate16453  (.A(g15143), .B(g28923), .Z(g29205) ) ;
INV     gate16454  (.A(g29205), .Z(II38924) ) ;
INV     gate16455  (.A(II38924), .Z(g29546) ) ;
NOR2    gate16456  (.A(g15196), .B(g28936), .Z(g29209) ) ;
INV     gate16457  (.A(g29209), .Z(II38931) ) ;
INV     gate16458  (.A(II38931), .Z(g29551) ) ;
NOR2    gate16459  (.A(g15219), .B(g28944), .Z(g29212) ) ;
INV     gate16460  (.A(g29212), .Z(II38936) ) ;
INV     gate16461  (.A(II38936), .Z(g29554) ) ;
NOR2    gate16462  (.A(g15235), .B(g28949), .Z(g29213) ) ;
INV     gate16463  (.A(g29213), .Z(II38940) ) ;
INV     gate16464  (.A(II38940), .Z(g29556) ) ;
NOR2    gate16465  (.A(g15282), .B(g28966), .Z(g29218) ) ;
INV     gate16466  (.A(g29218), .Z(II38947) ) ;
INV     gate16467  (.A(II38947), .Z(g29561) ) ;
NOR2    gate16468  (.A(g15305), .B(g28971), .Z(g29221) ) ;
INV     gate16469  (.A(g29221), .Z(II38951) ) ;
INV     gate16470  (.A(II38951), .Z(g29563) ) ;
NOR2    gate16471  (.A(g15374), .B(g28997), .Z(g29226) ) ;
INV     gate16472  (.A(g29226), .Z(II38958) ) ;
INV     gate16473  (.A(II38958), .Z(g29568) ) ;
OR3     gate16474  (.A(g1942), .B(g1939), .C(g29113), .Z(g29348) ) ;
INV     gate16475  (.A(g29348), .Z(II38975) ) ;
INV     gate16476  (.A(II38975), .Z(g29583) ) ;
INV     gate16477  (.A(g29496), .Z(II38999) ) ;
INV     gate16478  (.A(g29506), .Z(II39002) ) ;
INV     gate16479  (.A(g29507), .Z(II39005) ) ;
INV     gate16480  (.A(g29509), .Z(II39008) ) ;
INV     gate16481  (.A(g29530), .Z(II39011) ) ;
INV     gate16482  (.A(g29535), .Z(II39014) ) ;
INV     gate16483  (.A(g29542), .Z(II39017) ) ;
INV     gate16484  (.A(g29499), .Z(II39020) ) ;
INV     gate16485  (.A(g29508), .Z(II39023) ) ;
INV     gate16486  (.A(g29510), .Z(II39026) ) ;
INV     gate16487  (.A(g29512), .Z(II39029) ) ;
INV     gate16488  (.A(g29537), .Z(II39032) ) ;
INV     gate16489  (.A(g29544), .Z(II39035) ) ;
INV     gate16490  (.A(g29551), .Z(II39038) ) ;
INV     gate16491  (.A(g29501), .Z(II39041) ) ;
INV     gate16492  (.A(g29511), .Z(II39044) ) ;
INV     gate16493  (.A(g29513), .Z(II39047) ) ;
INV     gate16494  (.A(g29515), .Z(II39050) ) ;
INV     gate16495  (.A(g29546), .Z(II39053) ) ;
INV     gate16496  (.A(g29554), .Z(II39056) ) ;
INV     gate16497  (.A(g29561), .Z(II39059) ) ;
INV     gate16498  (.A(g29504), .Z(II39062) ) ;
INV     gate16499  (.A(g29514), .Z(II39065) ) ;
INV     gate16500  (.A(g29516), .Z(II39068) ) ;
INV     gate16501  (.A(g29517), .Z(II39071) ) ;
INV     gate16502  (.A(g29556), .Z(II39074) ) ;
INV     gate16503  (.A(g29563), .Z(II39077) ) ;
INV     gate16504  (.A(g29568), .Z(II39080) ) ;
INV     gate16505  (.A(g29519), .Z(II39083) ) ;
INV     gate16506  (.A(g29497), .Z(II39086) ) ;
INV     gate16507  (.A(g29495), .Z(II39089) ) ;
NOR2    gate16508  (.A(g28712), .B(g29180), .Z(g29574) ) ;
INV     gate16509  (.A(g29574), .Z(g29658) ) ;
NOR2    gate16510  (.A(g28710), .B(g29176), .Z(g29571) ) ;
INV     gate16511  (.A(g29571), .Z(g29659) ) ;
NOR2    gate16512  (.A(g28715), .B(g29188), .Z(g29578) ) ;
INV     gate16513  (.A(g29578), .Z(g29660) ) ;
NOR2    gate16514  (.A(g28713), .B(g29183), .Z(g29576) ) ;
INV     gate16515  (.A(g29576), .Z(g29661) ) ;
NOR2    gate16516  (.A(g28709), .B(g29175), .Z(g29570) ) ;
INV     gate16517  (.A(g29570), .Z(g29662) ) ;
NOR2    gate16518  (.A(g29130), .B(g29411), .Z(g29552) ) ;
INV     gate16519  (.A(g29552), .Z(g29664) ) ;
NOR2    gate16520  (.A(g28714), .B(g29186), .Z(g29577) ) ;
INV     gate16521  (.A(g29577), .Z(g29666) ) ;
NOR2    gate16522  (.A(g28708), .B(g29174), .Z(g29569) ) ;
INV     gate16523  (.A(g29569), .Z(g29668) ) ;
INV     gate16524  (.A(g29583), .Z(g29673) ) ;
NOR2    gate16525  (.A(g29399), .B(g17001), .Z(g29579) ) ;
INV     gate16526  (.A(g29579), .Z(II39121) ) ;
INV     gate16527  (.A(II39121), .Z(g29689) ) ;
NOR2    gate16528  (.A(g13878), .B(g29248), .Z(g29606) ) ;
INV     gate16529  (.A(g29606), .Z(II39124) ) ;
INV     gate16530  (.A(II39124), .Z(g29690) ) ;
NOR2    gate16531  (.A(g13892), .B(g29251), .Z(g29608) ) ;
INV     gate16532  (.A(g29608), .Z(II39127) ) ;
INV     gate16533  (.A(II39127), .Z(g29691) ) ;
NOR2    gate16534  (.A(g29403), .B(g17031), .Z(g29580) ) ;
INV     gate16535  (.A(g29580), .Z(II39130) ) ;
INV     gate16536  (.A(II39130), .Z(g29692) ) ;
NOR2    gate16537  (.A(g13900), .B(g29252), .Z(g29609) ) ;
INV     gate16538  (.A(g29609), .Z(II39133) ) ;
INV     gate16539  (.A(II39133), .Z(g29693) ) ;
NOR2    gate16540  (.A(g13913), .B(g29255), .Z(g29611) ) ;
INV     gate16541  (.A(g29611), .Z(II39136) ) ;
INV     gate16542  (.A(II39136), .Z(g29694) ) ;
NOR2    gate16543  (.A(g13933), .B(g29256), .Z(g29612) ) ;
INV     gate16544  (.A(g29612), .Z(II39139) ) ;
INV     gate16545  (.A(II39139), .Z(g29695) ) ;
NOR2    gate16546  (.A(g29406), .B(g17065), .Z(g29581) ) ;
INV     gate16547  (.A(g29581), .Z(II39142) ) ;
INV     gate16548  (.A(II39142), .Z(g29696) ) ;
NOR2    gate16549  (.A(g13941), .B(g29257), .Z(g29613) ) ;
INV     gate16550  (.A(g29613), .Z(II39145) ) ;
INV     gate16551  (.A(II39145), .Z(g29697) ) ;
NOR2    gate16552  (.A(g13969), .B(g29259), .Z(g29616) ) ;
INV     gate16553  (.A(g29616), .Z(II39148) ) ;
INV     gate16554  (.A(II39148), .Z(g29698) ) ;
NOR2    gate16555  (.A(g13989), .B(g29260), .Z(g29617) ) ;
INV     gate16556  (.A(g29617), .Z(II39151) ) ;
INV     gate16557  (.A(II39151), .Z(g29699) ) ;
NOR2    gate16558  (.A(g29409), .B(g17100), .Z(g29582) ) ;
INV     gate16559  (.A(g29582), .Z(II39154) ) ;
INV     gate16560  (.A(II39154), .Z(g29700) ) ;
NOR2    gate16561  (.A(g13997), .B(g29261), .Z(g29618) ) ;
INV     gate16562  (.A(g29618), .Z(II39157) ) ;
INV     gate16563  (.A(II39157), .Z(g29701) ) ;
NOR2    gate16564  (.A(g14039), .B(g29262), .Z(g29620) ) ;
INV     gate16565  (.A(g29620), .Z(II39160) ) ;
INV     gate16566  (.A(II39160), .Z(g29702) ) ;
NOR2    gate16567  (.A(g14059), .B(g29263), .Z(g29621) ) ;
INV     gate16568  (.A(g29621), .Z(II39164) ) ;
INV     gate16569  (.A(II39164), .Z(g29704) ) ;
NOR2    gate16570  (.A(g14130), .B(g29264), .Z(g29623) ) ;
INV     gate16571  (.A(g29623), .Z(II39168) ) ;
INV     gate16572  (.A(II39168), .Z(g29708) ) ;
NAND2   gate16573  (.A(II38811), .B(II38812), .Z(g29498) ) ;
INV     gate16574  (.A(g29498), .Z(g29716) ) ;
NAND2   gate16575  (.A(II38821), .B(II38822), .Z(g29500) ) ;
INV     gate16576  (.A(g29500), .Z(g29724) ) ;
NAND2   gate16577  (.A(II38832), .B(II38833), .Z(g29503) ) ;
INV     gate16578  (.A(g29503), .Z(g29726) ) ;
NAND2   gate16579  (.A(II38842), .B(II38843), .Z(g29505) ) ;
INV     gate16580  (.A(g29505), .Z(g29739) ) ;
INV     gate16581  (.A(g29689), .Z(II39234) ) ;
INV     gate16582  (.A(g29690), .Z(II39237) ) ;
INV     gate16583  (.A(g29691), .Z(II39240) ) ;
INV     gate16584  (.A(g29694), .Z(II39243) ) ;
INV     gate16585  (.A(g29692), .Z(II39246) ) ;
INV     gate16586  (.A(g29693), .Z(II39249) ) ;
INV     gate16587  (.A(g29695), .Z(II39252) ) ;
INV     gate16588  (.A(g29698), .Z(II39255) ) ;
INV     gate16589  (.A(g29696), .Z(II39258) ) ;
INV     gate16590  (.A(g29697), .Z(II39261) ) ;
INV     gate16591  (.A(g29699), .Z(II39264) ) ;
INV     gate16592  (.A(g29702), .Z(II39267) ) ;
INV     gate16593  (.A(g29700), .Z(II39270) ) ;
INV     gate16594  (.A(g29701), .Z(II39273) ) ;
INV     gate16595  (.A(g29704), .Z(II39276) ) ;
INV     gate16596  (.A(g29708), .Z(II39279) ) ;
NOR2    gate16597  (.A(g29518), .B(g29284), .Z(g29663) ) ;
INV     gate16598  (.A(g29663), .Z(g29823) ) ;
NOR2    gate16599  (.A(g29521), .B(g29289), .Z(g29665) ) ;
INV     gate16600  (.A(g29665), .Z(g29829) ) ;
NOR2    gate16601  (.A(g29524), .B(g29294), .Z(g29667) ) ;
INV     gate16602  (.A(g29667), .Z(g29835) ) ;
NOR2    gate16603  (.A(g29528), .B(g29300), .Z(g29669) ) ;
INV     gate16604  (.A(g29669), .Z(g29840) ) ;
NOR2    gate16605  (.A(g29529), .B(g29302), .Z(g29670) ) ;
INV     gate16606  (.A(g29670), .Z(g29844) ) ;
NOR3    gate16607  (.A(g28707), .B(g28711), .C(g29466), .Z(g29761) ) ;
INV     gate16608  (.A(g29761), .Z(g29848) ) ;
NOR2    gate16609  (.A(g29534), .B(g29310), .Z(g29671) ) ;
INV     gate16610  (.A(g29671), .Z(g29849) ) ;
NOR2    gate16611  (.A(g29536), .B(g29312), .Z(g29672) ) ;
INV     gate16612  (.A(g29672), .Z(g29853) ) ;
NOR2    gate16613  (.A(g29540), .B(g29320), .Z(g29676) ) ;
INV     gate16614  (.A(g29676), .Z(g29857) ) ;
NOR2    gate16615  (.A(g29543), .B(g29321), .Z(g29677) ) ;
INV     gate16616  (.A(g29677), .Z(g29861) ) ;
NOR2    gate16617  (.A(g29545), .B(g29323), .Z(g29678) ) ;
INV     gate16618  (.A(g29678), .Z(g29865) ) ;
NOR2    gate16619  (.A(g29549), .B(g29329), .Z(g29679) ) ;
INV     gate16620  (.A(g29679), .Z(g29869) ) ;
NOR2    gate16621  (.A(g29553), .B(g29330), .Z(g29680) ) ;
INV     gate16622  (.A(g29680), .Z(g29873) ) ;
NOR2    gate16623  (.A(g29555), .B(g29332), .Z(g29681) ) ;
INV     gate16624  (.A(g29681), .Z(g29877) ) ;
NOR2    gate16625  (.A(g29557), .B(g29336), .Z(g29682) ) ;
INV     gate16626  (.A(g29682), .Z(g29881) ) ;
NOR2    gate16627  (.A(g29559), .B(g29337), .Z(g29683) ) ;
INV     gate16628  (.A(g29683), .Z(g29885) ) ;
NOR2    gate16629  (.A(g29562), .B(g29338), .Z(g29684) ) ;
INV     gate16630  (.A(g29684), .Z(g29889) ) ;
NOR2    gate16631  (.A(g29564), .B(g29341), .Z(g29685) ) ;
INV     gate16632  (.A(g29685), .Z(g29893) ) ;
NOR2    gate16633  (.A(g29566), .B(g29342), .Z(g29686) ) ;
INV     gate16634  (.A(g29686), .Z(g29897) ) ;
NOR2    gate16635  (.A(g29572), .B(g29344), .Z(g29687) ) ;
INV     gate16636  (.A(g29687), .Z(g29901) ) ;
NOR2    gate16637  (.A(g29575), .B(g29346), .Z(g29688) ) ;
INV     gate16638  (.A(g29688), .Z(g29905) ) ;
INV     gate16639  (.A(g29664), .Z(II39398) ) ;
INV     gate16640  (.A(II39398), .Z(g29932) ) ;
INV     gate16641  (.A(g29662), .Z(II39401) ) ;
INV     gate16642  (.A(II39401), .Z(g29933) ) ;
INV     gate16643  (.A(g29661), .Z(II39404) ) ;
INV     gate16644  (.A(II39404), .Z(g29934) ) ;
INV     gate16645  (.A(g29660), .Z(II39407) ) ;
INV     gate16646  (.A(II39407), .Z(g29935) ) ;
INV     gate16647  (.A(g29659), .Z(II39411) ) ;
INV     gate16648  (.A(II39411), .Z(g29937) ) ;
INV     gate16649  (.A(g29658), .Z(II39414) ) ;
INV     gate16650  (.A(II39414), .Z(g29938) ) ;
INV     gate16651  (.A(g29668), .Z(II39418) ) ;
INV     gate16652  (.A(II39418), .Z(g29940) ) ;
INV     gate16653  (.A(g29666), .Z(II39423) ) ;
INV     gate16654  (.A(II39423), .Z(g29943) ) ;
INV     gate16655  (.A(g29940), .Z(II39454) ) ;
INV     gate16656  (.A(g29943), .Z(II39457) ) ;
INV     gate16657  (.A(g29932), .Z(II39460) ) ;
INV     gate16658  (.A(g29933), .Z(II39463) ) ;
INV     gate16659  (.A(g29934), .Z(II39466) ) ;
INV     gate16660  (.A(g29935), .Z(II39469) ) ;
INV     gate16661  (.A(g29937), .Z(II39472) ) ;
INV     gate16662  (.A(g29938), .Z(II39475) ) ;
NOR2    gate16663  (.A(g24676), .B(g29716), .Z(g29912) ) ;
INV     gate16664  (.A(g29912), .Z(g30036) ) ;
NOR2    gate16665  (.A(g24695), .B(g29724), .Z(g29914) ) ;
INV     gate16666  (.A(g29914), .Z(g30040) ) ;
NOR2    gate16667  (.A(g24712), .B(g29726), .Z(g29916) ) ;
INV     gate16668  (.A(g29916), .Z(g30044) ) ;
NOR2    gate16669  (.A(g24723), .B(g29739), .Z(g29920) ) ;
INV     gate16670  (.A(g29920), .Z(g30048) ) ;
INV     gate16671  (.A(g29848), .Z(II39550) ) ;
INV     gate16672  (.A(II39550), .Z(g30052) ) ;
NOR2    gate16673  (.A(g16049), .B(g29790), .Z(g29936) ) ;
INV     gate16674  (.A(g29936), .Z(II39573) ) ;
INV     gate16675  (.A(II39573), .Z(g30076) ) ;
NOR2    gate16676  (.A(g16102), .B(g29792), .Z(g29939) ) ;
INV     gate16677  (.A(g29939), .Z(II39577) ) ;
INV     gate16678  (.A(II39577), .Z(g30078) ) ;
NOR2    gate16679  (.A(g16182), .B(g29793), .Z(g29941) ) ;
INV     gate16680  (.A(g29941), .Z(II39585) ) ;
INV     gate16681  (.A(II39585), .Z(g30084) ) ;
INV     gate16682  (.A(g30052), .Z(II39622) ) ;
INV     gate16683  (.A(g30076), .Z(II39625) ) ;
INV     gate16684  (.A(g30078), .Z(II39628) ) ;
INV     gate16685  (.A(g30084), .Z(II39631) ) ;
NOR2    gate16686  (.A(g29965), .B(g13326), .Z(g30055) ) ;
INV     gate16687  (.A(g30055), .Z(II39635) ) ;
INV     gate16688  (.A(II39635), .Z(g30124) ) ;
NOR2    gate16689  (.A(g29966), .B(g13345), .Z(g30056) ) ;
INV     gate16690  (.A(g30056), .Z(II39638) ) ;
INV     gate16691  (.A(II39638), .Z(g30125) ) ;
NOR2    gate16692  (.A(g29967), .B(g13368), .Z(g30057) ) ;
INV     gate16693  (.A(g30057), .Z(II39641) ) ;
INV     gate16694  (.A(II39641), .Z(g30126) ) ;
NOR2    gate16695  (.A(g29968), .B(g13395), .Z(g30058) ) ;
INV     gate16696  (.A(g30058), .Z(II39647) ) ;
INV     gate16697  (.A(II39647), .Z(g30130) ) ;
NOR2    gate16698  (.A(g29520), .B(g29942), .Z(g30010) ) ;
INV     gate16699  (.A(g30010), .Z(g30134) ) ;
NOR2    gate16700  (.A(g29522), .B(g29944), .Z(g30011) ) ;
INV     gate16701  (.A(g30011), .Z(g30139) ) ;
NOR2    gate16702  (.A(g29523), .B(g29945), .Z(g30012) ) ;
INV     gate16703  (.A(g30012), .Z(g30143) ) ;
NOR2    gate16704  (.A(g29525), .B(g29946), .Z(g30013) ) ;
INV     gate16705  (.A(g30013), .Z(g30147) ) ;
NOR2    gate16706  (.A(g29526), .B(g29947), .Z(g30014) ) ;
INV     gate16707  (.A(g30014), .Z(g30151) ) ;
NOR2    gate16708  (.A(g29527), .B(g29948), .Z(g30015) ) ;
INV     gate16709  (.A(g30015), .Z(g30155) ) ;
NOR2    gate16710  (.A(g29531), .B(g29949), .Z(g30016) ) ;
INV     gate16711  (.A(g30016), .Z(g30159) ) ;
NOR2    gate16712  (.A(g29532), .B(g29950), .Z(g30017) ) ;
INV     gate16713  (.A(g30017), .Z(g30163) ) ;
NOR2    gate16714  (.A(g29533), .B(g29951), .Z(g30018) ) ;
INV     gate16715  (.A(g30018), .Z(g30167) ) ;
NOR2    gate16716  (.A(g29538), .B(g29952), .Z(g30019) ) ;
INV     gate16717  (.A(g30019), .Z(g30171) ) ;
NOR2    gate16718  (.A(g29539), .B(g29953), .Z(g30020) ) ;
INV     gate16719  (.A(g30020), .Z(g30175) ) ;
NOR2    gate16720  (.A(g29541), .B(g29954), .Z(g30021) ) ;
INV     gate16721  (.A(g30021), .Z(g30179) ) ;
NOR2    gate16722  (.A(g29547), .B(g29955), .Z(g30022) ) ;
INV     gate16723  (.A(g30022), .Z(g30183) ) ;
NOR2    gate16724  (.A(g29548), .B(g29956), .Z(g30023) ) ;
INV     gate16725  (.A(g30023), .Z(g30187) ) ;
NOR2    gate16726  (.A(g29550), .B(g29957), .Z(g30024) ) ;
INV     gate16727  (.A(g30024), .Z(g30191) ) ;
NOR2    gate16728  (.A(g29558), .B(g29958), .Z(g30025) ) ;
INV     gate16729  (.A(g30025), .Z(g30195) ) ;
NOR2    gate16730  (.A(g29560), .B(g29959), .Z(g30026) ) ;
INV     gate16731  (.A(g30026), .Z(g30199) ) ;
NOR2    gate16732  (.A(g29565), .B(g29960), .Z(g30027) ) ;
INV     gate16733  (.A(g30027), .Z(g30203) ) ;
NOR2    gate16734  (.A(g29567), .B(g29961), .Z(g30028) ) ;
INV     gate16735  (.A(g30028), .Z(g30207) ) ;
NOR2    gate16736  (.A(g29573), .B(g29962), .Z(g30029) ) ;
INV     gate16737  (.A(g30029), .Z(g30211) ) ;
NOR2    gate16738  (.A(g29910), .B(g8947), .Z(g30072) ) ;
INV     gate16739  (.A(g30072), .Z(II39674) ) ;
INV     gate16740  (.A(II39674), .Z(g30215) ) ;
NOR2    gate16741  (.A(g24676), .B(g29923), .Z(g30030) ) ;
INV     gate16742  (.A(g30030), .Z(g30229) ) ;
NOR2    gate16743  (.A(g24695), .B(g29925), .Z(g30031) ) ;
INV     gate16744  (.A(g30031), .Z(g30233) ) ;
NOR2    gate16745  (.A(g24712), .B(g29927), .Z(g30032) ) ;
INV     gate16746  (.A(g30032), .Z(g30237) ) ;
NOR2    gate16747  (.A(g24723), .B(g29931), .Z(g30033) ) ;
INV     gate16748  (.A(g30033), .Z(g30241) ) ;
INV     gate16749  (.A(g30072), .Z(II39761) ) ;
INV     gate16750  (.A(II39761), .Z(g30306) ) ;
NOR2    gate16751  (.A(g29970), .B(g11612), .Z(g30060) ) ;
INV     gate16752  (.A(g30060), .Z(II39764) ) ;
INV     gate16753  (.A(II39764), .Z(g30307) ) ;
NOR2    gate16754  (.A(g29971), .B(g13493), .Z(g30061) ) ;
INV     gate16755  (.A(g30061), .Z(II39767) ) ;
INV     gate16756  (.A(II39767), .Z(g30308) ) ;
NOR2    gate16757  (.A(g29812), .B(g11637), .Z(g30063) ) ;
INV     gate16758  (.A(g30063), .Z(II39770) ) ;
INV     gate16759  (.A(II39770), .Z(g30309) ) ;
NOR2    gate16760  (.A(g29813), .B(g13506), .Z(g30064) ) ;
INV     gate16761  (.A(g30064), .Z(II39773) ) ;
INV     gate16762  (.A(II39773), .Z(g30310) ) ;
NOR2    gate16763  (.A(g29816), .B(g13517), .Z(g30066) ) ;
INV     gate16764  (.A(g30066), .Z(II39776) ) ;
INV     gate16765  (.A(II39776), .Z(g30311) ) ;
NOR2    gate16766  (.A(g29963), .B(g16286), .Z(g30053) ) ;
INV     gate16767  (.A(g30053), .Z(II39779) ) ;
INV     gate16768  (.A(II39779), .Z(g30312) ) ;
NOR2    gate16769  (.A(g29964), .B(g16336), .Z(g30054) ) ;
INV     gate16770  (.A(g30054), .Z(II39782) ) ;
INV     gate16771  (.A(II39782), .Z(g30313) ) ;
INV     gate16772  (.A(g30124), .Z(II39785) ) ;
INV     gate16773  (.A(g30125), .Z(II39788) ) ;
INV     gate16774  (.A(g30126), .Z(II39791) ) ;
INV     gate16775  (.A(g30130), .Z(II39794) ) ;
INV     gate16776  (.A(g30307), .Z(II39797) ) ;
INV     gate16777  (.A(g30309), .Z(II39800) ) ;
INV     gate16778  (.A(g30308), .Z(II39803) ) ;
INV     gate16779  (.A(g30310), .Z(II39806) ) ;
INV     gate16780  (.A(g30311), .Z(II39809) ) ;
INV     gate16781  (.A(g30312), .Z(II39812) ) ;
INV     gate16782  (.A(g30313), .Z(II39815) ) ;
INV     gate16783  (.A(g30215), .Z(II39818) ) ;
NOR2    gate16784  (.A(g16380), .B(g30101), .Z(g30267) ) ;
INV     gate16785  (.A(g30267), .Z(II39821) ) ;
INV     gate16786  (.A(II39821), .Z(g30326) ) ;
NOR2    gate16787  (.A(g16382), .B(g30102), .Z(g30268) ) ;
INV     gate16788  (.A(g30268), .Z(II39825) ) ;
INV     gate16789  (.A(II39825), .Z(g30328) ) ;
NOR2    gate16790  (.A(g16386), .B(g30103), .Z(g30269) ) ;
INV     gate16791  (.A(g30269), .Z(II39828) ) ;
INV     gate16792  (.A(II39828), .Z(g30329) ) ;
NOR2    gate16793  (.A(g16387), .B(g30104), .Z(g30270) ) ;
INV     gate16794  (.A(g30270), .Z(II39832) ) ;
INV     gate16795  (.A(II39832), .Z(g30331) ) ;
NOR2    gate16796  (.A(g16388), .B(g30105), .Z(g30271) ) ;
INV     gate16797  (.A(g30271), .Z(II39835) ) ;
INV     gate16798  (.A(II39835), .Z(g30332) ) ;
NOR2    gate16799  (.A(g16392), .B(g30106), .Z(g30272) ) ;
INV     gate16800  (.A(g30272), .Z(II39840) ) ;
INV     gate16801  (.A(II39840), .Z(g30335) ) ;
NOR2    gate16802  (.A(g16393), .B(g30107), .Z(g30273) ) ;
INV     gate16803  (.A(g30273), .Z(II39843) ) ;
INV     gate16804  (.A(II39843), .Z(g30336) ) ;
NOR2    gate16805  (.A(g16403), .B(g30108), .Z(g30274) ) ;
INV     gate16806  (.A(g30274), .Z(II39848) ) ;
INV     gate16807  (.A(II39848), .Z(g30339) ) ;
NOR2    gate16808  (.A(g16413), .B(g30109), .Z(g30275) ) ;
INV     gate16809  (.A(g30275), .Z(II39853) ) ;
INV     gate16810  (.A(II39853), .Z(g30342) ) ;
NOR2    gate16811  (.A(g16415), .B(g30110), .Z(g30276) ) ;
INV     gate16812  (.A(g30276), .Z(II39856) ) ;
INV     gate16813  (.A(II39856), .Z(g30343) ) ;
NOR2    gate16814  (.A(g16418), .B(g30111), .Z(g30277) ) ;
INV     gate16815  (.A(g30277), .Z(II39859) ) ;
INV     gate16816  (.A(II39859), .Z(g30344) ) ;
NOR2    gate16817  (.A(g16420), .B(g30112), .Z(g30278) ) ;
INV     gate16818  (.A(g30278), .Z(II39863) ) ;
INV     gate16819  (.A(II39863), .Z(g30346) ) ;
NOR2    gate16820  (.A(g16424), .B(g30113), .Z(g30279) ) ;
INV     gate16821  (.A(g30279), .Z(II39866) ) ;
INV     gate16822  (.A(II39866), .Z(g30347) ) ;
NOR2    gate16823  (.A(g16425), .B(g30114), .Z(g30280) ) ;
INV     gate16824  (.A(g30280), .Z(II39870) ) ;
INV     gate16825  (.A(II39870), .Z(g30349) ) ;
NOR2    gate16826  (.A(g16426), .B(g30115), .Z(g30281) ) ;
INV     gate16827  (.A(g30281), .Z(II39873) ) ;
INV     gate16828  (.A(II39873), .Z(g30350) ) ;
NOR2    gate16829  (.A(g16430), .B(g30117), .Z(g30282) ) ;
INV     gate16830  (.A(g30282), .Z(II39878) ) ;
INV     gate16831  (.A(II39878), .Z(g30353) ) ;
NOR2    gate16832  (.A(g16431), .B(g30118), .Z(g30283) ) ;
INV     gate16833  (.A(g30283), .Z(II39881) ) ;
INV     gate16834  (.A(II39881), .Z(g30354) ) ;
NOR2    gate16835  (.A(g16444), .B(g29980), .Z(g30284) ) ;
INV     gate16836  (.A(g30284), .Z(II39886) ) ;
INV     gate16837  (.A(II39886), .Z(g30357) ) ;
NOR2    gate16838  (.A(g16447), .B(g29981), .Z(g30285) ) ;
INV     gate16839  (.A(g30285), .Z(II39889) ) ;
INV     gate16840  (.A(II39889), .Z(g30358) ) ;
NOR2    gate16841  (.A(g16449), .B(g29982), .Z(g30286) ) ;
INV     gate16842  (.A(g30286), .Z(II39892) ) ;
INV     gate16843  (.A(II39892), .Z(g30359) ) ;
NOR2    gate16844  (.A(g16452), .B(g29983), .Z(g30287) ) ;
INV     gate16845  (.A(g30287), .Z(II39895) ) ;
INV     gate16846  (.A(II39895), .Z(g30360) ) ;
NOR2    gate16847  (.A(g16454), .B(g29984), .Z(g30288) ) ;
INV     gate16848  (.A(g30288), .Z(II39899) ) ;
INV     gate16849  (.A(II39899), .Z(g30362) ) ;
NOR2    gate16850  (.A(g16458), .B(g29985), .Z(g30289) ) ;
INV     gate16851  (.A(g30289), .Z(II39902) ) ;
INV     gate16852  (.A(II39902), .Z(g30363) ) ;
NOR2    gate16853  (.A(g16459), .B(g29986), .Z(g30290) ) ;
INV     gate16854  (.A(g30290), .Z(II39906) ) ;
INV     gate16855  (.A(II39906), .Z(g30365) ) ;
NOR2    gate16856  (.A(g16460), .B(g29987), .Z(g30291) ) ;
INV     gate16857  (.A(g30291), .Z(II39909) ) ;
INV     gate16858  (.A(II39909), .Z(g30366) ) ;
NOR2    gate16859  (.A(g13477), .B(g29988), .Z(g30292) ) ;
INV     gate16860  (.A(g30292), .Z(II39913) ) ;
INV     gate16861  (.A(II39913), .Z(g30368) ) ;
NOR2    gate16862  (.A(g13480), .B(g29989), .Z(g30293) ) ;
INV     gate16863  (.A(g30293), .Z(II39916) ) ;
INV     gate16864  (.A(II39916), .Z(g30369) ) ;
NOR2    gate16865  (.A(g13483), .B(g29990), .Z(g30294) ) ;
INV     gate16866  (.A(g30294), .Z(II39919) ) ;
INV     gate16867  (.A(II39919), .Z(g30370) ) ;
NOR2    gate16868  (.A(g13485), .B(g29991), .Z(g30295) ) ;
INV     gate16869  (.A(g30295), .Z(II39922) ) ;
INV     gate16870  (.A(II39922), .Z(g30371) ) ;
NOR2    gate16871  (.A(g13488), .B(g29993), .Z(g30296) ) ;
INV     gate16872  (.A(g30296), .Z(II39926) ) ;
INV     gate16873  (.A(II39926), .Z(g30373) ) ;
NOR2    gate16874  (.A(g13490), .B(g29994), .Z(g30297) ) ;
INV     gate16875  (.A(g30297), .Z(II39930) ) ;
INV     gate16876  (.A(II39930), .Z(g30375) ) ;
NOR2    gate16877  (.A(g13496), .B(g29995), .Z(g30298) ) ;
INV     gate16878  (.A(g30298), .Z(II39933) ) ;
INV     gate16879  (.A(II39933), .Z(g30376) ) ;
NOR2    gate16880  (.A(g13499), .B(g29996), .Z(g30299) ) ;
INV     gate16881  (.A(g30299), .Z(II39936) ) ;
INV     gate16882  (.A(II39936), .Z(g30377) ) ;
NOR2    gate16883  (.A(g13502), .B(g30001), .Z(g30300) ) ;
INV     gate16884  (.A(g30300), .Z(II39939) ) ;
INV     gate16885  (.A(II39939), .Z(g30378) ) ;
NOR2    gate16886  (.A(g13504), .B(g30002), .Z(g30301) ) ;
INV     gate16887  (.A(g30301), .Z(II39942) ) ;
INV     gate16888  (.A(II39942), .Z(g30379) ) ;
NOR2    gate16889  (.A(g13513), .B(g30003), .Z(g30302) ) ;
INV     gate16890  (.A(g30302), .Z(II39945) ) ;
INV     gate16891  (.A(II39945), .Z(g30380) ) ;
NOR2    gate16892  (.A(g13516), .B(g30005), .Z(g30303) ) ;
INV     gate16893  (.A(g30303), .Z(II39948) ) ;
INV     gate16894  (.A(II39948), .Z(g30381) ) ;
NOR2    gate16895  (.A(g13527), .B(g30007), .Z(g30304) ) ;
INV     gate16896  (.A(g30304), .Z(II39951) ) ;
INV     gate16897  (.A(II39951), .Z(g30382) ) ;
INV     gate16898  (.A(g30306), .Z(g30383) ) ;
NOR2    gate16899  (.A(g16074), .B(g30077), .Z(g30245) ) ;
INV     gate16900  (.A(g30245), .Z(II39976) ) ;
INV     gate16901  (.A(II39976), .Z(g30408) ) ;
OR3     gate16902  (.A(g2636), .B(g2633), .C(g30072), .Z(g30305) ) ;
INV     gate16903  (.A(g30305), .Z(II39982) ) ;
INV     gate16904  (.A(II39982), .Z(g30412) ) ;
NOR2    gate16905  (.A(g16107), .B(g30079), .Z(g30246) ) ;
INV     gate16906  (.A(g30246), .Z(II39985) ) ;
INV     gate16907  (.A(II39985), .Z(g30435) ) ;
NOR2    gate16908  (.A(g16112), .B(g30080), .Z(g30247) ) ;
INV     gate16909  (.A(g30247), .Z(II39991) ) ;
INV     gate16910  (.A(II39991), .Z(g30439) ) ;
NOR2    gate16911  (.A(g16139), .B(g30081), .Z(g30248) ) ;
INV     gate16912  (.A(g30248), .Z(II39997) ) ;
INV     gate16913  (.A(II39997), .Z(g30443) ) ;
NOR2    gate16914  (.A(g16158), .B(g30082), .Z(g30249) ) ;
INV     gate16915  (.A(g30249), .Z(II40002) ) ;
INV     gate16916  (.A(II40002), .Z(g30446) ) ;
NOR2    gate16917  (.A(g16163), .B(g30083), .Z(g30250) ) ;
INV     gate16918  (.A(g30250), .Z(II40008) ) ;
INV     gate16919  (.A(II40008), .Z(g30450) ) ;
NOR2    gate16920  (.A(g16198), .B(g30085), .Z(g30251) ) ;
INV     gate16921  (.A(g30251), .Z(II40016) ) ;
INV     gate16922  (.A(II40016), .Z(g30456) ) ;
NOR2    gate16923  (.A(g16217), .B(g30086), .Z(g30252) ) ;
INV     gate16924  (.A(g30252), .Z(II40021) ) ;
INV     gate16925  (.A(II40021), .Z(g30459) ) ;
NOR2    gate16926  (.A(g16222), .B(g30087), .Z(g30253) ) ;
INV     gate16927  (.A(g30253), .Z(II40027) ) ;
INV     gate16928  (.A(II40027), .Z(g30463) ) ;
NOR2    gate16929  (.A(g16242), .B(g30088), .Z(g30254) ) ;
INV     gate16930  (.A(g30254), .Z(II40032) ) ;
INV     gate16931  (.A(II40032), .Z(g30466) ) ;
NOR2    gate16932  (.A(g16263), .B(g30089), .Z(g30255) ) ;
INV     gate16933  (.A(g30255), .Z(II40039) ) ;
INV     gate16934  (.A(II40039), .Z(g30471) ) ;
NOR2    gate16935  (.A(g16282), .B(g30090), .Z(g30256) ) ;
INV     gate16936  (.A(g30256), .Z(II40044) ) ;
INV     gate16937  (.A(II40044), .Z(g30474) ) ;
NOR2    gate16938  (.A(g16290), .B(g30091), .Z(g30257) ) ;
INV     gate16939  (.A(g30257), .Z(II40051) ) ;
INV     gate16940  (.A(II40051), .Z(g30479) ) ;
NOR2    gate16941  (.A(g16291), .B(g30092), .Z(g30258) ) ;
INV     gate16942  (.A(g30258), .Z(II40054) ) ;
INV     gate16943  (.A(II40054), .Z(g30480) ) ;
NOR2    gate16944  (.A(g16301), .B(g30093), .Z(g30259) ) ;
INV     gate16945  (.A(g30259), .Z(II40059) ) ;
INV     gate16946  (.A(II40059), .Z(g30483) ) ;
NOR2    gate16947  (.A(g16322), .B(g30094), .Z(g30260) ) ;
INV     gate16948  (.A(g30260), .Z(II40066) ) ;
INV     gate16949  (.A(II40066), .Z(g30488) ) ;
NOR2    gate16950  (.A(g16342), .B(g30095), .Z(g30261) ) ;
INV     gate16951  (.A(g30261), .Z(II40071) ) ;
INV     gate16952  (.A(II40071), .Z(g30491) ) ;
NOR2    gate16953  (.A(g16343), .B(g30096), .Z(g30262) ) ;
INV     gate16954  (.A(g30262), .Z(II40075) ) ;
INV     gate16955  (.A(II40075), .Z(g30493) ) ;
NOR2    gate16956  (.A(g16344), .B(g30097), .Z(g30263) ) ;
INV     gate16957  (.A(g30263), .Z(II40078) ) ;
INV     gate16958  (.A(II40078), .Z(g30494) ) ;
NOR2    gate16959  (.A(g16348), .B(g30098), .Z(g30264) ) ;
INV     gate16960  (.A(g30264), .Z(II40083) ) ;
INV     gate16961  (.A(II40083), .Z(g30497) ) ;
NOR2    gate16962  (.A(g16349), .B(g30099), .Z(g30265) ) ;
INV     gate16963  (.A(g30265), .Z(II40086) ) ;
INV     gate16964  (.A(II40086), .Z(g30498) ) ;
NOR2    gate16965  (.A(g16359), .B(g30100), .Z(g30266) ) ;
INV     gate16966  (.A(g30266), .Z(II40091) ) ;
INV     gate16967  (.A(II40091), .Z(g30501) ) ;
INV     gate16968  (.A(g30491), .Z(II40098) ) ;
INV     gate16969  (.A(g30326), .Z(II40101) ) ;
INV     gate16970  (.A(g30342), .Z(II40104) ) ;
INV     gate16971  (.A(g30343), .Z(II40107) ) ;
INV     gate16972  (.A(g30357), .Z(II40110) ) ;
INV     gate16973  (.A(g30368), .Z(II40113) ) ;
INV     gate16974  (.A(g30408), .Z(II40116) ) ;
INV     gate16975  (.A(g30435), .Z(II40119) ) ;
INV     gate16976  (.A(g30443), .Z(II40122) ) ;
INV     gate16977  (.A(g30466), .Z(II40125) ) ;
INV     gate16978  (.A(g30479), .Z(II40128) ) ;
INV     gate16979  (.A(g30493), .Z(II40131) ) ;
INV     gate16980  (.A(g30480), .Z(II40134) ) ;
INV     gate16981  (.A(g30494), .Z(II40137) ) ;
INV     gate16982  (.A(g30328), .Z(II40140) ) ;
INV     gate16983  (.A(g30329), .Z(II40143) ) ;
INV     gate16984  (.A(g30344), .Z(II40146) ) ;
INV     gate16985  (.A(g30358), .Z(II40149) ) ;
INV     gate16986  (.A(g30359), .Z(II40152) ) ;
INV     gate16987  (.A(g30369), .Z(II40155) ) ;
INV     gate16988  (.A(g30376), .Z(II40158) ) ;
INV     gate16989  (.A(g30439), .Z(II40161) ) ;
INV     gate16990  (.A(g30446), .Z(II40164) ) ;
INV     gate16991  (.A(g30456), .Z(II40167) ) ;
INV     gate16992  (.A(g30483), .Z(II40170) ) ;
INV     gate16993  (.A(g30497), .Z(II40173) ) ;
INV     gate16994  (.A(g30331), .Z(II40176) ) ;
INV     gate16995  (.A(g30498), .Z(II40179) ) ;
INV     gate16996  (.A(g30332), .Z(II40182) ) ;
INV     gate16997  (.A(g30346), .Z(II40185) ) ;
INV     gate16998  (.A(g30347), .Z(II40188) ) ;
INV     gate16999  (.A(g30360), .Z(II40191) ) ;
INV     gate17000  (.A(g30370), .Z(II40194) ) ;
INV     gate17001  (.A(g30371), .Z(II40197) ) ;
INV     gate17002  (.A(g30377), .Z(II40200) ) ;
INV     gate17003  (.A(g30380), .Z(II40203) ) ;
INV     gate17004  (.A(g30450), .Z(II40206) ) ;
INV     gate17005  (.A(g30459), .Z(II40209) ) ;
INV     gate17006  (.A(g30471), .Z(II40212) ) ;
INV     gate17007  (.A(g30501), .Z(II40215) ) ;
INV     gate17008  (.A(g30335), .Z(II40218) ) ;
INV     gate17009  (.A(g30349), .Z(II40221) ) ;
INV     gate17010  (.A(g30336), .Z(II40224) ) ;
INV     gate17011  (.A(g30350), .Z(II40227) ) ;
INV     gate17012  (.A(g30362), .Z(II40230) ) ;
INV     gate17013  (.A(g30363), .Z(II40233) ) ;
INV     gate17014  (.A(g30373), .Z(II40236) ) ;
INV     gate17015  (.A(g30378), .Z(II40239) ) ;
INV     gate17016  (.A(g30379), .Z(II40242) ) ;
INV     gate17017  (.A(g30381), .Z(II40245) ) ;
INV     gate17018  (.A(g30382), .Z(II40248) ) ;
INV     gate17019  (.A(g30463), .Z(II40251) ) ;
INV     gate17020  (.A(g30474), .Z(II40254) ) ;
INV     gate17021  (.A(g30488), .Z(II40257) ) ;
INV     gate17022  (.A(g30339), .Z(II40260) ) ;
INV     gate17023  (.A(g30353), .Z(II40263) ) ;
INV     gate17024  (.A(g30365), .Z(II40266) ) ;
INV     gate17025  (.A(g30354), .Z(II40269) ) ;
INV     gate17026  (.A(g30366), .Z(II40272) ) ;
INV     gate17027  (.A(g30375), .Z(II40275) ) ;
NOR2    gate17028  (.A(g30004), .B(g30131), .Z(g30403) ) ;
INV     gate17029  (.A(g30403), .Z(g30567) ) ;
NOR2    gate17030  (.A(g29999), .B(g30129), .Z(g30402) ) ;
INV     gate17031  (.A(g30402), .Z(g30568) ) ;
NOR2    gate17032  (.A(g30009), .B(g30138), .Z(g30406) ) ;
INV     gate17033  (.A(g30406), .Z(g30569) ) ;
NOR2    gate17034  (.A(g30006), .B(g30132), .Z(g30404) ) ;
INV     gate17035  (.A(g30404), .Z(g30570) ) ;
NOR2    gate17036  (.A(g29998), .B(g30128), .Z(g30401) ) ;
INV     gate17037  (.A(g30401), .Z(g30571) ) ;
NOR2    gate17038  (.A(g30116), .B(g30123), .Z(g30399) ) ;
INV     gate17039  (.A(g30399), .Z(g30572) ) ;
NOR2    gate17040  (.A(g30008), .B(g30133), .Z(g30405) ) ;
INV     gate17041  (.A(g30405), .Z(g30573) ) ;
NOR2    gate17042  (.A(g29997), .B(g30127), .Z(g30400) ) ;
INV     gate17043  (.A(g30400), .Z(g30574) ) ;
INV     gate17044  (.A(g30412), .Z(g30575) ) ;
NOR2    gate17045  (.A(g13953), .B(g30216), .Z(g30455) ) ;
INV     gate17046  (.A(g30455), .Z(II40288) ) ;
INV     gate17047  (.A(II40288), .Z(g30578) ) ;
NOR2    gate17048  (.A(g14007), .B(g30217), .Z(g30468) ) ;
INV     gate17049  (.A(g30468), .Z(II40291) ) ;
INV     gate17050  (.A(II40291), .Z(g30579) ) ;
NOR2    gate17051  (.A(g14023), .B(g30218), .Z(g30470) ) ;
INV     gate17052  (.A(g30470), .Z(II40294) ) ;
INV     gate17053  (.A(II40294), .Z(g30580) ) ;
NOR2    gate17054  (.A(g14067), .B(g30219), .Z(g30482) ) ;
INV     gate17055  (.A(g30482), .Z(II40297) ) ;
INV     gate17056  (.A(II40297), .Z(g30581) ) ;
NOR2    gate17057  (.A(g14098), .B(g30220), .Z(g30485) ) ;
INV     gate17058  (.A(g30485), .Z(II40300) ) ;
INV     gate17059  (.A(II40300), .Z(g30582) ) ;
NOR2    gate17060  (.A(g14114), .B(g30221), .Z(g30487) ) ;
INV     gate17061  (.A(g30487), .Z(II40303) ) ;
INV     gate17062  (.A(II40303), .Z(g30583) ) ;
NOR2    gate17063  (.A(g14182), .B(g30222), .Z(g30500) ) ;
INV     gate17064  (.A(g30500), .Z(II40307) ) ;
INV     gate17065  (.A(II40307), .Z(g30585) ) ;
NOR2    gate17066  (.A(g14213), .B(g30223), .Z(g30503) ) ;
INV     gate17067  (.A(g30503), .Z(II40310) ) ;
INV     gate17068  (.A(II40310), .Z(g30586) ) ;
NOR2    gate17069  (.A(g14229), .B(g30224), .Z(g30505) ) ;
INV     gate17070  (.A(g30505), .Z(II40313) ) ;
INV     gate17071  (.A(II40313), .Z(g30587) ) ;
NOR2    gate17072  (.A(g14297), .B(g30225), .Z(g30338) ) ;
INV     gate17073  (.A(g30338), .Z(II40317) ) ;
INV     gate17074  (.A(II40317), .Z(g30591) ) ;
NOR2    gate17075  (.A(g14328), .B(g30226), .Z(g30341) ) ;
INV     gate17076  (.A(g30341), .Z(II40320) ) ;
INV     gate17077  (.A(II40320), .Z(g30592) ) ;
NOR2    gate17078  (.A(g14419), .B(g30227), .Z(g30356) ) ;
INV     gate17079  (.A(g30356), .Z(II40326) ) ;
INV     gate17080  (.A(II40326), .Z(g30600) ) ;
INV     gate17081  (.A(g30578), .Z(II40420) ) ;
INV     gate17082  (.A(g30579), .Z(II40423) ) ;
INV     gate17083  (.A(g30581), .Z(II40426) ) ;
INV     gate17084  (.A(g30580), .Z(II40429) ) ;
INV     gate17085  (.A(g30582), .Z(II40432) ) ;
INV     gate17086  (.A(g30585), .Z(II40435) ) ;
INV     gate17087  (.A(g30583), .Z(II40438) ) ;
INV     gate17088  (.A(g30586), .Z(II40441) ) ;
INV     gate17089  (.A(g30591), .Z(II40444) ) ;
INV     gate17090  (.A(g30587), .Z(II40447) ) ;
INV     gate17091  (.A(g30592), .Z(II40450) ) ;
INV     gate17092  (.A(g30600), .Z(II40453) ) ;
NOR2    gate17093  (.A(g16381), .B(g30478), .Z(g30668) ) ;
INV     gate17094  (.A(g30668), .Z(II40456) ) ;
INV     gate17095  (.A(II40456), .Z(g30722) ) ;
NOR2    gate17096  (.A(g16383), .B(g30481), .Z(g30669) ) ;
INV     gate17097  (.A(g30669), .Z(II40459) ) ;
INV     gate17098  (.A(II40459), .Z(g30723) ) ;
NOR2    gate17099  (.A(g16389), .B(g30484), .Z(g30670) ) ;
INV     gate17100  (.A(g30670), .Z(II40462) ) ;
INV     gate17101  (.A(II40462), .Z(g30724) ) ;
NOR2    gate17102  (.A(g16391), .B(g30486), .Z(g30671) ) ;
INV     gate17103  (.A(g30671), .Z(II40465) ) ;
INV     gate17104  (.A(II40465), .Z(g30725) ) ;
NOR2    gate17105  (.A(g16401), .B(g30489), .Z(g30672) ) ;
INV     gate17106  (.A(g30672), .Z(II40468) ) ;
INV     gate17107  (.A(II40468), .Z(g30726) ) ;
NOR2    gate17108  (.A(g16402), .B(g30490), .Z(g30673) ) ;
INV     gate17109  (.A(g30673), .Z(II40471) ) ;
INV     gate17110  (.A(II40471), .Z(g30727) ) ;
NOR2    gate17111  (.A(g16414), .B(g30492), .Z(g30674) ) ;
INV     gate17112  (.A(g30674), .Z(II40475) ) ;
INV     gate17113  (.A(II40475), .Z(g30729) ) ;
NOR2    gate17114  (.A(g16416), .B(g30495), .Z(g30675) ) ;
INV     gate17115  (.A(g30675), .Z(II40478) ) ;
INV     gate17116  (.A(II40478), .Z(g30730) ) ;
NOR2    gate17117  (.A(g16419), .B(g30496), .Z(g30676) ) ;
INV     gate17118  (.A(g30676), .Z(II40481) ) ;
INV     gate17119  (.A(II40481), .Z(g30731) ) ;
NOR2    gate17120  (.A(g16421), .B(g30499), .Z(g30677) ) ;
INV     gate17121  (.A(g30677), .Z(II40484) ) ;
INV     gate17122  (.A(II40484), .Z(g30732) ) ;
NOR2    gate17123  (.A(g16427), .B(g30502), .Z(g30678) ) ;
INV     gate17124  (.A(g30678), .Z(II40487) ) ;
INV     gate17125  (.A(II40487), .Z(g30733) ) ;
NOR2    gate17126  (.A(g16429), .B(g30504), .Z(g30679) ) ;
INV     gate17127  (.A(g30679), .Z(II40490) ) ;
INV     gate17128  (.A(II40490), .Z(g30734) ) ;
NOR2    gate17129  (.A(g16443), .B(g30327), .Z(g30680) ) ;
INV     gate17130  (.A(g30680), .Z(II40495) ) ;
INV     gate17131  (.A(II40495), .Z(g30737) ) ;
NOR2    gate17132  (.A(g16448), .B(g30330), .Z(g30681) ) ;
INV     gate17133  (.A(g30681), .Z(II40498) ) ;
INV     gate17134  (.A(II40498), .Z(g30738) ) ;
NOR2    gate17135  (.A(g16450), .B(g30333), .Z(g30682) ) ;
INV     gate17136  (.A(g30682), .Z(II40501) ) ;
INV     gate17137  (.A(II40501), .Z(g30739) ) ;
NOR2    gate17138  (.A(g16453), .B(g30334), .Z(g30683) ) ;
INV     gate17139  (.A(g30683), .Z(II40504) ) ;
INV     gate17140  (.A(II40504), .Z(g30740) ) ;
NOR2    gate17141  (.A(g16455), .B(g30337), .Z(g30684) ) ;
INV     gate17142  (.A(g30684), .Z(II40507) ) ;
INV     gate17143  (.A(II40507), .Z(g30741) ) ;
NOR2    gate17144  (.A(g16461), .B(g30340), .Z(g30686) ) ;
INV     gate17145  (.A(g30686), .Z(II40510) ) ;
INV     gate17146  (.A(II40510), .Z(g30742) ) ;
NOR2    gate17147  (.A(g13479), .B(g30345), .Z(g30687) ) ;
INV     gate17148  (.A(g30687), .Z(II40515) ) ;
INV     gate17149  (.A(II40515), .Z(g30745) ) ;
NOR2    gate17150  (.A(g13484), .B(g30348), .Z(g30688) ) ;
INV     gate17151  (.A(g30688), .Z(II40518) ) ;
INV     gate17152  (.A(II40518), .Z(g30746) ) ;
NOR2    gate17153  (.A(g13486), .B(g30351), .Z(g30689) ) ;
INV     gate17154  (.A(g30689), .Z(II40521) ) ;
INV     gate17155  (.A(II40521), .Z(g30747) ) ;
NOR2    gate17156  (.A(g13489), .B(g30352), .Z(g30690) ) ;
INV     gate17157  (.A(g30690), .Z(II40524) ) ;
INV     gate17158  (.A(II40524), .Z(g30748) ) ;
NOR2    gate17159  (.A(g13491), .B(g30355), .Z(g30691) ) ;
INV     gate17160  (.A(g30691), .Z(II40527) ) ;
INV     gate17161  (.A(II40527), .Z(g30749) ) ;
NOR2    gate17162  (.A(g13498), .B(g30361), .Z(g30692) ) ;
INV     gate17163  (.A(g30692), .Z(II40531) ) ;
INV     gate17164  (.A(II40531), .Z(g30751) ) ;
NOR2    gate17165  (.A(g13503), .B(g30364), .Z(g30693) ) ;
INV     gate17166  (.A(g30693), .Z(II40534) ) ;
INV     gate17167  (.A(II40534), .Z(g30752) ) ;
NOR2    gate17168  (.A(g13505), .B(g30367), .Z(g30694) ) ;
INV     gate17169  (.A(g30694), .Z(II40537) ) ;
INV     gate17170  (.A(II40537), .Z(g30753) ) ;
NOR2    gate17171  (.A(g13515), .B(g30374), .Z(g30695) ) ;
INV     gate17172  (.A(g30695), .Z(II40542) ) ;
INV     gate17173  (.A(II40542), .Z(g30756) ) ;
NOR3    gate17174  (.A(g29992), .B(g30000), .C(g30372), .Z(g30685) ) ;
INV     gate17175  (.A(g30685), .Z(g30765) ) ;
NOR2    gate17176  (.A(g13914), .B(g30387), .Z(g30699) ) ;
INV     gate17177  (.A(g30699), .Z(II40555) ) ;
INV     gate17178  (.A(II40555), .Z(g30767) ) ;
NOR2    gate17179  (.A(g13952), .B(g30388), .Z(g30700) ) ;
INV     gate17180  (.A(g30700), .Z(II40565) ) ;
INV     gate17181  (.A(II40565), .Z(g30769) ) ;
NOR2    gate17182  (.A(g13970), .B(g30389), .Z(g30701) ) ;
INV     gate17183  (.A(g30701), .Z(II40568) ) ;
INV     gate17184  (.A(II40568), .Z(g30770) ) ;
NOR2    gate17185  (.A(g14006), .B(g30390), .Z(g30702) ) ;
INV     gate17186  (.A(g30702), .Z(II40578) ) ;
INV     gate17187  (.A(II40578), .Z(g30772) ) ;
NOR2    gate17188  (.A(g14022), .B(g30391), .Z(g30703) ) ;
INV     gate17189  (.A(g30703), .Z(II40581) ) ;
INV     gate17190  (.A(II40581), .Z(g30773) ) ;
NOR2    gate17191  (.A(g14040), .B(g30392), .Z(g30704) ) ;
INV     gate17192  (.A(g30704), .Z(II40584) ) ;
INV     gate17193  (.A(II40584), .Z(g30774) ) ;
NOR2    gate17194  (.A(g14097), .B(g30393), .Z(g30705) ) ;
INV     gate17195  (.A(g30705), .Z(II40594) ) ;
INV     gate17196  (.A(II40594), .Z(g30776) ) ;
NOR2    gate17197  (.A(g14113), .B(g30394), .Z(g30706) ) ;
INV     gate17198  (.A(g30706), .Z(II40597) ) ;
INV     gate17199  (.A(II40597), .Z(g30777) ) ;
NOR2    gate17200  (.A(g14131), .B(g30395), .Z(g30707) ) ;
INV     gate17201  (.A(g30707), .Z(II40600) ) ;
INV     gate17202  (.A(II40600), .Z(g30778) ) ;
NOR2    gate17203  (.A(g14212), .B(g30396), .Z(g30708) ) ;
INV     gate17204  (.A(g30708), .Z(II40611) ) ;
INV     gate17205  (.A(II40611), .Z(g30781) ) ;
NOR2    gate17206  (.A(g14228), .B(g30397), .Z(g30709) ) ;
INV     gate17207  (.A(g30709), .Z(II40614) ) ;
INV     gate17208  (.A(II40614), .Z(g30782) ) ;
NOR2    gate17209  (.A(g14327), .B(g30398), .Z(g30566) ) ;
INV     gate17210  (.A(g30566), .Z(II40618) ) ;
INV     gate17211  (.A(II40618), .Z(g30784) ) ;
INV     gate17212  (.A(g30571), .Z(II40634) ) ;
INV     gate17213  (.A(II40634), .Z(g30792) ) ;
INV     gate17214  (.A(g30570), .Z(II40637) ) ;
INV     gate17215  (.A(II40637), .Z(g30793) ) ;
INV     gate17216  (.A(g30569), .Z(II40640) ) ;
INV     gate17217  (.A(II40640), .Z(g30794) ) ;
INV     gate17218  (.A(g30568), .Z(II40643) ) ;
INV     gate17219  (.A(II40643), .Z(g30795) ) ;
INV     gate17220  (.A(g30567), .Z(II40647) ) ;
INV     gate17221  (.A(II40647), .Z(g30797) ) ;
INV     gate17222  (.A(g30574), .Z(II40651) ) ;
INV     gate17223  (.A(II40651), .Z(g30799) ) ;
INV     gate17224  (.A(g30573), .Z(II40654) ) ;
INV     gate17225  (.A(II40654), .Z(g30800) ) ;
INV     gate17226  (.A(g30572), .Z(II40658) ) ;
INV     gate17227  (.A(II40658), .Z(g30802) ) ;
NOR2    gate17228  (.A(g16108), .B(g30407), .Z(g30635) ) ;
INV     gate17229  (.A(g30635), .Z(II40661) ) ;
INV     gate17230  (.A(II40661), .Z(g30803) ) ;
NOR2    gate17231  (.A(g16140), .B(g30409), .Z(g30636) ) ;
INV     gate17232  (.A(g30636), .Z(II40664) ) ;
INV     gate17233  (.A(II40664), .Z(g30804) ) ;
NOR2    gate17234  (.A(g16141), .B(g30410), .Z(g30637) ) ;
INV     gate17235  (.A(g30637), .Z(II40667) ) ;
INV     gate17236  (.A(II40667), .Z(g30805) ) ;
NOR2    gate17237  (.A(g16159), .B(g30411), .Z(g30638) ) ;
INV     gate17238  (.A(g30638), .Z(II40670) ) ;
INV     gate17239  (.A(II40670), .Z(g30806) ) ;
NOR2    gate17240  (.A(g16186), .B(g30436), .Z(g30639) ) ;
INV     gate17241  (.A(g30639), .Z(II40673) ) ;
INV     gate17242  (.A(II40673), .Z(g30807) ) ;
NOR2    gate17243  (.A(g16187), .B(g30437), .Z(g30640) ) ;
INV     gate17244  (.A(g30640), .Z(II40676) ) ;
INV     gate17245  (.A(II40676), .Z(g30808) ) ;
NOR2    gate17246  (.A(g16188), .B(g30438), .Z(g30641) ) ;
INV     gate17247  (.A(g30641), .Z(II40679) ) ;
INV     gate17248  (.A(II40679), .Z(g30809) ) ;
NOR2    gate17249  (.A(g16199), .B(g30440), .Z(g30642) ) ;
INV     gate17250  (.A(g30642), .Z(II40682) ) ;
INV     gate17251  (.A(II40682), .Z(g30810) ) ;
NOR2    gate17252  (.A(g16200), .B(g30441), .Z(g30643) ) ;
INV     gate17253  (.A(g30643), .Z(II40685) ) ;
INV     gate17254  (.A(II40685), .Z(g30811) ) ;
NOR2    gate17255  (.A(g16218), .B(g30442), .Z(g30644) ) ;
INV     gate17256  (.A(g30644), .Z(II40688) ) ;
INV     gate17257  (.A(II40688), .Z(g30812) ) ;
NOR2    gate17258  (.A(g16240), .B(g30444), .Z(g30645) ) ;
INV     gate17259  (.A(g30645), .Z(II40691) ) ;
INV     gate17260  (.A(II40691), .Z(g30813) ) ;
NOR2    gate17261  (.A(g16241), .B(g30445), .Z(g30646) ) ;
INV     gate17262  (.A(g30646), .Z(II40694) ) ;
INV     gate17263  (.A(II40694), .Z(g30814) ) ;
NOR2    gate17264  (.A(g16251), .B(g30447), .Z(g30647) ) ;
INV     gate17265  (.A(g30647), .Z(II40697) ) ;
INV     gate17266  (.A(II40697), .Z(g30815) ) ;
NOR2    gate17267  (.A(g16252), .B(g30448), .Z(g30648) ) ;
INV     gate17268  (.A(g30648), .Z(II40700) ) ;
INV     gate17269  (.A(II40700), .Z(g30816) ) ;
NOR2    gate17270  (.A(g16253), .B(g30449), .Z(g30649) ) ;
INV     gate17271  (.A(g30649), .Z(II40703) ) ;
INV     gate17272  (.A(II40703), .Z(g30817) ) ;
NOR2    gate17273  (.A(g16264), .B(g30451), .Z(g30650) ) ;
INV     gate17274  (.A(g30650), .Z(II40706) ) ;
INV     gate17275  (.A(II40706), .Z(g30818) ) ;
NOR2    gate17276  (.A(g16265), .B(g30452), .Z(g30651) ) ;
INV     gate17277  (.A(g30651), .Z(II40709) ) ;
INV     gate17278  (.A(II40709), .Z(g30819) ) ;
NOR2    gate17279  (.A(g16283), .B(g30453), .Z(g30652) ) ;
INV     gate17280  (.A(g30652), .Z(II40712) ) ;
INV     gate17281  (.A(II40712), .Z(g30820) ) ;
NOR2    gate17282  (.A(g16289), .B(g30454), .Z(g30653) ) ;
INV     gate17283  (.A(g30653), .Z(II40715) ) ;
INV     gate17284  (.A(II40715), .Z(g30821) ) ;
NOR2    gate17285  (.A(g16299), .B(g30457), .Z(g30654) ) ;
INV     gate17286  (.A(g30654), .Z(II40718) ) ;
INV     gate17287  (.A(II40718), .Z(g30822) ) ;
NOR2    gate17288  (.A(g16300), .B(g30458), .Z(g30655) ) ;
INV     gate17289  (.A(g30655), .Z(II40721) ) ;
INV     gate17290  (.A(II40721), .Z(g30823) ) ;
NOR2    gate17291  (.A(g16310), .B(g30460), .Z(g30656) ) ;
INV     gate17292  (.A(g30656), .Z(II40724) ) ;
INV     gate17293  (.A(II40724), .Z(g30824) ) ;
NOR2    gate17294  (.A(g16311), .B(g30461), .Z(g30657) ) ;
INV     gate17295  (.A(g30657), .Z(II40727) ) ;
INV     gate17296  (.A(II40727), .Z(g30825) ) ;
NOR2    gate17297  (.A(g16312), .B(g30462), .Z(g30658) ) ;
INV     gate17298  (.A(g30658), .Z(II40730) ) ;
INV     gate17299  (.A(II40730), .Z(g30826) ) ;
NOR2    gate17300  (.A(g16323), .B(g30464), .Z(g30659) ) ;
INV     gate17301  (.A(g30659), .Z(II40733) ) ;
INV     gate17302  (.A(II40733), .Z(g30827) ) ;
NOR2    gate17303  (.A(g16324), .B(g30465), .Z(g30660) ) ;
INV     gate17304  (.A(g30660), .Z(II40736) ) ;
INV     gate17305  (.A(II40736), .Z(g30828) ) ;
NOR2    gate17306  (.A(g16345), .B(g30467), .Z(g30661) ) ;
INV     gate17307  (.A(g30661), .Z(II40739) ) ;
INV     gate17308  (.A(II40739), .Z(g30829) ) ;
NOR2    gate17309  (.A(g16347), .B(g30469), .Z(g30662) ) ;
INV     gate17310  (.A(g30662), .Z(II40742) ) ;
INV     gate17311  (.A(II40742), .Z(g30830) ) ;
NOR2    gate17312  (.A(g16357), .B(g30472), .Z(g30663) ) ;
INV     gate17313  (.A(g30663), .Z(II40745) ) ;
INV     gate17314  (.A(II40745), .Z(g30831) ) ;
NOR2    gate17315  (.A(g16358), .B(g30473), .Z(g30664) ) ;
INV     gate17316  (.A(g30664), .Z(II40748) ) ;
INV     gate17317  (.A(II40748), .Z(g30832) ) ;
NOR2    gate17318  (.A(g16368), .B(g30475), .Z(g30665) ) ;
INV     gate17319  (.A(g30665), .Z(II40751) ) ;
INV     gate17320  (.A(II40751), .Z(g30833) ) ;
NOR2    gate17321  (.A(g16369), .B(g30476), .Z(g30666) ) ;
INV     gate17322  (.A(g30666), .Z(II40754) ) ;
INV     gate17323  (.A(II40754), .Z(g30834) ) ;
NOR2    gate17324  (.A(g16370), .B(g30477), .Z(g30667) ) ;
INV     gate17325  (.A(g30667), .Z(II40757) ) ;
INV     gate17326  (.A(II40757), .Z(g30835) ) ;
INV     gate17327  (.A(g30722), .Z(II40760) ) ;
INV     gate17328  (.A(g30729), .Z(II40763) ) ;
INV     gate17329  (.A(g30737), .Z(II40766) ) ;
INV     gate17330  (.A(g30803), .Z(II40769) ) ;
INV     gate17331  (.A(g30804), .Z(II40772) ) ;
INV     gate17332  (.A(g30807), .Z(II40775) ) ;
INV     gate17333  (.A(g30805), .Z(II40778) ) ;
INV     gate17334  (.A(g30808), .Z(II40781) ) ;
INV     gate17335  (.A(g30813), .Z(II40784) ) ;
INV     gate17336  (.A(g30809), .Z(II40787) ) ;
INV     gate17337  (.A(g30814), .Z(II40790) ) ;
INV     gate17338  (.A(g30821), .Z(II40793) ) ;
INV     gate17339  (.A(g30829), .Z(II40796) ) ;
INV     gate17340  (.A(g30723), .Z(II40799) ) ;
INV     gate17341  (.A(g30730), .Z(II40802) ) ;
INV     gate17342  (.A(g30767), .Z(II40805) ) ;
INV     gate17343  (.A(g30769), .Z(II40808) ) ;
INV     gate17344  (.A(g30772), .Z(II40811) ) ;
INV     gate17345  (.A(g30731), .Z(II40814) ) ;
INV     gate17346  (.A(g30738), .Z(II40817) ) ;
INV     gate17347  (.A(g30745), .Z(II40820) ) ;
INV     gate17348  (.A(g30806), .Z(II40823) ) ;
INV     gate17349  (.A(g30810), .Z(II40826) ) ;
INV     gate17350  (.A(g30815), .Z(II40829) ) ;
INV     gate17351  (.A(g30811), .Z(II40832) ) ;
INV     gate17352  (.A(g30816), .Z(II40835) ) ;
INV     gate17353  (.A(g30822), .Z(II40838) ) ;
INV     gate17354  (.A(g30817), .Z(II40841) ) ;
INV     gate17355  (.A(g30823), .Z(II40844) ) ;
INV     gate17356  (.A(g30830), .Z(II40847) ) ;
INV     gate17357  (.A(g30724), .Z(II40850) ) ;
INV     gate17358  (.A(g30732), .Z(II40853) ) ;
INV     gate17359  (.A(g30739), .Z(II40856) ) ;
INV     gate17360  (.A(g30770), .Z(II40859) ) ;
INV     gate17361  (.A(g30773), .Z(II40862) ) ;
INV     gate17362  (.A(g30776), .Z(II40865) ) ;
INV     gate17363  (.A(g30740), .Z(II40868) ) ;
INV     gate17364  (.A(g30746), .Z(II40871) ) ;
INV     gate17365  (.A(g30751), .Z(II40874) ) ;
INV     gate17366  (.A(g30812), .Z(II40877) ) ;
INV     gate17367  (.A(g30818), .Z(II40880) ) ;
INV     gate17368  (.A(g30824), .Z(II40883) ) ;
INV     gate17369  (.A(g30819), .Z(II40886) ) ;
INV     gate17370  (.A(g30825), .Z(II40889) ) ;
INV     gate17371  (.A(g30831), .Z(II40892) ) ;
INV     gate17372  (.A(g30826), .Z(II40895) ) ;
INV     gate17373  (.A(g30832), .Z(II40898) ) ;
INV     gate17374  (.A(g30725), .Z(II40901) ) ;
INV     gate17375  (.A(g30733), .Z(II40904) ) ;
INV     gate17376  (.A(g30741), .Z(II40907) ) ;
INV     gate17377  (.A(g30747), .Z(II40910) ) ;
INV     gate17378  (.A(g30774), .Z(II40913) ) ;
INV     gate17379  (.A(g30777), .Z(II40916) ) ;
INV     gate17380  (.A(g30781), .Z(II40919) ) ;
INV     gate17381  (.A(g30748), .Z(II40922) ) ;
INV     gate17382  (.A(g30752), .Z(II40925) ) ;
INV     gate17383  (.A(g30756), .Z(II40928) ) ;
INV     gate17384  (.A(g30820), .Z(II40931) ) ;
INV     gate17385  (.A(g30827), .Z(II40934) ) ;
INV     gate17386  (.A(g30833), .Z(II40937) ) ;
INV     gate17387  (.A(g30828), .Z(II40940) ) ;
INV     gate17388  (.A(g30834), .Z(II40943) ) ;
INV     gate17389  (.A(g30726), .Z(II40946) ) ;
INV     gate17390  (.A(g30835), .Z(II40949) ) ;
INV     gate17391  (.A(g30727), .Z(II40952) ) ;
INV     gate17392  (.A(g30734), .Z(II40955) ) ;
INV     gate17393  (.A(g30742), .Z(II40958) ) ;
INV     gate17394  (.A(g30749), .Z(II40961) ) ;
INV     gate17395  (.A(g30753), .Z(II40964) ) ;
INV     gate17396  (.A(g30778), .Z(II40967) ) ;
INV     gate17397  (.A(g30782), .Z(II40970) ) ;
INV     gate17398  (.A(g30784), .Z(II40973) ) ;
INV     gate17399  (.A(g30799), .Z(II40976) ) ;
INV     gate17400  (.A(g30800), .Z(II40979) ) ;
INV     gate17401  (.A(g30802), .Z(II40982) ) ;
INV     gate17402  (.A(g30792), .Z(II40985) ) ;
INV     gate17403  (.A(g30793), .Z(II40988) ) ;
INV     gate17404  (.A(g30794), .Z(II40991) ) ;
INV     gate17405  (.A(g30795), .Z(II40994) ) ;
INV     gate17406  (.A(g30797), .Z(II40997) ) ;
INV     gate17407  (.A(g30765), .Z(II41024) ) ;
INV     gate17408  (.A(II41024), .Z(g30928) ) ;
NOR2    gate17409  (.A(g16069), .B(g30696), .Z(g30796) ) ;
INV     gate17410  (.A(g30796), .Z(II41035) ) ;
INV     gate17411  (.A(II41035), .Z(g30937) ) ;
NOR2    gate17412  (.A(g16134), .B(g30697), .Z(g30798) ) ;
INV     gate17413  (.A(g30798), .Z(II41038) ) ;
INV     gate17414  (.A(II41038), .Z(g30938) ) ;
NOR2    gate17415  (.A(g16237), .B(g30698), .Z(g30801) ) ;
INV     gate17416  (.A(g30801), .Z(II41041) ) ;
INV     gate17417  (.A(II41041), .Z(g30939) ) ;
INV     gate17418  (.A(g30928), .Z(II41044) ) ;
INV     gate17419  (.A(g30937), .Z(II41047) ) ;
INV     gate17420  (.A(g30938), .Z(II41050) ) ;
INV     gate17421  (.A(g30939), .Z(II41053) ) ;
NOR2    gate17422  (.A(g30922), .B(g30948), .Z(g30958) ) ;
INV     gate17423  (.A(g30958), .Z(g30962) ) ;
NOR2    gate17424  (.A(g30920), .B(g30947), .Z(g30957) ) ;
INV     gate17425  (.A(g30957), .Z(g30963) ) ;
NOR2    gate17426  (.A(g30925), .B(g30951), .Z(g30961) ) ;
INV     gate17427  (.A(g30961), .Z(g30964) ) ;
NOR2    gate17428  (.A(g30923), .B(g30949), .Z(g30959) ) ;
INV     gate17429  (.A(g30959), .Z(g30965) ) ;
NOR2    gate17430  (.A(g30919), .B(g30946), .Z(g30956) ) ;
INV     gate17431  (.A(g30956), .Z(g30966) ) ;
NOR2    gate17432  (.A(g30916), .B(g30944), .Z(g30954) ) ;
INV     gate17433  (.A(g30954), .Z(g30967) ) ;
NOR2    gate17434  (.A(g30924), .B(g30950), .Z(g30960) ) ;
INV     gate17435  (.A(g30960), .Z(g30968) ) ;
NOR2    gate17436  (.A(g30918), .B(g30945), .Z(g30955) ) ;
INV     gate17437  (.A(g30955), .Z(g30969) ) ;
NOR3    gate17438  (.A(g30917), .B(g30921), .C(g30953), .Z(g30970) ) ;
INV     gate17439  (.A(g30970), .Z(g30971) ) ;
INV     gate17440  (.A(g30965), .Z(II41090) ) ;
INV     gate17441  (.A(II41090), .Z(g30972) ) ;
INV     gate17442  (.A(g30964), .Z(II41093) ) ;
INV     gate17443  (.A(II41093), .Z(g30973) ) ;
INV     gate17444  (.A(g30963), .Z(II41096) ) ;
INV     gate17445  (.A(II41096), .Z(g30974) ) ;
INV     gate17446  (.A(g30962), .Z(II41099) ) ;
INV     gate17447  (.A(II41099), .Z(g30975) ) ;
INV     gate17448  (.A(g30969), .Z(II41102) ) ;
INV     gate17449  (.A(II41102), .Z(g30976) ) ;
INV     gate17450  (.A(g30968), .Z(II41105) ) ;
INV     gate17451  (.A(II41105), .Z(g30977) ) ;
INV     gate17452  (.A(g30967), .Z(II41108) ) ;
INV     gate17453  (.A(II41108), .Z(g30978) ) ;
INV     gate17454  (.A(g30966), .Z(II41111) ) ;
INV     gate17455  (.A(II41111), .Z(g30979) ) ;
INV     gate17456  (.A(g30976), .Z(II41114) ) ;
INV     gate17457  (.A(g30977), .Z(II41117) ) ;
INV     gate17458  (.A(g30978), .Z(II41120) ) ;
INV     gate17459  (.A(g30979), .Z(II41123) ) ;
INV     gate17460  (.A(g30972), .Z(II41126) ) ;
INV     gate17461  (.A(g30973), .Z(II41129) ) ;
INV     gate17462  (.A(g30974), .Z(II41132) ) ;
INV     gate17463  (.A(g30975), .Z(II41135) ) ;
INV     gate17464  (.A(g30971), .Z(II41138) ) ;
INV     gate17465  (.A(II41138), .Z(g30988) ) ;
INV     gate17466  (.A(g30988), .Z(II41141) ) ;
AND2    gate17467  (.A(g325), .B(g349), .Z(g5630) ) ;
AND2    gate17468  (.A(g331), .B(g351), .Z(g5649) ) ;
AND2    gate17469  (.A(g325), .B(g364), .Z(g5650) ) ;
AND2    gate17470  (.A(g1012), .B(g1036), .Z(g5658) ) ;
AND2    gate17471  (.A(g337), .B(g353), .Z(g5676) ) ;
AND2    gate17472  (.A(g331), .B(g366), .Z(g5677) ) ;
AND2    gate17473  (.A(g325), .B(g379), .Z(g5678) ) ;
AND2    gate17474  (.A(g1018), .B(g1038), .Z(g5687) ) ;
AND2    gate17475  (.A(g1012), .B(g1051), .Z(g5688) ) ;
AND2    gate17476  (.A(g1706), .B(g1730), .Z(g5696) ) ;
AND2    gate17477  (.A(g337), .B(g368), .Z(g5709) ) ;
AND2    gate17478  (.A(g331), .B(g381), .Z(g5710) ) ;
AND2    gate17479  (.A(g325), .B(g394), .Z(g5711) ) ;
AND2    gate17480  (.A(g1024), .B(g1040), .Z(g5728) ) ;
AND2    gate17481  (.A(g1018), .B(g1053), .Z(g5729) ) ;
AND2    gate17482  (.A(g1012), .B(g1066), .Z(g5730) ) ;
AND2    gate17483  (.A(g1712), .B(g1732), .Z(g5739) ) ;
AND2    gate17484  (.A(g1706), .B(g1745), .Z(g5740) ) ;
AND2    gate17485  (.A(g2400), .B(g2424), .Z(g5748) ) ;
AND2    gate17486  (.A(g337), .B(g383), .Z(g5757) ) ;
AND2    gate17487  (.A(g331), .B(g396), .Z(g5758) ) ;
AND2    gate17488  (.A(g1024), .B(g1055), .Z(g5767) ) ;
AND2    gate17489  (.A(g1018), .B(g1068), .Z(g5768) ) ;
AND2    gate17490  (.A(g1012), .B(g1081), .Z(g5769) ) ;
AND2    gate17491  (.A(g1718), .B(g1734), .Z(g5786) ) ;
AND2    gate17492  (.A(g1712), .B(g1747), .Z(g5787) ) ;
AND2    gate17493  (.A(g1706), .B(g1760), .Z(g5788) ) ;
AND2    gate17494  (.A(g2406), .B(g2426), .Z(g5797) ) ;
AND2    gate17495  (.A(g2400), .B(g2439), .Z(g5798) ) ;
AND2    gate17496  (.A(g337), .B(g324), .Z(g5807) ) ;
AND2    gate17497  (.A(g1024), .B(g1070), .Z(g5816) ) ;
AND2    gate17498  (.A(g1018), .B(g1083), .Z(g5817) ) ;
AND2    gate17499  (.A(g1718), .B(g1749), .Z(g5826) ) ;
AND2    gate17500  (.A(g1712), .B(g1762), .Z(g5827) ) ;
AND2    gate17501  (.A(g1706), .B(g1775), .Z(g5828) ) ;
AND2    gate17502  (.A(g2412), .B(g2428), .Z(g5845) ) ;
AND2    gate17503  (.A(g2406), .B(g2441), .Z(g5846) ) ;
AND2    gate17504  (.A(g2400), .B(g2454), .Z(g5847) ) ;
AND2    gate17505  (.A(g1024), .B(g1011), .Z(g5863) ) ;
AND2    gate17506  (.A(g1718), .B(g1764), .Z(g5872) ) ;
AND2    gate17507  (.A(g1712), .B(g1777), .Z(g5873) ) ;
AND2    gate17508  (.A(g2412), .B(g2443), .Z(g5882) ) ;
AND2    gate17509  (.A(g2406), .B(g2456), .Z(g5883) ) ;
AND2    gate17510  (.A(g2400), .B(g2469), .Z(g5884) ) ;
AND2    gate17511  (.A(g1718), .B(g1705), .Z(g5910) ) ;
AND2    gate17512  (.A(g2412), .B(g2458), .Z(g5919) ) ;
AND2    gate17513  (.A(g2406), .B(g2471), .Z(g5920) ) ;
AND2    gate17514  (.A(g2412), .B(g2399), .Z(g5949) ) ;
AND2    gate17515  (.A(g3254), .B(g219), .Z(g8327) ) ;
AND2    gate17516  (.A(g6314), .B(g225), .Z(g8328) ) ;
AND2    gate17517  (.A(g6232), .B(g231), .Z(g8329) ) ;
AND2    gate17518  (.A(g6519), .B(g903), .Z(g8339) ) ;
AND2    gate17519  (.A(g6369), .B(g909), .Z(g8340) ) ;
AND2    gate17520  (.A(g6574), .B(g1594), .Z(g8350) ) ;
AND2    gate17521  (.A(g3254), .B(g228), .Z(g8385) ) ;
AND2    gate17522  (.A(g6314), .B(g234), .Z(g8386) ) ;
AND2    gate17523  (.A(g6232), .B(g240), .Z(g8387) ) ;
AND2    gate17524  (.A(g3410), .B(g906), .Z(g8394) ) ;
AND2    gate17525  (.A(g6519), .B(g912), .Z(g8395) ) ;
AND2    gate17526  (.A(g6369), .B(g918), .Z(g8396) ) ;
AND2    gate17527  (.A(g6783), .B(g1597), .Z(g8406) ) ;
AND2    gate17528  (.A(g6574), .B(g1603), .Z(g8407) ) ;
AND2    gate17529  (.A(g6838), .B(g2288), .Z(g8417) ) ;
AND2    gate17530  (.A(g3254), .B(g237), .Z(g8431) ) ;
AND2    gate17531  (.A(g6314), .B(g243), .Z(g8432) ) ;
AND2    gate17532  (.A(g6232), .B(g249), .Z(g8433) ) ;
AND2    gate17533  (.A(g3410), .B(g915), .Z(g8437) ) ;
AND2    gate17534  (.A(g6519), .B(g921), .Z(g8438) ) ;
AND2    gate17535  (.A(g6369), .B(g927), .Z(g8439) ) ;
AND2    gate17536  (.A(g3566), .B(g1600), .Z(g8446) ) ;
AND2    gate17537  (.A(g6783), .B(g1606), .Z(g8447) ) ;
AND2    gate17538  (.A(g6574), .B(g1612), .Z(g8448) ) ;
AND2    gate17539  (.A(g7085), .B(g2291), .Z(g8458) ) ;
AND2    gate17540  (.A(g6838), .B(g2297), .Z(g8459) ) ;
AND2    gate17541  (.A(g3254), .B(g246), .Z(g8463) ) ;
AND2    gate17542  (.A(g6314), .B(g252), .Z(g8464) ) ;
AND2    gate17543  (.A(g6232), .B(g258), .Z(g8465) ) ;
AND2    gate17544  (.A(g3410), .B(g924), .Z(g8466) ) ;
AND2    gate17545  (.A(g6519), .B(g930), .Z(g8467) ) ;
AND2    gate17546  (.A(g6369), .B(g936), .Z(g8468) ) ;
AND2    gate17547  (.A(g3566), .B(g1609), .Z(g8472) ) ;
AND2    gate17548  (.A(g6783), .B(g1615), .Z(g8473) ) ;
AND2    gate17549  (.A(g6574), .B(g1621), .Z(g8474) ) ;
AND2    gate17550  (.A(g3722), .B(g2294), .Z(g8481) ) ;
AND2    gate17551  (.A(g7085), .B(g2300), .Z(g8482) ) ;
AND2    gate17552  (.A(g6838), .B(g2306), .Z(g8483) ) ;
AND2    gate17553  (.A(g6232), .B(g186), .Z(g8484) ) ;
AND2    gate17554  (.A(g3254), .B(g255), .Z(g8485) ) ;
AND2    gate17555  (.A(g6314), .B(g261), .Z(g8486) ) ;
AND2    gate17556  (.A(g6232), .B(g267), .Z(g8487) ) ;
AND2    gate17557  (.A(g3410), .B(g933), .Z(g8488) ) ;
AND2    gate17558  (.A(g6519), .B(g939), .Z(g8489) ) ;
AND2    gate17559  (.A(g6369), .B(g945), .Z(g8490) ) ;
AND2    gate17560  (.A(g3566), .B(g1618), .Z(g8491) ) ;
AND2    gate17561  (.A(g6783), .B(g1624), .Z(g8492) ) ;
AND2    gate17562  (.A(g6574), .B(g1630), .Z(g8493) ) ;
AND2    gate17563  (.A(g3722), .B(g2303), .Z(g8497) ) ;
AND2    gate17564  (.A(g7085), .B(g2309), .Z(g8498) ) ;
AND2    gate17565  (.A(g6838), .B(g2315), .Z(g8499) ) ;
AND2    gate17566  (.A(g6314), .B(g189), .Z(g8500) ) ;
AND2    gate17567  (.A(g6232), .B(g195), .Z(g8501) ) ;
AND2    gate17568  (.A(g3254), .B(g264), .Z(g8502) ) ;
AND2    gate17569  (.A(g6314), .B(g270), .Z(g8503) ) ;
AND2    gate17570  (.A(g6369), .B(g873), .Z(g8504) ) ;
AND2    gate17571  (.A(g3410), .B(g942), .Z(g8505) ) ;
AND2    gate17572  (.A(g6519), .B(g948), .Z(g8506) ) ;
AND2    gate17573  (.A(g6369), .B(g954), .Z(g8507) ) ;
AND2    gate17574  (.A(g3566), .B(g1627), .Z(g8508) ) ;
AND2    gate17575  (.A(g6783), .B(g1633), .Z(g8509) ) ;
AND2    gate17576  (.A(g6574), .B(g1639), .Z(g8510) ) ;
AND2    gate17577  (.A(g3722), .B(g2312), .Z(g8511) ) ;
AND2    gate17578  (.A(g7085), .B(g2318), .Z(g8512) ) ;
AND2    gate17579  (.A(g6838), .B(g2324), .Z(g8513) ) ;
AND2    gate17580  (.A(g3254), .B(g192), .Z(g8515) ) ;
AND2    gate17581  (.A(g6314), .B(g198), .Z(g8516) ) ;
AND2    gate17582  (.A(g6232), .B(g204), .Z(g8517) ) ;
AND2    gate17583  (.A(g3254), .B(g273), .Z(g8518) ) ;
AND2    gate17584  (.A(g6519), .B(g876), .Z(g8519) ) ;
AND2    gate17585  (.A(g6369), .B(g882), .Z(g8520) ) ;
AND2    gate17586  (.A(g3410), .B(g951), .Z(g8521) ) ;
AND2    gate17587  (.A(g6519), .B(g957), .Z(g8522) ) ;
AND2    gate17588  (.A(g6574), .B(g1567), .Z(g8523) ) ;
AND2    gate17589  (.A(g3566), .B(g1636), .Z(g8524) ) ;
AND2    gate17590  (.A(g6783), .B(g1642), .Z(g8525) ) ;
AND2    gate17591  (.A(g6574), .B(g1648), .Z(g8526) ) ;
AND2    gate17592  (.A(g3722), .B(g2321), .Z(g8527) ) ;
AND2    gate17593  (.A(g7085), .B(g2327), .Z(g8528) ) ;
AND2    gate17594  (.A(g6838), .B(g2333), .Z(g8529) ) ;
AND2    gate17595  (.A(g3254), .B(g201), .Z(g8531) ) ;
AND2    gate17596  (.A(g6314), .B(g207), .Z(g8532) ) ;
AND2    gate17597  (.A(g3410), .B(g879), .Z(g8534) ) ;
AND2    gate17598  (.A(g6519), .B(g885), .Z(g8535) ) ;
AND2    gate17599  (.A(g6369), .B(g891), .Z(g8536) ) ;
AND2    gate17600  (.A(g3410), .B(g960), .Z(g8537) ) ;
AND2    gate17601  (.A(g6783), .B(g1570), .Z(g8538) ) ;
AND2    gate17602  (.A(g6574), .B(g1576), .Z(g8539) ) ;
AND2    gate17603  (.A(g3566), .B(g1645), .Z(g8540) ) ;
AND2    gate17604  (.A(g6783), .B(g1651), .Z(g8541) ) ;
AND2    gate17605  (.A(g6838), .B(g2261), .Z(g8542) ) ;
AND2    gate17606  (.A(g3722), .B(g2330), .Z(g8543) ) ;
AND2    gate17607  (.A(g7085), .B(g2336), .Z(g8544) ) ;
AND2    gate17608  (.A(g6838), .B(g2342), .Z(g8545) ) ;
AND2    gate17609  (.A(g3254), .B(g210), .Z(g8546) ) ;
AND2    gate17610  (.A(g3410), .B(g888), .Z(g8548) ) ;
AND2    gate17611  (.A(g6519), .B(g894), .Z(g8549) ) ;
AND2    gate17612  (.A(g3566), .B(g1573), .Z(g8551) ) ;
AND2    gate17613  (.A(g6783), .B(g1579), .Z(g8552) ) ;
AND2    gate17614  (.A(g6574), .B(g1585), .Z(g8553) ) ;
AND2    gate17615  (.A(g3566), .B(g1654), .Z(g8554) ) ;
AND2    gate17616  (.A(g7085), .B(g2264), .Z(g8555) ) ;
AND2    gate17617  (.A(g6838), .B(g2270), .Z(g8556) ) ;
AND2    gate17618  (.A(g3722), .B(g2339), .Z(g8557) ) ;
AND2    gate17619  (.A(g7085), .B(g2345), .Z(g8558) ) ;
AND2    gate17620  (.A(g3410), .B(g897), .Z(g8559) ) ;
AND2    gate17621  (.A(g3566), .B(g1582), .Z(g8561) ) ;
AND2    gate17622  (.A(g6783), .B(g1588), .Z(g8562) ) ;
AND2    gate17623  (.A(g3722), .B(g2267), .Z(g8564) ) ;
AND2    gate17624  (.A(g7085), .B(g2273), .Z(g8565) ) ;
AND2    gate17625  (.A(g6838), .B(g2279), .Z(g8566) ) ;
AND2    gate17626  (.A(g3722), .B(g2348), .Z(g8567) ) ;
AND2    gate17627  (.A(g3566), .B(g1591), .Z(g8570) ) ;
AND2    gate17628  (.A(g3722), .B(g2276), .Z(g8572) ) ;
AND2    gate17629  (.A(g7085), .B(g2282), .Z(g8573) ) ;
AND2    gate17630  (.A(g3722), .B(g2285), .Z(g8576) ) ;
AND2    gate17631  (.A(g6643), .B(g7153), .Z(g8601) ) ;
AND2    gate17632  (.A(g3338), .B(g6908), .Z(g8612) ) ;
AND2    gate17633  (.A(g6945), .B(g7349), .Z(g8613) ) ;
AND2    gate17634  (.A(g6486), .B(g6672), .Z(g8621) ) ;
AND2    gate17635  (.A(g3494), .B(g7158), .Z(g8625) ) ;
AND2    gate17636  (.A(g7195), .B(g7479), .Z(g8626) ) ;
AND2    gate17637  (.A(g6751), .B(g6974), .Z(g8631) ) ;
AND2    gate17638  (.A(g3650), .B(g7354), .Z(g8635) ) ;
AND2    gate17639  (.A(g7391), .B(g7535), .Z(g8636) ) ;
AND2    gate17640  (.A(g7053), .B(g7224), .Z(g8650) ) ;
AND2    gate17641  (.A(g3806), .B(g7484), .Z(g8654) ) ;
AND2    gate17642  (.A(g7303), .B(g7420), .Z(g8666) ) ;
AND2    gate17643  (.A(g6643), .B(g7838), .Z(g8676) ) ;
AND2    gate17644  (.A(g3338), .B(g7827), .Z(g8687) ) ;
AND2    gate17645  (.A(g6945), .B(g7858), .Z(g8688) ) ;
AND2    gate17646  (.A(g6486), .B(g7819), .Z(g8703) ) ;
AND2    gate17647  (.A(g6643), .B(g7996), .Z(g8704) ) ;
AND2    gate17648  (.A(g3494), .B(g7842), .Z(g8705) ) ;
AND2    gate17649  (.A(g7195), .B(g7888), .Z(g8706) ) ;
AND2    gate17650  (.A(g3338), .B(g7953), .Z(g8717) ) ;
AND2    gate17651  (.A(g6751), .B(g7830), .Z(g8722) ) ;
AND2    gate17652  (.A(g6945), .B(g8071), .Z(g8723) ) ;
AND2    gate17653  (.A(g3650), .B(g7862), .Z(g8724) ) ;
AND2    gate17654  (.A(g7391), .B(g7912), .Z(g8725) ) ;
AND2    gate17655  (.A(g6486), .B(g7906), .Z(g8751) ) ;
AND2    gate17656  (.A(g3494), .B(g8004), .Z(g8755) ) ;
AND2    gate17657  (.A(g7053), .B(g7845), .Z(g8760) ) ;
AND2    gate17658  (.A(g7195), .B(g8156), .Z(g8761) ) ;
AND2    gate17659  (.A(g3806), .B(g7892), .Z(g8762) ) ;
AND2    gate17660  (.A(g6751), .B(g7958), .Z(g8774) ) ;
AND2    gate17661  (.A(g3650), .B(g8079), .Z(g8778) ) ;
AND2    gate17662  (.A(g7303), .B(g7865), .Z(g8783) ) ;
AND2    gate17663  (.A(g7391), .B(g8242), .Z(g8784) ) ;
AND2    gate17664  (.A(g7053), .B(g8009), .Z(g8797) ) ;
AND2    gate17665  (.A(g3806), .B(g8164), .Z(g8801) ) ;
AND2    gate17666  (.A(g7303), .B(g8084), .Z(g8816) ) ;
AND2    gate17667  (.A(g6486), .B(g490), .Z(g8841) ) ;
AND2    gate17668  (.A(g6512), .B(g5508), .Z(g8842) ) ;
AND2    gate17669  (.A(g6643), .B(g493), .Z(g8861) ) ;
AND2    gate17670  (.A(g6751), .B(g1177), .Z(g8868) ) ;
AND2    gate17671  (.A(g6776), .B(g5552), .Z(g8869) ) ;
AND2    gate17672  (.A(g3338), .B(g496), .Z(g8892) ) ;
AND2    gate17673  (.A(g6945), .B(g1180), .Z(g8899) ) ;
AND2    gate17674  (.A(g7053), .B(g1871), .Z(g8906) ) ;
AND2    gate17675  (.A(g7078), .B(g5598), .Z(g8907) ) ;
AND2    gate17676  (.A(g3494), .B(g1183), .Z(g8932) ) ;
AND2    gate17677  (.A(g7195), .B(g1874), .Z(g8939) ) ;
AND2    gate17678  (.A(g7303), .B(g2565), .Z(g8946) ) ;
AND2    gate17679  (.A(g7328), .B(g5615), .Z(g8947) ) ;
AND2    gate17680  (.A(g3650), .B(g1877), .Z(g8972) ) ;
AND2    gate17681  (.A(g7391), .B(g2568), .Z(g8979) ) ;
AND2    gate17682  (.A(g3806), .B(g2571), .Z(g9004) ) ;
AND2    gate17683  (.A(g6486), .B(g565), .Z(g9009) ) ;
AND2    gate17684  (.A(g5438), .B(g7610), .Z(g9026) ) ;
AND2    gate17685  (.A(g6643), .B(g567), .Z(g9033) ) ;
AND2    gate17686  (.A(g6751), .B(g1251), .Z(g9034) ) ;
AND2    gate17687  (.A(g6448), .B(g7616), .Z(g9047) ) ;
AND2    gate17688  (.A(g3338), .B(g489), .Z(g9048) ) ;
AND2    gate17689  (.A(g5473), .B(g7619), .Z(g9049) ) ;
AND2    gate17690  (.A(g6945), .B(g1253), .Z(g9056) ) ;
AND2    gate17691  (.A(g7053), .B(g1945), .Z(g9057) ) ;
AND2    gate17692  (.A(g3306), .B(g7623), .Z(g9061) ) ;
AND2    gate17693  (.A(g5438), .B(g7626), .Z(g9062) ) ;
AND2    gate17694  (.A(g5438), .B(g7629), .Z(g9063) ) ;
AND2    gate17695  (.A(g6713), .B(g7632), .Z(g9064) ) ;
AND2    gate17696  (.A(g3494), .B(g1176), .Z(g9065) ) ;
AND2    gate17697  (.A(g5512), .B(g7635), .Z(g9066) ) ;
AND2    gate17698  (.A(g7195), .B(g1947), .Z(g9073) ) ;
AND2    gate17699  (.A(g7303), .B(g2639), .Z(g9074) ) ;
AND2    gate17700  (.A(g6448), .B(g7643), .Z(g9075) ) ;
AND2    gate17701  (.A(g5438), .B(g7646), .Z(g9076) ) ;
AND2    gate17702  (.A(g6448), .B(g7649), .Z(g9077) ) ;
AND2    gate17703  (.A(g3462), .B(g7652), .Z(g9078) ) ;
AND2    gate17704  (.A(g5473), .B(g7655), .Z(g9079) ) ;
AND2    gate17705  (.A(g5473), .B(g7658), .Z(g9080) ) ;
AND2    gate17706  (.A(g7015), .B(g7661), .Z(g9081) ) ;
AND2    gate17707  (.A(g3650), .B(g1870), .Z(g9082) ) ;
AND2    gate17708  (.A(g5556), .B(g7664), .Z(g9083) ) ;
AND2    gate17709  (.A(g7391), .B(g2641), .Z(g9090) ) ;
AND2    gate17710  (.A(g3306), .B(g7670), .Z(g9091) ) ;
AND2    gate17711  (.A(g6448), .B(g7673), .Z(g9092) ) ;
AND2    gate17712  (.A(g3306), .B(g7676), .Z(g9093) ) ;
AND2    gate17713  (.A(g6713), .B(g7679), .Z(g9094) ) ;
AND2    gate17714  (.A(g5473), .B(g7682), .Z(g9095) ) ;
AND2    gate17715  (.A(g6713), .B(g7685), .Z(g9096) ) ;
AND2    gate17716  (.A(g3618), .B(g7688), .Z(g9097) ) ;
AND2    gate17717  (.A(g5512), .B(g7691), .Z(g9098) ) ;
AND2    gate17718  (.A(g5512), .B(g7694), .Z(g9099) ) ;
AND2    gate17719  (.A(g7265), .B(g7697), .Z(g9100) ) ;
AND2    gate17720  (.A(g3806), .B(g2564), .Z(g9101) ) ;
AND2    gate17721  (.A(g3306), .B(g7703), .Z(g9102) ) ;
AND2    gate17722  (.A(g3462), .B(g7706), .Z(g9103) ) ;
AND2    gate17723  (.A(g6713), .B(g7709), .Z(g9104) ) ;
AND2    gate17724  (.A(g3462), .B(g7712), .Z(g9105) ) ;
AND2    gate17725  (.A(g7015), .B(g7715), .Z(g9106) ) ;
AND2    gate17726  (.A(g5512), .B(g7718), .Z(g9107) ) ;
AND2    gate17727  (.A(g7015), .B(g7721), .Z(g9108) ) ;
AND2    gate17728  (.A(g3774), .B(g7724), .Z(g9109) ) ;
AND2    gate17729  (.A(g5556), .B(g7727), .Z(g9110) ) ;
AND2    gate17730  (.A(g5556), .B(g7730), .Z(g9111) ) ;
AND2    gate17731  (.A(g3462), .B(g7733), .Z(g9112) ) ;
AND2    gate17732  (.A(g3618), .B(g7736), .Z(g9113) ) ;
AND2    gate17733  (.A(g7015), .B(g7739), .Z(g9114) ) ;
AND2    gate17734  (.A(g3618), .B(g7742), .Z(g9115) ) ;
AND2    gate17735  (.A(g7265), .B(g7745), .Z(g9116) ) ;
AND2    gate17736  (.A(g5556), .B(g7748), .Z(g9117) ) ;
AND2    gate17737  (.A(g7265), .B(g7751), .Z(g9118) ) ;
AND2    gate17738  (.A(g5438), .B(g7754), .Z(g9119) ) ;
AND2    gate17739  (.A(g3618), .B(g7757), .Z(g9120) ) ;
AND2    gate17740  (.A(g3774), .B(g7760), .Z(g9121) ) ;
AND2    gate17741  (.A(g7265), .B(g7763), .Z(g9122) ) ;
AND2    gate17742  (.A(g3774), .B(g7766), .Z(g9123) ) ;
AND2    gate17743  (.A(g6448), .B(g7769), .Z(g9124) ) ;
AND2    gate17744  (.A(g5473), .B(g7776), .Z(g9125) ) ;
AND2    gate17745  (.A(g3774), .B(g7779), .Z(g9126) ) ;
AND2    gate17746  (.A(g3306), .B(g7782), .Z(g9127) ) ;
AND2    gate17747  (.A(g6713), .B(g7785), .Z(g9131) ) ;
AND2    gate17748  (.A(g5512), .B(g7792), .Z(g9132) ) ;
AND2    gate17749  (.A(g3462), .B(g7796), .Z(g9133) ) ;
AND2    gate17750  (.A(g7015), .B(g7799), .Z(g9137) ) ;
AND2    gate17751  (.A(g5556), .B(g7806), .Z(g9138) ) ;
AND2    gate17752  (.A(g3618), .B(g7809), .Z(g9139) ) ;
AND2    gate17753  (.A(g7265), .B(g7812), .Z(g9143) ) ;
AND2    gate17754  (.A(g3774), .B(g7823), .Z(g9145) ) ;
AND2    gate17755  (.A(g6232), .B(g7950), .Z(g9241) ) ;
AND2    gate17756  (.A(g6314), .B(g7990), .Z(g9301) ) ;
AND2    gate17757  (.A(g6232), .B(g7993), .Z(g9302) ) ;
AND2    gate17758  (.A(g6369), .B(g8001), .Z(g9319) ) ;
AND2    gate17759  (.A(g3254), .B(g8053), .Z(g9364) ) ;
AND2    gate17760  (.A(g6314), .B(g8056), .Z(g9365) ) ;
AND2    gate17761  (.A(g6232), .B(g8059), .Z(g9366) ) ;
AND2    gate17762  (.A(g6232), .B(g8062), .Z(g9367) ) ;
AND2    gate17763  (.A(g6519), .B(g8065), .Z(g9382) ) ;
AND2    gate17764  (.A(g6369), .B(g8068), .Z(g9383) ) ;
AND2    gate17765  (.A(g6574), .B(g8076), .Z(g9400) ) ;
AND2    gate17766  (.A(g3254), .B(g8123), .Z(g9438) ) ;
AND2    gate17767  (.A(g6314), .B(g8126), .Z(g9439) ) ;
AND2    gate17768  (.A(g6232), .B(g8129), .Z(g9440) ) ;
AND2    gate17769  (.A(g6314), .B(g8132), .Z(g9441) ) ;
AND2    gate17770  (.A(g6232), .B(g8135), .Z(g9442) ) ;
AND2    gate17771  (.A(g3410), .B(g8138), .Z(g9461) ) ;
AND2    gate17772  (.A(g6519), .B(g8141), .Z(g9462) ) ;
AND2    gate17773  (.A(g6369), .B(g8144), .Z(g9463) ) ;
AND2    gate17774  (.A(g6369), .B(g8147), .Z(g9464) ) ;
AND2    gate17775  (.A(g6783), .B(g8150), .Z(g9479) ) ;
AND2    gate17776  (.A(g6574), .B(g8153), .Z(g9480) ) ;
AND2    gate17777  (.A(g6838), .B(g8161), .Z(g9497) ) ;
AND2    gate17778  (.A(g3254), .B(g8191), .Z(g9518) ) ;
AND2    gate17779  (.A(g6314), .B(g8194), .Z(g9519) ) ;
AND2    gate17780  (.A(g6232), .B(g8197), .Z(g9520) ) ;
AND2    gate17781  (.A(g3254), .B(g8200), .Z(g9521) ) ;
AND2    gate17782  (.A(g6314), .B(g8203), .Z(g9522) ) ;
AND2    gate17783  (.A(g6232), .B(g8206), .Z(g9523) ) ;
AND3    gate17784  (.A(g7772), .B(g6135), .C(g538), .Z(g9534) ) ;
AND2    gate17785  (.A(g3410), .B(g8209), .Z(g9580) ) ;
AND2    gate17786  (.A(g6519), .B(g8212), .Z(g9581) ) ;
AND2    gate17787  (.A(g6369), .B(g8215), .Z(g9582) ) ;
AND2    gate17788  (.A(g6519), .B(g8218), .Z(g9583) ) ;
AND2    gate17789  (.A(g6369), .B(g8221), .Z(g9584) ) ;
AND2    gate17790  (.A(g3566), .B(g8224), .Z(g9603) ) ;
AND2    gate17791  (.A(g6783), .B(g8227), .Z(g9604) ) ;
AND2    gate17792  (.A(g6574), .B(g8230), .Z(g9605) ) ;
AND2    gate17793  (.A(g6574), .B(g8233), .Z(g9606) ) ;
AND2    gate17794  (.A(g7085), .B(g8236), .Z(g9621) ) ;
AND2    gate17795  (.A(g6838), .B(g8239), .Z(g9622) ) ;
AND2    gate17796  (.A(g3254), .B(g3922), .Z(g9630) ) ;
AND2    gate17797  (.A(g6314), .B(g3925), .Z(g9631) ) ;
AND2    gate17798  (.A(g6232), .B(g3928), .Z(g9632) ) ;
AND2    gate17799  (.A(g3254), .B(g3931), .Z(g9633) ) ;
AND2    gate17800  (.A(g6314), .B(g3934), .Z(g9634) ) ;
AND2    gate17801  (.A(g6232), .B(g3937), .Z(g9635) ) ;
AND4    gate17802  (.A(g5856), .B(g4338), .C(g4339), .D(g5141), .Z(II16735) ) ;
AND4    gate17803  (.A(g5713), .B(g5958), .C(g4735), .D(g4736), .Z(II16736) ) ;
AND2    gate17804  (.A(II16735), .B(II16736), .Z(g9636) ) ;
AND2    gate17805  (.A(g5438), .B(g408), .Z(g9639) ) ;
AND2    gate17806  (.A(g6678), .B(g3942), .Z(g9647) ) ;
AND2    gate17807  (.A(g6678), .B(g3945), .Z(g9648) ) ;
AND2    gate17808  (.A(g3410), .B(g3948), .Z(g9660) ) ;
AND2    gate17809  (.A(g6519), .B(g3951), .Z(g9661) ) ;
AND2    gate17810  (.A(g6369), .B(g3954), .Z(g9662) ) ;
AND2    gate17811  (.A(g3410), .B(g3957), .Z(g9663) ) ;
AND2    gate17812  (.A(g6519), .B(g3960), .Z(g9664) ) ;
AND2    gate17813  (.A(g6369), .B(g3963), .Z(g9665) ) ;
AND3    gate17814  (.A(g7788), .B(g6145), .C(g1224), .Z(g9676) ) ;
AND2    gate17815  (.A(g3566), .B(g3966), .Z(g9722) ) ;
AND2    gate17816  (.A(g6783), .B(g3969), .Z(g9723) ) ;
AND2    gate17817  (.A(g6574), .B(g3972), .Z(g9724) ) ;
AND2    gate17818  (.A(g6783), .B(g3975), .Z(g9725) ) ;
AND2    gate17819  (.A(g6574), .B(g3978), .Z(g9726) ) ;
AND2    gate17820  (.A(g3722), .B(g3981), .Z(g9745) ) ;
AND2    gate17821  (.A(g7085), .B(g3984), .Z(g9746) ) ;
AND2    gate17822  (.A(g6838), .B(g3987), .Z(g9747) ) ;
AND2    gate17823  (.A(g6838), .B(g3990), .Z(g9748) ) ;
AND2    gate17824  (.A(g3254), .B(g4000), .Z(g9759) ) ;
AND2    gate17825  (.A(g6314), .B(g4003), .Z(g9760) ) ;
AND2    gate17826  (.A(g6232), .B(g4006), .Z(g9761) ) ;
AND2    gate17827  (.A(g3254), .B(g4009), .Z(g9762) ) ;
AND2    gate17828  (.A(g6314), .B(g4012), .Z(g9763) ) ;
AND2    gate17829  (.A(g6448), .B(g411), .Z(g9764) ) ;
AND2    gate17830  (.A(g5438), .B(g417), .Z(g9765) ) ;
AND2    gate17831  (.A(g5438), .B(g4017), .Z(g9766) ) ;
AND2    gate17832  (.A(g6912), .B(g4020), .Z(g9773) ) ;
AND2    gate17833  (.A(g6678), .B(g4023), .Z(g9774) ) ;
AND2    gate17834  (.A(g6912), .B(g4026), .Z(g9775) ) ;
AND2    gate17835  (.A(g3410), .B(g4029), .Z(g9776) ) ;
AND2    gate17836  (.A(g6519), .B(g4032), .Z(g9777) ) ;
AND2    gate17837  (.A(g6369), .B(g4035), .Z(g9778) ) ;
AND2    gate17838  (.A(g3410), .B(g4038), .Z(g9779) ) ;
AND2    gate17839  (.A(g6519), .B(g4041), .Z(g9780) ) ;
AND2    gate17840  (.A(g6369), .B(g4044), .Z(g9781) ) ;
AND4    gate17841  (.A(g5903), .B(g4507), .C(g4508), .D(g5234), .Z(II16826) ) ;
AND4    gate17842  (.A(g5771), .B(g5987), .C(g4911), .D(g4912), .Z(II16827) ) ;
AND2    gate17843  (.A(II16826), .B(II16827), .Z(g9782) ) ;
AND2    gate17844  (.A(g5473), .B(g1095), .Z(g9785) ) ;
AND2    gate17845  (.A(g6980), .B(g4049), .Z(g9793) ) ;
AND2    gate17846  (.A(g6980), .B(g4052), .Z(g9794) ) ;
AND2    gate17847  (.A(g3566), .B(g4055), .Z(g9806) ) ;
AND2    gate17848  (.A(g6783), .B(g4058), .Z(g9807) ) ;
AND2    gate17849  (.A(g6574), .B(g4061), .Z(g9808) ) ;
AND2    gate17850  (.A(g3566), .B(g4064), .Z(g9809) ) ;
AND2    gate17851  (.A(g6783), .B(g4067), .Z(g9810) ) ;
AND2    gate17852  (.A(g6574), .B(g4070), .Z(g9811) ) ;
AND3    gate17853  (.A(g7802), .B(g6166), .C(g1918), .Z(g9822) ) ;
AND2    gate17854  (.A(g3722), .B(g4073), .Z(g9868) ) ;
AND2    gate17855  (.A(g7085), .B(g4076), .Z(g9869) ) ;
AND2    gate17856  (.A(g6838), .B(g4079), .Z(g9870) ) ;
AND2    gate17857  (.A(g7085), .B(g4082), .Z(g9871) ) ;
AND2    gate17858  (.A(g6838), .B(g4085), .Z(g9872) ) ;
AND2    gate17859  (.A(g6232), .B(g4095), .Z(g9887) ) ;
AND2    gate17860  (.A(g3254), .B(g4098), .Z(g9888) ) ;
AND2    gate17861  (.A(g6314), .B(g4101), .Z(g9889) ) ;
AND2    gate17862  (.A(g6232), .B(g4104), .Z(g9890) ) ;
AND2    gate17863  (.A(g3254), .B(g4107), .Z(g9891) ) ;
AND2    gate17864  (.A(g3306), .B(g414), .Z(g9892) ) ;
AND2    gate17865  (.A(g6448), .B(g420), .Z(g9893) ) ;
AND2    gate17866  (.A(g6448), .B(g4112), .Z(g9894) ) ;
AND2    gate17867  (.A(g3366), .B(g4115), .Z(g9901) ) ;
AND2    gate17868  (.A(g6912), .B(g4118), .Z(g9902) ) ;
AND2    gate17869  (.A(g6678), .B(g4121), .Z(g9903) ) ;
AND2    gate17870  (.A(g3366), .B(g4124), .Z(g9904) ) ;
AND2    gate17871  (.A(g3410), .B(g4127), .Z(g9905) ) ;
AND2    gate17872  (.A(g6519), .B(g4130), .Z(g9906) ) ;
AND2    gate17873  (.A(g6369), .B(g4133), .Z(g9907) ) ;
AND2    gate17874  (.A(g3410), .B(g4136), .Z(g9908) ) ;
AND2    gate17875  (.A(g6519), .B(g4139), .Z(g9909) ) ;
AND2    gate17876  (.A(g6713), .B(g1098), .Z(g9910) ) ;
AND2    gate17877  (.A(g5473), .B(g1104), .Z(g9911) ) ;
AND2    gate17878  (.A(g5473), .B(g4144), .Z(g9912) ) ;
AND2    gate17879  (.A(g7162), .B(g4147), .Z(g9919) ) ;
AND2    gate17880  (.A(g6980), .B(g4150), .Z(g9920) ) ;
AND2    gate17881  (.A(g7162), .B(g4153), .Z(g9921) ) ;
AND2    gate17882  (.A(g3566), .B(g4156), .Z(g9922) ) ;
AND2    gate17883  (.A(g6783), .B(g4159), .Z(g9923) ) ;
AND2    gate17884  (.A(g6574), .B(g4162), .Z(g9924) ) ;
AND2    gate17885  (.A(g3566), .B(g4165), .Z(g9925) ) ;
AND2    gate17886  (.A(g6783), .B(g4168), .Z(g9926) ) ;
AND2    gate17887  (.A(g6574), .B(g4171), .Z(g9927) ) ;
AND4    gate17888  (.A(g5942), .B(g4683), .C(g4684), .D(g5297), .Z(II16930) ) ;
AND4    gate17889  (.A(g5830), .B(g6024), .C(g5070), .D(g5071), .Z(II16931) ) ;
AND2    gate17890  (.A(II16930), .B(II16931), .Z(g9928) ) ;
AND2    gate17891  (.A(g5512), .B(g1789), .Z(g9931) ) ;
AND2    gate17892  (.A(g7230), .B(g4176), .Z(g9939) ) ;
AND2    gate17893  (.A(g7230), .B(g4179), .Z(g9940) ) ;
AND2    gate17894  (.A(g3722), .B(g4182), .Z(g9952) ) ;
AND2    gate17895  (.A(g7085), .B(g4185), .Z(g9953) ) ;
AND2    gate17896  (.A(g6838), .B(g4188), .Z(g9954) ) ;
AND2    gate17897  (.A(g3722), .B(g4191), .Z(g9955) ) ;
AND2    gate17898  (.A(g7085), .B(g4194), .Z(g9956) ) ;
AND2    gate17899  (.A(g6838), .B(g4197), .Z(g9957) ) ;
AND3    gate17900  (.A(g7815), .B(g6193), .C(g2612), .Z(g9968) ) ;
AND2    gate17901  (.A(g6314), .B(g4205), .Z(g10007) ) ;
AND2    gate17902  (.A(g6232), .B(g4208), .Z(g10008) ) ;
AND2    gate17903  (.A(g3254), .B(g4211), .Z(g10009) ) ;
AND2    gate17904  (.A(g6314), .B(g4214), .Z(g10010) ) ;
AND2    gate17905  (.A(g5438), .B(g4217), .Z(g10011) ) ;
AND2    gate17906  (.A(g3306), .B(g423), .Z(g10012) ) ;
AND2    gate17907  (.A(g3306), .B(g4221), .Z(g10013) ) ;
AND2    gate17908  (.A(g5438), .B(g429), .Z(g10014) ) ;
AND2    gate17909  (.A(g3398), .B(g6912), .Z(g10024) ) ;
AND2    gate17910  (.A(g3366), .B(g4225), .Z(g10035) ) ;
AND2    gate17911  (.A(g6912), .B(g4228), .Z(g10036) ) ;
AND2    gate17912  (.A(g6678), .B(g4231), .Z(g10037) ) ;
AND2    gate17913  (.A(g6369), .B(g4234), .Z(g10041) ) ;
AND2    gate17914  (.A(g3410), .B(g4237), .Z(g10042) ) ;
AND2    gate17915  (.A(g6519), .B(g4240), .Z(g10043) ) ;
AND2    gate17916  (.A(g6369), .B(g4243), .Z(g10044) ) ;
AND2    gate17917  (.A(g3410), .B(g4246), .Z(g10045) ) ;
AND2    gate17918  (.A(g3462), .B(g1101), .Z(g10046) ) ;
AND2    gate17919  (.A(g6713), .B(g1107), .Z(g10047) ) ;
AND2    gate17920  (.A(g6713), .B(g4251), .Z(g10048) ) ;
AND2    gate17921  (.A(g3522), .B(g4254), .Z(g10055) ) ;
AND2    gate17922  (.A(g7162), .B(g4257), .Z(g10056) ) ;
AND2    gate17923  (.A(g6980), .B(g4260), .Z(g10057) ) ;
AND2    gate17924  (.A(g3522), .B(g4263), .Z(g10058) ) ;
AND2    gate17925  (.A(g3566), .B(g4266), .Z(g10059) ) ;
AND2    gate17926  (.A(g6783), .B(g4269), .Z(g10060) ) ;
AND2    gate17927  (.A(g6574), .B(g4272), .Z(g10061) ) ;
AND2    gate17928  (.A(g3566), .B(g4275), .Z(g10062) ) ;
AND2    gate17929  (.A(g6783), .B(g4278), .Z(g10063) ) ;
AND2    gate17930  (.A(g7015), .B(g1792), .Z(g10064) ) ;
AND2    gate17931  (.A(g5512), .B(g1798), .Z(g10065) ) ;
AND2    gate17932  (.A(g5512), .B(g4283), .Z(g10066) ) ;
AND2    gate17933  (.A(g7358), .B(g4286), .Z(g10073) ) ;
AND2    gate17934  (.A(g7230), .B(g4289), .Z(g10074) ) ;
AND2    gate17935  (.A(g7358), .B(g4292), .Z(g10075) ) ;
AND2    gate17936  (.A(g3722), .B(g4295), .Z(g10076) ) ;
AND2    gate17937  (.A(g7085), .B(g4298), .Z(g10077) ) ;
AND2    gate17938  (.A(g6838), .B(g4301), .Z(g10078) ) ;
AND2    gate17939  (.A(g3722), .B(g4304), .Z(g10079) ) ;
AND2    gate17940  (.A(g7085), .B(g4307), .Z(g10080) ) ;
AND2    gate17941  (.A(g6838), .B(g4310), .Z(g10081) ) ;
AND4    gate17942  (.A(g5976), .B(g4860), .C(g4861), .D(g5334), .Z(II17042) ) ;
AND4    gate17943  (.A(g5886), .B(g6040), .C(g5199), .D(g5200), .Z(II17043) ) ;
AND2    gate17944  (.A(II17042), .B(II17043), .Z(g10082) ) ;
AND2    gate17945  (.A(g5556), .B(g2483), .Z(g10085) ) ;
AND2    gate17946  (.A(g7426), .B(g4315), .Z(g10093) ) ;
AND2    gate17947  (.A(g7426), .B(g4318), .Z(g10094) ) ;
AND2    gate17948  (.A(g3254), .B(g4329), .Z(g10101) ) ;
AND2    gate17949  (.A(g6314), .B(g4332), .Z(g10102) ) ;
AND2    gate17950  (.A(g3254), .B(g4335), .Z(g10103) ) ;
AND2    gate17951  (.A(g6448), .B(g4340), .Z(g10104) ) ;
AND2    gate17952  (.A(g5438), .B(g4343), .Z(g10105) ) ;
AND2    gate17953  (.A(g6448), .B(g432), .Z(g10106) ) ;
AND2    gate17954  (.A(g5438), .B(g438), .Z(g10107) ) ;
AND2    gate17955  (.A(g6486), .B(g569), .Z(g10108) ) ;
AND2    gate17956  (.A(g3366), .B(g4348), .Z(g10112) ) ;
AND2    gate17957  (.A(g6912), .B(g4351), .Z(g10113) ) ;
AND2    gate17958  (.A(g6678), .B(g4354), .Z(g10114) ) ;
AND2    gate17959  (.A(g6678), .B(g4357), .Z(g10115) ) ;
AND2    gate17960  (.A(g6519), .B(g4360), .Z(g10116) ) ;
AND2    gate17961  (.A(g6369), .B(g4363), .Z(g10117) ) ;
AND2    gate17962  (.A(g3410), .B(g4366), .Z(g10118) ) ;
AND2    gate17963  (.A(g6519), .B(g4369), .Z(g10119) ) ;
AND2    gate17964  (.A(g5473), .B(g4372), .Z(g10120) ) ;
AND2    gate17965  (.A(g3462), .B(g1110), .Z(g10121) ) ;
AND2    gate17966  (.A(g3462), .B(g4376), .Z(g10122) ) ;
AND2    gate17967  (.A(g5473), .B(g1116), .Z(g10123) ) ;
AND2    gate17968  (.A(g3554), .B(g7162), .Z(g10133) ) ;
AND2    gate17969  (.A(g3522), .B(g4380), .Z(g10144) ) ;
AND2    gate17970  (.A(g7162), .B(g4383), .Z(g10145) ) ;
AND2    gate17971  (.A(g6980), .B(g4386), .Z(g10146) ) ;
AND2    gate17972  (.A(g6574), .B(g4389), .Z(g10150) ) ;
AND2    gate17973  (.A(g3566), .B(g4392), .Z(g10151) ) ;
AND2    gate17974  (.A(g6783), .B(g4395), .Z(g10152) ) ;
AND2    gate17975  (.A(g6574), .B(g4398), .Z(g10153) ) ;
AND2    gate17976  (.A(g3566), .B(g4401), .Z(g10154) ) ;
AND2    gate17977  (.A(g3618), .B(g1795), .Z(g10155) ) ;
AND2    gate17978  (.A(g7015), .B(g1801), .Z(g10156) ) ;
AND2    gate17979  (.A(g7015), .B(g4406), .Z(g10157) ) ;
AND2    gate17980  (.A(g3678), .B(g4409), .Z(g10164) ) ;
AND2    gate17981  (.A(g7358), .B(g4412), .Z(g10165) ) ;
AND2    gate17982  (.A(g7230), .B(g4415), .Z(g10166) ) ;
AND2    gate17983  (.A(g3678), .B(g4418), .Z(g10167) ) ;
AND2    gate17984  (.A(g3722), .B(g4421), .Z(g10168) ) ;
AND2    gate17985  (.A(g7085), .B(g4424), .Z(g10169) ) ;
AND2    gate17986  (.A(g6838), .B(g4427), .Z(g10170) ) ;
AND2    gate17987  (.A(g3722), .B(g4430), .Z(g10171) ) ;
AND2    gate17988  (.A(g7085), .B(g4433), .Z(g10172) ) ;
AND2    gate17989  (.A(g7265), .B(g2486), .Z(g10173) ) ;
AND2    gate17990  (.A(g5556), .B(g2492), .Z(g10174) ) ;
AND2    gate17991  (.A(g5556), .B(g4438), .Z(g10175) ) ;
AND2    gate17992  (.A(g7488), .B(g4441), .Z(g10182) ) ;
AND2    gate17993  (.A(g7426), .B(g4444), .Z(g10183) ) ;
AND2    gate17994  (.A(g7488), .B(g4447), .Z(g10184) ) ;
AND4    gate17995  (.A(g6898), .B(g2998), .C(g6901), .D(g3002), .Z(II17156) ) ;
AND4    gate17996  (.A(g3013), .B(g7466), .C(g3024), .D(II17156), .Z(g10186) ) ;
AND2    gate17997  (.A(g3254), .B(g4453), .Z(g10192) ) ;
AND2    gate17998  (.A(g3306), .B(g4465), .Z(g10193) ) ;
AND2    gate17999  (.A(g6448), .B(g4468), .Z(g10194) ) ;
AND2    gate18000  (.A(g5438), .B(g4471), .Z(g10195) ) ;
AND2    gate18001  (.A(g3306), .B(g435), .Z(g10196) ) ;
AND2    gate18002  (.A(g6448), .B(g441), .Z(g10197) ) ;
AND2    gate18003  (.A(g6643), .B(g571), .Z(g10198) ) ;
AND2    gate18004  (.A(g6486), .B(g4476), .Z(g10199) ) ;
AND2    gate18005  (.A(g6486), .B(g587), .Z(g10200) ) ;
AND2    gate18006  (.A(g3366), .B(g4480), .Z(g10201) ) ;
AND2    gate18007  (.A(g6912), .B(g4483), .Z(g10202) ) ;
AND2    gate18008  (.A(g6678), .B(g4486), .Z(g10203) ) ;
AND2    gate18009  (.A(g6912), .B(g4489), .Z(g10204) ) ;
AND2    gate18010  (.A(g6678), .B(g4492), .Z(g10205) ) ;
AND2    gate18011  (.A(g3410), .B(g4498), .Z(g10206) ) ;
AND2    gate18012  (.A(g6519), .B(g4501), .Z(g10207) ) ;
AND2    gate18013  (.A(g3410), .B(g4504), .Z(g10208) ) ;
AND2    gate18014  (.A(g6713), .B(g4509), .Z(g10209) ) ;
AND2    gate18015  (.A(g5473), .B(g4512), .Z(g10210) ) ;
AND2    gate18016  (.A(g6713), .B(g1119), .Z(g10211) ) ;
AND2    gate18017  (.A(g5473), .B(g1125), .Z(g10212) ) ;
AND2    gate18018  (.A(g6751), .B(g1255), .Z(g10213) ) ;
AND2    gate18019  (.A(g3522), .B(g4517), .Z(g10217) ) ;
AND2    gate18020  (.A(g7162), .B(g4520), .Z(g10218) ) ;
AND2    gate18021  (.A(g6980), .B(g4523), .Z(g10219) ) ;
AND2    gate18022  (.A(g6980), .B(g4526), .Z(g10220) ) ;
AND2    gate18023  (.A(g6783), .B(g4529), .Z(g10221) ) ;
AND2    gate18024  (.A(g6574), .B(g4532), .Z(g10222) ) ;
AND2    gate18025  (.A(g3566), .B(g4535), .Z(g10223) ) ;
AND2    gate18026  (.A(g6783), .B(g4538), .Z(g10224) ) ;
AND2    gate18027  (.A(g5512), .B(g4541), .Z(g10225) ) ;
AND2    gate18028  (.A(g3618), .B(g1804), .Z(g10226) ) ;
AND2    gate18029  (.A(g3618), .B(g4545), .Z(g10227) ) ;
AND2    gate18030  (.A(g5512), .B(g1810), .Z(g10228) ) ;
AND2    gate18031  (.A(g3710), .B(g7358), .Z(g10238) ) ;
AND2    gate18032  (.A(g3678), .B(g4549), .Z(g10249) ) ;
AND2    gate18033  (.A(g7358), .B(g4552), .Z(g10250) ) ;
AND2    gate18034  (.A(g7230), .B(g4555), .Z(g10251) ) ;
AND2    gate18035  (.A(g6838), .B(g4558), .Z(g10255) ) ;
AND2    gate18036  (.A(g3722), .B(g4561), .Z(g10256) ) ;
AND2    gate18037  (.A(g7085), .B(g4564), .Z(g10257) ) ;
AND2    gate18038  (.A(g6838), .B(g4567), .Z(g10258) ) ;
AND2    gate18039  (.A(g3722), .B(g4570), .Z(g10259) ) ;
AND2    gate18040  (.A(g3774), .B(g2489), .Z(g10260) ) ;
AND2    gate18041  (.A(g7265), .B(g2495), .Z(g10261) ) ;
AND2    gate18042  (.A(g7265), .B(g4575), .Z(g10262) ) ;
AND2    gate18043  (.A(g3834), .B(g4578), .Z(g10269) ) ;
AND2    gate18044  (.A(g7488), .B(g4581), .Z(g10270) ) ;
AND2    gate18045  (.A(g7426), .B(g4584), .Z(g10271) ) ;
AND2    gate18046  (.A(g3834), .B(g4587), .Z(g10272) ) ;
AND2    gate18047  (.A(g3306), .B(g4592), .Z(g10279) ) ;
AND2    gate18048  (.A(g6448), .B(g4595), .Z(g10280) ) ;
AND2    gate18049  (.A(g5438), .B(g4598), .Z(g10281) ) ;
AND2    gate18050  (.A(g3306), .B(g444), .Z(g10282) ) ;
AND2    gate18051  (.A(g3338), .B(g573), .Z(g10283) ) ;
AND2    gate18052  (.A(g6643), .B(g4603), .Z(g10284) ) ;
AND2    gate18053  (.A(g6486), .B(g4606), .Z(g10285) ) ;
AND2    gate18054  (.A(g6643), .B(g590), .Z(g10286) ) ;
AND2    gate18055  (.A(g6486), .B(g596), .Z(g10287) ) ;
AND2    gate18056  (.A(g3366), .B(g4611), .Z(g10288) ) ;
AND2    gate18057  (.A(g6912), .B(g4614), .Z(g10289) ) ;
AND2    gate18058  (.A(g6678), .B(g4617), .Z(g10290) ) ;
AND2    gate18059  (.A(g3366), .B(g4620), .Z(g10291) ) ;
AND2    gate18060  (.A(g6912), .B(g4623), .Z(g10292) ) ;
AND2    gate18061  (.A(g6678), .B(g4626), .Z(g10293) ) ;
AND2    gate18062  (.A(g3410), .B(g4629), .Z(g10294) ) ;
AND2    gate18063  (.A(g3462), .B(g4641), .Z(g10295) ) ;
AND2    gate18064  (.A(g6713), .B(g4644), .Z(g10296) ) ;
AND2    gate18065  (.A(g5473), .B(g4647), .Z(g10297) ) ;
AND2    gate18066  (.A(g3462), .B(g1122), .Z(g10298) ) ;
AND2    gate18067  (.A(g6713), .B(g1128), .Z(g10299) ) ;
AND2    gate18068  (.A(g6945), .B(g1257), .Z(g10300) ) ;
AND2    gate18069  (.A(g6751), .B(g4652), .Z(g10301) ) ;
AND2    gate18070  (.A(g6751), .B(g1273), .Z(g10302) ) ;
AND2    gate18071  (.A(g3522), .B(g4656), .Z(g10303) ) ;
AND2    gate18072  (.A(g7162), .B(g4659), .Z(g10304) ) ;
AND2    gate18073  (.A(g6980), .B(g4662), .Z(g10305) ) ;
AND2    gate18074  (.A(g7162), .B(g4665), .Z(g10306) ) ;
AND2    gate18075  (.A(g6980), .B(g4668), .Z(g10307) ) ;
AND2    gate18076  (.A(g3566), .B(g4674), .Z(g10308) ) ;
AND2    gate18077  (.A(g6783), .B(g4677), .Z(g10309) ) ;
AND2    gate18078  (.A(g3566), .B(g4680), .Z(g10310) ) ;
AND2    gate18079  (.A(g7015), .B(g4685), .Z(g10311) ) ;
AND2    gate18080  (.A(g5512), .B(g4688), .Z(g10312) ) ;
AND2    gate18081  (.A(g7015), .B(g1813), .Z(g10313) ) ;
AND2    gate18082  (.A(g5512), .B(g1819), .Z(g10314) ) ;
AND2    gate18083  (.A(g7053), .B(g1949), .Z(g10315) ) ;
AND2    gate18084  (.A(g3678), .B(g4693), .Z(g10319) ) ;
AND2    gate18085  (.A(g7358), .B(g4696), .Z(g10320) ) ;
AND2    gate18086  (.A(g7230), .B(g4699), .Z(g10321) ) ;
AND2    gate18087  (.A(g7230), .B(g4702), .Z(g10322) ) ;
AND2    gate18088  (.A(g7085), .B(g4705), .Z(g10323) ) ;
AND2    gate18089  (.A(g6838), .B(g4708), .Z(g10324) ) ;
AND2    gate18090  (.A(g3722), .B(g4711), .Z(g10325) ) ;
AND2    gate18091  (.A(g7085), .B(g4714), .Z(g10326) ) ;
AND2    gate18092  (.A(g5556), .B(g4717), .Z(g10327) ) ;
AND2    gate18093  (.A(g3774), .B(g2498), .Z(g10328) ) ;
AND2    gate18094  (.A(g3774), .B(g4721), .Z(g10329) ) ;
AND2    gate18095  (.A(g5556), .B(g2504), .Z(g10330) ) ;
AND2    gate18096  (.A(g3866), .B(g7488), .Z(g10340) ) ;
AND2    gate18097  (.A(g3834), .B(g4725), .Z(g10351) ) ;
AND2    gate18098  (.A(g7488), .B(g4728), .Z(g10352) ) ;
AND2    gate18099  (.A(g7426), .B(g4731), .Z(g10353) ) ;
AND2    gate18100  (.A(g3306), .B(g4737), .Z(g10360) ) ;
AND2    gate18101  (.A(g6448), .B(g4740), .Z(g10361) ) ;
AND2    gate18102  (.A(g3338), .B(g4743), .Z(g10362) ) ;
AND2    gate18103  (.A(g6643), .B(g4746), .Z(g10363) ) ;
AND2    gate18104  (.A(g6486), .B(g4749), .Z(g10364) ) ;
AND2    gate18105  (.A(g3338), .B(g593), .Z(g10365) ) ;
AND2    gate18106  (.A(g6643), .B(g599), .Z(g10366) ) ;
AND2    gate18107  (.A(g3366), .B(g4754), .Z(g10367) ) ;
AND2    gate18108  (.A(g6912), .B(g4757), .Z(g10368) ) ;
AND2    gate18109  (.A(g6678), .B(g4760), .Z(g10369) ) ;
AND2    gate18110  (.A(g3366), .B(g4763), .Z(g10370) ) ;
AND2    gate18111  (.A(g6912), .B(g4766), .Z(g10371) ) ;
AND2    gate18112  (.A(g3462), .B(g4769), .Z(g10372) ) ;
AND2    gate18113  (.A(g6713), .B(g4772), .Z(g10373) ) ;
AND2    gate18114  (.A(g5473), .B(g4775), .Z(g10374) ) ;
AND2    gate18115  (.A(g3462), .B(g1131), .Z(g10375) ) ;
AND2    gate18116  (.A(g3494), .B(g1259), .Z(g10376) ) ;
AND2    gate18117  (.A(g6945), .B(g4780), .Z(g10377) ) ;
AND2    gate18118  (.A(g6751), .B(g4783), .Z(g10378) ) ;
AND2    gate18119  (.A(g6945), .B(g1276), .Z(g10379) ) ;
AND2    gate18120  (.A(g6751), .B(g1282), .Z(g10380) ) ;
AND2    gate18121  (.A(g3522), .B(g4788), .Z(g10381) ) ;
AND2    gate18122  (.A(g7162), .B(g4791), .Z(g10382) ) ;
AND2    gate18123  (.A(g6980), .B(g4794), .Z(g10383) ) ;
AND2    gate18124  (.A(g3522), .B(g4797), .Z(g10384) ) ;
AND2    gate18125  (.A(g7162), .B(g4800), .Z(g10385) ) ;
AND2    gate18126  (.A(g6980), .B(g4803), .Z(g10386) ) ;
AND2    gate18127  (.A(g3566), .B(g4806), .Z(g10387) ) ;
AND2    gate18128  (.A(g3618), .B(g4818), .Z(g10388) ) ;
AND2    gate18129  (.A(g7015), .B(g4821), .Z(g10389) ) ;
AND2    gate18130  (.A(g5512), .B(g4824), .Z(g10390) ) ;
AND2    gate18131  (.A(g3618), .B(g1816), .Z(g10391) ) ;
AND2    gate18132  (.A(g7015), .B(g1822), .Z(g10392) ) ;
AND2    gate18133  (.A(g7195), .B(g1951), .Z(g10393) ) ;
AND2    gate18134  (.A(g7053), .B(g4829), .Z(g10394) ) ;
AND2    gate18135  (.A(g7053), .B(g1967), .Z(g10395) ) ;
AND2    gate18136  (.A(g3678), .B(g4833), .Z(g10396) ) ;
AND2    gate18137  (.A(g7358), .B(g4836), .Z(g10397) ) ;
AND2    gate18138  (.A(g7230), .B(g4839), .Z(g10398) ) ;
AND2    gate18139  (.A(g7358), .B(g4842), .Z(g10399) ) ;
AND2    gate18140  (.A(g7230), .B(g4845), .Z(g10400) ) ;
AND2    gate18141  (.A(g3722), .B(g4851), .Z(g10401) ) ;
AND2    gate18142  (.A(g7085), .B(g4854), .Z(g10402) ) ;
AND2    gate18143  (.A(g3722), .B(g4857), .Z(g10403) ) ;
AND2    gate18144  (.A(g7265), .B(g4862), .Z(g10404) ) ;
AND2    gate18145  (.A(g5556), .B(g4865), .Z(g10405) ) ;
AND2    gate18146  (.A(g7265), .B(g2507), .Z(g10406) ) ;
AND2    gate18147  (.A(g5556), .B(g2513), .Z(g10407) ) ;
AND2    gate18148  (.A(g7303), .B(g2643), .Z(g10408) ) ;
AND2    gate18149  (.A(g3834), .B(g4870), .Z(g10412) ) ;
AND2    gate18150  (.A(g7488), .B(g4873), .Z(g10413) ) ;
AND2    gate18151  (.A(g7426), .B(g4876), .Z(g10414) ) ;
AND2    gate18152  (.A(g7426), .B(g4879), .Z(g10415) ) ;
AND2    gate18153  (.A(g3306), .B(g4882), .Z(g10422) ) ;
AND2    gate18154  (.A(g5438), .B(g4885), .Z(g10423) ) ;
AND2    gate18155  (.A(g3338), .B(g4888), .Z(g10430) ) ;
AND2    gate18156  (.A(g6643), .B(g4891), .Z(g10431) ) ;
AND2    gate18157  (.A(g6486), .B(g4894), .Z(g10432) ) ;
AND2    gate18158  (.A(g3338), .B(g602), .Z(g10433) ) ;
AND2    gate18159  (.A(g6486), .B(g605), .Z(g10434) ) ;
AND2    gate18160  (.A(g3366), .B(g4899), .Z(g10435) ) ;
AND2    gate18161  (.A(g6912), .B(g4902), .Z(g10436) ) ;
AND2    gate18162  (.A(g6678), .B(g4905), .Z(g10437) ) ;
AND2    gate18163  (.A(g3366), .B(g4908), .Z(g10438) ) ;
AND2    gate18164  (.A(g3462), .B(g4913), .Z(g10439) ) ;
AND2    gate18165  (.A(g6713), .B(g4916), .Z(g10440) ) ;
AND2    gate18166  (.A(g3494), .B(g4919), .Z(g10441) ) ;
AND2    gate18167  (.A(g6945), .B(g4922), .Z(g10442) ) ;
AND2    gate18168  (.A(g6751), .B(g4925), .Z(g10443) ) ;
AND2    gate18169  (.A(g3494), .B(g1279), .Z(g10444) ) ;
AND2    gate18170  (.A(g6945), .B(g1285), .Z(g10445) ) ;
AND2    gate18171  (.A(g3522), .B(g4930), .Z(g10446) ) ;
AND2    gate18172  (.A(g7162), .B(g4933), .Z(g10447) ) ;
AND2    gate18173  (.A(g6980), .B(g4936), .Z(g10448) ) ;
AND2    gate18174  (.A(g3522), .B(g4939), .Z(g10449) ) ;
AND2    gate18175  (.A(g7162), .B(g4942), .Z(g10450) ) ;
AND2    gate18176  (.A(g3618), .B(g4945), .Z(g10451) ) ;
AND2    gate18177  (.A(g7015), .B(g4948), .Z(g10452) ) ;
AND2    gate18178  (.A(g5512), .B(g4951), .Z(g10453) ) ;
AND2    gate18179  (.A(g3618), .B(g1825), .Z(g10454) ) ;
AND2    gate18180  (.A(g3650), .B(g1953), .Z(g10455) ) ;
AND2    gate18181  (.A(g7195), .B(g4956), .Z(g10456) ) ;
AND2    gate18182  (.A(g7053), .B(g4959), .Z(g10457) ) ;
AND2    gate18183  (.A(g7195), .B(g1970), .Z(g10458) ) ;
AND2    gate18184  (.A(g7053), .B(g1976), .Z(g10459) ) ;
AND2    gate18185  (.A(g3678), .B(g4964), .Z(g10460) ) ;
AND2    gate18186  (.A(g7358), .B(g4967), .Z(g10461) ) ;
AND2    gate18187  (.A(g7230), .B(g4970), .Z(g10462) ) ;
AND2    gate18188  (.A(g3678), .B(g4973), .Z(g10463) ) ;
AND2    gate18189  (.A(g7358), .B(g4976), .Z(g10464) ) ;
AND2    gate18190  (.A(g7230), .B(g4979), .Z(g10465) ) ;
AND2    gate18191  (.A(g3722), .B(g4982), .Z(g10466) ) ;
AND2    gate18192  (.A(g3774), .B(g4994), .Z(g10467) ) ;
AND2    gate18193  (.A(g7265), .B(g4997), .Z(g10468) ) ;
AND2    gate18194  (.A(g5556), .B(g5000), .Z(g10469) ) ;
AND2    gate18195  (.A(g3774), .B(g2510), .Z(g10470) ) ;
AND2    gate18196  (.A(g7265), .B(g2516), .Z(g10471) ) ;
AND2    gate18197  (.A(g7391), .B(g2645), .Z(g10472) ) ;
AND2    gate18198  (.A(g7303), .B(g5005), .Z(g10473) ) ;
AND2    gate18199  (.A(g7303), .B(g2661), .Z(g10474) ) ;
AND2    gate18200  (.A(g3834), .B(g5009), .Z(g10475) ) ;
AND2    gate18201  (.A(g7488), .B(g5012), .Z(g10476) ) ;
AND2    gate18202  (.A(g7426), .B(g5015), .Z(g10477) ) ;
AND2    gate18203  (.A(g7488), .B(g5018), .Z(g10478) ) ;
AND2    gate18204  (.A(g7426), .B(g5021), .Z(g10479) ) ;
AND3    gate18205  (.A(g6901), .B(g7338), .C(g7146), .Z(II17429) ) ;
AND2    gate18206  (.A(g6448), .B(g5024), .Z(g10485) ) ;
AND2    gate18207  (.A(g3338), .B(g5027), .Z(g10492) ) ;
AND2    gate18208  (.A(g6643), .B(g5030), .Z(g10493) ) ;
AND2    gate18209  (.A(g6643), .B(g608), .Z(g10494) ) ;
AND2    gate18210  (.A(g6486), .B(g614), .Z(g10495) ) ;
AND2    gate18211  (.A(g3366), .B(g5035), .Z(g10496) ) ;
AND2    gate18212  (.A(g6912), .B(g5038), .Z(g10497) ) ;
AND2    gate18213  (.A(g3462), .B(g5041), .Z(g10498) ) ;
AND2    gate18214  (.A(g5473), .B(g5044), .Z(g10499) ) ;
AND2    gate18215  (.A(g3494), .B(g5047), .Z(g10506) ) ;
AND2    gate18216  (.A(g6945), .B(g5050), .Z(g10507) ) ;
AND2    gate18217  (.A(g6751), .B(g5053), .Z(g10508) ) ;
AND2    gate18218  (.A(g3494), .B(g1288), .Z(g10509) ) ;
AND2    gate18219  (.A(g6751), .B(g1291), .Z(g10510) ) ;
AND2    gate18220  (.A(g3522), .B(g5058), .Z(g10511) ) ;
AND2    gate18221  (.A(g7162), .B(g5061), .Z(g10512) ) ;
AND2    gate18222  (.A(g6980), .B(g5064), .Z(g10513) ) ;
AND2    gate18223  (.A(g3522), .B(g5067), .Z(g10514) ) ;
AND2    gate18224  (.A(g3618), .B(g5072), .Z(g10515) ) ;
AND2    gate18225  (.A(g7015), .B(g5075), .Z(g10516) ) ;
AND2    gate18226  (.A(g3650), .B(g5078), .Z(g10517) ) ;
AND2    gate18227  (.A(g7195), .B(g5081), .Z(g10518) ) ;
AND2    gate18228  (.A(g7053), .B(g5084), .Z(g10519) ) ;
AND2    gate18229  (.A(g3650), .B(g1973), .Z(g10520) ) ;
AND2    gate18230  (.A(g7195), .B(g1979), .Z(g10521) ) ;
AND2    gate18231  (.A(g3678), .B(g5089), .Z(g10522) ) ;
AND2    gate18232  (.A(g7358), .B(g5092), .Z(g10523) ) ;
AND2    gate18233  (.A(g7230), .B(g5095), .Z(g10524) ) ;
AND2    gate18234  (.A(g3678), .B(g5098), .Z(g10525) ) ;
AND2    gate18235  (.A(g7358), .B(g5101), .Z(g10526) ) ;
AND2    gate18236  (.A(g3774), .B(g5104), .Z(g10527) ) ;
AND2    gate18237  (.A(g7265), .B(g5107), .Z(g10528) ) ;
AND2    gate18238  (.A(g5556), .B(g5110), .Z(g10529) ) ;
AND2    gate18239  (.A(g3774), .B(g2519), .Z(g10530) ) ;
AND2    gate18240  (.A(g3806), .B(g2647), .Z(g10531) ) ;
AND2    gate18241  (.A(g7391), .B(g5115), .Z(g10532) ) ;
AND2    gate18242  (.A(g7303), .B(g5118), .Z(g10533) ) ;
AND2    gate18243  (.A(g7391), .B(g2664), .Z(g10534) ) ;
AND2    gate18244  (.A(g7303), .B(g2670), .Z(g10535) ) ;
AND2    gate18245  (.A(g3834), .B(g5123), .Z(g10536) ) ;
AND2    gate18246  (.A(g7488), .B(g5126), .Z(g10537) ) ;
AND2    gate18247  (.A(g7426), .B(g5129), .Z(g10538) ) ;
AND2    gate18248  (.A(g3834), .B(g5132), .Z(g10539) ) ;
AND2    gate18249  (.A(g7488), .B(g5135), .Z(g10540) ) ;
AND2    gate18250  (.A(g7426), .B(g5138), .Z(g10541) ) ;
AND2    gate18251  (.A(g3306), .B(g5142), .Z(g10548) ) ;
AND2    gate18252  (.A(g3338), .B(g5145), .Z(g10555) ) ;
AND2    gate18253  (.A(g3338), .B(g611), .Z(g10556) ) ;
AND2    gate18254  (.A(g6643), .B(g617), .Z(g10557) ) ;
AND2    gate18255  (.A(g3366), .B(g5150), .Z(g10558) ) ;
AND2    gate18256  (.A(g6713), .B(g5153), .Z(g10559) ) ;
AND2    gate18257  (.A(g3494), .B(g5156), .Z(g10566) ) ;
AND2    gate18258  (.A(g6945), .B(g5159), .Z(g10567) ) ;
AND2    gate18259  (.A(g6945), .B(g1294), .Z(g10568) ) ;
AND2    gate18260  (.A(g6751), .B(g1300), .Z(g10569) ) ;
AND2    gate18261  (.A(g3522), .B(g5164), .Z(g10570) ) ;
AND2    gate18262  (.A(g7162), .B(g5167), .Z(g10571) ) ;
AND2    gate18263  (.A(g3618), .B(g5170), .Z(g10572) ) ;
AND2    gate18264  (.A(g5512), .B(g5173), .Z(g10573) ) ;
AND2    gate18265  (.A(g3650), .B(g5176), .Z(g10580) ) ;
AND2    gate18266  (.A(g7195), .B(g5179), .Z(g10581) ) ;
AND2    gate18267  (.A(g7053), .B(g5182), .Z(g10582) ) ;
AND2    gate18268  (.A(g3650), .B(g1982), .Z(g10583) ) ;
AND2    gate18269  (.A(g7053), .B(g1985), .Z(g10584) ) ;
AND2    gate18270  (.A(g3678), .B(g5187), .Z(g10585) ) ;
AND2    gate18271  (.A(g7358), .B(g5190), .Z(g10586) ) ;
AND2    gate18272  (.A(g7230), .B(g5193), .Z(g10587) ) ;
AND2    gate18273  (.A(g3678), .B(g5196), .Z(g10588) ) ;
AND2    gate18274  (.A(g3774), .B(g5201), .Z(g10589) ) ;
AND2    gate18275  (.A(g7265), .B(g5204), .Z(g10590) ) ;
AND2    gate18276  (.A(g3806), .B(g5207), .Z(g10591) ) ;
AND2    gate18277  (.A(g7391), .B(g5210), .Z(g10592) ) ;
AND2    gate18278  (.A(g7303), .B(g5213), .Z(g10593) ) ;
AND2    gate18279  (.A(g3806), .B(g2667), .Z(g10594) ) ;
AND2    gate18280  (.A(g7391), .B(g2673), .Z(g10595) ) ;
AND2    gate18281  (.A(g3834), .B(g5218), .Z(g10596) ) ;
AND2    gate18282  (.A(g7488), .B(g5221), .Z(g10597) ) ;
AND2    gate18283  (.A(g7426), .B(g5224), .Z(g10598) ) ;
AND2    gate18284  (.A(g3834), .B(g5227), .Z(g10599) ) ;
AND2    gate18285  (.A(g7488), .B(g5230), .Z(g10600) ) ;
AND2    gate18286  (.A(g3338), .B(g620), .Z(g10604) ) ;
AND2    gate18287  (.A(g3462), .B(g5235), .Z(g10605) ) ;
AND2    gate18288  (.A(g3494), .B(g5238), .Z(g10612) ) ;
AND2    gate18289  (.A(g3494), .B(g1297), .Z(g10613) ) ;
AND2    gate18290  (.A(g6945), .B(g1303), .Z(g10614) ) ;
AND2    gate18291  (.A(g3522), .B(g5243), .Z(g10615) ) ;
AND2    gate18292  (.A(g7015), .B(g5246), .Z(g10616) ) ;
AND2    gate18293  (.A(g3650), .B(g5249), .Z(g10623) ) ;
AND2    gate18294  (.A(g7195), .B(g5252), .Z(g10624) ) ;
AND2    gate18295  (.A(g7195), .B(g1988), .Z(g10625) ) ;
AND2    gate18296  (.A(g7053), .B(g1994), .Z(g10626) ) ;
AND2    gate18297  (.A(g3678), .B(g5257), .Z(g10627) ) ;
AND2    gate18298  (.A(g7358), .B(g5260), .Z(g10628) ) ;
AND2    gate18299  (.A(g3774), .B(g5263), .Z(g10629) ) ;
AND2    gate18300  (.A(g5556), .B(g5266), .Z(g10630) ) ;
AND2    gate18301  (.A(g3806), .B(g5269), .Z(g10637) ) ;
AND2    gate18302  (.A(g7391), .B(g5272), .Z(g10638) ) ;
AND2    gate18303  (.A(g7303), .B(g5275), .Z(g10639) ) ;
AND2    gate18304  (.A(g3806), .B(g2676), .Z(g10640) ) ;
AND2    gate18305  (.A(g7303), .B(g2679), .Z(g10641) ) ;
AND2    gate18306  (.A(g3834), .B(g5280), .Z(g10642) ) ;
AND2    gate18307  (.A(g7488), .B(g5283), .Z(g10643) ) ;
AND2    gate18308  (.A(g7426), .B(g5286), .Z(g10644) ) ;
AND2    gate18309  (.A(g3834), .B(g5289), .Z(g10645) ) ;
AND2    gate18310  (.A(g6678), .B(g5293), .Z(g10650) ) ;
AND2    gate18311  (.A(g3494), .B(g1306), .Z(g10651) ) ;
AND2    gate18312  (.A(g3618), .B(g5298), .Z(g10652) ) ;
AND2    gate18313  (.A(g3650), .B(g5301), .Z(g10659) ) ;
AND2    gate18314  (.A(g3650), .B(g1991), .Z(g10660) ) ;
AND2    gate18315  (.A(g7195), .B(g1997), .Z(g10661) ) ;
AND2    gate18316  (.A(g3678), .B(g5306), .Z(g10662) ) ;
AND2    gate18317  (.A(g7265), .B(g5309), .Z(g10663) ) ;
AND2    gate18318  (.A(g3806), .B(g5312), .Z(g10670) ) ;
AND2    gate18319  (.A(g7391), .B(g5315), .Z(g10671) ) ;
AND2    gate18320  (.A(g7391), .B(g2682), .Z(g10672) ) ;
AND2    gate18321  (.A(g7303), .B(g2688), .Z(g10673) ) ;
AND2    gate18322  (.A(g3834), .B(g5320), .Z(g10674) ) ;
AND2    gate18323  (.A(g7488), .B(g5323), .Z(g10675) ) ;
AND2    gate18324  (.A(g6912), .B(g5327), .Z(g10678) ) ;
AND2    gate18325  (.A(g6980), .B(g5330), .Z(g10680) ) ;
AND2    gate18326  (.A(g3650), .B(g2000), .Z(g10681) ) ;
AND2    gate18327  (.A(g3774), .B(g5335), .Z(g10682) ) ;
AND2    gate18328  (.A(g3806), .B(g5338), .Z(g10689) ) ;
AND2    gate18329  (.A(g3806), .B(g2685), .Z(g10690) ) ;
AND2    gate18330  (.A(g7391), .B(g2691), .Z(g10691) ) ;
AND2    gate18331  (.A(g3834), .B(g5343), .Z(g10692) ) ;
AND4    gate18332  (.A(g7462), .B(g7522), .C(g2924), .D(g7545), .Z(g10693) ) ;
AND2    gate18333  (.A(g3366), .B(g5352), .Z(g10704) ) ;
AND2    gate18334  (.A(g7162), .B(g5355), .Z(g10707) ) ;
AND2    gate18335  (.A(g7230), .B(g5358), .Z(g10709) ) ;
AND2    gate18336  (.A(g3806), .B(g2694), .Z(g10710) ) ;
AND3    gate18337  (.A(g7566), .B(g7583), .C(g7587), .Z(II17599) ) ;
AND2    gate18338  (.A(g3522), .B(g5369), .Z(g10724) ) ;
AND2    gate18339  (.A(g7358), .B(g5372), .Z(g10727) ) ;
AND2    gate18340  (.A(g7426), .B(g5375), .Z(g10729) ) ;
AND2    gate18341  (.A(g3678), .B(g5382), .Z(g10745) ) ;
AND2    gate18342  (.A(g7488), .B(g5385), .Z(g10748) ) ;
AND2    gate18343  (.A(g3834), .B(g5391), .Z(g10764) ) ;
AND2    gate18344  (.A(g6232), .B(g213), .Z(g11347) ) ;
AND2    gate18345  (.A(g6314), .B(g216), .Z(g11420) ) ;
AND2    gate18346  (.A(g6232), .B(g222), .Z(g11421) ) ;
AND2    gate18347  (.A(g6369), .B(g900), .Z(g11431) ) ;
AND2    gate18348  (.A(g5871), .B(g8360), .Z(g11607) ) ;
AND2    gate18349  (.A(g5881), .B(g8378), .Z(g11612) ) ;
AND2    gate18350  (.A(g5918), .B(g8427), .Z(g11637) ) ;
AND2    gate18351  (.A(g554), .B(g8622), .Z(g11771) ) ;
AND2    gate18352  (.A(g1240), .B(g8632), .Z(g11788) ) ;
AND2    gate18353  (.A(g6173), .B(g8643), .Z(g11805) ) ;
AND2    gate18354  (.A(g1934), .B(g8651), .Z(g11814) ) ;
AND2    gate18355  (.A(g7869), .B(g8655), .Z(g11816) ) ;
AND2    gate18356  (.A(g6205), .B(g8659), .Z(g11838) ) ;
AND2    gate18357  (.A(g2628), .B(g8667), .Z(g11847) ) ;
AND2    gate18358  (.A(g7849), .B(g8670), .Z(g11851) ) ;
AND2    gate18359  (.A(g6294), .B(g8678), .Z(g11880) ) ;
AND2    gate18360  (.A(g7834), .B(g8684), .Z(g11885) ) ;
AND2    gate18361  (.A(g6431), .B(g8690), .Z(g11922) ) ;
AND2    gate18362  (.A(g8169), .B(g8696), .Z(g11926) ) ;
AND2    gate18363  (.A(g8090), .B(g8708), .Z(g11966) ) ;
AND2    gate18364  (.A(g7967), .B(g8711), .Z(g11967) ) ;
AND2    gate18365  (.A(g8015), .B(g8745), .Z(g12012) ) ;
AND2    gate18366  (.A(g7964), .B(g8763), .Z(g12069) ) ;
AND2    gate18367  (.A(g8018), .B(g8766), .Z(g12070) ) ;
AND2    gate18368  (.A(g7916), .B(g8785), .Z(g12128) ) ;
AND2    gate18369  (.A(g7872), .B(g8788), .Z(g12129) ) ;
AND2    gate18370  (.A(g8093), .B(g8805), .Z(g12186) ) ;
AND2    gate18371  (.A(g8172), .B(g8829), .Z(g12273) ) ;
AND2    gate18372  (.A(g7900), .B(g8832), .Z(g12274) ) ;
AND2    gate18373  (.A(g7919), .B(g8853), .Z(g12307) ) ;
AND2    gate18374  (.A(g8246), .B(g8879), .Z(g12330) ) ;
AND2    gate18375  (.A(g7927), .B(g8882), .Z(g12331) ) ;
AND2    gate18376  (.A(g7852), .B(g8915), .Z(g12353) ) ;
AND2    gate18377  (.A(g7974), .B(g8949), .Z(g12376) ) ;
AND2    gate18378  (.A(g8028), .B(g9006), .Z(g12419) ) ;
AND2    gate18379  (.A(g8101), .B(g9044), .Z(g12429) ) ;
AND2    gate18380  (.A(g7822), .B(g9128), .Z(g12477) ) ;
AND2    gate18381  (.A(g7833), .B(g9134), .Z(g12494) ) ;
AND2    gate18382  (.A(g7848), .B(g9140), .Z(g12514) ) ;
AND2    gate18383  (.A(g7868), .B(g9146), .Z(g12531) ) ;
AND2    gate18384  (.A(g6149), .B(g9290), .Z(g12650) ) ;
AND4    gate18385  (.A(g9507), .B(g9427), .C(g9356), .D(g9293), .Z(II19937) ) ;
AND4    gate18386  (.A(g9232), .B(g9187), .C(g9161), .D(g9150), .Z(II19938) ) ;
AND2    gate18387  (.A(II19937), .B(II19938), .Z(g12876) ) ;
AND2    gate18388  (.A(g7899), .B(g10004), .Z(g12908) ) ;
AND4    gate18389  (.A(g9649), .B(g9569), .C(g9453), .D(g9374), .Z(II19971) ) ;
AND4    gate18390  (.A(g9310), .B(g9248), .C(g9203), .D(g9174), .Z(II19972) ) ;
AND2    gate18391  (.A(II19971), .B(II19972), .Z(g12916) ) ;
AND2    gate18392  (.A(g8179), .B(g10096), .Z(g12938) ) ;
AND4    gate18393  (.A(g9795), .B(g9711), .C(g9595), .D(g9471), .Z(II19996) ) ;
AND4    gate18394  (.A(g9391), .B(g9326), .C(g9264), .D(g9216), .Z(II19997) ) ;
AND2    gate18395  (.A(II19996), .B(II19997), .Z(g12945) ) ;
AND2    gate18396  (.A(g7926), .B(g10189), .Z(g12966) ) ;
AND4    gate18397  (.A(g9941), .B(g9857), .C(g9737), .D(g9613), .Z(II20021) ) ;
AND4    gate18398  (.A(g9488), .B(g9407), .C(g9342), .D(g9277), .Z(II20022) ) ;
AND2    gate18399  (.A(II20021), .B(II20022), .Z(g12974) ) ;
AND2    gate18400  (.A(g8254), .B(g10273), .Z(g12989) ) ;
AND2    gate18401  (.A(g8180), .B(g10276), .Z(g12990) ) ;
AND2    gate18402  (.A(g7973), .B(g10357), .Z(g13000) ) ;
AND2    gate18403  (.A(g3995), .B(g10416), .Z(g13009) ) ;
AND2    gate18404  (.A(g8255), .B(g10419), .Z(g13010) ) ;
AND2    gate18405  (.A(g8027), .B(g10482), .Z(g13023) ) ;
AND2    gate18406  (.A(g7879), .B(g10542), .Z(g13031) ) ;
AND2    gate18407  (.A(g3996), .B(g10545), .Z(g13032) ) ;
AND2    gate18408  (.A(g8100), .B(g10601), .Z(g13042) ) ;
AND3    gate18409  (.A(g10186), .B(g3018), .C(g3028), .Z(II20100) ) ;
AND2    gate18410  (.A(g4092), .B(g10646), .Z(g13056) ) ;
AND4    gate18411  (.A(g8313), .B(g7542), .C(g2888), .D(g7566), .Z(II20131) ) ;
AND4    gate18412  (.A(g2892), .B(g2903), .C(g7595), .D(g2908), .Z(II20132) ) ;
AND2    gate18413  (.A(g298), .B(g11032), .Z(g13247) ) ;
AND2    gate18414  (.A(g5628), .B(g11088), .Z(g13266) ) ;
AND2    gate18415  (.A(g985), .B(g11102), .Z(g13270) ) ;
AND2    gate18416  (.A(g5647), .B(g11141), .Z(g13289) ) ;
AND2    gate18417  (.A(g5656), .B(g11154), .Z(g13291) ) ;
AND2    gate18418  (.A(g1679), .B(g11170), .Z(g13295) ) ;
AND2    gate18419  (.A(g5675), .B(g11210), .Z(g13316) ) ;
AND2    gate18420  (.A(g5685), .B(g11225), .Z(g13320) ) ;
AND2    gate18421  (.A(g5694), .B(g11240), .Z(g13322) ) ;
AND2    gate18422  (.A(g2373), .B(g11256), .Z(g13326) ) ;
AND2    gate18423  (.A(g5708), .B(g11278), .Z(g13335) ) ;
AND2    gate18424  (.A(g5727), .B(g11294), .Z(g13340) ) ;
AND2    gate18425  (.A(g5737), .B(g11309), .Z(g13343) ) ;
AND2    gate18426  (.A(g5746), .B(g11324), .Z(g13345) ) ;
AND2    gate18427  (.A(g5756), .B(g11355), .Z(g13355) ) ;
AND2    gate18428  (.A(g5766), .B(g11373), .Z(g13360) ) ;
AND2    gate18429  (.A(g5785), .B(g11389), .Z(g13365) ) ;
AND2    gate18430  (.A(g5795), .B(g11404), .Z(g13368) ) ;
AND2    gate18431  (.A(g5815), .B(g11441), .Z(g13385) ) ;
AND2    gate18432  (.A(g5825), .B(g11459), .Z(g13390) ) ;
AND2    gate18433  (.A(g5844), .B(g11475), .Z(g13395) ) ;
AND2    gate18434  (.A(g6016), .B(g12191), .Z(g13477) ) ;
AND2    gate18435  (.A(g6017), .B(g12196), .Z(g13479) ) ;
AND2    gate18436  (.A(g6018), .B(g12197), .Z(g13480) ) ;
AND2    gate18437  (.A(g5864), .B(g11603), .Z(g13481) ) ;
AND2    gate18438  (.A(g6020), .B(g12209), .Z(g13483) ) ;
AND2    gate18439  (.A(g6021), .B(g12210), .Z(g13484) ) ;
AND2    gate18440  (.A(g6022), .B(g12211), .Z(g13485) ) ;
AND2    gate18441  (.A(g6023), .B(g12212), .Z(g13486) ) ;
AND2    gate18442  (.A(g5874), .B(g11608), .Z(g13487) ) ;
AND2    gate18443  (.A(g6025), .B(g12218), .Z(g13488) ) ;
AND2    gate18444  (.A(g6026), .B(g12219), .Z(g13489) ) ;
AND2    gate18445  (.A(g6027), .B(g12220), .Z(g13490) ) ;
AND2    gate18446  (.A(g6028), .B(g12221), .Z(g13491) ) ;
AND2    gate18447  (.A(g2371), .B(g12222), .Z(g13492) ) ;
AND2    gate18448  (.A(g5887), .B(g11613), .Z(g13493) ) ;
AND2    gate18449  (.A(g6032), .B(g12246), .Z(g13496) ) ;
AND2    gate18450  (.A(g6033), .B(g12251), .Z(g13498) ) ;
AND2    gate18451  (.A(g6034), .B(g12252), .Z(g13499) ) ;
AND2    gate18452  (.A(g5911), .B(g11633), .Z(g13500) ) ;
AND2    gate18453  (.A(g6036), .B(g12264), .Z(g13502) ) ;
AND2    gate18454  (.A(g6037), .B(g12265), .Z(g13503) ) ;
AND2    gate18455  (.A(g6038), .B(g12266), .Z(g13504) ) ;
AND2    gate18456  (.A(g6039), .B(g12267), .Z(g13505) ) ;
AND2    gate18457  (.A(g5921), .B(g11638), .Z(g13506) ) ;
AND2    gate18458  (.A(g6043), .B(g12289), .Z(g13513) ) ;
AND2    gate18459  (.A(g6044), .B(g12294), .Z(g13515) ) ;
AND2    gate18460  (.A(g6045), .B(g12295), .Z(g13516) ) ;
AND2    gate18461  (.A(g5950), .B(g11656), .Z(g13517) ) ;
AND2    gate18462  (.A(g6047), .B(g12325), .Z(g13527) ) ;
AND2    gate18463  (.A(g6141), .B(g12456), .Z(g13609) ) ;
AND2    gate18464  (.A(g6162), .B(g12466), .Z(g13619) ) ;
AND2    gate18465  (.A(g5428), .B(g12472), .Z(g13623) ) ;
AND2    gate18466  (.A(g6173), .B(g12476), .Z(g13625) ) ;
AND2    gate18467  (.A(g6189), .B(g12481), .Z(g13631) ) ;
AND2    gate18468  (.A(g12776), .B(g8617), .Z(g13634) ) ;
AND2    gate18469  (.A(g6205), .B(g12493), .Z(g13636) ) ;
AND2    gate18470  (.A(g6221), .B(g12498), .Z(g13642) ) ;
AND2    gate18471  (.A(g5431), .B(g12502), .Z(g13643) ) ;
AND2    gate18472  (.A(g6281), .B(g12504), .Z(g13645) ) ;
AND2    gate18473  (.A(g7772), .B(g12505), .Z(g13646) ) ;
AND2    gate18474  (.A(g6294), .B(g12513), .Z(g13648) ) ;
AND2    gate18475  (.A(g8093), .B(g11791), .Z(g13654) ) ;
AND2    gate18476  (.A(g7540), .B(g12518), .Z(g13655) ) ;
AND2    gate18477  (.A(g12776), .B(g8640), .Z(g13656) ) ;
AND2    gate18478  (.A(g6418), .B(g12521), .Z(g13671) ) ;
AND2    gate18479  (.A(g7788), .B(g12522), .Z(g13672) ) ;
AND2    gate18480  (.A(g6431), .B(g12530), .Z(g13674) ) ;
AND2    gate18481  (.A(g7561), .B(g12532), .Z(g13675) ) ;
AND2    gate18482  (.A(g5434), .B(g12533), .Z(g13676) ) ;
AND2    gate18483  (.A(g6623), .B(g12536), .Z(g13701) ) ;
AND2    gate18484  (.A(g7802), .B(g12537), .Z(g13702) ) ;
AND2    gate18485  (.A(g8018), .B(g11848), .Z(g13703) ) ;
AND2    gate18486  (.A(g7581), .B(g12542), .Z(g13704) ) ;
AND2    gate18487  (.A(g12776), .B(g8673), .Z(g13705) ) ;
AND2    gate18488  (.A(g6887), .B(g12545), .Z(g13738) ) ;
AND2    gate18489  (.A(g7815), .B(g12546), .Z(g13739) ) ;
AND2    gate18490  (.A(g6636), .B(g12547), .Z(g13740) ) ;
AND2    gate18491  (.A(g7347), .B(g12551), .Z(g13755) ) ;
AND2    gate18492  (.A(g7967), .B(g11923), .Z(g13787) ) ;
AND2    gate18493  (.A(g6897), .B(g12553), .Z(g13788) ) ;
AND2    gate18494  (.A(g7140), .B(g12554), .Z(g13789) ) ;
AND2    gate18495  (.A(g7475), .B(g12558), .Z(g13790) ) ;
AND2    gate18496  (.A(g7477), .B(g12559), .Z(g13796) ) ;
AND2    gate18497  (.A(g7139), .B(g12560), .Z(g13815) ) ;
AND2    gate18498  (.A(g7530), .B(g12596), .Z(g13816) ) ;
AND2    gate18499  (.A(g7531), .B(g12597), .Z(g13818) ) ;
AND2    gate18500  (.A(g7533), .B(g12598), .Z(g13824) ) ;
AND2    gate18501  (.A(g7919), .B(g12009), .Z(g13833) ) ;
AND2    gate18502  (.A(g7336), .B(g12599), .Z(g13834) ) ;
AND2    gate18503  (.A(g7461), .B(g12600), .Z(g13835) ) ;
AND2    gate18504  (.A(g7556), .B(g12642), .Z(g13837) ) ;
AND2    gate18505  (.A(g7557), .B(g12643), .Z(g13839) ) ;
AND2    gate18506  (.A(g7559), .B(g12644), .Z(g13845) ) ;
AND2    gate18507  (.A(g7460), .B(g12645), .Z(g13846) ) ;
AND2    gate18508  (.A(g7521), .B(g12646), .Z(g13847) ) ;
AND2    gate18509  (.A(g7579), .B(g12688), .Z(g13851) ) ;
AND2    gate18510  (.A(g7580), .B(g12689), .Z(g13853) ) ;
AND2    gate18511  (.A(g5349), .B(g12690), .Z(g13854) ) ;
AND2    gate18512  (.A(g7541), .B(g12691), .Z(g13855) ) ;
AND2    gate18513  (.A(g7593), .B(g12742), .Z(g13860) ) ;
AND2    gate18514  (.A(g5366), .B(g12743), .Z(g13862) ) ;
AND2    gate18515  (.A(g7582), .B(g12768), .Z(g13870) ) ;
AND2    gate18516  (.A(g7898), .B(g12775), .Z(g13871) ) ;
AND2    gate18517  (.A(g7610), .B(g12782), .Z(g13878) ) ;
AND2    gate18518  (.A(g1234), .B(g12790), .Z(g13880) ) ;
AND2    gate18519  (.A(g7594), .B(g12807), .Z(g13884) ) ;
AND2    gate18520  (.A(g7616), .B(g12815), .Z(g13892) ) ;
AND2    gate18521  (.A(g7619), .B(g12821), .Z(g13900) ) ;
AND2    gate18522  (.A(g1928), .B(g12829), .Z(g13902) ) ;
AND2    gate18523  (.A(g7337), .B(g12843), .Z(g13904) ) ;
AND2    gate18524  (.A(g7925), .B(g12847), .Z(g13905) ) ;
AND2    gate18525  (.A(g7623), .B(g12850), .Z(g13913) ) ;
AND2    gate18526  (.A(g7626), .B(g12851), .Z(g13914) ) ;
AND2    gate18527  (.A(g7632), .B(g12853), .Z(g13933) ) ;
AND2    gate18528  (.A(g7635), .B(g12859), .Z(g13941) ) ;
AND2    gate18529  (.A(g2622), .B(g12867), .Z(g13943) ) ;
AND2    gate18530  (.A(g7141), .B(g12874), .Z(g13944) ) ;
AND2    gate18531  (.A(g7643), .B(g12881), .Z(g13952) ) ;
AND2    gate18532  (.A(g7646), .B(g12882), .Z(g13953) ) ;
AND2    gate18533  (.A(g7652), .B(g12891), .Z(g13969) ) ;
AND2    gate18534  (.A(g7655), .B(g12892), .Z(g13970) ) ;
AND2    gate18535  (.A(g7661), .B(g12894), .Z(g13989) ) ;
AND2    gate18536  (.A(g7664), .B(g12900), .Z(g13997) ) ;
AND2    gate18537  (.A(g7972), .B(g12907), .Z(g13998) ) ;
AND2    gate18538  (.A(g7670), .B(g12914), .Z(g14006) ) ;
AND2    gate18539  (.A(g7673), .B(g12915), .Z(g14007) ) ;
AND2    gate18540  (.A(g7679), .B(g12921), .Z(g14022) ) ;
AND2    gate18541  (.A(g7682), .B(g12922), .Z(g14023) ) ;
AND2    gate18542  (.A(g7688), .B(g12931), .Z(g14039) ) ;
AND2    gate18543  (.A(g7691), .B(g12932), .Z(g14040) ) ;
AND2    gate18544  (.A(g7697), .B(g12934), .Z(g14059) ) ;
AND2    gate18545  (.A(g7703), .B(g12940), .Z(g14067) ) ;
AND2    gate18546  (.A(g7706), .B(g12943), .Z(g14097) ) ;
AND2    gate18547  (.A(g7709), .B(g12944), .Z(g14098) ) ;
AND2    gate18548  (.A(g7715), .B(g12950), .Z(g14113) ) ;
AND2    gate18549  (.A(g7718), .B(g12951), .Z(g14114) ) ;
AND2    gate18550  (.A(g7724), .B(g12960), .Z(g14130) ) ;
AND2    gate18551  (.A(g7727), .B(g12961), .Z(g14131) ) ;
AND2    gate18552  (.A(g8026), .B(g12965), .Z(g14143) ) ;
AND2    gate18553  (.A(g7733), .B(g12969), .Z(g14182) ) ;
AND2    gate18554  (.A(g7736), .B(g12972), .Z(g14212) ) ;
AND2    gate18555  (.A(g7739), .B(g12973), .Z(g14213) ) ;
AND2    gate18556  (.A(g7745), .B(g12979), .Z(g14228) ) ;
AND2    gate18557  (.A(g7748), .B(g12980), .Z(g14229) ) ;
AND2    gate18558  (.A(g7757), .B(g12993), .Z(g14297) ) ;
AND2    gate18559  (.A(g7760), .B(g12996), .Z(g14327) ) ;
AND2    gate18560  (.A(g7763), .B(g12997), .Z(g14328) ) ;
AND2    gate18561  (.A(g8099), .B(g12998), .Z(g14336) ) ;
AND2    gate18562  (.A(g7779), .B(g13003), .Z(g14419) ) ;
AND2    gate18563  (.A(g7841), .B(g13101), .Z(g14690) ) ;
AND2    gate18564  (.A(g7861), .B(g13117), .Z(g14724) ) ;
AND2    gate18565  (.A(g7891), .B(g13130), .Z(g14752) ) ;
NAND2   gate18566  (.A(g10779), .B(g7901), .Z(g13245) ) ;
AND2    gate18567  (.A(g13245), .B(g10765), .Z(g14767) ) ;
AND2    gate18568  (.A(g7915), .B(g13141), .Z(g14773) ) ;
AND2    gate18569  (.A(g8169), .B(g12548), .Z(g14884) ) ;
AND2    gate18570  (.A(g3940), .B(g13148), .Z(g14894) ) ;
AND2    gate18571  (.A(g11059), .B(g13151), .Z(g14956) ) ;
AND2    gate18572  (.A(g4015), .B(g13152), .Z(g14957) ) ;
AND2    gate18573  (.A(g4016), .B(g13153), .Z(g14958) ) ;
AND2    gate18574  (.A(g4047), .B(g13154), .Z(g14975) ) ;
AND2    gate18575  (.A(g8090), .B(g12561), .Z(g15020) ) ;
AND2    gate18576  (.A(g4110), .B(g13158), .Z(g15030) ) ;
AND2    gate18577  (.A(g4111), .B(g13159), .Z(g15031) ) ;
AND2    gate18578  (.A(g4142), .B(g13161), .Z(g15046) ) ;
AND2    gate18579  (.A(g4143), .B(g13162), .Z(g15047) ) ;
AND2    gate18580  (.A(g4174), .B(g13163), .Z(g15064) ) ;
AND2    gate18581  (.A(g7869), .B(g12601), .Z(g15093) ) ;
AND2    gate18582  (.A(g7872), .B(g12604), .Z(g15094) ) ;
AND2    gate18583  (.A(g4220), .B(g13167), .Z(g15104) ) ;
AND2    gate18584  (.A(g4224), .B(g13168), .Z(g15105) ) ;
AND2    gate18585  (.A(g4249), .B(g13169), .Z(g15126) ) ;
AND2    gate18586  (.A(g4250), .B(g13170), .Z(g15127) ) ;
AND2    gate18587  (.A(g4281), .B(g13172), .Z(g15142) ) ;
AND2    gate18588  (.A(g4282), .B(g13173), .Z(g15143) ) ;
AND2    gate18589  (.A(g4313), .B(g13174), .Z(g15160) ) ;
AND2    gate18590  (.A(g8015), .B(g12647), .Z(g15171) ) ;
AND2    gate18591  (.A(g4346), .B(g13176), .Z(g15172) ) ;
AND2    gate18592  (.A(g4347), .B(g13177), .Z(g15173) ) ;
AND2    gate18593  (.A(g640), .B(g12651), .Z(g15178) ) ;
AND2    gate18594  (.A(g4375), .B(g13178), .Z(g15196) ) ;
AND2    gate18595  (.A(g4379), .B(g13179), .Z(g15197) ) ;
AND2    gate18596  (.A(g4404), .B(g13180), .Z(g15218) ) ;
AND2    gate18597  (.A(g4405), .B(g13181), .Z(g15219) ) ;
AND2    gate18598  (.A(g4436), .B(g13183), .Z(g15234) ) ;
AND2    gate18599  (.A(g4437), .B(g13184), .Z(g15235) ) ;
AND2    gate18600  (.A(g7849), .B(g12692), .Z(g15243) ) ;
AND2    gate18601  (.A(g7852), .B(g12695), .Z(g15244) ) ;
AND2    gate18602  (.A(g4474), .B(g13185), .Z(g15245) ) ;
AND2    gate18603  (.A(g4475), .B(g13186), .Z(g15246) ) ;
AND2    gate18604  (.A(g4479), .B(g13187), .Z(g15247) ) ;
AND2    gate18605  (.A(g4357), .B(g12702), .Z(g15257) ) ;
AND2    gate18606  (.A(g4515), .B(g13188), .Z(g15258) ) ;
AND2    gate18607  (.A(g4516), .B(g13189), .Z(g15259) ) ;
AND2    gate18608  (.A(g1326), .B(g12705), .Z(g15264) ) ;
AND2    gate18609  (.A(g4544), .B(g13190), .Z(g15282) ) ;
AND2    gate18610  (.A(g4548), .B(g13191), .Z(g15283) ) ;
AND2    gate18611  (.A(g4573), .B(g13192), .Z(g15304) ) ;
AND2    gate18612  (.A(g4574), .B(g13193), .Z(g15305) ) ;
AND2    gate18613  (.A(g7964), .B(g12744), .Z(g15320) ) ;
AND2    gate18614  (.A(g4601), .B(g13195), .Z(g15321) ) ;
AND2    gate18615  (.A(g4609), .B(g13196), .Z(g15324) ) ;
AND2    gate18616  (.A(g4610), .B(g13197), .Z(g15325) ) ;
AND2    gate18617  (.A(g4489), .B(g12749), .Z(g15335) ) ;
AND2    gate18618  (.A(g4492), .B(g12752), .Z(g15336) ) ;
AND2    gate18619  (.A(g4650), .B(g13198), .Z(g15337) ) ;
AND2    gate18620  (.A(g4651), .B(g13199), .Z(g15338) ) ;
AND2    gate18621  (.A(g4655), .B(g13200), .Z(g15339) ) ;
AND2    gate18622  (.A(g4526), .B(g12759), .Z(g15349) ) ;
AND2    gate18623  (.A(g4691), .B(g13201), .Z(g15350) ) ;
AND2    gate18624  (.A(g4692), .B(g13202), .Z(g15351) ) ;
AND2    gate18625  (.A(g2020), .B(g12762), .Z(g15356) ) ;
AND2    gate18626  (.A(g4720), .B(g13203), .Z(g15374) ) ;
AND2    gate18627  (.A(g4724), .B(g13204), .Z(g15375) ) ;
AND2    gate18628  (.A(g7834), .B(g12769), .Z(g15388) ) ;
AND2    gate18629  (.A(g8246), .B(g12772), .Z(g15389) ) ;
AND2    gate18630  (.A(g4752), .B(g13205), .Z(g15391) ) ;
AND2    gate18631  (.A(g4753), .B(g13206), .Z(g15392) ) ;
AND2    gate18632  (.A(g4620), .B(g12783), .Z(g15402) ) ;
AND2    gate18633  (.A(g4623), .B(g12786), .Z(g15403) ) ;
AND2    gate18634  (.A(g4778), .B(g13207), .Z(g15407) ) ;
AND2    gate18635  (.A(g4786), .B(g13208), .Z(g15410) ) ;
AND2    gate18636  (.A(g4787), .B(g13209), .Z(g15411) ) ;
AND2    gate18637  (.A(g4665), .B(g12791), .Z(g15421) ) ;
AND2    gate18638  (.A(g4668), .B(g12794), .Z(g15422) ) ;
AND2    gate18639  (.A(g4827), .B(g13210), .Z(g15423) ) ;
AND2    gate18640  (.A(g4828), .B(g13211), .Z(g15424) ) ;
AND2    gate18641  (.A(g4832), .B(g13212), .Z(g15425) ) ;
AND2    gate18642  (.A(g4702), .B(g12801), .Z(g15435) ) ;
AND2    gate18643  (.A(g4868), .B(g13213), .Z(g15436) ) ;
AND2    gate18644  (.A(g4869), .B(g13214), .Z(g15437) ) ;
AND2    gate18645  (.A(g2714), .B(g12804), .Z(g15442) ) ;
AND2    gate18646  (.A(g7916), .B(g12808), .Z(g15452) ) ;
AND2    gate18647  (.A(g6898), .B(g12811), .Z(g15453) ) ;
AND2    gate18648  (.A(g4897), .B(g13218), .Z(g15459) ) ;
AND2    gate18649  (.A(g4898), .B(g13219), .Z(g15460) ) ;
AND2    gate18650  (.A(g4763), .B(g12816), .Z(g15470) ) ;
AND2    gate18651  (.A(g4928), .B(g13220), .Z(g15475) ) ;
AND2    gate18652  (.A(g4929), .B(g13221), .Z(g15476) ) ;
AND2    gate18653  (.A(g4797), .B(g12822), .Z(g15486) ) ;
AND2    gate18654  (.A(g4800), .B(g12825), .Z(g15487) ) ;
AND2    gate18655  (.A(g4954), .B(g13222), .Z(g15491) ) ;
AND2    gate18656  (.A(g4962), .B(g13223), .Z(g15494) ) ;
AND2    gate18657  (.A(g4963), .B(g13224), .Z(g15495) ) ;
AND2    gate18658  (.A(g4842), .B(g12830), .Z(g15505) ) ;
AND2    gate18659  (.A(g4845), .B(g12833), .Z(g15506) ) ;
AND2    gate18660  (.A(g5003), .B(g13225), .Z(g15507) ) ;
AND2    gate18661  (.A(g5004), .B(g13226), .Z(g15508) ) ;
AND2    gate18662  (.A(g5008), .B(g13227), .Z(g15509) ) ;
AND2    gate18663  (.A(g4879), .B(g12840), .Z(g15519) ) ;
AND2    gate18664  (.A(g8172), .B(g12844), .Z(g15520) ) ;
AND2    gate18665  (.A(g5033), .B(g13232), .Z(g15526) ) ;
AND2    gate18666  (.A(g5034), .B(g13233), .Z(g15527) ) ;
AND2    gate18667  (.A(g5056), .B(g13237), .Z(g15545) ) ;
AND2    gate18668  (.A(g5057), .B(g13238), .Z(g15546) ) ;
AND2    gate18669  (.A(g4939), .B(g12854), .Z(g15556) ) ;
AND2    gate18670  (.A(g5087), .B(g13239), .Z(g15561) ) ;
AND2    gate18671  (.A(g5088), .B(g13240), .Z(g15562) ) ;
AND2    gate18672  (.A(g4973), .B(g12860), .Z(g15572) ) ;
AND2    gate18673  (.A(g4976), .B(g12863), .Z(g15573) ) ;
AND2    gate18674  (.A(g5113), .B(g13241), .Z(g15577) ) ;
AND2    gate18675  (.A(g5121), .B(g13242), .Z(g15580) ) ;
AND2    gate18676  (.A(g5122), .B(g13243), .Z(g15581) ) ;
AND2    gate18677  (.A(g5018), .B(g12868), .Z(g15591) ) ;
AND2    gate18678  (.A(g5021), .B(g12871), .Z(g15592) ) ;
AND2    gate18679  (.A(g7897), .B(g13244), .Z(g15593) ) ;
AND2    gate18680  (.A(g5148), .B(g13249), .Z(g15594) ) ;
AND2    gate18681  (.A(g5149), .B(g13250), .Z(g15595) ) ;
AND2    gate18682  (.A(g5162), .B(g13255), .Z(g15604) ) ;
AND2    gate18683  (.A(g5163), .B(g13256), .Z(g15605) ) ;
AND2    gate18684  (.A(g5185), .B(g13260), .Z(g15623) ) ;
AND2    gate18685  (.A(g5186), .B(g13261), .Z(g15624) ) ;
AND2    gate18686  (.A(g5098), .B(g12895), .Z(g15634) ) ;
AND2    gate18687  (.A(g5216), .B(g13262), .Z(g15639) ) ;
AND2    gate18688  (.A(g5217), .B(g13263), .Z(g15640) ) ;
AND2    gate18689  (.A(g5132), .B(g12901), .Z(g15650) ) ;
AND2    gate18690  (.A(g5135), .B(g12904), .Z(g15651) ) ;
AND2    gate18691  (.A(g8177), .B(g13264), .Z(g15658) ) ;
AND2    gate18692  (.A(g5233), .B(g13268), .Z(g15666) ) ;
AND2    gate18693  (.A(g5241), .B(g13272), .Z(g15670) ) ;
AND2    gate18694  (.A(g5242), .B(g13273), .Z(g15671) ) ;
AND2    gate18695  (.A(g5255), .B(g13278), .Z(g15680) ) ;
AND2    gate18696  (.A(g5256), .B(g13279), .Z(g15681) ) ;
AND2    gate18697  (.A(g5278), .B(g13283), .Z(g15699) ) ;
AND2    gate18698  (.A(g5279), .B(g13284), .Z(g15700) ) ;
AND2    gate18699  (.A(g5227), .B(g12935), .Z(g15710) ) ;
AND2    gate18700  (.A(g7924), .B(g13285), .Z(g15717) ) ;
AND2    gate18701  (.A(g5296), .B(g13293), .Z(g15725) ) ;
AND2    gate18702  (.A(g5304), .B(g13297), .Z(g15729) ) ;
AND2    gate18703  (.A(g5305), .B(g13298), .Z(g15730) ) ;
AND2    gate18704  (.A(g5318), .B(g13303), .Z(g15739) ) ;
AND2    gate18705  (.A(g5319), .B(g13304), .Z(g15740) ) ;
AND2    gate18706  (.A(g7542), .B(g12962), .Z(g15753) ) ;
AND2    gate18707  (.A(g7837), .B(g13308), .Z(g15754) ) ;
AND2    gate18708  (.A(g8178), .B(g13309), .Z(g15755) ) ;
AND2    gate18709  (.A(g5333), .B(g13324), .Z(g15765) ) ;
AND2    gate18710  (.A(g5341), .B(g13328), .Z(g15769) ) ;
AND2    gate18711  (.A(g5342), .B(g13329), .Z(g15770) ) ;
AND3    gate18712  (.A(g13004), .B(g3018), .C(g7549), .Z(II22028) ) ;
AND3    gate18713  (.A(g7471), .B(g3032), .C(II22028), .Z(g15780) ) ;
AND2    gate18714  (.A(g7971), .B(g13330), .Z(g15781) ) ;
AND2    gate18715  (.A(g5361), .B(g13347), .Z(g15793) ) ;
AND2    gate18716  (.A(g7856), .B(g13351), .Z(g15801) ) ;
AND2    gate18717  (.A(g8253), .B(g13352), .Z(g15802) ) ;
AND2    gate18718  (.A(g8025), .B(g13373), .Z(g15817) ) ;
AND2    gate18719  (.A(g7877), .B(g13398), .Z(g15828) ) ;
AND2    gate18720  (.A(g7857), .B(g13400), .Z(g15829) ) ;
AND2    gate18721  (.A(g8098), .B(g11620), .Z(g15840) ) ;
AND2    gate18722  (.A(g7878), .B(g11642), .Z(g15852) ) ;
AND3    gate18723  (.A(g13082), .B(g2912), .C(g7522), .Z(II22136) ) ;
AND3    gate18724  (.A(g7607), .B(g2920), .C(II22136), .Z(g15902) ) ;
AND2    gate18725  (.A(g5469), .B(g11732), .Z(g15998) ) ;
AND2    gate18726  (.A(g12013), .B(g10826), .Z(g16003) ) ;
AND2    gate18727  (.A(g5587), .B(g11734), .Z(g16004) ) ;
AND2    gate18728  (.A(g5504), .B(g11735), .Z(g16008) ) ;
AND2    gate18729  (.A(g12071), .B(g10843), .Z(g16009) ) ;
AND2    gate18730  (.A(g7639), .B(g11736), .Z(g16010) ) ;
AND2    gate18731  (.A(g12013), .B(g10859), .Z(g16015) ) ;
AND2    gate18732  (.A(g5601), .B(g11740), .Z(g16016) ) ;
AND2    gate18733  (.A(g12130), .B(g10862), .Z(g16017) ) ;
AND2    gate18734  (.A(g6149), .B(g11741), .Z(g16018) ) ;
AND2    gate18735  (.A(g5507), .B(g11742), .Z(g16019) ) ;
AND2    gate18736  (.A(g5543), .B(g11745), .Z(g16028) ) ;
AND2    gate18737  (.A(g12071), .B(g10877), .Z(g16029) ) ;
AND2    gate18738  (.A(g7667), .B(g11746), .Z(g16030) ) ;
AND2    gate18739  (.A(g6227), .B(g11747), .Z(g16031) ) ;
AND2    gate18740  (.A(g12187), .B(g10883), .Z(g16032) ) ;
AND2    gate18741  (.A(g5546), .B(g11748), .Z(g16033) ) ;
AND2    gate18742  (.A(g12013), .B(g10892), .Z(g16045) ) ;
AND2    gate18743  (.A(g5618), .B(g11761), .Z(g16046) ) ;
AND2    gate18744  (.A(g12130), .B(g10895), .Z(g16047) ) ;
AND2    gate18745  (.A(g6170), .B(g11762), .Z(g16048) ) ;
AND2    gate18746  (.A(g6638), .B(g11763), .Z(g16049) ) ;
AND2    gate18747  (.A(g5590), .B(g11764), .Z(g16050) ) ;
AND2    gate18748  (.A(g12235), .B(g10901), .Z(g16051) ) ;
AND2    gate18749  (.A(g5591), .B(g11765), .Z(g16052) ) ;
AND2    gate18750  (.A(g12071), .B(g10912), .Z(g16066) ) ;
AND2    gate18751  (.A(g7700), .B(g11774), .Z(g16067) ) ;
AND2    gate18752  (.A(g6310), .B(g11775), .Z(g16068) ) ;
AND2    gate18753  (.A(g5346), .B(g11776), .Z(g16069) ) ;
AND2    gate18754  (.A(g12187), .B(g10921), .Z(g16070) ) ;
AND2    gate18755  (.A(g5604), .B(g11777), .Z(g16071) ) ;
AND2    gate18756  (.A(g12275), .B(g10924), .Z(g16072) ) ;
AND2    gate18757  (.A(g5605), .B(g11778), .Z(g16073) ) ;
AND2    gate18758  (.A(g5646), .B(g11782), .Z(g16074) ) ;
AND2    gate18759  (.A(g984), .B(g11787), .Z(g16089) ) ;
AND2    gate18760  (.A(g12130), .B(g10937), .Z(g16100) ) ;
AND2    gate18761  (.A(g6197), .B(g11794), .Z(g16101) ) ;
AND2    gate18762  (.A(g6905), .B(g11795), .Z(g16102) ) ;
AND2    gate18763  (.A(g5621), .B(g11796), .Z(g16103) ) ;
AND2    gate18764  (.A(g12235), .B(g10946), .Z(g16104) ) ;
AND2    gate18765  (.A(g5622), .B(g11797), .Z(g16105) ) ;
AND2    gate18766  (.A(g12308), .B(g10949), .Z(g16106) ) ;
AND2    gate18767  (.A(g5666), .B(g11801), .Z(g16107) ) ;
AND2    gate18768  (.A(g5667), .B(g11802), .Z(g16108) ) ;
AND2    gate18769  (.A(g5551), .B(g13215), .Z(g16111) ) ;
AND2    gate18770  (.A(g5684), .B(g11808), .Z(g16112) ) ;
AND2    gate18771  (.A(g3460), .B(g11809), .Z(g16119) ) ;
AND2    gate18772  (.A(g1678), .B(g11813), .Z(g16127) ) ;
AND2    gate18773  (.A(g6444), .B(g11817), .Z(g16133) ) ;
AND2    gate18774  (.A(g5363), .B(g11818), .Z(g16134) ) ;
AND2    gate18775  (.A(g12187), .B(g10980), .Z(g16135) ) ;
AND2    gate18776  (.A(g5640), .B(g11819), .Z(g16136) ) ;
AND2    gate18777  (.A(g12275), .B(g10983), .Z(g16137) ) ;
AND2    gate18778  (.A(g5641), .B(g11820), .Z(g16138) ) ;
AND2    gate18779  (.A(g5704), .B(g11824), .Z(g16139) ) ;
AND2    gate18780  (.A(g5705), .B(g11825), .Z(g16140) ) ;
AND2    gate18781  (.A(g5706), .B(g11826), .Z(g16141) ) ;
AND2    gate18782  (.A(g5592), .B(g13229), .Z(g16153) ) ;
AND2    gate18783  (.A(g5718), .B(g11834), .Z(g16158) ) ;
AND2    gate18784  (.A(g5719), .B(g11835), .Z(g16159) ) ;
AND2    gate18785  (.A(g8286), .B(g11836), .Z(g16160) ) ;
AND2    gate18786  (.A(g1202), .B(g11837), .Z(g16161) ) ;
AND2    gate18787  (.A(g5597), .B(g13234), .Z(g16162) ) ;
AND2    gate18788  (.A(g5736), .B(g11841), .Z(g16163) ) ;
AND2    gate18789  (.A(g3616), .B(g11842), .Z(g16170) ) ;
AND2    gate18790  (.A(g2372), .B(g11846), .Z(g16178) ) ;
AND2    gate18791  (.A(g7149), .B(g11852), .Z(g16182) ) ;
AND2    gate18792  (.A(g12235), .B(g11014), .Z(g16183) ) ;
AND2    gate18793  (.A(g5663), .B(g11853), .Z(g16184) ) ;
AND2    gate18794  (.A(g12308), .B(g11017), .Z(g16185) ) ;
AND2    gate18795  (.A(g5753), .B(g11856), .Z(g16186) ) ;
AND2    gate18796  (.A(g5754), .B(g11857), .Z(g16187) ) ;
AND2    gate18797  (.A(g5755), .B(g11858), .Z(g16188) ) ;
AND2    gate18798  (.A(g5762), .B(g11866), .Z(g16198) ) ;
AND2    gate18799  (.A(g5763), .B(g11867), .Z(g16199) ) ;
AND2    gate18800  (.A(g5764), .B(g11868), .Z(g16200) ) ;
AND2    gate18801  (.A(g1203), .B(g11871), .Z(g16211) ) ;
AND2    gate18802  (.A(g5609), .B(g13252), .Z(g16212) ) ;
AND2    gate18803  (.A(g5776), .B(g11876), .Z(g16217) ) ;
AND2    gate18804  (.A(g5777), .B(g11877), .Z(g16218) ) ;
AND2    gate18805  (.A(g8295), .B(g11878), .Z(g16219) ) ;
AND2    gate18806  (.A(g1896), .B(g11879), .Z(g16220) ) ;
AND2    gate18807  (.A(g5614), .B(g13257), .Z(g16221) ) ;
AND2    gate18808  (.A(g5794), .B(g11883), .Z(g16222) ) ;
AND2    gate18809  (.A(g3772), .B(g11884), .Z(g16229) ) ;
AND2    gate18810  (.A(g5379), .B(g11886), .Z(g16237) ) ;
AND2    gate18811  (.A(g12275), .B(g11066), .Z(g16238) ) ;
AND2    gate18812  (.A(g5700), .B(g11887), .Z(g16239) ) ;
AND2    gate18813  (.A(g5804), .B(g11891), .Z(g16240) ) ;
AND2    gate18814  (.A(g5805), .B(g11892), .Z(g16241) ) ;
AND2    gate18815  (.A(g5806), .B(g11893), .Z(g16242) ) ;
AND2    gate18816  (.A(g5812), .B(g11898), .Z(g16251) ) ;
AND2    gate18817  (.A(g5813), .B(g11899), .Z(g16252) ) ;
AND2    gate18818  (.A(g5814), .B(g11900), .Z(g16253) ) ;
AND2    gate18819  (.A(g1204), .B(g11904), .Z(g16262) ) ;
AND2    gate18820  (.A(g5821), .B(g11908), .Z(g16263) ) ;
AND2    gate18821  (.A(g5822), .B(g11909), .Z(g16264) ) ;
AND2    gate18822  (.A(g5823), .B(g11910), .Z(g16265) ) ;
AND2    gate18823  (.A(g1897), .B(g11913), .Z(g16276) ) ;
AND2    gate18824  (.A(g5634), .B(g13275), .Z(g16277) ) ;
AND2    gate18825  (.A(g5835), .B(g11918), .Z(g16282) ) ;
AND2    gate18826  (.A(g5836), .B(g11919), .Z(g16283) ) ;
AND2    gate18827  (.A(g8304), .B(g11920), .Z(g16284) ) ;
AND2    gate18828  (.A(g2590), .B(g11921), .Z(g16285) ) ;
AND2    gate18829  (.A(g5639), .B(g13280), .Z(g16286) ) ;
AND2    gate18830  (.A(g12308), .B(g11129), .Z(g16288) ) ;
AND2    gate18831  (.A(g5853), .B(g11929), .Z(g16289) ) ;
AND2    gate18832  (.A(g5854), .B(g11930), .Z(g16290) ) ;
AND2    gate18833  (.A(g5855), .B(g11931), .Z(g16291) ) ;
AND2    gate18834  (.A(g520), .B(g11936), .Z(g16298) ) ;
AND2    gate18835  (.A(g5860), .B(g11941), .Z(g16299) ) ;
AND2    gate18836  (.A(g5861), .B(g11942), .Z(g16300) ) ;
AND2    gate18837  (.A(g5862), .B(g11943), .Z(g16301) ) ;
AND2    gate18838  (.A(g1205), .B(g11945), .Z(g16309) ) ;
AND2    gate18839  (.A(g5868), .B(g11948), .Z(g16310) ) ;
AND2    gate18840  (.A(g5869), .B(g11949), .Z(g16311) ) ;
AND2    gate18841  (.A(g5870), .B(g11950), .Z(g16312) ) ;
AND2    gate18842  (.A(g1898), .B(g11954), .Z(g16321) ) ;
AND2    gate18843  (.A(g5877), .B(g11958), .Z(g16322) ) ;
AND2    gate18844  (.A(g5878), .B(g11959), .Z(g16323) ) ;
AND2    gate18845  (.A(g5879), .B(g11960), .Z(g16324) ) ;
AND2    gate18846  (.A(g2591), .B(g11963), .Z(g16335) ) ;
AND2    gate18847  (.A(g5662), .B(g13300), .Z(g16336) ) ;
AND2    gate18848  (.A(g5894), .B(g11968), .Z(g16342) ) ;
AND2    gate18849  (.A(g5895), .B(g11969), .Z(g16343) ) ;
AND2    gate18850  (.A(g5896), .B(g11970), .Z(g16344) ) ;
AND2    gate18851  (.A(g5897), .B(g11971), .Z(g16345) ) ;
AND2    gate18852  (.A(g5900), .B(g11982), .Z(g16347) ) ;
AND2    gate18853  (.A(g5901), .B(g11983), .Z(g16348) ) ;
AND2    gate18854  (.A(g5902), .B(g11984), .Z(g16349) ) ;
AND2    gate18855  (.A(g981), .B(g11985), .Z(g16350) ) ;
AND2    gate18856  (.A(g1206), .B(g11989), .Z(g16356) ) ;
AND2    gate18857  (.A(g5907), .B(g11994), .Z(g16357) ) ;
AND2    gate18858  (.A(g5908), .B(g11995), .Z(g16358) ) ;
AND2    gate18859  (.A(g5909), .B(g11996), .Z(g16359) ) ;
AND2    gate18860  (.A(g1899), .B(g11998), .Z(g16367) ) ;
AND2    gate18861  (.A(g5915), .B(g12001), .Z(g16368) ) ;
AND2    gate18862  (.A(g5916), .B(g12002), .Z(g16369) ) ;
AND2    gate18863  (.A(g5917), .B(g12003), .Z(g16370) ) ;
AND2    gate18864  (.A(g2592), .B(g12007), .Z(g16379) ) ;
AND2    gate18865  (.A(g5925), .B(g12020), .Z(g16380) ) ;
AND2    gate18866  (.A(g5926), .B(g12021), .Z(g16381) ) ;
AND2    gate18867  (.A(g5927), .B(g12022), .Z(g16382) ) ;
AND2    gate18868  (.A(g5928), .B(g12023), .Z(g16383) ) ;
AND2    gate18869  (.A(g5714), .B(g13336), .Z(g16385) ) ;
AND2    gate18870  (.A(g5933), .B(g12037), .Z(g16386) ) ;
AND2    gate18871  (.A(g5934), .B(g12038), .Z(g16387) ) ;
AND2    gate18872  (.A(g5935), .B(g12039), .Z(g16388) ) ;
AND2    gate18873  (.A(g5936), .B(g12040), .Z(g16389) ) ;
AND2    gate18874  (.A(g982), .B(g12041), .Z(g16390) ) ;
AND2    gate18875  (.A(g5939), .B(g12051), .Z(g16391) ) ;
AND2    gate18876  (.A(g5940), .B(g12052), .Z(g16392) ) ;
AND2    gate18877  (.A(g5941), .B(g12053), .Z(g16393) ) ;
AND2    gate18878  (.A(g1675), .B(g12054), .Z(g16394) ) ;
AND2    gate18879  (.A(g1900), .B(g12058), .Z(g16400) ) ;
AND2    gate18880  (.A(g5946), .B(g12063), .Z(g16401) ) ;
AND2    gate18881  (.A(g5947), .B(g12064), .Z(g16402) ) ;
AND2    gate18882  (.A(g5948), .B(g12065), .Z(g16403) ) ;
AND2    gate18883  (.A(g2593), .B(g12067), .Z(g16411) ) ;
AND2    gate18884  (.A(g5954), .B(g12075), .Z(g16413) ) ;
AND2    gate18885  (.A(g5955), .B(g12076), .Z(g16414) ) ;
AND2    gate18886  (.A(g5956), .B(g12077), .Z(g16415) ) ;
AND2    gate18887  (.A(g5957), .B(g12078), .Z(g16416) ) ;
AND2    gate18888  (.A(g5759), .B(g13356), .Z(g16417) ) ;
AND2    gate18889  (.A(g5959), .B(g12084), .Z(g16418) ) ;
AND2    gate18890  (.A(g5960), .B(g12085), .Z(g16419) ) ;
AND2    gate18891  (.A(g5961), .B(g12086), .Z(g16420) ) ;
AND2    gate18892  (.A(g5962), .B(g12087), .Z(g16421) ) ;
AND2    gate18893  (.A(g983), .B(g12088), .Z(g16422) ) ;
AND2    gate18894  (.A(g5772), .B(g13361), .Z(g16423) ) ;
AND2    gate18895  (.A(g5967), .B(g12101), .Z(g16424) ) ;
AND2    gate18896  (.A(g5968), .B(g12102), .Z(g16425) ) ;
AND2    gate18897  (.A(g5969), .B(g12103), .Z(g16426) ) ;
AND2    gate18898  (.A(g5970), .B(g12104), .Z(g16427) ) ;
AND2    gate18899  (.A(g1676), .B(g12105), .Z(g16428) ) ;
AND2    gate18900  (.A(g5973), .B(g12115), .Z(g16429) ) ;
AND2    gate18901  (.A(g5974), .B(g12116), .Z(g16430) ) ;
AND2    gate18902  (.A(g5975), .B(g12117), .Z(g16431) ) ;
AND2    gate18903  (.A(g2369), .B(g12118), .Z(g16432) ) ;
AND2    gate18904  (.A(g2594), .B(g12122), .Z(g16438) ) ;
AND2    gate18905  (.A(g5980), .B(g12134), .Z(g16443) ) ;
AND2    gate18906  (.A(g5981), .B(g12135), .Z(g16444) ) ;
AND2    gate18907  (.A(g5808), .B(g13381), .Z(g16445) ) ;
AND2    gate18908  (.A(g5983), .B(g12147), .Z(g16447) ) ;
AND2    gate18909  (.A(g5984), .B(g12148), .Z(g16448) ) ;
AND2    gate18910  (.A(g5985), .B(g12149), .Z(g16449) ) ;
AND2    gate18911  (.A(g5986), .B(g12150), .Z(g16450) ) ;
AND2    gate18912  (.A(g5818), .B(g13386), .Z(g16451) ) ;
AND2    gate18913  (.A(g5988), .B(g12156), .Z(g16452) ) ;
AND2    gate18914  (.A(g5989), .B(g12157), .Z(g16453) ) ;
AND2    gate18915  (.A(g5990), .B(g12158), .Z(g16454) ) ;
AND2    gate18916  (.A(g5991), .B(g12159), .Z(g16455) ) ;
AND2    gate18917  (.A(g1677), .B(g12160), .Z(g16456) ) ;
AND2    gate18918  (.A(g5831), .B(g13391), .Z(g16457) ) ;
AND2    gate18919  (.A(g5996), .B(g12173), .Z(g16458) ) ;
AND2    gate18920  (.A(g5997), .B(g12174), .Z(g16459) ) ;
AND2    gate18921  (.A(g5998), .B(g12175), .Z(g16460) ) ;
AND2    gate18922  (.A(g5999), .B(g12176), .Z(g16461) ) ;
AND2    gate18923  (.A(g2370), .B(g12177), .Z(g16462) ) ;
AND4    gate18924  (.A(g14776), .B(g14797), .C(g16142), .D(g16243), .Z(g16505) ) ;
AND4    gate18925  (.A(g15065), .B(g13724), .C(g13764), .D(g13797), .Z(g16513) ) ;
AND4    gate18926  (.A(g14811), .B(g14849), .C(g16201), .D(g16302), .Z(g16527) ) ;
AND4    gate18927  (.A(g15161), .B(g13774), .C(g13805), .D(g13825), .Z(g16535) ) ;
AND4    gate18928  (.A(g14863), .B(g14922), .C(g16266), .D(g16360), .Z(g16558) ) ;
AND4    gate18929  (.A(g14936), .B(g15003), .C(g16325), .D(g16404), .Z(g16590) ) ;
AND2    gate18930  (.A(g15022), .B(g15096), .Z(g16607) ) ;
AND2    gate18931  (.A(g15118), .B(g15188), .Z(g16625) ) ;
AND2    gate18932  (.A(g15210), .B(g15274), .Z(g16639) ) ;
AND2    gate18933  (.A(g15296), .B(g15366), .Z(g16650) ) ;
AND2    gate18934  (.A(g6226), .B(g14764), .Z(g16850) ) ;
AND2    gate18935  (.A(g15722), .B(g8646), .Z(g16855) ) ;
AND2    gate18936  (.A(g6443), .B(g14794), .Z(g16856) ) ;
AND2    gate18937  (.A(g15762), .B(g8662), .Z(g16859) ) ;
AND2    gate18938  (.A(g15790), .B(g8681), .Z(g16864) ) ;
AND2    gate18939  (.A(g6896), .B(g14881), .Z(g16865) ) ;
AND2    gate18940  (.A(g15813), .B(g8693), .Z(g16879) ) ;
AND2    gate18941  (.A(g7156), .B(g14959), .Z(g16894) ) ;
AND2    gate18942  (.A(g7335), .B(g15017), .Z(g16907) ) ;
AND2    gate18943  (.A(g7838), .B(g15032), .Z(g16908) ) ;
AND2    gate18944  (.A(g6908), .B(g15033), .Z(g16909) ) ;
AND2    gate18945  (.A(g7352), .B(g15048), .Z(g16923) ) ;
AND2    gate18946  (.A(g7858), .B(g15128), .Z(g16938) ) ;
AND2    gate18947  (.A(g7158), .B(g15129), .Z(g16939) ) ;
AND2    gate18948  (.A(g7482), .B(g15144), .Z(g16953) ) ;
AND2    gate18949  (.A(g7520), .B(g15170), .Z(g16964) ) ;
AND2    gate18950  (.A(g7529), .B(g15174), .Z(g16966) ) ;
AND2    gate18951  (.A(g7827), .B(g15175), .Z(g16967) ) ;
AND2    gate18952  (.A(g6672), .B(g15176), .Z(g16968) ) ;
AND2    gate18953  (.A(g7888), .B(g15220), .Z(g16969) ) ;
AND2    gate18954  (.A(g7354), .B(g15221), .Z(g16970) ) ;
AND2    gate18955  (.A(g7538), .B(g15236), .Z(g16984) ) ;
AND2    gate18956  (.A(g7555), .B(g15260), .Z(g16987) ) ;
AND2    gate18957  (.A(g7842), .B(g15261), .Z(g16988) ) ;
AND2    gate18958  (.A(g6974), .B(g15262), .Z(g16989) ) ;
AND2    gate18959  (.A(g7912), .B(g15306), .Z(g16990) ) ;
AND2    gate18960  (.A(g7484), .B(g15307), .Z(g16991) ) ;
AND2    gate18961  (.A(g7576), .B(g15322), .Z(g16993) ) ;
AND2    gate18962  (.A(g7819), .B(g15323), .Z(g16994) ) ;
AND2    gate18963  (.A(g7578), .B(g15352), .Z(g16997) ) ;
AND2    gate18964  (.A(g7862), .B(g15353), .Z(g16998) ) ;
AND2    gate18965  (.A(g7224), .B(g15354), .Z(g16999) ) ;
AND3    gate18966  (.A(g3254), .B(g10694), .C(g14144), .Z(g17001) ) ;
AND2    gate18967  (.A(g7996), .B(g15390), .Z(g17015) ) ;
AND2    gate18968  (.A(g7590), .B(g15408), .Z(g17017) ) ;
AND2    gate18969  (.A(g7830), .B(g15409), .Z(g17018) ) ;
AND2    gate18970  (.A(g7592), .B(g15438), .Z(g17021) ) ;
AND2    gate18971  (.A(g7892), .B(g15439), .Z(g17022) ) ;
AND2    gate18972  (.A(g7420), .B(g15440), .Z(g17023) ) ;
AND2    gate18973  (.A(g7604), .B(g15458), .Z(g17028) ) ;
AND3    gate18974  (.A(g3410), .B(g10714), .C(g14259), .Z(g17031) ) ;
AND2    gate18975  (.A(g8071), .B(g15474), .Z(g17045) ) ;
AND2    gate18976  (.A(g7605), .B(g15492), .Z(g17047) ) ;
AND2    gate18977  (.A(g7845), .B(g15493), .Z(g17048) ) ;
AND2    gate18978  (.A(g7153), .B(g15524), .Z(g17055) ) ;
AND2    gate18979  (.A(g7953), .B(g15525), .Z(g17056) ) ;
AND2    gate18980  (.A(g7613), .B(g15544), .Z(g17062) ) ;
AND3    gate18981  (.A(g3566), .B(g10735), .C(g14381), .Z(g17065) ) ;
AND2    gate18982  (.A(g8156), .B(g15560), .Z(g17079) ) ;
AND2    gate18983  (.A(g7614), .B(g15578), .Z(g17081) ) ;
AND2    gate18984  (.A(g7865), .B(g15579), .Z(g17082) ) ;
AND2    gate18985  (.A(g7629), .B(g13954), .Z(g17084) ) ;
AND2    gate18986  (.A(g7349), .B(g15602), .Z(g17090) ) ;
AND2    gate18987  (.A(g8004), .B(g15603), .Z(g17091) ) ;
AND2    gate18988  (.A(g7622), .B(g15622), .Z(g17097) ) ;
AND3    gate18989  (.A(g3722), .B(g10754), .C(g14493), .Z(g17100) ) ;
AND2    gate18990  (.A(g8242), .B(g15638), .Z(g17114) ) ;
AND2    gate18991  (.A(g7649), .B(g14008), .Z(g17116) ) ;
AND2    gate18992  (.A(g7906), .B(g15665), .Z(g17117) ) ;
AND2    gate18993  (.A(g7658), .B(g14024), .Z(g17122) ) ;
AND2    gate18994  (.A(g7479), .B(g15678), .Z(g17128) ) ;
AND2    gate18995  (.A(g8079), .B(g15679), .Z(g17129) ) ;
AND2    gate18996  (.A(g7638), .B(g15698), .Z(g17135) ) ;
AND2    gate18997  (.A(g7676), .B(g14068), .Z(g17138) ) ;
AND2    gate18998  (.A(g7685), .B(g14099), .Z(g17143) ) ;
AND2    gate18999  (.A(g7958), .B(g15724), .Z(g17144) ) ;
AND2    gate19000  (.A(g7694), .B(g14115), .Z(g17149) ) ;
AND2    gate19001  (.A(g7535), .B(g15737), .Z(g17155) ) ;
AND2    gate19002  (.A(g8164), .B(g15738), .Z(g17156) ) ;
AND2    gate19003  (.A(g7712), .B(g14183), .Z(g17161) ) ;
AND2    gate19004  (.A(g7721), .B(g14214), .Z(g17166) ) ;
AND2    gate19005  (.A(g8009), .B(g15764), .Z(g17167) ) ;
AND2    gate19006  (.A(g7730), .B(g14230), .Z(g17172) ) ;
AND2    gate19007  (.A(g7742), .B(g14298), .Z(g17176) ) ;
AND2    gate19008  (.A(g7751), .B(g14329), .Z(g17181) ) ;
AND2    gate19009  (.A(g8084), .B(g15792), .Z(g17182) ) ;
AND2    gate19010  (.A(g7766), .B(g14420), .Z(g17193) ) ;
AND2    gate19011  (.A(g8024), .B(g15991), .Z(g17268) ) ;
AND2    gate19012  (.A(g8097), .B(g15994), .Z(g17301) ) ;
AND2    gate19013  (.A(g8176), .B(g15997), .Z(g17339) ) ;
AND2    gate19014  (.A(g3942), .B(g14960), .Z(g17352) ) ;
AND2    gate19015  (.A(g3945), .B(g14963), .Z(g17353) ) ;
AND2    gate19016  (.A(g8250), .B(g16001), .Z(g17381) ) ;
AND2    gate19017  (.A(g8252), .B(g16002), .Z(g17382) ) ;
AND2    gate19018  (.A(g3941), .B(g16005), .Z(g17393) ) ;
AND2    gate19019  (.A(g6177), .B(g15034), .Z(g17395) ) ;
AND2    gate19020  (.A(g4020), .B(g15037), .Z(g17396) ) ;
AND2    gate19021  (.A(g4023), .B(g15040), .Z(g17397) ) ;
AND2    gate19022  (.A(g4026), .B(g15043), .Z(g17398) ) ;
AND2    gate19023  (.A(g4049), .B(g15049), .Z(g17408) ) ;
AND2    gate19024  (.A(g4052), .B(g15052), .Z(g17409) ) ;
AND2    gate19025  (.A(g3994), .B(g16007), .Z(g17428) ) ;
AND2    gate19026  (.A(g6284), .B(g16011), .Z(g17446) ) ;
AND2    gate19027  (.A(g4115), .B(g15106), .Z(g17447) ) ;
AND2    gate19028  (.A(g4118), .B(g15109), .Z(g17448) ) ;
AND2    gate19029  (.A(g4121), .B(g15112), .Z(g17449) ) ;
AND2    gate19030  (.A(g4124), .B(g15115), .Z(g17450) ) ;
AND2    gate19031  (.A(g4048), .B(g16012), .Z(g17460) ) ;
AND2    gate19032  (.A(g6209), .B(g15130), .Z(g17461) ) ;
AND2    gate19033  (.A(g4147), .B(g15133), .Z(g17462) ) ;
AND2    gate19034  (.A(g4150), .B(g15136), .Z(g17463) ) ;
AND2    gate19035  (.A(g4153), .B(g15139), .Z(g17464) ) ;
AND2    gate19036  (.A(g4176), .B(g15145), .Z(g17474) ) ;
AND2    gate19037  (.A(g4179), .B(g15148), .Z(g17475) ) ;
AND2    gate19038  (.A(g4089), .B(g16013), .Z(g17485) ) ;
AND2    gate19039  (.A(g4091), .B(g16014), .Z(g17486) ) ;
AND2    gate19040  (.A(g6675), .B(g16023), .Z(g17506) ) ;
AND2    gate19041  (.A(g4225), .B(g15179), .Z(g17508) ) ;
AND2    gate19042  (.A(g4228), .B(g15182), .Z(g17509) ) ;
AND2    gate19043  (.A(g4231), .B(g15185), .Z(g17510) ) ;
AND2    gate19044  (.A(g6421), .B(g16025), .Z(g17526) ) ;
AND2    gate19045  (.A(g4254), .B(g15198), .Z(g17527) ) ;
AND2    gate19046  (.A(g4257), .B(g15201), .Z(g17528) ) ;
AND2    gate19047  (.A(g4260), .B(g15204), .Z(g17529) ) ;
AND2    gate19048  (.A(g4263), .B(g15207), .Z(g17530) ) ;
AND2    gate19049  (.A(g4175), .B(g16026), .Z(g17540) ) ;
AND2    gate19050  (.A(g6298), .B(g15222), .Z(g17541) ) ;
AND2    gate19051  (.A(g4286), .B(g15225), .Z(g17542) ) ;
AND2    gate19052  (.A(g4289), .B(g15228), .Z(g17543) ) ;
AND2    gate19053  (.A(g4292), .B(g15231), .Z(g17544) ) ;
AND2    gate19054  (.A(g4315), .B(g15237), .Z(g17554) ) ;
AND2    gate19055  (.A(g4318), .B(g15240), .Z(g17555) ) ;
AND2    gate19056  (.A(g4201), .B(g16027), .Z(g17556) ) ;
AND2    gate19057  (.A(g4348), .B(g15248), .Z(g17576) ) ;
AND2    gate19058  (.A(g4351), .B(g15251), .Z(g17577) ) ;
AND2    gate19059  (.A(g4354), .B(g15254), .Z(g17578) ) ;
AND2    gate19060  (.A(g6977), .B(g16039), .Z(g17597) ) ;
AND2    gate19061  (.A(g4380), .B(g15265), .Z(g17598) ) ;
AND2    gate19062  (.A(g4383), .B(g15268), .Z(g17599) ) ;
AND2    gate19063  (.A(g4386), .B(g15271), .Z(g17600) ) ;
AND2    gate19064  (.A(g6626), .B(g16041), .Z(g17616) ) ;
AND2    gate19065  (.A(g4409), .B(g15284), .Z(g17617) ) ;
AND2    gate19066  (.A(g4412), .B(g15287), .Z(g17618) ) ;
AND2    gate19067  (.A(g4415), .B(g15290), .Z(g17619) ) ;
AND2    gate19068  (.A(g4418), .B(g15293), .Z(g17620) ) ;
AND2    gate19069  (.A(g4314), .B(g16042), .Z(g17630) ) ;
AND2    gate19070  (.A(g6435), .B(g15308), .Z(g17631) ) ;
AND2    gate19071  (.A(g4441), .B(g15311), .Z(g17632) ) ;
AND2    gate19072  (.A(g4444), .B(g15314), .Z(g17633) ) ;
AND2    gate19073  (.A(g4447), .B(g15317), .Z(g17634) ) ;
AND2    gate19074  (.A(g4322), .B(g16043), .Z(g17635) ) ;
AND2    gate19075  (.A(g4324), .B(g16044), .Z(g17636) ) ;
AND2    gate19076  (.A(g4480), .B(g15326), .Z(g17652) ) ;
AND2    gate19077  (.A(g4483), .B(g15329), .Z(g17653) ) ;
AND2    gate19078  (.A(g4486), .B(g15332), .Z(g17654) ) ;
AND2    gate19079  (.A(g4517), .B(g15340), .Z(g17673) ) ;
AND2    gate19080  (.A(g4520), .B(g15343), .Z(g17674) ) ;
AND2    gate19081  (.A(g4523), .B(g15346), .Z(g17675) ) ;
AND2    gate19082  (.A(g7227), .B(g16061), .Z(g17694) ) ;
AND2    gate19083  (.A(g4549), .B(g15357), .Z(g17695) ) ;
AND2    gate19084  (.A(g4552), .B(g15360), .Z(g17696) ) ;
AND2    gate19085  (.A(g4555), .B(g15363), .Z(g17697) ) ;
AND2    gate19086  (.A(g6890), .B(g16063), .Z(g17713) ) ;
AND2    gate19087  (.A(g4578), .B(g15376), .Z(g17714) ) ;
AND2    gate19088  (.A(g4581), .B(g15379), .Z(g17715) ) ;
AND2    gate19089  (.A(g4584), .B(g15382), .Z(g17716) ) ;
AND2    gate19090  (.A(g4587), .B(g15385), .Z(g17717) ) ;
AND2    gate19091  (.A(g4451), .B(g16064), .Z(g17718) ) ;
AND2    gate19092  (.A(g2993), .B(g16065), .Z(g17719) ) ;
AND2    gate19093  (.A(g4611), .B(g15393), .Z(g17734) ) ;
AND2    gate19094  (.A(g4614), .B(g15396), .Z(g17735) ) ;
AND2    gate19095  (.A(g4617), .B(g15399), .Z(g17736) ) ;
AND2    gate19096  (.A(g4626), .B(g15404), .Z(g17737) ) ;
AND2    gate19097  (.A(g4656), .B(g15412), .Z(g17752) ) ;
AND2    gate19098  (.A(g4659), .B(g15415), .Z(g17753) ) ;
AND2    gate19099  (.A(g4662), .B(g15418), .Z(g17754) ) ;
AND2    gate19100  (.A(g4693), .B(g15426), .Z(g17773) ) ;
AND2    gate19101  (.A(g4696), .B(g15429), .Z(g17774) ) ;
AND2    gate19102  (.A(g4699), .B(g15432), .Z(g17775) ) ;
AND2    gate19103  (.A(g7423), .B(g16097), .Z(g17794) ) ;
AND2    gate19104  (.A(g4725), .B(g15443), .Z(g17795) ) ;
AND2    gate19105  (.A(g4728), .B(g15446), .Z(g17796) ) ;
AND2    gate19106  (.A(g4731), .B(g15449), .Z(g17797) ) ;
AND2    gate19107  (.A(g4591), .B(g16099), .Z(g17798) ) ;
AND2    gate19108  (.A(g4754), .B(g15461), .Z(g17812) ) ;
AND2    gate19109  (.A(g4757), .B(g15464), .Z(g17813) ) ;
AND2    gate19110  (.A(g4760), .B(g15467), .Z(g17814) ) ;
AND2    gate19111  (.A(g4766), .B(g15471), .Z(g17824) ) ;
AND2    gate19112  (.A(g4788), .B(g15477), .Z(g17835) ) ;
AND2    gate19113  (.A(g4791), .B(g15480), .Z(g17836) ) ;
AND2    gate19114  (.A(g4794), .B(g15483), .Z(g17837) ) ;
AND2    gate19115  (.A(g4803), .B(g15488), .Z(g17838) ) ;
AND2    gate19116  (.A(g4833), .B(g15496), .Z(g17853) ) ;
AND2    gate19117  (.A(g4836), .B(g15499), .Z(g17854) ) ;
AND2    gate19118  (.A(g4839), .B(g15502), .Z(g17855) ) ;
AND2    gate19119  (.A(g4870), .B(g15510), .Z(g17874) ) ;
AND2    gate19120  (.A(g4873), .B(g15513), .Z(g17875) ) ;
AND2    gate19121  (.A(g4876), .B(g15516), .Z(g17876) ) ;
AND2    gate19122  (.A(g2998), .B(g15521), .Z(g17877) ) ;
AND2    gate19123  (.A(g4899), .B(g15528), .Z(g17900) ) ;
AND2    gate19124  (.A(g4902), .B(g15531), .Z(g17901) ) ;
AND2    gate19125  (.A(g4905), .B(g15534), .Z(g17902) ) ;
AND2    gate19126  (.A(g4908), .B(g15537), .Z(g17912) ) ;
AND2    gate19127  (.A(g4930), .B(g15547), .Z(g17924) ) ;
AND2    gate19128  (.A(g4933), .B(g15550), .Z(g17925) ) ;
AND2    gate19129  (.A(g4936), .B(g15553), .Z(g17926) ) ;
AND2    gate19130  (.A(g4942), .B(g15557), .Z(g17936) ) ;
AND2    gate19131  (.A(g4964), .B(g15563), .Z(g17947) ) ;
AND2    gate19132  (.A(g4967), .B(g15566), .Z(g17948) ) ;
AND2    gate19133  (.A(g4970), .B(g15569), .Z(g17949) ) ;
AND2    gate19134  (.A(g4979), .B(g15574), .Z(g17950) ) ;
AND2    gate19135  (.A(g5009), .B(g15582), .Z(g17965) ) ;
AND2    gate19136  (.A(g5012), .B(g15585), .Z(g17966) ) ;
AND2    gate19137  (.A(g5015), .B(g15588), .Z(g17967) ) ;
AND2    gate19138  (.A(g5035), .B(g15596), .Z(g17989) ) ;
AND2    gate19139  (.A(g5038), .B(g15599), .Z(g17990) ) ;
AND2    gate19140  (.A(g5058), .B(g15606), .Z(g18011) ) ;
AND2    gate19141  (.A(g5061), .B(g15609), .Z(g18012) ) ;
AND2    gate19142  (.A(g5064), .B(g15612), .Z(g18013) ) ;
AND2    gate19143  (.A(g5067), .B(g15615), .Z(g18023) ) ;
AND2    gate19144  (.A(g5089), .B(g15625), .Z(g18035) ) ;
AND2    gate19145  (.A(g5092), .B(g15628), .Z(g18036) ) ;
AND2    gate19146  (.A(g5095), .B(g15631), .Z(g18037) ) ;
AND2    gate19147  (.A(g5101), .B(g15635), .Z(g18047) ) ;
AND2    gate19148  (.A(g5123), .B(g15641), .Z(g18058) ) ;
AND2    gate19149  (.A(g5126), .B(g15644), .Z(g18059) ) ;
AND2    gate19150  (.A(g5129), .B(g15647), .Z(g18060) ) ;
AND2    gate19151  (.A(g5138), .B(g15652), .Z(g18061) ) ;
AND2    gate19152  (.A(g7462), .B(g15655), .Z(g18062) ) ;
AND2    gate19153  (.A(g5150), .B(g15667), .Z(g18088) ) ;
AND2    gate19154  (.A(g5164), .B(g15672), .Z(g18106) ) ;
AND2    gate19155  (.A(g5167), .B(g15675), .Z(g18107) ) ;
AND2    gate19156  (.A(g5187), .B(g15682), .Z(g18128) ) ;
AND2    gate19157  (.A(g5190), .B(g15685), .Z(g18129) ) ;
AND2    gate19158  (.A(g5193), .B(g15688), .Z(g18130) ) ;
AND2    gate19159  (.A(g5196), .B(g15691), .Z(g18140) ) ;
AND2    gate19160  (.A(g5218), .B(g15701), .Z(g18152) ) ;
AND2    gate19161  (.A(g5221), .B(g15704), .Z(g18153) ) ;
AND2    gate19162  (.A(g5224), .B(g15707), .Z(g18154) ) ;
AND2    gate19163  (.A(g5230), .B(g15711), .Z(g18164) ) ;
AND2    gate19164  (.A(g2883), .B(g16287), .Z(g18165) ) ;
AND2    gate19165  (.A(g7527), .B(g15714), .Z(g18169) ) ;
AND2    gate19166  (.A(g5243), .B(g15726), .Z(g18204) ) ;
AND2    gate19167  (.A(g5257), .B(g15731), .Z(g18222) ) ;
AND2    gate19168  (.A(g5260), .B(g15734), .Z(g18223) ) ;
AND2    gate19169  (.A(g5280), .B(g15741), .Z(g18244) ) ;
AND2    gate19170  (.A(g5283), .B(g15744), .Z(g18245) ) ;
AND2    gate19171  (.A(g5286), .B(g15747), .Z(g18246) ) ;
AND2    gate19172  (.A(g5289), .B(g15750), .Z(g18256) ) ;
AND2    gate19173  (.A(g5306), .B(g15766), .Z(g18311) ) ;
AND2    gate19174  (.A(g5320), .B(g15771), .Z(g18329) ) ;
AND2    gate19175  (.A(g5323), .B(g15774), .Z(g18330) ) ;
AND2    gate19176  (.A(g2888), .B(g15777), .Z(g18333) ) ;
AND2    gate19177  (.A(g5343), .B(g15794), .Z(g18404) ) ;
AND3    gate19178  (.A(g14776), .B(g14837), .C(g16142), .Z(II24619) ) ;
AND3    gate19179  (.A(g13677), .B(g13750), .C(II24619), .Z(g18547) ) ;
AND3    gate19180  (.A(g14811), .B(g14910), .C(g16201), .Z(II24689) ) ;
AND3    gate19181  (.A(g13714), .B(g13791), .C(II24689), .Z(g18597) ) ;
AND3    gate19182  (.A(g14863), .B(g14991), .C(g16266), .Z(II24738) ) ;
AND3    gate19183  (.A(g13764), .B(g13819), .C(II24738), .Z(g18629) ) ;
AND3    gate19184  (.A(g14936), .B(g15080), .C(g16325), .Z(II24758) ) ;
AND3    gate19185  (.A(g13805), .B(g13840), .C(II24758), .Z(g18638) ) ;
AND4    gate19186  (.A(g14776), .B(g14895), .C(g16142), .D(g13750), .Z(g18645) ) ;
AND3    gate19187  (.A(g14895), .B(g16142), .C(g16243), .Z(g18647) ) ;
AND4    gate19188  (.A(g14811), .B(g14976), .C(g16201), .D(g13791), .Z(g18648) ) ;
AND4    gate19189  (.A(g14776), .B(g14837), .C(g13657), .D(g16189), .Z(g18649) ) ;
AND3    gate19190  (.A(g14976), .B(g16201), .C(g16302), .Z(g18650) ) ;
AND4    gate19191  (.A(g14863), .B(g15065), .C(g16266), .D(g13819), .Z(g18651) ) ;
AND4    gate19192  (.A(g14797), .B(g13657), .C(g13677), .D(g16243), .Z(g18652) ) ;
AND4    gate19193  (.A(g14811), .B(g14910), .C(g13687), .D(g16254), .Z(g18653) ) ;
AND3    gate19194  (.A(g15065), .B(g16266), .C(g16360), .Z(g18654) ) ;
AND4    gate19195  (.A(g14936), .B(g15161), .C(g16325), .D(g13840), .Z(g18655) ) ;
AND4    gate19196  (.A(g14776), .B(g14837), .C(g16189), .D(g13706), .Z(g18665) ) ;
AND4    gate19197  (.A(g14849), .B(g13687), .C(g13714), .D(g16302), .Z(g18666) ) ;
AND4    gate19198  (.A(g14863), .B(g14991), .C(g13724), .D(g16313), .Z(g18667) ) ;
AND3    gate19199  (.A(g15161), .B(g16325), .C(g16404), .Z(g18668) ) ;
AND4    gate19200  (.A(g14811), .B(g14910), .C(g16254), .D(g13756), .Z(g18688) ) ;
AND4    gate19201  (.A(g14922), .B(g13724), .C(g13764), .D(g16360), .Z(g18689) ) ;
AND4    gate19202  (.A(g14936), .B(g15080), .C(g13774), .D(g16371), .Z(g18690) ) ;
AND4    gate19203  (.A(g14863), .B(g14991), .C(g16313), .D(g13797), .Z(g18717) ) ;
AND4    gate19204  (.A(g15003), .B(g13774), .C(g13805), .D(g16404), .Z(g18718) ) ;
AND4    gate19205  (.A(g14936), .B(g15080), .C(g16371), .D(g13825), .Z(g18753) ) ;
AND2    gate19206  (.A(g13519), .B(g16154), .Z(g18982) ) ;
AND2    gate19207  (.A(g13530), .B(g16213), .Z(g18990) ) ;
AND4    gate19208  (.A(g14895), .B(g13657), .C(g13677), .D(g13706), .Z(g18994) ) ;
AND2    gate19209  (.A(g13541), .B(g16278), .Z(g18997) ) ;
AND4    gate19210  (.A(g14976), .B(g13687), .C(g13714), .D(g13756), .Z(g19007) ) ;
AND2    gate19211  (.A(g13552), .B(g16337), .Z(g19010) ) ;
AND4    gate19212  (.A(g18679), .B(g14910), .C(g13687), .D(g16254), .Z(g19063) ) ;
AND4    gate19213  (.A(g14797), .B(g18692), .C(g16142), .D(g16189), .Z(g19079) ) ;
AND4    gate19214  (.A(g18708), .B(g14991), .C(g13724), .D(g16313), .Z(g19080) ) ;
NOR2    gate19215  (.A(g15904), .B(g14642), .Z(g17215) ) ;
AND2    gate19216  (.A(g17215), .B(g16540), .Z(g19087) ) ;
AND4    gate19217  (.A(g18656), .B(g14797), .C(g16189), .D(g13706), .Z(g19088) ) ;
AND4    gate19218  (.A(g14849), .B(g18728), .C(g16201), .D(g16254), .Z(g19089) ) ;
AND4    gate19219  (.A(g18744), .B(g15080), .C(g13774), .D(g16371), .Z(g19090) ) ;
AND4    gate19220  (.A(g14776), .B(g18670), .C(g18692), .D(g16293), .Z(g19092) ) ;
NOR2    gate19221  (.A(g15933), .B(g14669), .Z(g17218) ) ;
AND2    gate19222  (.A(g17218), .B(g16572), .Z(g19093) ) ;
AND4    gate19223  (.A(g18679), .B(g14849), .C(g16254), .D(g13756), .Z(g19094) ) ;
AND4    gate19224  (.A(g14922), .B(g18765), .C(g16266), .D(g16313), .Z(g19095) ) ;
AND3    gate19225  (.A(g18656), .B(g18670), .C(g18720), .Z(II25280) ) ;
AND3    gate19226  (.A(g13657), .B(g16243), .C(II25280), .Z(g19097) ) ;
AND4    gate19227  (.A(g14811), .B(g18699), .C(g18728), .D(g16351), .Z(g19099) ) ;
NOR2    gate19228  (.A(g15962), .B(g14703), .Z(g17220) ) ;
AND2    gate19229  (.A(g17220), .B(g16596), .Z(g19100) ) ;
AND4    gate19230  (.A(g18708), .B(g14922), .C(g16313), .D(g13797), .Z(g19101) ) ;
AND4    gate19231  (.A(g15003), .B(g18796), .C(g16325), .D(g16371), .Z(g19102) ) ;
AND3    gate19232  (.A(g18679), .B(g18699), .C(g18758), .Z(II25291) ) ;
AND3    gate19233  (.A(g13687), .B(g16302), .C(II25291), .Z(g19104) ) ;
AND4    gate19234  (.A(g14863), .B(g18735), .C(g18765), .D(g16395), .Z(g19106) ) ;
NOR2    gate19235  (.A(g15981), .B(g14737), .Z(g17223) ) ;
AND2    gate19236  (.A(g17223), .B(g16616), .Z(g19107) ) ;
AND4    gate19237  (.A(g18744), .B(g15003), .C(g16371), .D(g13825), .Z(g19108) ) ;
AND3    gate19238  (.A(g18708), .B(g18735), .C(g18789), .Z(II25300) ) ;
AND3    gate19239  (.A(g13724), .B(g16360), .C(II25300), .Z(g19109) ) ;
AND4    gate19240  (.A(g14936), .B(g18772), .C(g18796), .D(g16433), .Z(g19111) ) ;
AND2    gate19241  (.A(g14657), .B(g16633), .Z(g19112) ) ;
AND3    gate19242  (.A(g18744), .B(g18772), .C(g18815), .Z(II25311) ) ;
AND3    gate19243  (.A(g13774), .B(g16404), .C(II25311), .Z(g19116) ) ;
AND2    gate19244  (.A(g14691), .B(g16644), .Z(g19117) ) ;
AND2    gate19245  (.A(g14725), .B(g16656), .Z(g19124) ) ;
AND2    gate19246  (.A(g14753), .B(g16673), .Z(g19131) ) ;
NAND2   gate19247  (.A(g14642), .B(g14657), .Z(g17159) ) ;
AND2    gate19248  (.A(g17159), .B(g16719), .Z(g19142) ) ;
NAND2   gate19249  (.A(g14669), .B(g14691), .Z(g17174) ) ;
AND2    gate19250  (.A(g17174), .B(g16761), .Z(g19143) ) ;
NAND2   gate19251  (.A(g14703), .B(g14725), .Z(g17191) ) ;
AND2    gate19252  (.A(g17191), .B(g16788), .Z(g19146) ) ;
NAND2   gate19253  (.A(g14737), .B(g14753), .Z(g17202) ) ;
AND2    gate19254  (.A(g17202), .B(g16817), .Z(g19148) ) ;
AND2    gate19255  (.A(g17189), .B(g8602), .Z(g19150) ) ;
AND2    gate19256  (.A(g17200), .B(g8614), .Z(g19155) ) ;
AND2    gate19257  (.A(g17207), .B(g8627), .Z(g19161) ) ;
AND2    gate19258  (.A(g17212), .B(g8637), .Z(g19166) ) ;
NAND2   gate19259  (.A(II22706), .B(II22707), .Z(g16662) ) ;
AND2    gate19260  (.A(g16662), .B(g12125), .Z(g19228) ) ;
NAND2   gate19261  (.A(II22885), .B(II22886), .Z(g16935) ) ;
AND2    gate19262  (.A(g16935), .B(g8802), .Z(g19236) ) ;
AND3    gate19263  (.A(g16867), .B(g14158), .C(g14071), .Z(g19241) ) ;
AND2    gate19264  (.A(g16662), .B(g8817), .Z(g19248) ) ;
AND2    gate19265  (.A(g18725), .B(g9527), .Z(g19252) ) ;
AND3    gate19266  (.A(g16895), .B(g14273), .C(g14186), .Z(g19254) ) ;
AND2    gate19267  (.A(g16749), .B(g3124), .Z(g19260) ) ;
AND3    gate19268  (.A(g16924), .B(g14395), .C(g14301), .Z(g19267) ) ;
AND3    gate19269  (.A(g16954), .B(g14507), .C(g14423), .Z(g19282) ) ;
AND2    gate19270  (.A(g18063), .B(g3111), .Z(g19284) ) ;
AND2    gate19271  (.A(g16749), .B(g7642), .Z(g19285) ) ;
AND2    gate19272  (.A(g17029), .B(g8580), .Z(g19289) ) ;
AND3    gate19273  (.A(g16867), .B(g16543), .C(g14071), .Z(g19303) ) ;
AND2    gate19274  (.A(g17063), .B(g8587), .Z(g19307) ) ;
AND2    gate19275  (.A(g18063), .B(g3110), .Z(g19316) ) ;
AND2    gate19276  (.A(g16749), .B(g3126), .Z(g19317) ) ;
AND3    gate19277  (.A(g16867), .B(g16515), .C(g14158), .Z(g19320) ) ;
AND3    gate19278  (.A(g16895), .B(g16575), .C(g14186), .Z(g19324) ) ;
AND2    gate19279  (.A(g17098), .B(g8594), .Z(g19328) ) ;
AND3    gate19280  (.A(g16895), .B(g16546), .C(g14273), .Z(g19347) ) ;
AND3    gate19281  (.A(g16924), .B(g16599), .C(g14301), .Z(g19351) ) ;
AND2    gate19282  (.A(g17136), .B(g8605), .Z(g19355) ) ;
AND2    gate19283  (.A(g18063), .B(g3112), .Z(g19356) ) ;
AND3    gate19284  (.A(g16924), .B(g16578), .C(g14395), .Z(g19381) ) ;
AND3    gate19285  (.A(g16954), .B(g16619), .C(g14423), .Z(g19385) ) ;
AND3    gate19286  (.A(g16954), .B(g16602), .C(g14507), .Z(g19413) ) ;
AND3    gate19287  (.A(g16884), .B(g14797), .C(g14776), .Z(g19449) ) ;
AND3    gate19288  (.A(g16913), .B(g14849), .C(g14811), .Z(g19476) ) ;
AND3    gate19289  (.A(g16943), .B(g14922), .C(g14863), .Z(g19499) ) ;
AND3    gate19290  (.A(g16974), .B(g15003), .C(g14936), .Z(g19520) ) ;
AND3    gate19291  (.A(g16884), .B(g16722), .C(g14776), .Z(g19531) ) ;
AND3    gate19292  (.A(g16884), .B(g16697), .C(g14797), .Z(g19540) ) ;
AND3    gate19293  (.A(g16913), .B(g16764), .C(g14811), .Z(g19541) ) ;
AND3    gate19294  (.A(g16913), .B(g16728), .C(g14849), .Z(g19544) ) ;
AND3    gate19295  (.A(g16943), .B(g16791), .C(g14863), .Z(g19545) ) ;
AND3    gate19296  (.A(g16943), .B(g16770), .C(g14922), .Z(g19547) ) ;
AND3    gate19297  (.A(g16974), .B(g16820), .C(g14936), .Z(g19548) ) ;
AND2    gate19298  (.A(g7950), .B(g17230), .Z(g19549) ) ;
AND3    gate19299  (.A(g16974), .B(g16797), .C(g15003), .Z(g19551) ) ;
NOR2    gate19300  (.A(g14956), .B(g12564), .Z(g16829) ) ;
AND2    gate19301  (.A(g16829), .B(g6048), .Z(g19552) ) ;
AND2    gate19302  (.A(g7990), .B(g17237), .Z(g19553) ) ;
AND2    gate19303  (.A(g7993), .B(g17240), .Z(g19554) ) ;
AND2    gate19304  (.A(g8001), .B(g17243), .Z(g19555) ) ;
AND2    gate19305  (.A(g8053), .B(g17249), .Z(g19557) ) ;
AND2    gate19306  (.A(g8056), .B(g17252), .Z(g19558) ) ;
AND2    gate19307  (.A(g8059), .B(g17255), .Z(g19559) ) ;
AND2    gate19308  (.A(g8065), .B(g17259), .Z(g19560) ) ;
AND2    gate19309  (.A(g8068), .B(g17262), .Z(g19561) ) ;
AND2    gate19310  (.A(g8076), .B(g17265), .Z(g19562) ) ;
AND2    gate19311  (.A(g8123), .B(g17272), .Z(g19564) ) ;
AND2    gate19312  (.A(g8126), .B(g17275), .Z(g19565) ) ;
AND2    gate19313  (.A(g8129), .B(g17278), .Z(g19566) ) ;
AND2    gate19314  (.A(g8138), .B(g17282), .Z(g19567) ) ;
AND2    gate19315  (.A(g8141), .B(g17285), .Z(g19568) ) ;
AND2    gate19316  (.A(g8144), .B(g17288), .Z(g19569) ) ;
AND2    gate19317  (.A(g8150), .B(g17291), .Z(g19570) ) ;
AND2    gate19318  (.A(g8153), .B(g17294), .Z(g19571) ) ;
AND2    gate19319  (.A(g8161), .B(g17297), .Z(g19572) ) ;
AND2    gate19320  (.A(g8191), .B(g17304), .Z(g19574) ) ;
AND2    gate19321  (.A(g8194), .B(g17307), .Z(g19575) ) ;
AND2    gate19322  (.A(g8197), .B(g17310), .Z(g19576) ) ;
AND2    gate19323  (.A(g640), .B(g18756), .Z(g19584) ) ;
AND2    gate19324  (.A(g692), .B(g18757), .Z(g19585) ) ;
AND2    gate19325  (.A(g8209), .B(g17315), .Z(g19586) ) ;
AND2    gate19326  (.A(g8212), .B(g17318), .Z(g19587) ) ;
AND2    gate19327  (.A(g8215), .B(g17321), .Z(g19588) ) ;
AND2    gate19328  (.A(g8224), .B(g17324), .Z(g19589) ) ;
AND2    gate19329  (.A(g8227), .B(g17327), .Z(g19590) ) ;
AND2    gate19330  (.A(g8230), .B(g17330), .Z(g19591) ) ;
AND2    gate19331  (.A(g8236), .B(g17333), .Z(g19592) ) ;
AND2    gate19332  (.A(g8239), .B(g17336), .Z(g19593) ) ;
AND2    gate19333  (.A(g16935), .B(g12555), .Z(g19594) ) ;
AND2    gate19334  (.A(g3922), .B(g17342), .Z(g19597) ) ;
AND2    gate19335  (.A(g3925), .B(g17345), .Z(g19598) ) ;
AND2    gate19336  (.A(g3928), .B(g17348), .Z(g19599) ) ;
AND2    gate19337  (.A(g633), .B(g18783), .Z(g19600) ) ;
AND2    gate19338  (.A(g640), .B(g18784), .Z(g19601) ) ;
AND2    gate19339  (.A(g633), .B(g18785), .Z(g19602) ) ;
AND2    gate19340  (.A(g692), .B(g18786), .Z(g19603) ) ;
AND2    gate19341  (.A(g3948), .B(g17354), .Z(g19604) ) ;
AND2    gate19342  (.A(g3951), .B(g17357), .Z(g19605) ) ;
AND2    gate19343  (.A(g3954), .B(g17360), .Z(g19606) ) ;
AND2    gate19344  (.A(g1326), .B(g18787), .Z(g19614) ) ;
AND2    gate19345  (.A(g1378), .B(g18788), .Z(g19615) ) ;
AND2    gate19346  (.A(g3966), .B(g17363), .Z(g19616) ) ;
AND2    gate19347  (.A(g3969), .B(g17366), .Z(g19617) ) ;
AND2    gate19348  (.A(g3972), .B(g17369), .Z(g19618) ) ;
AND2    gate19349  (.A(g3981), .B(g17372), .Z(g19619) ) ;
AND2    gate19350  (.A(g3984), .B(g17375), .Z(g19620) ) ;
AND2    gate19351  (.A(g3987), .B(g17378), .Z(g19621) ) ;
AND2    gate19352  (.A(g4000), .B(g17384), .Z(g19623) ) ;
AND2    gate19353  (.A(g4003), .B(g17387), .Z(g19624) ) ;
AND2    gate19354  (.A(g4006), .B(g17390), .Z(g19625) ) ;
AND2    gate19355  (.A(g640), .B(g18805), .Z(g19626) ) ;
AND2    gate19356  (.A(g633), .B(g18806), .Z(g19627) ) ;
AND2    gate19357  (.A(g653), .B(g18807), .Z(g19628) ) ;
AND2    gate19358  (.A(g692), .B(g18808), .Z(g19629) ) ;
AND2    gate19359  (.A(g4029), .B(g17399), .Z(g19630) ) ;
AND2    gate19360  (.A(g4032), .B(g17402), .Z(g19631) ) ;
AND2    gate19361  (.A(g4035), .B(g17405), .Z(g19632) ) ;
AND2    gate19362  (.A(g1319), .B(g18809), .Z(g19633) ) ;
AND2    gate19363  (.A(g1326), .B(g18810), .Z(g19634) ) ;
AND2    gate19364  (.A(g1319), .B(g18811), .Z(g19635) ) ;
AND2    gate19365  (.A(g1378), .B(g18812), .Z(g19636) ) ;
AND2    gate19366  (.A(g4055), .B(g17410), .Z(g19637) ) ;
AND2    gate19367  (.A(g4058), .B(g17413), .Z(g19638) ) ;
AND2    gate19368  (.A(g4061), .B(g17416), .Z(g19639) ) ;
AND2    gate19369  (.A(g2020), .B(g18813), .Z(g19647) ) ;
AND2    gate19370  (.A(g2072), .B(g18814), .Z(g19648) ) ;
AND2    gate19371  (.A(g4073), .B(g17419), .Z(g19649) ) ;
AND2    gate19372  (.A(g4076), .B(g17422), .Z(g19650) ) ;
AND2    gate19373  (.A(g4079), .B(g17425), .Z(g19651) ) ;
AND2    gate19374  (.A(g4095), .B(g17430), .Z(g19653) ) ;
AND2    gate19375  (.A(g4098), .B(g17433), .Z(g19654) ) ;
AND2    gate19376  (.A(g4101), .B(g17436), .Z(g19655) ) ;
AND2    gate19377  (.A(g4104), .B(g17439), .Z(g19656) ) ;
AND2    gate19378  (.A(g633), .B(g18822), .Z(g19660) ) ;
AND2    gate19379  (.A(g653), .B(g18823), .Z(g19661) ) ;
AND2    gate19380  (.A(g646), .B(g18824), .Z(g19662) ) ;
AND2    gate19381  (.A(g4127), .B(g17451), .Z(g19663) ) ;
AND2    gate19382  (.A(g4130), .B(g17454), .Z(g19664) ) ;
AND2    gate19383  (.A(g4133), .B(g17457), .Z(g19665) ) ;
AND2    gate19384  (.A(g1326), .B(g18825), .Z(g19666) ) ;
AND2    gate19385  (.A(g1319), .B(g18826), .Z(g19667) ) ;
AND2    gate19386  (.A(g1339), .B(g18827), .Z(g19668) ) ;
AND2    gate19387  (.A(g1378), .B(g18828), .Z(g19669) ) ;
AND2    gate19388  (.A(g4156), .B(g17465), .Z(g19670) ) ;
AND2    gate19389  (.A(g4159), .B(g17468), .Z(g19671) ) ;
AND2    gate19390  (.A(g4162), .B(g17471), .Z(g19672) ) ;
AND2    gate19391  (.A(g2013), .B(g18829), .Z(g19673) ) ;
AND2    gate19392  (.A(g2020), .B(g18830), .Z(g19674) ) ;
AND2    gate19393  (.A(g2013), .B(g18831), .Z(g19675) ) ;
AND2    gate19394  (.A(g2072), .B(g18832), .Z(g19676) ) ;
AND2    gate19395  (.A(g4182), .B(g17476), .Z(g19677) ) ;
AND2    gate19396  (.A(g4185), .B(g17479), .Z(g19678) ) ;
AND2    gate19397  (.A(g4188), .B(g17482), .Z(g19679) ) ;
AND2    gate19398  (.A(g2714), .B(g18833), .Z(g19687) ) ;
AND2    gate19399  (.A(g2766), .B(g18834), .Z(g19688) ) ;
NOR2    gate19400  (.A(g15021), .B(g12607), .Z(g16841) ) ;
AND2    gate19401  (.A(g16841), .B(g10865), .Z(g19691) ) ;
AND2    gate19402  (.A(g4205), .B(g17487), .Z(g19692) ) ;
AND2    gate19403  (.A(g4208), .B(g17490), .Z(g19693) ) ;
AND2    gate19404  (.A(g4211), .B(g17493), .Z(g19694) ) ;
AND2    gate19405  (.A(g4214), .B(g17496), .Z(g19695) ) ;
AND2    gate19406  (.A(g653), .B(g18838), .Z(g19697) ) ;
AND2    gate19407  (.A(g646), .B(g18839), .Z(g19698) ) ;
AND2    gate19408  (.A(g660), .B(g18840), .Z(g19699) ) ;
AND2    gate19409  (.A(g17815), .B(g16024), .Z(g19700) ) ;
AND2    gate19410  (.A(g4234), .B(g17511), .Z(g19701) ) ;
AND2    gate19411  (.A(g4237), .B(g17514), .Z(g19702) ) ;
AND2    gate19412  (.A(g4240), .B(g17517), .Z(g19703) ) ;
AND2    gate19413  (.A(g4243), .B(g17520), .Z(g19704) ) ;
AND2    gate19414  (.A(g1319), .B(g18841), .Z(g19708) ) ;
AND2    gate19415  (.A(g1339), .B(g18842), .Z(g19709) ) ;
AND2    gate19416  (.A(g1332), .B(g18843), .Z(g19710) ) ;
AND2    gate19417  (.A(g4266), .B(g17531), .Z(g19711) ) ;
AND2    gate19418  (.A(g4269), .B(g17534), .Z(g19712) ) ;
AND2    gate19419  (.A(g4272), .B(g17537), .Z(g19713) ) ;
AND2    gate19420  (.A(g2020), .B(g18844), .Z(g19714) ) ;
AND2    gate19421  (.A(g2013), .B(g18845), .Z(g19715) ) ;
AND2    gate19422  (.A(g2033), .B(g18846), .Z(g19716) ) ;
AND2    gate19423  (.A(g2072), .B(g18847), .Z(g19717) ) ;
AND2    gate19424  (.A(g4295), .B(g17545), .Z(g19718) ) ;
AND2    gate19425  (.A(g4298), .B(g17548), .Z(g19719) ) ;
AND2    gate19426  (.A(g4301), .B(g17551), .Z(g19720) ) ;
AND2    gate19427  (.A(g2707), .B(g18848), .Z(g19721) ) ;
AND2    gate19428  (.A(g2714), .B(g18849), .Z(g19722) ) ;
AND2    gate19429  (.A(g2707), .B(g18850), .Z(g19723) ) ;
AND2    gate19430  (.A(g2766), .B(g18851), .Z(g19724) ) ;
NOR2    gate19431  (.A(g15095), .B(g12650), .Z(g16847) ) ;
AND2    gate19432  (.A(g16847), .B(g6131), .Z(g19726) ) ;
AND2    gate19433  (.A(g4329), .B(g17557), .Z(g19727) ) ;
AND2    gate19434  (.A(g4332), .B(g17560), .Z(g19728) ) ;
AND2    gate19435  (.A(g4335), .B(g17563), .Z(g19729) ) ;
AND2    gate19436  (.A(g653), .B(g17573), .Z(g19730) ) ;
AND2    gate19437  (.A(g646), .B(g18853), .Z(g19731) ) ;
AND2    gate19438  (.A(g660), .B(g18854), .Z(g19732) ) ;
AND2    gate19439  (.A(g672), .B(g18855), .Z(g19733) ) ;
AND2    gate19440  (.A(g17815), .B(g16034), .Z(g19734) ) ;
AND2    gate19441  (.A(g17903), .B(g16035), .Z(g19735) ) ;
AND2    gate19442  (.A(g4360), .B(g17579), .Z(g19736) ) ;
AND2    gate19443  (.A(g4363), .B(g17582), .Z(g19737) ) ;
AND2    gate19444  (.A(g4366), .B(g17585), .Z(g19738) ) ;
AND2    gate19445  (.A(g4369), .B(g17588), .Z(g19739) ) ;
AND2    gate19446  (.A(g1339), .B(g18856), .Z(g19741) ) ;
AND2    gate19447  (.A(g1332), .B(g18857), .Z(g19742) ) ;
AND2    gate19448  (.A(g1346), .B(g18858), .Z(g19743) ) ;
AND2    gate19449  (.A(g17927), .B(g16040), .Z(g19744) ) ;
AND2    gate19450  (.A(g4389), .B(g17601), .Z(g19745) ) ;
AND2    gate19451  (.A(g4392), .B(g17604), .Z(g19746) ) ;
AND2    gate19452  (.A(g4395), .B(g17607), .Z(g19747) ) ;
AND2    gate19453  (.A(g4398), .B(g17610), .Z(g19748) ) ;
AND2    gate19454  (.A(g2013), .B(g18859), .Z(g19752) ) ;
AND2    gate19455  (.A(g2033), .B(g18860), .Z(g19753) ) ;
AND2    gate19456  (.A(g2026), .B(g18861), .Z(g19754) ) ;
AND2    gate19457  (.A(g4421), .B(g17621), .Z(g19755) ) ;
AND2    gate19458  (.A(g4424), .B(g17624), .Z(g19756) ) ;
AND2    gate19459  (.A(g4427), .B(g17627), .Z(g19757) ) ;
AND2    gate19460  (.A(g2714), .B(g18862), .Z(g19758) ) ;
AND2    gate19461  (.A(g2707), .B(g18863), .Z(g19759) ) ;
AND2    gate19462  (.A(g2727), .B(g18864), .Z(g19760) ) ;
AND2    gate19463  (.A(g2766), .B(g18865), .Z(g19761) ) ;
AND2    gate19464  (.A(g4453), .B(g17637), .Z(g19764) ) ;
AND2    gate19465  (.A(g660), .B(g18870), .Z(g19765) ) ;
AND2    gate19466  (.A(g672), .B(g18871), .Z(g19766) ) ;
AND2    gate19467  (.A(g666), .B(g18872), .Z(g19767) ) ;
AND2    gate19468  (.A(g17815), .B(g16054), .Z(g19768) ) ;
AND2    gate19469  (.A(g17903), .B(g16055), .Z(g19769) ) ;
AND2    gate19470  (.A(g4498), .B(g17655), .Z(g19770) ) ;
AND2    gate19471  (.A(g4501), .B(g17658), .Z(g19771) ) ;
AND2    gate19472  (.A(g4504), .B(g17661), .Z(g19772) ) ;
AND2    gate19473  (.A(g1339), .B(g17670), .Z(g19773) ) ;
AND2    gate19474  (.A(g1332), .B(g18874), .Z(g19774) ) ;
AND2    gate19475  (.A(g1346), .B(g18875), .Z(g19775) ) ;
AND2    gate19476  (.A(g1358), .B(g18876), .Z(g19776) ) ;
AND2    gate19477  (.A(g17927), .B(g16056), .Z(g19777) ) ;
AND2    gate19478  (.A(g18014), .B(g16057), .Z(g19778) ) ;
AND2    gate19479  (.A(g4529), .B(g17676), .Z(g19779) ) ;
AND2    gate19480  (.A(g4532), .B(g17679), .Z(g19780) ) ;
AND2    gate19481  (.A(g4535), .B(g17682), .Z(g19781) ) ;
AND2    gate19482  (.A(g4538), .B(g17685), .Z(g19782) ) ;
AND2    gate19483  (.A(g2033), .B(g18877), .Z(g19784) ) ;
AND2    gate19484  (.A(g2026), .B(g18878), .Z(g19785) ) ;
AND2    gate19485  (.A(g2040), .B(g18879), .Z(g19786) ) ;
AND2    gate19486  (.A(g18038), .B(g16062), .Z(g19787) ) ;
AND2    gate19487  (.A(g4558), .B(g17698), .Z(g19788) ) ;
AND2    gate19488  (.A(g4561), .B(g17701), .Z(g19789) ) ;
AND2    gate19489  (.A(g4564), .B(g17704), .Z(g19790) ) ;
AND2    gate19490  (.A(g4567), .B(g17707), .Z(g19791) ) ;
AND2    gate19491  (.A(g2707), .B(g18880), .Z(g19795) ) ;
AND2    gate19492  (.A(g2727), .B(g18881), .Z(g19796) ) ;
AND2    gate19493  (.A(g2720), .B(g18882), .Z(g19797) ) ;
AND3    gate19494  (.A(g18174), .B(g18341), .C(g17974), .Z(II26240) ) ;
AND3    gate19495  (.A(g17640), .B(g18074), .C(II26240), .Z(g19799) ) ;
AND2    gate19496  (.A(g672), .B(g18891), .Z(g19802) ) ;
AND2    gate19497  (.A(g666), .B(g18892), .Z(g19803) ) ;
AND2    gate19498  (.A(g679), .B(g18893), .Z(g19804) ) ;
AND2    gate19499  (.A(g17903), .B(g16088), .Z(g19805) ) ;
AND2    gate19500  (.A(g4629), .B(g17738), .Z(g19806) ) ;
AND2    gate19501  (.A(g1346), .B(g18896), .Z(g19807) ) ;
AND2    gate19502  (.A(g1358), .B(g18897), .Z(g19808) ) ;
AND2    gate19503  (.A(g1352), .B(g18898), .Z(g19809) ) ;
AND2    gate19504  (.A(g17927), .B(g16090), .Z(g19810) ) ;
AND2    gate19505  (.A(g18014), .B(g16091), .Z(g19811) ) ;
AND2    gate19506  (.A(g4674), .B(g17755), .Z(g19812) ) ;
AND2    gate19507  (.A(g4677), .B(g17758), .Z(g19813) ) ;
AND2    gate19508  (.A(g4680), .B(g17761), .Z(g19814) ) ;
AND2    gate19509  (.A(g2033), .B(g17770), .Z(g19815) ) ;
AND2    gate19510  (.A(g2026), .B(g18900), .Z(g19816) ) ;
AND2    gate19511  (.A(g2040), .B(g18901), .Z(g19817) ) ;
AND2    gate19512  (.A(g2052), .B(g18902), .Z(g19818) ) ;
AND2    gate19513  (.A(g18038), .B(g16092), .Z(g19819) ) ;
AND2    gate19514  (.A(g18131), .B(g16093), .Z(g19820) ) ;
AND2    gate19515  (.A(g4705), .B(g17776), .Z(g19821) ) ;
AND2    gate19516  (.A(g4708), .B(g17779), .Z(g19822) ) ;
AND2    gate19517  (.A(g4711), .B(g17782), .Z(g19823) ) ;
AND2    gate19518  (.A(g4714), .B(g17785), .Z(g19824) ) ;
AND2    gate19519  (.A(g2727), .B(g18903), .Z(g19826) ) ;
AND2    gate19520  (.A(g2720), .B(g18904), .Z(g19827) ) ;
AND2    gate19521  (.A(g2734), .B(g18905), .Z(g19828) ) ;
AND2    gate19522  (.A(g18155), .B(g16098), .Z(g19829) ) ;
AND2    gate19523  (.A(g7143), .B(g18908), .Z(g19836) ) ;
AND2    gate19524  (.A(g6901), .B(g17799), .Z(g19837) ) ;
AND2    gate19525  (.A(g666), .B(g18909), .Z(g19839) ) ;
AND2    gate19526  (.A(g679), .B(g18910), .Z(g19840) ) ;
AND2    gate19527  (.A(g686), .B(g18911), .Z(g19841) ) ;
AND3    gate19528  (.A(g18188), .B(g18089), .C(g17991), .Z(II26282) ) ;
AND3    gate19529  (.A(g14525), .B(g13922), .C(II26282), .Z(g19842) ) ;
AND3    gate19530  (.A(g18281), .B(g18436), .C(g18091), .Z(II26285) ) ;
AND3    gate19531  (.A(g17741), .B(g18190), .C(II26285), .Z(g19843) ) ;
AND2    gate19532  (.A(g1358), .B(g18914), .Z(g19846) ) ;
AND2    gate19533  (.A(g1352), .B(g18915), .Z(g19847) ) ;
AND2    gate19534  (.A(g1365), .B(g18916), .Z(g19848) ) ;
AND2    gate19535  (.A(g18014), .B(g16126), .Z(g19849) ) ;
AND2    gate19536  (.A(g4806), .B(g17839), .Z(g19850) ) ;
AND2    gate19537  (.A(g2040), .B(g18919), .Z(g19851) ) ;
AND2    gate19538  (.A(g2052), .B(g18920), .Z(g19852) ) ;
AND2    gate19539  (.A(g2046), .B(g18921), .Z(g19853) ) ;
AND2    gate19540  (.A(g18038), .B(g16128), .Z(g19854) ) ;
AND2    gate19541  (.A(g18131), .B(g16129), .Z(g19855) ) ;
AND2    gate19542  (.A(g4851), .B(g17856), .Z(g19856) ) ;
AND2    gate19543  (.A(g4854), .B(g17859), .Z(g19857) ) ;
AND2    gate19544  (.A(g4857), .B(g17862), .Z(g19858) ) ;
AND2    gate19545  (.A(g2727), .B(g17871), .Z(g19859) ) ;
AND2    gate19546  (.A(g2720), .B(g18923), .Z(g19860) ) ;
AND2    gate19547  (.A(g2734), .B(g18924), .Z(g19861) ) ;
AND2    gate19548  (.A(g2746), .B(g18925), .Z(g19862) ) ;
AND2    gate19549  (.A(g18155), .B(g16130), .Z(g19863) ) ;
AND2    gate19550  (.A(g18247), .B(g16131), .Z(g19864) ) ;
NOR2    gate19551  (.A(g14158), .B(g14347), .Z(g16498) ) ;
AND3    gate19552  (.A(g16498), .B(g16867), .C(g19001), .Z(g19868) ) ;
AND2    gate19553  (.A(g679), .B(g18926), .Z(g19869) ) ;
AND2    gate19554  (.A(g686), .B(g18927), .Z(g19870) ) ;
AND3    gate19555  (.A(g18353), .B(g13958), .C(g14011), .Z(II26311) ) ;
AND3    gate19556  (.A(g14086), .B(g18275), .C(II26311), .Z(g19871) ) ;
AND2    gate19557  (.A(g1352), .B(g18928), .Z(g19872) ) ;
AND2    gate19558  (.A(g1365), .B(g18929), .Z(g19873) ) ;
AND2    gate19559  (.A(g1372), .B(g18930), .Z(g19874) ) ;
AND3    gate19560  (.A(g18295), .B(g18205), .C(g18108), .Z(II26317) ) ;
AND3    gate19561  (.A(g14580), .B(g13978), .C(II26317), .Z(g19875) ) ;
AND3    gate19562  (.A(g18374), .B(g18509), .C(g18207), .Z(II26320) ) ;
AND3    gate19563  (.A(g17842), .B(g18297), .C(II26320), .Z(g19876) ) ;
AND2    gate19564  (.A(g2052), .B(g18933), .Z(g19879) ) ;
AND2    gate19565  (.A(g2046), .B(g18934), .Z(g19880) ) ;
AND2    gate19566  (.A(g2059), .B(g18935), .Z(g19881) ) ;
AND2    gate19567  (.A(g18131), .B(g16177), .Z(g19882) ) ;
AND2    gate19568  (.A(g4982), .B(g17951), .Z(g19883) ) ;
AND2    gate19569  (.A(g2734), .B(g18938), .Z(g19884) ) ;
AND2    gate19570  (.A(g2746), .B(g18939), .Z(g19885) ) ;
AND2    gate19571  (.A(g2740), .B(g18940), .Z(g19886) ) ;
AND2    gate19572  (.A(g18155), .B(g16179), .Z(g19887) ) ;
AND2    gate19573  (.A(g18247), .B(g16180), .Z(g19888) ) ;
AND2    gate19574  (.A(g2912), .B(g18943), .Z(g19889) ) ;
AND2    gate19575  (.A(g686), .B(g18945), .Z(g19895) ) ;
NOR2    gate19576  (.A(g14273), .B(g14459), .Z(g16520) ) ;
AND3    gate19577  (.A(g16520), .B(g16895), .C(g16507), .Z(g19899) ) ;
AND2    gate19578  (.A(g1365), .B(g18946), .Z(g19900) ) ;
AND2    gate19579  (.A(g1372), .B(g18947), .Z(g19901) ) ;
AND3    gate19580  (.A(g18448), .B(g14028), .C(g14102), .Z(II26348) ) ;
AND3    gate19581  (.A(g14201), .B(g18368), .C(II26348), .Z(g19902) ) ;
AND2    gate19582  (.A(g2046), .B(g18948), .Z(g19903) ) ;
AND2    gate19583  (.A(g2059), .B(g18949), .Z(g19904) ) ;
AND2    gate19584  (.A(g2066), .B(g18950), .Z(g19905) ) ;
AND3    gate19585  (.A(g18388), .B(g18312), .C(g18224), .Z(II26354) ) ;
AND3    gate19586  (.A(g14614), .B(g14048), .C(II26354), .Z(g19906) ) ;
AND3    gate19587  (.A(g18469), .B(g18573), .C(g18314), .Z(II26357) ) ;
AND3    gate19588  (.A(g17954), .B(g18390), .C(II26357), .Z(g19907) ) ;
AND2    gate19589  (.A(g2746), .B(g18953), .Z(g19910) ) ;
AND2    gate19590  (.A(g2740), .B(g18954), .Z(g19911) ) ;
AND2    gate19591  (.A(g2753), .B(g18955), .Z(g19912) ) ;
AND2    gate19592  (.A(g18247), .B(g16236), .Z(g19913) ) ;
AND2    gate19593  (.A(g3018), .B(g18958), .Z(g19914) ) ;
AND2    gate19594  (.A(g1372), .B(g18961), .Z(g19920) ) ;
NOR2    gate19595  (.A(g14395), .B(g14546), .Z(g16551) ) ;
AND3    gate19596  (.A(g16551), .B(g16924), .C(g16529), .Z(g19924) ) ;
AND2    gate19597  (.A(g2059), .B(g18962), .Z(g19925) ) ;
AND2    gate19598  (.A(g2066), .B(g18963), .Z(g19926) ) ;
AND3    gate19599  (.A(g18521), .B(g14119), .C(g14217), .Z(II26377) ) ;
AND3    gate19600  (.A(g14316), .B(g18463), .C(II26377), .Z(g19927) ) ;
AND2    gate19601  (.A(g2740), .B(g18964), .Z(g19928) ) ;
AND2    gate19602  (.A(g2753), .B(g18965), .Z(g19929) ) ;
AND2    gate19603  (.A(g2760), .B(g18966), .Z(g19930) ) ;
AND3    gate19604  (.A(g18483), .B(g18405), .C(g18331), .Z(II26383) ) ;
AND3    gate19605  (.A(g14637), .B(g14139), .C(II26383), .Z(g19931) ) ;
AND2    gate19606  (.A(g2917), .B(g18166), .Z(g19932) ) ;
AND2    gate19607  (.A(g2066), .B(g18972), .Z(g19935) ) ;
NOR2    gate19608  (.A(g14507), .B(g14601), .Z(g16583) ) ;
AND3    gate19609  (.A(g16583), .B(g16954), .C(g16560), .Z(g19939) ) ;
AND2    gate19610  (.A(g2753), .B(g18973), .Z(g19940) ) ;
AND2    gate19611  (.A(g2760), .B(g18974), .Z(g19941) ) ;
AND3    gate19612  (.A(g18585), .B(g14234), .C(g14332), .Z(II26396) ) ;
AND3    gate19613  (.A(g14438), .B(g18536), .C(II26396), .Z(g19942) ) ;
AND2    gate19614  (.A(g7562), .B(g18976), .Z(g19943) ) ;
AND2    gate19615  (.A(g3028), .B(g18258), .Z(g19944) ) ;
AND2    gate19616  (.A(g5293), .B(g18278), .Z(g19949) ) ;
AND2    gate19617  (.A(g2760), .B(g18987), .Z(g19952) ) ;
AND2    gate19618  (.A(g7566), .B(g18334), .Z(g19953) ) ;
NAND2   gate19619  (.A(II24625), .B(II24626), .Z(g18553) ) ;
NAND2   gate19620  (.A(II24531), .B(II24532), .Z(g18491) ) ;
NAND2   gate19621  (.A(II24453), .B(II24454), .Z(g18431) ) ;
AND3    gate19622  (.A(g18553), .B(g18491), .C(g18431), .Z(II26416) ) ;
NAND2   gate19623  (.A(II24362), .B(II24363), .Z(g18354) ) ;
NAND2   gate19624  (.A(II24272), .B(II24273), .Z(g18276) ) ;
AND3    gate19625  (.A(g18354), .B(g18276), .C(II26416), .Z(g19970) ) ;
AND2    gate19626  (.A(g5327), .B(g18355), .Z(g19971) ) ;
AND2    gate19627  (.A(g5330), .B(g18371), .Z(g19976) ) ;
NAND2   gate19628  (.A(II24279), .B(II24280), .Z(g18277) ) ;
NAND2   gate19629  (.A(II24187), .B(II24188), .Z(g18189) ) ;
NAND2   gate19630  (.A(II24103), .B(II24104), .Z(g18090) ) ;
AND3    gate19631  (.A(g18277), .B(g18189), .C(g18090), .Z(II26432) ) ;
NAND2   gate19632  (.A(II24029), .B(II24030), .Z(g17992) ) ;
NAND2   gate19633  (.A(II23959), .B(II23960), .Z(g17913) ) ;
AND3    gate19634  (.A(g17992), .B(g17913), .C(II26432), .Z(g19982) ) ;
AND2    gate19635  (.A(g5352), .B(g18432), .Z(g19983) ) ;
NAND2   gate19636  (.A(II24695), .B(II24696), .Z(g18603) ) ;
NAND2   gate19637  (.A(II24633), .B(II24634), .Z(g18555) ) ;
NAND2   gate19638  (.A(II24554), .B(II24555), .Z(g18504) ) ;
AND3    gate19639  (.A(g18603), .B(g18555), .C(g18504), .Z(II26440) ) ;
NAND2   gate19640  (.A(II24475), .B(II24476), .Z(g18449) ) ;
NAND2   gate19641  (.A(II24381), .B(II24382), .Z(g18369) ) ;
AND3    gate19642  (.A(g18449), .B(g18369), .C(II26440), .Z(g20000) ) ;
AND2    gate19643  (.A(g5355), .B(g18450), .Z(g20001) ) ;
AND2    gate19644  (.A(g5358), .B(g18466), .Z(g20006) ) ;
AND2    gate19645  (.A(g18063), .B(g3113), .Z(g20011) ) ;
AND2    gate19646  (.A(g16804), .B(g3135), .Z(g20012) ) ;
AND2    gate19647  (.A(g17720), .B(g12848), .Z(g20013) ) ;
AND2    gate19648  (.A(g7615), .B(g16749), .Z(g20014) ) ;
NAND2   gate19649  (.A(II24388), .B(II24389), .Z(g18370) ) ;
NAND2   gate19650  (.A(II24299), .B(II24300), .Z(g18296) ) ;
NAND2   gate19651  (.A(II24206), .B(II24207), .Z(g18206) ) ;
AND3    gate19652  (.A(g18370), .B(g18296), .C(g18206), .Z(II26464) ) ;
NAND2   gate19653  (.A(II24124), .B(II24125), .Z(g18109) ) ;
NAND2   gate19654  (.A(II24054), .B(II24055), .Z(g18024) ) ;
AND3    gate19655  (.A(g18109), .B(g18024), .C(II26464), .Z(g20020) ) ;
AND2    gate19656  (.A(g5369), .B(g18505), .Z(g20021) ) ;
NAND2   gate19657  (.A(II24744), .B(II24745), .Z(g18635) ) ;
NAND2   gate19658  (.A(II24703), .B(II24704), .Z(g18605) ) ;
NAND2   gate19659  (.A(II24656), .B(II24657), .Z(g18568) ) ;
AND3    gate19660  (.A(g18635), .B(g18605), .C(g18568), .Z(II26472) ) ;
NAND2   gate19661  (.A(II24576), .B(II24577), .Z(g18522) ) ;
NAND2   gate19662  (.A(II24494), .B(II24495), .Z(g18464) ) ;
AND3    gate19663  (.A(g18522), .B(g18464), .C(II26472), .Z(g20038) ) ;
AND2    gate19664  (.A(g5372), .B(g18523), .Z(g20039) ) ;
AND2    gate19665  (.A(g5375), .B(g18539), .Z(g20044) ) ;
AND2    gate19666  (.A(g16749), .B(g3127), .Z(g20048) ) ;
AND2    gate19667  (.A(g17878), .B(g3155), .Z(g20049) ) ;
AND2    gate19668  (.A(g18070), .B(g3161), .Z(g20050) ) ;
AND2    gate19669  (.A(g18063), .B(g3114), .Z(g20051) ) ;
AND2    gate19670  (.A(g16804), .B(g3134), .Z(g20052) ) ;
AND2    gate19671  (.A(g17720), .B(g12875), .Z(g20053) ) ;
NAND2   gate19672  (.A(II24501), .B(II24502), .Z(g18465) ) ;
NAND2   gate19673  (.A(II24408), .B(II24409), .Z(g18389) ) ;
NAND2   gate19674  (.A(II24318), .B(II24319), .Z(g18313) ) ;
AND3    gate19675  (.A(g18465), .B(g18389), .C(g18313), .Z(II26500) ) ;
NAND2   gate19676  (.A(II24227), .B(II24228), .Z(g18225) ) ;
NAND2   gate19677  (.A(II24149), .B(II24150), .Z(g18141) ) ;
AND3    gate19678  (.A(g18225), .B(g18141), .C(II26500), .Z(g20062) ) ;
AND2    gate19679  (.A(g5382), .B(g18569), .Z(g20063) ) ;
NAND2   gate19680  (.A(II24764), .B(II24765), .Z(g18644) ) ;
NAND2   gate19681  (.A(II24752), .B(II24753), .Z(g18637) ) ;
NAND2   gate19682  (.A(II24726), .B(II24727), .Z(g18618) ) ;
AND3    gate19683  (.A(g18644), .B(g18637), .C(g18618), .Z(II26508) ) ;
NAND2   gate19684  (.A(II24678), .B(II24679), .Z(g18586) ) ;
NAND2   gate19685  (.A(II24595), .B(II24596), .Z(g18537) ) ;
AND3    gate19686  (.A(g18586), .B(g18537), .C(II26508), .Z(g20080) ) ;
AND2    gate19687  (.A(g5385), .B(g18587), .Z(g20081) ) ;
AND2    gate19688  (.A(g17969), .B(g3158), .Z(g20084) ) ;
AND2    gate19689  (.A(g18170), .B(g3164), .Z(g20085) ) ;
AND2    gate19690  (.A(g18337), .B(g3170), .Z(g20086) ) ;
AND2    gate19691  (.A(g16749), .B(g7574), .Z(g20087) ) ;
AND2    gate19692  (.A(g16836), .B(g3147), .Z(g20088) ) ;
AND2    gate19693  (.A(g17969), .B(g9160), .Z(g20089) ) ;
AND2    gate19694  (.A(g18063), .B(g3120), .Z(g20090) ) ;
AND2    gate19695  (.A(g16804), .B(g3136), .Z(g20091) ) ;
AND2    gate19696  (.A(g16749), .B(g7603), .Z(g20092) ) ;
AND3    gate19697  (.A(g18656), .B(g18670), .C(g18692), .Z(II26525) ) ;
AND4    gate19698  (.A(g13657), .B(g13677), .C(g13750), .D(II26525), .Z(g20093) ) ;
AND3    gate19699  (.A(g18656), .B(g14837), .C(g13657), .Z(II26528) ) ;
AND3    gate19700  (.A(g13677), .B(g13706), .C(II26528), .Z(g20094) ) ;
NAND2   gate19701  (.A(II24602), .B(II24603), .Z(g18538) ) ;
NAND2   gate19702  (.A(II24521), .B(II24522), .Z(g18484) ) ;
NAND2   gate19703  (.A(II24427), .B(II24428), .Z(g18406) ) ;
AND3    gate19704  (.A(g18538), .B(g18484), .C(g18406), .Z(II26541) ) ;
NAND2   gate19705  (.A(II24339), .B(II24340), .Z(g18332) ) ;
NAND2   gate19706  (.A(II24252), .B(II24253), .Z(g18257) ) ;
AND3    gate19707  (.A(g18332), .B(g18257), .C(II26541), .Z(g20103) ) ;
AND2    gate19708  (.A(g5391), .B(g18619), .Z(g20104) ) ;
AND2    gate19709  (.A(g18261), .B(g3167), .Z(g20106) ) ;
AND2    gate19710  (.A(g18415), .B(g3173), .Z(g20107) ) ;
AND2    gate19711  (.A(g18543), .B(g3179), .Z(g20108) ) ;
AND2    gate19712  (.A(g17878), .B(g9504), .Z(g20109) ) ;
AND2    gate19713  (.A(g18070), .B(g9286), .Z(g20110) ) ;
AND2    gate19714  (.A(g18261), .B(g9884), .Z(g20111) ) ;
AND2    gate19715  (.A(g16749), .B(g3132), .Z(g20112) ) ;
AND2    gate19716  (.A(g16836), .B(g3142), .Z(g20113) ) ;
AND2    gate19717  (.A(g17969), .B(g9755), .Z(g20114) ) ;
AND2    gate19718  (.A(g16804), .B(g3139), .Z(g20115) ) ;
AND3    gate19719  (.A(g14776), .B(g18670), .C(g18720), .Z(II26558) ) ;
AND4    gate19720  (.A(g16142), .B(g13677), .C(g13706), .D(II26558), .Z(g20116) ) ;
AND3    gate19721  (.A(g14776), .B(g18720), .C(g13657), .Z(II26561) ) ;
AND3    gate19722  (.A(g16189), .B(g13706), .C(II26561), .Z(g20117) ) ;
AND3    gate19723  (.A(g18679), .B(g18699), .C(g18728), .Z(II26564) ) ;
AND4    gate19724  (.A(g13687), .B(g13714), .C(g13791), .D(II26564), .Z(g20118) ) ;
AND3    gate19725  (.A(g18679), .B(g14910), .C(g13687), .Z(II26567) ) ;
AND3    gate19726  (.A(g13714), .B(g13756), .C(II26567), .Z(g20119) ) ;
AND2    gate19727  (.A(g18486), .B(g3176), .Z(g20131) ) ;
AND2    gate19728  (.A(g18593), .B(g3182), .Z(g20132) ) ;
AND2    gate19729  (.A(g18170), .B(g9505), .Z(g20133) ) ;
AND2    gate19730  (.A(g18337), .B(g9506), .Z(g20134) ) ;
AND2    gate19731  (.A(g18486), .B(g9885), .Z(g20135) ) ;
AND2    gate19732  (.A(g17878), .B(g9423), .Z(g20136) ) ;
AND2    gate19733  (.A(g18070), .B(g9226), .Z(g20137) ) ;
AND2    gate19734  (.A(g18261), .B(g9756), .Z(g20138) ) ;
AND2    gate19735  (.A(g16836), .B(g3151), .Z(g20139) ) ;
NOR2    gate19736  (.A(g14797), .B(g14895), .Z(g16679) ) ;
AND3    gate19737  (.A(g16679), .B(g16884), .C(g16665), .Z(g20144) ) ;
AND4    gate19738  (.A(g14776), .B(g18670), .C(g16142), .D(g16189), .Z(g20145) ) ;
AND3    gate19739  (.A(g14811), .B(g18699), .C(g18758), .Z(II26590) ) ;
AND4    gate19740  (.A(g16201), .B(g13714), .C(g13756), .D(II26590), .Z(g20146) ) ;
AND3    gate19741  (.A(g14811), .B(g18758), .C(g13687), .Z(II26593) ) ;
AND3    gate19742  (.A(g16254), .B(g13756), .C(II26593), .Z(g20147) ) ;
AND3    gate19743  (.A(g18708), .B(g18735), .C(g18765), .Z(II26596) ) ;
AND4    gate19744  (.A(g13724), .B(g13764), .C(g13819), .D(II26596), .Z(g20148) ) ;
AND3    gate19745  (.A(g18708), .B(g14991), .C(g13724), .Z(II26599) ) ;
AND3    gate19746  (.A(g13764), .B(g13797), .C(II26599), .Z(g20149) ) ;
AND2    gate19747  (.A(g16809), .B(g3185), .Z(g20156) ) ;
AND2    gate19748  (.A(g18415), .B(g9287), .Z(g20157) ) ;
AND2    gate19749  (.A(g18543), .B(g9886), .Z(g20158) ) ;
AND2    gate19750  (.A(g16809), .B(g9288), .Z(g20159) ) ;
AND2    gate19751  (.A(g18170), .B(g9424), .Z(g20160) ) ;
AND2    gate19752  (.A(g18337), .B(g9426), .Z(g20161) ) ;
AND2    gate19753  (.A(g18486), .B(g9757), .Z(g20162) ) ;
AND3    gate19754  (.A(g14797), .B(g18692), .C(g13657), .Z(II26615) ) ;
AND3    gate19755  (.A(g13677), .B(g13750), .C(II26615), .Z(g20177) ) ;
NOR2    gate19756  (.A(g14849), .B(g14976), .Z(g16705) ) ;
AND3    gate19757  (.A(g16705), .B(g16913), .C(g16686), .Z(g20182) ) ;
AND4    gate19758  (.A(g14811), .B(g18699), .C(g16201), .D(g16254), .Z(g20183) ) ;
AND3    gate19759  (.A(g14863), .B(g18735), .C(g18789), .Z(II26621) ) ;
AND4    gate19760  (.A(g16266), .B(g13764), .C(g13797), .D(II26621), .Z(g20184) ) ;
AND3    gate19761  (.A(g14863), .B(g18789), .C(g13724), .Z(II26624) ) ;
AND3    gate19762  (.A(g16313), .B(g13797), .C(II26624), .Z(g20185) ) ;
AND3    gate19763  (.A(g18744), .B(g18772), .C(g18796), .Z(II26627) ) ;
AND4    gate19764  (.A(g13774), .B(g13805), .C(g13840), .D(II26627), .Z(g20186) ) ;
AND3    gate19765  (.A(g18744), .B(g15080), .C(g13774), .Z(II26630) ) ;
AND3    gate19766  (.A(g13805), .B(g13825), .C(II26630), .Z(g20187) ) ;
AND2    gate19767  (.A(g18593), .B(g9425), .Z(g20188) ) ;
AND2    gate19768  (.A(g16825), .B(g9289), .Z(g20189) ) ;
AND2    gate19769  (.A(g18415), .B(g9227), .Z(g20190) ) ;
AND2    gate19770  (.A(g18543), .B(g9758), .Z(g20191) ) ;
AND2    gate19771  (.A(g16809), .B(g9228), .Z(g20192) ) ;
AND3    gate19772  (.A(g18656), .B(g18670), .C(g16142), .Z(II26639) ) ;
AND3    gate19773  (.A(g13677), .B(g13706), .C(II26639), .Z(g20197) ) ;
AND3    gate19774  (.A(g14849), .B(g18728), .C(g13687), .Z(II26645) ) ;
AND3    gate19775  (.A(g13714), .B(g13791), .C(II26645), .Z(g20211) ) ;
NOR2    gate19776  (.A(g14922), .B(g15065), .Z(g16736) ) ;
AND3    gate19777  (.A(g16736), .B(g16943), .C(g16712), .Z(g20216) ) ;
AND4    gate19778  (.A(g14863), .B(g18735), .C(g16266), .D(g16313), .Z(g20217) ) ;
AND3    gate19779  (.A(g14936), .B(g18772), .C(g18815), .Z(II26651) ) ;
AND4    gate19780  (.A(g16325), .B(g13805), .C(g13825), .D(II26651), .Z(g20218) ) ;
AND3    gate19781  (.A(g14936), .B(g18815), .C(g13774), .Z(II26654) ) ;
AND3    gate19782  (.A(g16371), .B(g13825), .C(II26654), .Z(g20219) ) ;
AND2    gate19783  (.A(g18593), .B(g9355), .Z(g20220) ) ;
AND2    gate19784  (.A(g16825), .B(g10099), .Z(g20221) ) ;
AND4    gate19785  (.A(g18656), .B(g18720), .C(g13657), .D(g16293), .Z(g20222) ) ;
AND3    gate19786  (.A(g18679), .B(g18699), .C(g16201), .Z(II26661) ) ;
AND3    gate19787  (.A(g13714), .B(g13756), .C(II26661), .Z(g20227) ) ;
AND3    gate19788  (.A(g14922), .B(g18765), .C(g13724), .Z(II26667) ) ;
AND3    gate19789  (.A(g13764), .B(g13819), .C(II26667), .Z(g20241) ) ;
NOR2    gate19790  (.A(g15003), .B(g15161), .Z(g16778) ) ;
AND3    gate19791  (.A(g16778), .B(g16974), .C(g16743), .Z(g20246) ) ;
AND4    gate19792  (.A(g14936), .B(g18772), .C(g16325), .D(g16371), .Z(g20247) ) ;
AND3    gate19793  (.A(g18656), .B(g14837), .C(g16293), .Z(g20248) ) ;
AND4    gate19794  (.A(g18679), .B(g18758), .C(g13687), .D(g16351), .Z(g20249) ) ;
AND3    gate19795  (.A(g18708), .B(g18735), .C(g16266), .Z(II26676) ) ;
AND3    gate19796  (.A(g13764), .B(g13797), .C(II26676), .Z(g20254) ) ;
AND3    gate19797  (.A(g15003), .B(g18796), .C(g13774), .Z(II26682) ) ;
AND3    gate19798  (.A(g13805), .B(g13840), .C(II26682), .Z(g20268) ) ;
AND4    gate19799  (.A(g14797), .B(g18692), .C(g13657), .D(g16243), .Z(g20270) ) ;
AND3    gate19800  (.A(g18679), .B(g14910), .C(g16351), .Z(g20271) ) ;
AND4    gate19801  (.A(g18708), .B(g18789), .C(g13724), .D(g16395), .Z(g20272) ) ;
AND3    gate19802  (.A(g18744), .B(g18772), .C(g16325), .Z(II26690) ) ;
AND3    gate19803  (.A(g13805), .B(g13825), .C(II26690), .Z(g20277) ) ;
AND3    gate19804  (.A(g18670), .B(g18692), .C(g16142), .Z(II26695) ) ;
AND3    gate19805  (.A(g13677), .B(g16243), .C(II26695), .Z(g20280) ) ;
AND4    gate19806  (.A(g14849), .B(g18728), .C(g13687), .D(g16302), .Z(g20282) ) ;
AND3    gate19807  (.A(g18708), .B(g14991), .C(g16395), .Z(g20283) ) ;
AND4    gate19808  (.A(g18744), .B(g18815), .C(g13774), .D(g16433), .Z(g20284) ) ;
AND2    gate19809  (.A(g16846), .B(g8103), .Z(g20285) ) ;
AND3    gate19810  (.A(g18699), .B(g18728), .C(g16201), .Z(II26708) ) ;
AND3    gate19811  (.A(g13714), .B(g16302), .C(II26708), .Z(g20291) ) ;
AND4    gate19812  (.A(g14922), .B(g18765), .C(g13724), .D(g16360), .Z(g20293) ) ;
AND3    gate19813  (.A(g18744), .B(g15080), .C(g16433), .Z(g20294) ) ;
AND3    gate19814  (.A(g18735), .B(g18765), .C(g16266), .Z(II26726) ) ;
AND3    gate19815  (.A(g13764), .B(g16360), .C(II26726), .Z(g20307) ) ;
AND4    gate19816  (.A(g15003), .B(g18796), .C(g13774), .D(g16404), .Z(g20309) ) ;
AND3    gate19817  (.A(g18772), .B(g18796), .C(g16325), .Z(II26745) ) ;
AND3    gate19818  (.A(g13805), .B(g16404), .C(II26745), .Z(g20326) ) ;
AND2    gate19819  (.A(g17351), .B(g13644), .Z(g20460) ) ;
AND2    gate19820  (.A(g17314), .B(g13669), .Z(g20472) ) ;
AND2    gate19821  (.A(g17313), .B(g11827), .Z(g20480) ) ;
AND2    gate19822  (.A(g17281), .B(g11859), .Z(g20486) ) ;
AND2    gate19823  (.A(g17258), .B(g11894), .Z(g20492) ) ;
AND2    gate19824  (.A(g17648), .B(g11933), .Z(g20499) ) ;
AND2    gate19825  (.A(g17566), .B(g11973), .Z(g20502) ) ;
NOR2    gate19826  (.A(g16298), .B(g13318), .Z(g17507) ) ;
AND2    gate19827  (.A(g17507), .B(g13817), .Z(g20503) ) ;
AND2    gate19828  (.A(g17499), .B(g12025), .Z(g20506) ) ;
AND2    gate19829  (.A(g17445), .B(g13836), .Z(g20512) ) ;
AND2    gate19830  (.A(g17394), .B(g13849), .Z(g20525) ) ;
AND4    gate19831  (.A(g18656), .B(g14837), .C(g13657), .D(g16189), .Z(g20538) ) ;
AND2    gate19832  (.A(g4809), .B(g19064), .Z(g20640) ) ;
AND2    gate19833  (.A(g5888), .B(g19075), .Z(g20647) ) ;
AND2    gate19834  (.A(g4985), .B(g19081), .Z(g20665) ) ;
AND2    gate19835  (.A(g5712), .B(g19113), .Z(g20809) ) ;
AND2    gate19836  (.A(g5770), .B(g19118), .Z(g20826) ) ;
AND2    gate19837  (.A(g5829), .B(g19125), .Z(g20836) ) ;
AND2    gate19838  (.A(g5885), .B(g19132), .Z(g20840) ) ;
AND3    gate19839  (.A(g20016), .B(g14079), .C(g14165), .Z(g21049) ) ;
AND2    gate19840  (.A(g20193), .B(g12030), .Z(g21067) ) ;
AND3    gate19841  (.A(g20058), .B(g14194), .C(g14280), .Z(g21068) ) ;
AND2    gate19842  (.A(g20223), .B(g12094), .Z(g21077) ) ;
AND3    gate19843  (.A(g20099), .B(g14309), .C(g14402), .Z(g21078) ) ;
AND3    gate19844  (.A(g19484), .B(g14158), .C(g19001), .Z(g21085) ) ;
AND2    gate19845  (.A(g20193), .B(g12142), .Z(g21086) ) ;
AND2    gate19846  (.A(g20250), .B(g12166), .Z(g21091) ) ;
AND3    gate19847  (.A(g20124), .B(g14431), .C(g14514), .Z(g21092) ) ;
AND3    gate19848  (.A(g19505), .B(g14273), .C(g16507), .Z(g21097) ) ;
AND2    gate19849  (.A(g20223), .B(g12204), .Z(g21098) ) ;
AND2    gate19850  (.A(g20273), .B(g12228), .Z(g21103) ) ;
AND3    gate19851  (.A(g19444), .B(g17893), .C(g14079), .Z(g21107) ) ;
AND3    gate19852  (.A(g19524), .B(g14395), .C(g16529), .Z(g21111) ) ;
AND2    gate19853  (.A(g20250), .B(g12259), .Z(g21112) ) ;
NOR2    gate19854  (.A(g19001), .B(g16867), .Z(g20054) ) ;
AND2    gate19855  (.A(g20054), .B(g14244), .Z(g21121) ) ;
AND2    gate19856  (.A(g20140), .B(g12279), .Z(g21122) ) ;
AND2    gate19857  (.A(g19970), .B(g19982), .Z(g21123) ) ;
AND3    gate19858  (.A(g19471), .B(g18004), .C(g14194), .Z(g21124) ) ;
AND3    gate19859  (.A(g19534), .B(g14507), .C(g16560), .Z(g21128) ) ;
AND2    gate19860  (.A(g20273), .B(g12302), .Z(g21129) ) ;
NAND2   gate19861  (.A(II25682), .B(II25683), .Z(g19318) ) ;
NAND2   gate19862  (.A(II25634), .B(II25635), .Z(g19300) ) ;
NAND2   gate19863  (.A(II25596), .B(II25597), .Z(g19286) ) ;
AND3    gate19864  (.A(g19318), .B(g19300), .C(g19286), .Z(II27695) ) ;
NAND2   gate19865  (.A(II25561), .B(II25562), .Z(g19271) ) ;
NAND2   gate19866  (.A(II25533), .B(II25534), .Z(g19261) ) ;
AND3    gate19867  (.A(g19271), .B(g19261), .C(II27695), .Z(g21136) ) ;
AND2    gate19868  (.A(g5750), .B(g19272), .Z(g21137) ) ;
AND2    gate19869  (.A(g19484), .B(g14347), .Z(g21138) ) ;
NOR2    gate19870  (.A(g16507), .B(g16895), .Z(g20095) ) ;
AND2    gate19871  (.A(g20095), .B(g14366), .Z(g21140) ) ;
AND2    gate19872  (.A(g20178), .B(g12315), .Z(g21141) ) ;
AND2    gate19873  (.A(g20000), .B(g20020), .Z(g21142) ) ;
AND3    gate19874  (.A(g19494), .B(g18121), .C(g14309), .Z(g21143) ) ;
NAND2   gate19875  (.A(II25540), .B(II25541), .Z(g19262) ) ;
NAND2   gate19876  (.A(II25839), .B(II25840), .Z(g19414) ) ;
NAND2   gate19877  (.A(II25801), .B(II25802), .Z(g19386) ) ;
AND3    gate19878  (.A(g19262), .B(g19414), .C(g19386), .Z(II27711) ) ;
NAND2   gate19879  (.A(II25762), .B(II25763), .Z(g19357) ) ;
NAND2   gate19880  (.A(II25722), .B(II25723), .Z(g19334) ) ;
AND3    gate19881  (.A(g19357), .B(g19334), .C(II27711), .Z(g21152) ) ;
AND3    gate19882  (.A(g20054), .B(g16543), .C(g16501), .Z(g21153) ) ;
AND2    gate19883  (.A(g20193), .B(g12333), .Z(g21154) ) ;
AND2    gate19884  (.A(g20140), .B(g12336), .Z(g21155) ) ;
NAND2   gate19885  (.A(II25732), .B(II25733), .Z(g19345) ) ;
NAND2   gate19886  (.A(II25691), .B(II25692), .Z(g19321) ) ;
NAND2   gate19887  (.A(II25644), .B(II25645), .Z(g19304) ) ;
AND3    gate19888  (.A(g19345), .B(g19321), .C(g19304), .Z(II27717) ) ;
NAND2   gate19889  (.A(II25606), .B(II25607), .Z(g19290) ) ;
NAND2   gate19890  (.A(II25572), .B(II25573), .Z(g19276) ) ;
AND3    gate19891  (.A(g19290), .B(g19276), .C(II27717), .Z(g21156) ) ;
AND2    gate19892  (.A(g5809), .B(g19291), .Z(g21157) ) ;
AND2    gate19893  (.A(g19505), .B(g14459), .Z(g21158) ) ;
NOR2    gate19894  (.A(g16529), .B(g16924), .Z(g20120) ) ;
AND2    gate19895  (.A(g20120), .B(g14478), .Z(g21160) ) ;
AND2    gate19896  (.A(g20212), .B(g12343), .Z(g21161) ) ;
AND2    gate19897  (.A(g20038), .B(g20062), .Z(g21162) ) ;
AND3    gate19898  (.A(g19515), .B(g18237), .C(g14431), .Z(g21163) ) ;
NAND2   gate19899  (.A(II25579), .B(II25580), .Z(g19277) ) ;
NAND2   gate19900  (.A(II25881), .B(II25882), .Z(g19451) ) ;
NAND2   gate19901  (.A(II25847), .B(II25848), .Z(g19416) ) ;
AND3    gate19902  (.A(g19277), .B(g19451), .C(g19416), .Z(II27733) ) ;
NAND2   gate19903  (.A(II25810), .B(II25811), .Z(g19389) ) ;
NAND2   gate19904  (.A(II25772), .B(II25773), .Z(g19368) ) ;
AND3    gate19905  (.A(g19389), .B(g19368), .C(II27733), .Z(g21172) ) ;
AND3    gate19906  (.A(g20095), .B(g16575), .C(g16523), .Z(g21173) ) ;
AND2    gate19907  (.A(g20223), .B(g12363), .Z(g21174) ) ;
AND2    gate19908  (.A(g20178), .B(g12366), .Z(g21175) ) ;
NAND2   gate19909  (.A(II25782), .B(II25783), .Z(g19379) ) ;
NAND2   gate19910  (.A(II25741), .B(II25742), .Z(g19348) ) ;
NAND2   gate19911  (.A(II25701), .B(II25702), .Z(g19325) ) ;
AND3    gate19912  (.A(g19379), .B(g19348), .C(g19325), .Z(II27739) ) ;
NAND2   gate19913  (.A(II25654), .B(II25655), .Z(g19308) ) ;
NAND2   gate19914  (.A(II25617), .B(II25618), .Z(g19295) ) ;
AND3    gate19915  (.A(g19308), .B(g19295), .C(II27739), .Z(g21176) ) ;
AND2    gate19916  (.A(g5865), .B(g19309), .Z(g21177) ) ;
AND2    gate19917  (.A(g19524), .B(g14546), .Z(g21178) ) ;
NOR2    gate19918  (.A(g16560), .B(g16954), .Z(g20150) ) ;
AND2    gate19919  (.A(g20150), .B(g14565), .Z(g21180) ) ;
AND2    gate19920  (.A(g20242), .B(g12373), .Z(g21181) ) ;
AND2    gate19921  (.A(g20080), .B(g20103), .Z(g21182) ) ;
AND2    gate19922  (.A(g20140), .B(g12379), .Z(g21188) ) ;
NAND2   gate19923  (.A(II25624), .B(II25625), .Z(g19296) ) ;
NAND2   gate19924  (.A(II25914), .B(II25915), .Z(g19478) ) ;
NAND2   gate19925  (.A(II25889), .B(II25890), .Z(g19453) ) ;
AND3    gate19926  (.A(g19296), .B(g19478), .C(g19453), .Z(II27755) ) ;
NAND2   gate19927  (.A(II25856), .B(II25857), .Z(g19419) ) ;
NAND2   gate19928  (.A(II25820), .B(II25821), .Z(g19400) ) ;
AND3    gate19929  (.A(g19419), .B(g19400), .C(II27755), .Z(g21192) ) ;
AND3    gate19930  (.A(g20120), .B(g16599), .C(g16554), .Z(g21193) ) ;
AND2    gate19931  (.A(g20250), .B(g12382), .Z(g21194) ) ;
AND2    gate19932  (.A(g20212), .B(g12385), .Z(g21195) ) ;
NAND2   gate19933  (.A(II25830), .B(II25831), .Z(g19411) ) ;
NAND2   gate19934  (.A(II25791), .B(II25792), .Z(g19382) ) ;
NAND2   gate19935  (.A(II25751), .B(II25752), .Z(g19352) ) ;
AND3    gate19936  (.A(g19411), .B(g19382), .C(g19352), .Z(II27761) ) ;
NAND2   gate19937  (.A(II25711), .B(II25712), .Z(g19329) ) ;
NAND2   gate19938  (.A(II25665), .B(II25666), .Z(g19313) ) ;
AND3    gate19939  (.A(g19329), .B(g19313), .C(II27761), .Z(g21196) ) ;
AND2    gate19940  (.A(g5912), .B(g19330), .Z(g21197) ) ;
AND2    gate19941  (.A(g19534), .B(g14601), .Z(g21198) ) ;
AND2    gate19942  (.A(g20178), .B(g12409), .Z(g21203) ) ;
NAND2   gate19943  (.A(II25672), .B(II25673), .Z(g19314) ) ;
NAND2   gate19944  (.A(II25939), .B(II25940), .Z(g19501) ) ;
NAND2   gate19945  (.A(II25922), .B(II25923), .Z(g19480) ) ;
AND3    gate19946  (.A(g19314), .B(g19501), .C(g19480), .Z(II27772) ) ;
NAND2   gate19947  (.A(II25898), .B(II25899), .Z(g19456) ) ;
NAND2   gate19948  (.A(II25866), .B(II25867), .Z(g19430) ) ;
AND3    gate19949  (.A(g19456), .B(g19430), .C(II27772), .Z(g21207) ) ;
AND3    gate19950  (.A(g20150), .B(g16619), .C(g16586), .Z(g21208) ) ;
AND2    gate19951  (.A(g20273), .B(g12412), .Z(g21209) ) ;
AND2    gate19952  (.A(g20242), .B(g12415), .Z(g21210) ) ;
AND2    gate19953  (.A(g20212), .B(g12421), .Z(g21218) ) ;
AND2    gate19954  (.A(g20242), .B(g12426), .Z(g21226) ) ;
AND3    gate19955  (.A(g19578), .B(g14797), .C(g16665), .Z(g21229) ) ;
AND3    gate19956  (.A(g19608), .B(g14849), .C(g16686), .Z(g21234) ) ;
AND3    gate19957  (.A(g19641), .B(g14922), .C(g16712), .Z(g21243) ) ;
NOR2    gate19958  (.A(g16665), .B(g16884), .Z(g20299) ) ;
AND2    gate19959  (.A(g20299), .B(g14837), .Z(g21245) ) ;
AND3    gate19960  (.A(g19681), .B(g15003), .C(g16743), .Z(g21251) ) ;
AND2    gate19961  (.A(g19578), .B(g14895), .Z(g21252) ) ;
NOR2    gate19962  (.A(g16686), .B(g16913), .Z(g20318) ) ;
AND2    gate19963  (.A(g20318), .B(g14910), .Z(g21254) ) ;
AND3    gate19964  (.A(g20299), .B(g16722), .C(g16682), .Z(g21259) ) ;
AND2    gate19965  (.A(g19608), .B(g14976), .Z(g21260) ) ;
NOR2    gate19966  (.A(g16712), .B(g16943), .Z(g20337) ) ;
AND2    gate19967  (.A(g20337), .B(g14991), .Z(g21262) ) ;
AND3    gate19968  (.A(g20318), .B(g16764), .C(g16708), .Z(g21267) ) ;
AND2    gate19969  (.A(g19641), .B(g15065), .Z(g21268) ) ;
NOR2    gate19970  (.A(g16743), .B(g16974), .Z(g20357) ) ;
AND2    gate19971  (.A(g20357), .B(g15080), .Z(g21270) ) ;
AND3    gate19972  (.A(g20337), .B(g16791), .C(g16739), .Z(g21276) ) ;
AND2    gate19973  (.A(g19681), .B(g15161), .Z(g21277) ) ;
AND3    gate19974  (.A(g20357), .B(g16820), .C(g16781), .Z(g21283) ) ;
AND2    gate19975  (.A(g9356), .B(g20269), .Z(g21284) ) ;
AND2    gate19976  (.A(g9356), .B(g20278), .Z(g21290) ) ;
AND2    gate19977  (.A(g9293), .B(g20279), .Z(g21291) ) ;
AND2    gate19978  (.A(g9453), .B(g20281), .Z(g21292) ) ;
AND2    gate19979  (.A(g9356), .B(g20286), .Z(g21298) ) ;
AND2    gate19980  (.A(g9293), .B(g20287), .Z(g21299) ) ;
AND2    gate19981  (.A(g9232), .B(g20288), .Z(g21300) ) ;
AND2    gate19982  (.A(g9453), .B(g20289), .Z(g21301) ) ;
AND2    gate19983  (.A(g9374), .B(g20290), .Z(g21302) ) ;
AND2    gate19984  (.A(g9595), .B(g20292), .Z(g21303) ) ;
AND2    gate19985  (.A(g9293), .B(g20296), .Z(g21304) ) ;
AND2    gate19986  (.A(g9232), .B(g20297), .Z(g21305) ) ;
AND2    gate19987  (.A(g9187), .B(g20298), .Z(g21306) ) ;
AND2    gate19988  (.A(g9453), .B(g20302), .Z(g21307) ) ;
AND2    gate19989  (.A(g9374), .B(g20303), .Z(g21308) ) ;
AND2    gate19990  (.A(g9310), .B(g20304), .Z(g21309) ) ;
AND2    gate19991  (.A(g9595), .B(g20305), .Z(g21310) ) ;
AND2    gate19992  (.A(g9471), .B(g20306), .Z(g21311) ) ;
AND2    gate19993  (.A(g9737), .B(g20308), .Z(g21312) ) ;
AND2    gate19994  (.A(g9232), .B(g20311), .Z(g21313) ) ;
AND2    gate19995  (.A(g9187), .B(g20312), .Z(g21314) ) ;
AND2    gate19996  (.A(g9161), .B(g20313), .Z(g21315) ) ;
AND2    gate19997  (.A(g9374), .B(g20315), .Z(g21319) ) ;
AND2    gate19998  (.A(g9310), .B(g20316), .Z(g21320) ) ;
AND2    gate19999  (.A(g9248), .B(g20317), .Z(g21321) ) ;
AND2    gate20000  (.A(g9595), .B(g20321), .Z(g21322) ) ;
AND2    gate20001  (.A(g9471), .B(g20322), .Z(g21323) ) ;
AND2    gate20002  (.A(g9391), .B(g20323), .Z(g21324) ) ;
AND2    gate20003  (.A(g9737), .B(g20324), .Z(g21325) ) ;
AND2    gate20004  (.A(g9613), .B(g20325), .Z(g21326) ) ;
AND2    gate20005  (.A(g9187), .B(g20327), .Z(g21328) ) ;
AND2    gate20006  (.A(g9161), .B(g20328), .Z(g21329) ) ;
AND2    gate20007  (.A(g9150), .B(g20329), .Z(g21330) ) ;
AND2    gate20008  (.A(g9310), .B(g20330), .Z(g21334) ) ;
AND2    gate20009  (.A(g9248), .B(g20331), .Z(g21335) ) ;
AND2    gate20010  (.A(g9203), .B(g20332), .Z(g21336) ) ;
AND2    gate20011  (.A(g9471), .B(g20334), .Z(g21337) ) ;
AND2    gate20012  (.A(g9391), .B(g20335), .Z(g21338) ) ;
AND2    gate20013  (.A(g9326), .B(g20336), .Z(g21339) ) ;
AND2    gate20014  (.A(g9737), .B(g20340), .Z(g21340) ) ;
AND2    gate20015  (.A(g9613), .B(g20341), .Z(g21341) ) ;
AND2    gate20016  (.A(g9488), .B(g20342), .Z(g21342) ) ;
AND2    gate20017  (.A(g9161), .B(g20344), .Z(g21343) ) ;
AND2    gate20018  (.A(g9150), .B(g20345), .Z(g21344) ) ;
AND2    gate20019  (.A(g15096), .B(g20346), .Z(g21345) ) ;
AND2    gate20020  (.A(g9248), .B(g20347), .Z(g21349) ) ;
AND2    gate20021  (.A(g9203), .B(g20348), .Z(g21350) ) ;
AND2    gate20022  (.A(g9174), .B(g20349), .Z(g21351) ) ;
AND2    gate20023  (.A(g9391), .B(g20350), .Z(g21352) ) ;
AND2    gate20024  (.A(g9326), .B(g20351), .Z(g21353) ) ;
AND2    gate20025  (.A(g9264), .B(g20352), .Z(g21354) ) ;
AND2    gate20026  (.A(g9613), .B(g20354), .Z(g21355) ) ;
AND2    gate20027  (.A(g9488), .B(g20355), .Z(g21356) ) ;
AND2    gate20028  (.A(g9407), .B(g20356), .Z(g21357) ) ;
AND2    gate20029  (.A(g9507), .B(g20361), .Z(g21360) ) ;
AND2    gate20030  (.A(g9150), .B(g20362), .Z(g21361) ) ;
AND2    gate20031  (.A(g15096), .B(g20363), .Z(g21362) ) ;
AND2    gate20032  (.A(g15022), .B(g20364), .Z(g21363) ) ;
AND2    gate20033  (.A(g9203), .B(g20366), .Z(g21367) ) ;
AND2    gate20034  (.A(g9174), .B(g20367), .Z(g21368) ) ;
AND2    gate20035  (.A(g15188), .B(g20368), .Z(g21369) ) ;
AND2    gate20036  (.A(g9326), .B(g20369), .Z(g21370) ) ;
AND2    gate20037  (.A(g9264), .B(g20370), .Z(g21371) ) ;
AND2    gate20038  (.A(g9216), .B(g20371), .Z(g21372) ) ;
AND2    gate20039  (.A(g9488), .B(g20372), .Z(g21373) ) ;
AND2    gate20040  (.A(g9407), .B(g20373), .Z(g21374) ) ;
AND2    gate20041  (.A(g9342), .B(g20374), .Z(g21375) ) ;
AND2    gate20042  (.A(g9507), .B(g20378), .Z(g21378) ) ;
AND2    gate20043  (.A(g9427), .B(g20379), .Z(g21379) ) ;
AND2    gate20044  (.A(g15096), .B(g20380), .Z(g21380) ) ;
AND2    gate20045  (.A(g15022), .B(g20381), .Z(g21381) ) ;
AND2    gate20046  (.A(g6201), .B(g19657), .Z(g21388) ) ;
AND2    gate20047  (.A(g9649), .B(g20384), .Z(g21389) ) ;
AND2    gate20048  (.A(g9174), .B(g20385), .Z(g21390) ) ;
AND2    gate20049  (.A(g15188), .B(g20386), .Z(g21391) ) ;
AND2    gate20050  (.A(g15118), .B(g20387), .Z(g21392) ) ;
AND2    gate20051  (.A(g9264), .B(g20389), .Z(g21393) ) ;
AND2    gate20052  (.A(g9216), .B(g20390), .Z(g21394) ) ;
AND2    gate20053  (.A(g15274), .B(g20391), .Z(g21395) ) ;
AND2    gate20054  (.A(g9407), .B(g20392), .Z(g21396) ) ;
AND2    gate20055  (.A(g9342), .B(g20393), .Z(g21397) ) ;
AND2    gate20056  (.A(g9277), .B(g20394), .Z(g21398) ) ;
AND2    gate20057  (.A(g9507), .B(g20397), .Z(g21401) ) ;
AND2    gate20058  (.A(g9427), .B(g20398), .Z(g21402) ) ;
AND2    gate20059  (.A(g15022), .B(g20399), .Z(g21403) ) ;
AND2    gate20060  (.A(g6363), .B(g20402), .Z(g21410) ) ;
AND2    gate20061  (.A(g9649), .B(g20403), .Z(g21411) ) ;
AND2    gate20062  (.A(g9569), .B(g20404), .Z(g21412) ) ;
AND2    gate20063  (.A(g15188), .B(g20405), .Z(g21413) ) ;
AND2    gate20064  (.A(g15118), .B(g20406), .Z(g21414) ) ;
AND2    gate20065  (.A(g6290), .B(g19705), .Z(g21418) ) ;
AND2    gate20066  (.A(g9795), .B(g20409), .Z(g21419) ) ;
AND2    gate20067  (.A(g9216), .B(g20410), .Z(g21420) ) ;
AND2    gate20068  (.A(g15274), .B(g20411), .Z(g21421) ) ;
AND2    gate20069  (.A(g15210), .B(g20412), .Z(g21422) ) ;
AND2    gate20070  (.A(g9342), .B(g20414), .Z(g21423) ) ;
AND2    gate20071  (.A(g9277), .B(g20415), .Z(g21424) ) ;
AND2    gate20072  (.A(g15366), .B(g20416), .Z(g21425) ) ;
AND2    gate20073  (.A(g9427), .B(g20420), .Z(g21428) ) ;
AND2    gate20074  (.A(g9649), .B(g20422), .Z(g21438) ) ;
AND2    gate20075  (.A(g9569), .B(g20423), .Z(g21439) ) ;
AND2    gate20076  (.A(g15118), .B(g20424), .Z(g21440) ) ;
AND2    gate20077  (.A(g6568), .B(g20427), .Z(g21444) ) ;
AND2    gate20078  (.A(g9795), .B(g20428), .Z(g21445) ) ;
AND2    gate20079  (.A(g9711), .B(g20429), .Z(g21446) ) ;
AND2    gate20080  (.A(g15274), .B(g20430), .Z(g21447) ) ;
AND2    gate20081  (.A(g15210), .B(g20431), .Z(g21448) ) ;
AND2    gate20082  (.A(g6427), .B(g19749), .Z(g21452) ) ;
AND2    gate20083  (.A(g9941), .B(g20434), .Z(g21453) ) ;
AND2    gate20084  (.A(g9277), .B(g20435), .Z(g21454) ) ;
AND2    gate20085  (.A(g15366), .B(g20436), .Z(g21455) ) ;
AND2    gate20086  (.A(g15296), .B(g20437), .Z(g21456) ) ;
AND2    gate20087  (.A(g9569), .B(g20442), .Z(g21476) ) ;
AND2    gate20088  (.A(g9795), .B(g20444), .Z(g21480) ) ;
AND2    gate20089  (.A(g9711), .B(g20445), .Z(g21481) ) ;
AND2    gate20090  (.A(g15210), .B(g20446), .Z(g21482) ) ;
AND2    gate20091  (.A(g6832), .B(g20449), .Z(g21486) ) ;
AND2    gate20092  (.A(g9941), .B(g20450), .Z(g21487) ) ;
AND2    gate20093  (.A(g9857), .B(g20451), .Z(g21488) ) ;
AND2    gate20094  (.A(g15366), .B(g20452), .Z(g21489) ) ;
AND2    gate20095  (.A(g15296), .B(g20453), .Z(g21490) ) ;
AND2    gate20096  (.A(g6632), .B(g19792), .Z(g21494) ) ;
AND2    gate20097  (.A(g3006), .B(g20456), .Z(g21497) ) ;
AND2    gate20098  (.A(g9711), .B(g20461), .Z(g21517) ) ;
AND2    gate20099  (.A(g9941), .B(g20463), .Z(g21521) ) ;
AND2    gate20100  (.A(g9857), .B(g20464), .Z(g21522) ) ;
AND2    gate20101  (.A(g15296), .B(g20465), .Z(g21523) ) ;
AND2    gate20102  (.A(g7134), .B(g20468), .Z(g21527) ) ;
AND3    gate20103  (.A(g17802), .B(g18265), .C(g17882), .Z(II28068) ) ;
AND2    gate20104  (.A(g9857), .B(g20476), .Z(g21553) ) ;
AND3    gate20105  (.A(g13907), .B(g14238), .C(g13946), .Z(II28096) ) ;
AND4    gate20106  (.A(g13886), .B(g14153), .C(g19799), .D(II28096), .Z(g21564) ) ;
AND3    gate20107  (.A(g17914), .B(g18358), .C(g17993), .Z(II28103) ) ;
AND2    gate20108  (.A(g3002), .B(g19890), .Z(g21589) ) ;
AND3    gate20109  (.A(g16498), .B(g19484), .C(g14071), .Z(g21593) ) ;
AND3    gate20110  (.A(g13963), .B(g14360), .C(g14016), .Z(II28126) ) ;
AND4    gate20111  (.A(g13927), .B(g14268), .C(g19843), .D(II28126), .Z(g21597) ) ;
AND3    gate20112  (.A(g18025), .B(g18453), .C(g18110), .Z(II28133) ) ;
AND2    gate20113  (.A(g7522), .B(g20490), .Z(g21610) ) ;
AND2    gate20114  (.A(g7471), .B(g19915), .Z(g21611) ) ;
AND3    gate20115  (.A(g16520), .B(g19505), .C(g14186), .Z(g21622) ) ;
AND3    gate20116  (.A(g14033), .B(g14472), .C(g14107), .Z(II28155) ) ;
AND4    gate20117  (.A(g13983), .B(g14390), .C(g19876), .D(II28155), .Z(g21626) ) ;
AND3    gate20118  (.A(g18142), .B(g18526), .C(g18226), .Z(II28162) ) ;
AND2    gate20119  (.A(g7549), .B(g20496), .Z(g21635) ) ;
AND2    gate20120  (.A(g3398), .B(g20500), .Z(g21639) ) ;
AND3    gate20121  (.A(g16551), .B(g19524), .C(g14301), .Z(g21650) ) ;
AND3    gate20122  (.A(g14124), .B(g14559), .C(g14222), .Z(II28181) ) ;
AND4    gate20123  (.A(g14053), .B(g14502), .C(g19907), .D(II28181), .Z(g21654) ) ;
AND2    gate20124  (.A(g2896), .B(g20501), .Z(g21658) ) ;
AND2    gate20125  (.A(g3398), .B(g20504), .Z(g21666) ) ;
AND2    gate20126  (.A(g3554), .B(g20505), .Z(g21670) ) ;
AND3    gate20127  (.A(g16583), .B(g19534), .C(g14423), .Z(g21681) ) ;
AND2    gate20128  (.A(g3398), .B(g20516), .Z(g21687) ) ;
AND2    gate20129  (.A(g3554), .B(g20517), .Z(g21695) ) ;
AND2    gate20130  (.A(g3710), .B(g20518), .Z(g21699) ) ;
AND2    gate20131  (.A(g2892), .B(g19978), .Z(g21707) ) ;
AND2    gate20132  (.A(g3554), .B(g20534), .Z(g21723) ) ;
AND2    gate20133  (.A(g3710), .B(g20535), .Z(g21731) ) ;
AND2    gate20134  (.A(g3866), .B(g20536), .Z(g21735) ) ;
AND2    gate20135  (.A(g3710), .B(g20553), .Z(g21749) ) ;
AND2    gate20136  (.A(g3866), .B(g20554), .Z(g21757) ) ;
AND2    gate20137  (.A(g7607), .B(g20045), .Z(g21758) ) ;
AND2    gate20138  (.A(g3866), .B(g19078), .Z(g21773) ) ;
AND3    gate20139  (.A(g16679), .B(g19578), .C(g14776), .Z(g21805) ) ;
AND3    gate20140  (.A(g16705), .B(g19608), .C(g14811), .Z(g21812) ) ;
AND3    gate20141  (.A(g16736), .B(g19641), .C(g14863), .Z(g21818) ) ;
AND3    gate20142  (.A(g16778), .B(g19681), .C(g14936), .Z(g21822) ) ;
AND2    gate20143  (.A(g19302), .B(g11749), .Z(g21891) ) ;
NAND3   gate20144  (.A(g14685), .B(g8580), .C(g17057), .Z(g19288) ) ;
AND2    gate20145  (.A(g19288), .B(g13011), .Z(g21892) ) ;
AND2    gate20146  (.A(g19323), .B(g11749), .Z(g21899) ) ;
NAND3   gate20147  (.A(g14719), .B(g8587), .C(g17092), .Z(g19306) ) ;
AND2    gate20148  (.A(g19306), .B(g13011), .Z(g21900) ) ;
AND2    gate20149  (.A(g5715), .B(g20513), .Z(g21906) ) ;
AND2    gate20150  (.A(g19350), .B(g11749), .Z(g21911) ) ;
NAND3   gate20151  (.A(g14747), .B(g8594), .C(g17130), .Z(g19327) ) ;
AND2    gate20152  (.A(g19327), .B(g13011), .Z(g21912) ) ;
AND2    gate20153  (.A(g4456), .B(g20519), .Z(g21913) ) ;
AND2    gate20154  (.A(g5773), .B(g20531), .Z(g21920) ) ;
AND2    gate20155  (.A(g19384), .B(g11749), .Z(g21925) ) ;
NAND3   gate20156  (.A(g14768), .B(g8605), .C(g17157), .Z(g19354) ) ;
AND2    gate20157  (.A(g19354), .B(g13011), .Z(g21926) ) ;
AND2    gate20158  (.A(g4632), .B(g20539), .Z(g21931) ) ;
AND2    gate20159  (.A(g5832), .B(g20550), .Z(g21938) ) ;
AND2    gate20160  (.A(g291), .B(g21187), .Z(g21990) ) ;
AND2    gate20161  (.A(g978), .B(g21202), .Z(g22004) ) ;
AND2    gate20162  (.A(g1672), .B(g21217), .Z(g22015) ) ;
AND2    gate20163  (.A(g2366), .B(g21225), .Z(g22020) ) ;
NAND2   gate20164  (.A(g3088), .B(g16825), .Z(g19141) ) ;
NOR3    gate20165  (.A(g20108), .B(g20132), .C(g20156), .Z(g21133) ) ;
NOR3    gate20166  (.A(g20086), .B(g20107), .C(g20131), .Z(g21116) ) ;
AND3    gate20167  (.A(g19141), .B(g21133), .C(g21116), .Z(II28582) ) ;
NOR3    gate20168  (.A(g20050), .B(g20085), .C(g20106), .Z(g21104) ) ;
NOR3    gate20169  (.A(g20012), .B(g20049), .C(g20084), .Z(g21095) ) ;
NOR2    gate20170  (.A(g20011), .B(g20048), .Z(g21084) ) ;
NOR2    gate20171  (.A(g20159), .B(g20189), .Z(g21167) ) ;
NOR3    gate20172  (.A(g20135), .B(g20158), .C(g20188), .Z(g21147) ) ;
NOR3    gate20173  (.A(g20111), .B(g20134), .C(g20157), .Z(g21134) ) ;
AND3    gate20174  (.A(g21167), .B(g21147), .C(g21134), .Z(II28594) ) ;
NOR3    gate20175  (.A(g20089), .B(g20110), .C(g20133), .Z(g21117) ) ;
NOR3    gate20176  (.A(g20052), .B(g20088), .C(g20109), .Z(g21105) ) ;
NOR3    gate20177  (.A(g20013), .B(g20051), .C(g20087), .Z(g21096) ) ;
NOR2    gate20178  (.A(g20192), .B(g20221), .Z(g21183) ) ;
NOR3    gate20179  (.A(g20162), .B(g20191), .C(g20220), .Z(g21168) ) ;
NOR3    gate20180  (.A(g20138), .B(g20161), .C(g20190), .Z(g21148) ) ;
AND3    gate20181  (.A(g21183), .B(g21168), .C(g21148), .Z(II28609) ) ;
NOR3    gate20182  (.A(g20114), .B(g20137), .C(g20160), .Z(g21135) ) ;
NOR3    gate20183  (.A(g20091), .B(g20113), .C(g20136), .Z(g21118) ) ;
NOR3    gate20184  (.A(g20053), .B(g20090), .C(g20112), .Z(g21106) ) ;
AND2    gate20185  (.A(g21564), .B(g20986), .Z(g22187) ) ;
AND2    gate20186  (.A(g21597), .B(g21012), .Z(g22196) ) ;
AND2    gate20187  (.A(g21271), .B(g16881), .Z(g22201) ) ;
AND2    gate20188  (.A(g21626), .B(g21036), .Z(g22202) ) ;
AND2    gate20189  (.A(g21895), .B(g11976), .Z(g22206) ) ;
AND2    gate20190  (.A(g21278), .B(g16910), .Z(g22207) ) ;
AND2    gate20191  (.A(g21654), .B(g21057), .Z(g22208) ) ;
AND2    gate20192  (.A(g21661), .B(g12027), .Z(g22211) ) ;
AND2    gate20193  (.A(g21907), .B(g12045), .Z(g22214) ) ;
AND2    gate20194  (.A(g21285), .B(g16940), .Z(g22215) ) ;
AND2    gate20195  (.A(g21690), .B(g12091), .Z(g22220) ) ;
AND2    gate20196  (.A(g21921), .B(g12109), .Z(g22223) ) ;
AND2    gate20197  (.A(g21293), .B(g16971), .Z(g22224) ) ;
AND2    gate20198  (.A(g21716), .B(g12136), .Z(g22228) ) ;
AND2    gate20199  (.A(g21661), .B(g12139), .Z(g22229) ) ;
AND2    gate20200  (.A(g21726), .B(g12163), .Z(g22235) ) ;
AND2    gate20201  (.A(g21939), .B(g12181), .Z(g22238) ) ;
AND2    gate20202  (.A(g21742), .B(g12198), .Z(g22244) ) ;
AND2    gate20203  (.A(g21690), .B(g12201), .Z(g22245) ) ;
AND2    gate20204  (.A(g21752), .B(g12225), .Z(g22250) ) ;
AND2    gate20205  (.A(g21716), .B(g12239), .Z(g22254) ) ;
AND2    gate20206  (.A(g21661), .B(g12242), .Z(g22255) ) ;
AND2    gate20207  (.A(g21766), .B(g12253), .Z(g22264) ) ;
AND2    gate20208  (.A(g21726), .B(g12256), .Z(g22265) ) ;
AND2    gate20209  (.A(g92), .B(g21529), .Z(g22270) ) ;
AND2    gate20210  (.A(g21742), .B(g12282), .Z(g22272) ) ;
AND2    gate20211  (.A(g21690), .B(g12285), .Z(g22273) ) ;
AND2    gate20212  (.A(g21782), .B(g12296), .Z(g22281) ) ;
AND2    gate20213  (.A(g21752), .B(g12299), .Z(g22282) ) ;
AND2    gate20214  (.A(g21716), .B(g12312), .Z(g22285) ) ;
AND2    gate20215  (.A(g780), .B(g21565), .Z(g22289) ) ;
AND2    gate20216  (.A(g21766), .B(g12318), .Z(g22291) ) ;
AND2    gate20217  (.A(g21726), .B(g12321), .Z(g22292) ) ;
AND2    gate20218  (.A(g21742), .B(g12340), .Z(g22305) ) ;
AND2    gate20219  (.A(g1466), .B(g21598), .Z(g22309) ) ;
AND2    gate20220  (.A(g21782), .B(g12346), .Z(g22311) ) ;
AND2    gate20221  (.A(g21752), .B(g12349), .Z(g22312) ) ;
AND2    gate20222  (.A(g21766), .B(g12370), .Z(g22333) ) ;
AND2    gate20223  (.A(g2160), .B(g21627), .Z(g22337) ) ;
AND2    gate20224  (.A(g88), .B(g21184), .Z(g22340) ) ;
AND2    gate20225  (.A(g21782), .B(g12389), .Z(g22358) ) ;
AND2    gate20226  (.A(g776), .B(g21199), .Z(g22363) ) ;
AND2    gate20227  (.A(g1462), .B(g21214), .Z(g22383) ) ;
AND2    gate20228  (.A(g2156), .B(g21222), .Z(g22398) ) ;
AND2    gate20229  (.A(g646), .B(g21861), .Z(g22483) ) ;
AND2    gate20230  (.A(g13873), .B(g21382), .Z(g22515) ) ;
AND2    gate20231  (.A(g20885), .B(g17442), .Z(g22516) ) ;
AND2    gate20232  (.A(g21895), .B(g12608), .Z(g22517) ) ;
AND2    gate20233  (.A(g1332), .B(g21867), .Z(g22526) ) ;
AND2    gate20234  (.A(g13886), .B(g21404), .Z(g22546) ) ;
AND2    gate20235  (.A(g13895), .B(g21415), .Z(g22555) ) ;
AND2    gate20236  (.A(g20904), .B(g17523), .Z(g22556) ) ;
AND2    gate20237  (.A(g21907), .B(g12654), .Z(g22557) ) ;
AND2    gate20238  (.A(g2026), .B(g21872), .Z(g22566) ) ;
AND2    gate20239  (.A(g13907), .B(g21429), .Z(g22577) ) ;
AND2    gate20240  (.A(g21895), .B(g12699), .Z(g22581) ) ;
AND2    gate20241  (.A(g13927), .B(g21441), .Z(g22587) ) ;
AND2    gate20242  (.A(g13936), .B(g21449), .Z(g22595) ) ;
AND2    gate20243  (.A(g20928), .B(g17613), .Z(g22596) ) ;
AND2    gate20244  (.A(g21921), .B(g12708), .Z(g22597) ) ;
AND2    gate20245  (.A(g2720), .B(g21876), .Z(g22606) ) ;
AND2    gate20246  (.A(g13946), .B(g21458), .Z(g22607) ) ;
AND2    gate20247  (.A(g660), .B(g21473), .Z(g22610) ) ;
AND2    gate20248  (.A(g13963), .B(g21477), .Z(g22614) ) ;
AND2    gate20249  (.A(g21907), .B(g12756), .Z(g22618) ) ;
AND2    gate20250  (.A(g13983), .B(g21483), .Z(g22624) ) ;
AND2    gate20251  (.A(g13992), .B(g21491), .Z(g22632) ) ;
AND2    gate20252  (.A(g20956), .B(g17710), .Z(g22633) ) ;
AND2    gate20253  (.A(g21939), .B(g12765), .Z(g22634) ) ;
NOR2    gate20254  (.A(g14767), .B(g19552), .Z(g20841) ) ;
AND2    gate20255  (.A(g20841), .B(g10927), .Z(g22637) ) ;
AND2    gate20256  (.A(g14001), .B(g21498), .Z(g22638) ) ;
AND2    gate20257  (.A(g14016), .B(g21505), .Z(g22643) ) ;
AND2    gate20258  (.A(g1346), .B(g21514), .Z(g22646) ) ;
AND2    gate20259  (.A(g14033), .B(g21518), .Z(g22650) ) ;
AND2    gate20260  (.A(g21921), .B(g12798), .Z(g22654) ) ;
AND2    gate20261  (.A(g14053), .B(g21524), .Z(g22660) ) ;
NOR2    gate20262  (.A(g19691), .B(g19726), .Z(g20920) ) ;
AND2    gate20263  (.A(g20920), .B(g6153), .Z(g22665) ) ;
AND2    gate20264  (.A(g21825), .B(g20014), .Z(g22666) ) ;
AND2    gate20265  (.A(g14062), .B(g21530), .Z(g22667) ) ;
AND2    gate20266  (.A(g14092), .B(g21537), .Z(g22674) ) ;
AND2    gate20267  (.A(g14107), .B(g21541), .Z(g22679) ) ;
AND2    gate20268  (.A(g2040), .B(g21550), .Z(g22682) ) ;
AND2    gate20269  (.A(g14124), .B(g21554), .Z(g22686) ) ;
AND2    gate20270  (.A(g21939), .B(g12837), .Z(g22690) ) ;
AND2    gate20271  (.A(g7338), .B(g21883), .Z(g22699) ) ;
AND2    gate20272  (.A(g7146), .B(g21558), .Z(g22700) ) ;
AND2    gate20273  (.A(g18174), .B(g21561), .Z(g22701) ) ;
AND2    gate20274  (.A(g14177), .B(g21566), .Z(g22707) ) ;
AND2    gate20275  (.A(g14207), .B(g21573), .Z(g22714) ) ;
AND2    gate20276  (.A(g14222), .B(g21577), .Z(g22719) ) ;
AND2    gate20277  (.A(g2734), .B(g21586), .Z(g22722) ) ;
AND2    gate20278  (.A(g3036), .B(g21886), .Z(g22726) ) ;
AND2    gate20279  (.A(g14238), .B(g21590), .Z(g22727) ) ;
AND2    gate20280  (.A(g18281), .B(g21594), .Z(g22732) ) ;
AND2    gate20281  (.A(g14292), .B(g21599), .Z(g22738) ) ;
AND2    gate20282  (.A(g14322), .B(g21606), .Z(g22745) ) ;
AND2    gate20283  (.A(g14342), .B(g21612), .Z(g22754) ) ;
AND2    gate20284  (.A(g14360), .B(g21619), .Z(g22759) ) ;
AND2    gate20285  (.A(g18374), .B(g21623), .Z(g22764) ) ;
AND2    gate20286  (.A(g14414), .B(g21628), .Z(g22770) ) ;
AND2    gate20287  (.A(g14454), .B(g21640), .Z(g22788) ) ;
AND2    gate20288  (.A(g14472), .B(g21647), .Z(g22793) ) ;
AND2    gate20289  (.A(g18469), .B(g21651), .Z(g22798) ) ;
AND2    gate20290  (.A(g2920), .B(g21655), .Z(g22804) ) ;
AND2    gate20291  (.A(g14541), .B(g21671), .Z(g22830) ) ;
AND2    gate20292  (.A(g14559), .B(g21678), .Z(g22835) ) ;
AND2    gate20293  (.A(g7583), .B(g21902), .Z(g22841) ) ;
AND2    gate20294  (.A(g3032), .B(g21682), .Z(g22842) ) ;
AND2    gate20295  (.A(g14596), .B(g21700), .Z(g22869) ) ;
AND2    gate20296  (.A(g7587), .B(g21708), .Z(g22874) ) ;
AND2    gate20297  (.A(g2924), .B(g21927), .Z(g22906) ) ;
AND2    gate20298  (.A(g16840), .B(g21400), .Z(g22984) ) ;
AND2    gate20299  (.A(g20842), .B(g15859), .Z(g23104) ) ;
AND2    gate20300  (.A(g5857), .B(g21050), .Z(g23106) ) ;
AND2    gate20301  (.A(g20850), .B(g15890), .Z(g23118) ) ;
AND2    gate20302  (.A(g5904), .B(g21069), .Z(g23119) ) ;
AND2    gate20303  (.A(g20858), .B(g15923), .Z(g23127) ) ;
AND2    gate20304  (.A(g5943), .B(g21079), .Z(g23128) ) ;
AND2    gate20305  (.A(g20866), .B(g15952), .Z(g23138) ) ;
AND2    gate20306  (.A(g5977), .B(g21093), .Z(g23139) ) ;
AND2    gate20307  (.A(g21533), .B(g22408), .Z(g23409) ) ;
AND2    gate20308  (.A(g21569), .B(g22421), .Z(g23414) ) ;
NOR2    gate20309  (.A(g21271), .B(g20842), .Z(g22755) ) ;
AND2    gate20310  (.A(g22755), .B(g19577), .Z(g23419) ) ;
AND2    gate20311  (.A(g21602), .B(g22443), .Z(g23423) ) ;
NOR2    gate20312  (.A(g21278), .B(g20850), .Z(g22789) ) ;
AND2    gate20313  (.A(g22789), .B(g19607), .Z(g23428) ) ;
AND2    gate20314  (.A(g21631), .B(g22476), .Z(g23432) ) ;
NOR2    gate20315  (.A(g21285), .B(g20858), .Z(g22831) ) ;
AND2    gate20316  (.A(g22831), .B(g19640), .Z(g23434) ) ;
NOR2    gate20317  (.A(g21293), .B(g20866), .Z(g22870) ) ;
AND2    gate20318  (.A(g22870), .B(g19680), .Z(g23440) ) ;
AND2    gate20319  (.A(g18552), .B(g22547), .Z(g23451) ) ;
AND2    gate20320  (.A(g18602), .B(g22588), .Z(g23458) ) ;
AND2    gate20321  (.A(g17988), .B(g22609), .Z(g23462) ) ;
AND2    gate20322  (.A(g18634), .B(g22625), .Z(g23467) ) ;
AND2    gate20323  (.A(g18105), .B(g22645), .Z(g23471) ) ;
AND2    gate20324  (.A(g18643), .B(g22661), .Z(g23476) ) ;
AND2    gate20325  (.A(g22945), .B(g8847), .Z(g23483) ) ;
AND2    gate20326  (.A(g18221), .B(g22681), .Z(g23484) ) ;
AND2    gate20327  (.A(g18328), .B(g22721), .Z(g23494) ) ;
AND2    gate20328  (.A(g5802), .B(g22300), .Z(g23496) ) ;
AND2    gate20329  (.A(g5890), .B(g22753), .Z(g23510) ) ;
AND2    gate20330  (.A(g5858), .B(g22328), .Z(g23512) ) ;
AND2    gate20331  (.A(g5929), .B(g22787), .Z(g23525) ) ;
AND2    gate20332  (.A(g5905), .B(g22353), .Z(g23527) ) ;
AND2    gate20333  (.A(g5963), .B(g22829), .Z(g23536) ) ;
AND2    gate20334  (.A(g5944), .B(g22376), .Z(g23538) ) ;
AND2    gate20335  (.A(g5992), .B(g22868), .Z(g23544) ) ;
AND2    gate20336  (.A(g8062), .B(g22405), .Z(g23547) ) ;
AND2    gate20337  (.A(g8132), .B(g22409), .Z(g23550) ) ;
AND2    gate20338  (.A(g8135), .B(g22412), .Z(g23551) ) ;
AND2    gate20339  (.A(g6136), .B(g22415), .Z(g23552) ) ;
AND2    gate20340  (.A(g8147), .B(g22418), .Z(g23554) ) ;
AND2    gate20341  (.A(g8200), .B(g22422), .Z(g23558) ) ;
AND2    gate20342  (.A(g8203), .B(g22425), .Z(g23559) ) ;
AND2    gate20343  (.A(g8206), .B(g22428), .Z(g23560) ) ;
AND2    gate20344  (.A(g8218), .B(g22431), .Z(g23563) ) ;
AND2    gate20345  (.A(g8221), .B(g22434), .Z(g23564) ) ;
AND2    gate20346  (.A(g6146), .B(g22437), .Z(g23565) ) ;
AND2    gate20347  (.A(g8233), .B(g22440), .Z(g23567) ) ;
AND2    gate20348  (.A(g3931), .B(g22445), .Z(g23571) ) ;
AND2    gate20349  (.A(g3934), .B(g22448), .Z(g23572) ) ;
AND2    gate20350  (.A(g3937), .B(g22451), .Z(g23573) ) ;
AND2    gate20351  (.A(g3957), .B(g22455), .Z(g23577) ) ;
AND2    gate20352  (.A(g3960), .B(g22458), .Z(g23578) ) ;
AND2    gate20353  (.A(g3963), .B(g22461), .Z(g23579) ) ;
AND2    gate20354  (.A(g3975), .B(g22464), .Z(g23582) ) ;
AND2    gate20355  (.A(g3978), .B(g22467), .Z(g23583) ) ;
AND2    gate20356  (.A(g6167), .B(g22470), .Z(g23584) ) ;
AND2    gate20357  (.A(g3990), .B(g22473), .Z(g23586) ) ;
AND2    gate20358  (.A(g4009), .B(g22477), .Z(g23590) ) ;
AND2    gate20359  (.A(g4012), .B(g22480), .Z(g23591) ) ;
AND2    gate20360  (.A(g17640), .B(g22986), .Z(g23592) ) ;
NAND2   gate20361  (.A(g19441), .B(g20885), .Z(g22845) ) ;
AND2    gate20362  (.A(g22845), .B(g20365), .Z(g23593) ) ;
AND2    gate20363  (.A(g4038), .B(g22484), .Z(g23598) ) ;
AND2    gate20364  (.A(g4041), .B(g22487), .Z(g23599) ) ;
AND2    gate20365  (.A(g4044), .B(g22490), .Z(g23600) ) ;
AND2    gate20366  (.A(g4064), .B(g22494), .Z(g23604) ) ;
AND2    gate20367  (.A(g4067), .B(g22497), .Z(g23605) ) ;
AND2    gate20368  (.A(g4070), .B(g22500), .Z(g23606) ) ;
AND2    gate20369  (.A(g4082), .B(g22503), .Z(g23609) ) ;
AND2    gate20370  (.A(g4085), .B(g22506), .Z(g23610) ) ;
AND2    gate20371  (.A(g6194), .B(g22509), .Z(g23611) ) ;
AND2    gate20372  (.A(g4107), .B(g22512), .Z(g23615) ) ;
AND2    gate20373  (.A(g17724), .B(g22988), .Z(g23616) ) ;
NOR3    gate20374  (.A(g16075), .B(g20842), .C(g21271), .Z(g22810) ) ;
AND2    gate20375  (.A(g22810), .B(g20382), .Z(g23617) ) ;
NAND2   gate20376  (.A(g20842), .B(g20885), .Z(g22608) ) ;
AND2    gate20377  (.A(g22608), .B(g20383), .Z(g23618) ) ;
AND2    gate20378  (.A(g4136), .B(g22520), .Z(g23622) ) ;
AND2    gate20379  (.A(g4139), .B(g22523), .Z(g23623) ) ;
AND2    gate20380  (.A(g17741), .B(g22989), .Z(g23624) ) ;
NAND2   gate20381  (.A(g19468), .B(g20904), .Z(g22880) ) ;
AND2    gate20382  (.A(g22880), .B(g20388), .Z(g23625) ) ;
AND2    gate20383  (.A(g4165), .B(g22527), .Z(g23630) ) ;
AND2    gate20384  (.A(g4168), .B(g22530), .Z(g23631) ) ;
AND2    gate20385  (.A(g4171), .B(g22533), .Z(g23632) ) ;
AND2    gate20386  (.A(g4191), .B(g22537), .Z(g23636) ) ;
AND2    gate20387  (.A(g4194), .B(g22540), .Z(g23637) ) ;
AND2    gate20388  (.A(g4197), .B(g22543), .Z(g23638) ) ;
AND2    gate20389  (.A(g21825), .B(g22805), .Z(g23639) ) ;
AND2    gate20390  (.A(g17802), .B(g22991), .Z(g23643) ) ;
NOR2    gate20391  (.A(g16075), .B(g20885), .Z(g22784) ) ;
AND2    gate20392  (.A(g22784), .B(g17500), .Z(g23659) ) ;
AND2    gate20393  (.A(g4246), .B(g22552), .Z(g23664) ) ;
AND2    gate20394  (.A(g17825), .B(g22995), .Z(g23665) ) ;
NOR3    gate20395  (.A(g16113), .B(g20850), .C(g21278), .Z(g22851) ) ;
AND2    gate20396  (.A(g22851), .B(g20407), .Z(g23666) ) ;
NAND2   gate20397  (.A(g20850), .B(g20904), .Z(g22644) ) ;
AND2    gate20398  (.A(g22644), .B(g20408), .Z(g23667) ) ;
AND2    gate20399  (.A(g4275), .B(g22560), .Z(g23671) ) ;
AND2    gate20400  (.A(g4278), .B(g22563), .Z(g23672) ) ;
AND2    gate20401  (.A(g17842), .B(g22996), .Z(g23673) ) ;
NAND2   gate20402  (.A(g19491), .B(g20928), .Z(g22915) ) ;
AND2    gate20403  (.A(g22915), .B(g20413), .Z(g23674) ) ;
AND2    gate20404  (.A(g4304), .B(g22567), .Z(g23679) ) ;
AND2    gate20405  (.A(g4307), .B(g22570), .Z(g23680) ) ;
AND2    gate20406  (.A(g4310), .B(g22573), .Z(g23681) ) ;
AND2    gate20407  (.A(g17882), .B(g22998), .Z(g23686) ) ;
NAND2   gate20408  (.A(g16075), .B(g21271), .Z(g22668) ) ;
AND2    gate20409  (.A(g22668), .B(g17570), .Z(g23687) ) ;
AND2    gate20410  (.A(g6513), .B(g23001), .Z(g23689) ) ;
AND2    gate20411  (.A(g17914), .B(g23002), .Z(g23693) ) ;
NOR2    gate20412  (.A(g16113), .B(g20904), .Z(g22826) ) ;
AND2    gate20413  (.A(g22826), .B(g17591), .Z(g23709) ) ;
AND2    gate20414  (.A(g4401), .B(g22592), .Z(g23714) ) ;
AND2    gate20415  (.A(g17937), .B(g23006), .Z(g23715) ) ;
NOR3    gate20416  (.A(g16164), .B(g20858), .C(g21285), .Z(g22886) ) ;
AND2    gate20417  (.A(g22886), .B(g20432), .Z(g23716) ) ;
NAND2   gate20418  (.A(g20858), .B(g20928), .Z(g22680) ) ;
AND2    gate20419  (.A(g22680), .B(g20433), .Z(g23717) ) ;
AND2    gate20420  (.A(g4430), .B(g22600), .Z(g23721) ) ;
AND2    gate20421  (.A(g4433), .B(g22603), .Z(g23722) ) ;
AND2    gate20422  (.A(g17954), .B(g23007), .Z(g23723) ) ;
NAND2   gate20423  (.A(g19512), .B(g20956), .Z(g22940) ) ;
AND2    gate20424  (.A(g22940), .B(g20438), .Z(g23724) ) ;
AND2    gate20425  (.A(g21825), .B(g22843), .Z(g23726) ) ;
AND2    gate20426  (.A(g17974), .B(g23008), .Z(g23734) ) ;
AND2    gate20427  (.A(g22949), .B(g9450), .Z(g23735) ) ;
AND2    gate20428  (.A(g17993), .B(g23012), .Z(g23740) ) ;
NAND2   gate20429  (.A(g16113), .B(g21278), .Z(g22708) ) ;
AND2    gate20430  (.A(g22708), .B(g17667), .Z(g23741) ) ;
AND2    gate20431  (.A(g6777), .B(g23015), .Z(g23743) ) ;
AND2    gate20432  (.A(g18025), .B(g23016), .Z(g23747) ) ;
NOR2    gate20433  (.A(g16164), .B(g20928), .Z(g22865) ) ;
AND2    gate20434  (.A(g22865), .B(g17688), .Z(g23763) ) ;
AND2    gate20435  (.A(g4570), .B(g22629), .Z(g23768) ) ;
AND2    gate20436  (.A(g18048), .B(g23020), .Z(g23769) ) ;
NOR3    gate20437  (.A(g16223), .B(g20866), .C(g21293), .Z(g22921) ) ;
AND2    gate20438  (.A(g22921), .B(g20454), .Z(g23770) ) ;
NAND2   gate20439  (.A(g20866), .B(g20956), .Z(g22720) ) ;
AND2    gate20440  (.A(g22720), .B(g20455), .Z(g23771) ) ;
AND2    gate20441  (.A(g21825), .B(g22875), .Z(g23772) ) ;
AND2    gate20442  (.A(g18074), .B(g23021), .Z(g23776) ) ;
AND2    gate20443  (.A(g22949), .B(g9528), .Z(g23777) ) ;
AND2    gate20444  (.A(g22954), .B(g9531), .Z(g23778) ) ;
AND2    gate20445  (.A(g18091), .B(g23024), .Z(g23789) ) ;
AND2    gate20446  (.A(g22958), .B(g9592), .Z(g23790) ) ;
AND2    gate20447  (.A(g18110), .B(g23028), .Z(g23795) ) ;
NAND2   gate20448  (.A(g16164), .B(g21285), .Z(g22739) ) ;
AND2    gate20449  (.A(g22739), .B(g17767), .Z(g23796) ) ;
AND2    gate20450  (.A(g7079), .B(g23031), .Z(g23798) ) ;
AND2    gate20451  (.A(g18142), .B(g23032), .Z(g23802) ) ;
NOR2    gate20452  (.A(g16223), .B(g20956), .Z(g22900) ) ;
AND2    gate20453  (.A(g22900), .B(g17788), .Z(g23818) ) ;
AND2    gate20454  (.A(g3013), .B(g23036), .Z(g23820) ) ;
AND2    gate20455  (.A(g14148), .B(g23037), .Z(g23822) ) ;
AND2    gate20456  (.A(g22949), .B(g9641), .Z(g23824) ) ;
AND2    gate20457  (.A(g22954), .B(g9644), .Z(g23825) ) ;
AND2    gate20458  (.A(g18190), .B(g23038), .Z(g23829) ) ;
AND2    gate20459  (.A(g22958), .B(g9670), .Z(g23830) ) ;
AND2    gate20460  (.A(g22962), .B(g9673), .Z(g23831) ) ;
AND2    gate20461  (.A(g18207), .B(g23041), .Z(g23842) ) ;
AND2    gate20462  (.A(g22966), .B(g9734), .Z(g23843) ) ;
AND2    gate20463  (.A(g18226), .B(g23045), .Z(g23848) ) ;
NAND2   gate20464  (.A(g16223), .B(g21293), .Z(g22771) ) ;
AND2    gate20465  (.A(g22771), .B(g17868), .Z(g23849) ) ;
AND2    gate20466  (.A(g7329), .B(g23048), .Z(g23851) ) ;
NOR2    gate20467  (.A(g17719), .B(g15453), .Z(g19179) ) ;
AND2    gate20468  (.A(g19179), .B(g22696), .Z(g23852) ) ;
AND2    gate20469  (.A(g18265), .B(g23049), .Z(g23854) ) ;
AND2    gate20470  (.A(g22954), .B(g9767), .Z(g23855) ) ;
AND2    gate20471  (.A(g14263), .B(g23056), .Z(g23857) ) ;
AND2    gate20472  (.A(g22958), .B(g9787), .Z(g23859) ) ;
AND2    gate20473  (.A(g22962), .B(g9790), .Z(g23860) ) ;
AND2    gate20474  (.A(g18297), .B(g23057), .Z(g23864) ) ;
AND2    gate20475  (.A(g22966), .B(g9816), .Z(g23865) ) ;
AND2    gate20476  (.A(g22971), .B(g9819), .Z(g23866) ) ;
AND2    gate20477  (.A(g18314), .B(g23060), .Z(g23877) ) ;
AND2    gate20478  (.A(g22975), .B(g9880), .Z(g23878) ) ;
AND2    gate20479  (.A(g18341), .B(g23064), .Z(g23886) ) ;
AND2    gate20480  (.A(g18358), .B(g23069), .Z(g23888) ) ;
AND2    gate20481  (.A(g22962), .B(g9913), .Z(g23889) ) ;
AND2    gate20482  (.A(g14385), .B(g23074), .Z(g23891) ) ;
AND2    gate20483  (.A(g22966), .B(g9933), .Z(g23893) ) ;
AND2    gate20484  (.A(g22971), .B(g9936), .Z(g23894) ) ;
AND2    gate20485  (.A(g18390), .B(g23075), .Z(g23898) ) ;
AND2    gate20486  (.A(g22975), .B(g9962), .Z(g23899) ) ;
AND2    gate20487  (.A(g22980), .B(g9965), .Z(g23900) ) ;
AND2    gate20488  (.A(g3010), .B(g22750), .Z(g23904) ) ;
AND2    gate20489  (.A(g18436), .B(g23079), .Z(g23907) ) ;
AND2    gate20490  (.A(g18453), .B(g23082), .Z(g23909) ) ;
AND2    gate20491  (.A(g22971), .B(g10067), .Z(g23910) ) ;
AND2    gate20492  (.A(g14497), .B(g23087), .Z(g23912) ) ;
AND2    gate20493  (.A(g22975), .B(g10087), .Z(g23914) ) ;
AND2    gate20494  (.A(g22980), .B(g10090), .Z(g23915) ) ;
AND2    gate20495  (.A(g7545), .B(g23088), .Z(g23917) ) ;
AND2    gate20496  (.A(g18509), .B(g23095), .Z(g23939) ) ;
AND2    gate20497  (.A(g18526), .B(g23098), .Z(g23941) ) ;
AND2    gate20498  (.A(g22980), .B(g10176), .Z(g23942) ) ;
AND2    gate20499  (.A(g7570), .B(g23103), .Z(g23944) ) ;
AND2    gate20500  (.A(g18573), .B(g23112), .Z(g23971) ) ;
AND2    gate20501  (.A(g2903), .B(g23115), .Z(g23972) ) ;
AND2    gate20502  (.A(g2900), .B(g22903), .Z(g24029) ) ;
AND2    gate20503  (.A(g22014), .B(g10969), .Z(g24211) ) ;
AND2    gate20504  (.A(g22825), .B(g10999), .Z(g24217) ) ;
AND2    gate20505  (.A(g22979), .B(g11042), .Z(g24221) ) ;
AND2    gate20506  (.A(g22219), .B(g11045), .Z(g24224) ) ;
AND2    gate20507  (.A(g22232), .B(g11105), .Z(g24229) ) ;
AND2    gate20508  (.A(g22243), .B(g11157), .Z(g24236) ) ;
AND2    gate20509  (.A(g22259), .B(g11228), .Z(g24241) ) ;
AND2    gate20510  (.A(g21982), .B(g11291), .Z(g24246) ) ;
AND2    gate20511  (.A(g22551), .B(g11297), .Z(g24247) ) ;
AND2    gate20512  (.A(g21995), .B(g11370), .Z(g24253) ) ;
AND2    gate20513  (.A(g22003), .B(g11438), .Z(g24256) ) ;
AND3    gate20514  (.A(g17086), .B(g24134), .C(g13626), .Z(g24427) ) ;
AND2    gate20515  (.A(g24115), .B(g13614), .Z(g24429) ) ;
AND3    gate20516  (.A(g17124), .B(g24153), .C(g13637), .Z(g24431) ) ;
AND3    gate20517  (.A(g14642), .B(g15904), .C(g24115), .Z(g24432) ) ;
AND2    gate20518  (.A(g24134), .B(g13626), .Z(g24433) ) ;
AND3    gate20519  (.A(g17151), .B(g24168), .C(g13649), .Z(g24435) ) ;
AND3    gate20520  (.A(g14669), .B(g15933), .C(g24134), .Z(g24436) ) ;
AND2    gate20521  (.A(g24153), .B(g13637), .Z(g24437) ) ;
AND3    gate20522  (.A(g14703), .B(g15962), .C(g24153), .Z(g24439) ) ;
AND2    gate20523  (.A(g24168), .B(g13649), .Z(g24440) ) ;
AND3    gate20524  (.A(g14737), .B(g15981), .C(g24168), .Z(g24441) ) ;
NOR2    gate20525  (.A(g22984), .B(g20285), .Z(g23545) ) ;
NOR3    gate20526  (.A(g20092), .B(g20115), .C(g20139), .Z(g21119) ) ;
NOR3    gate20527  (.A(g18414), .B(g18485), .C(g20295), .Z(g21227) ) ;
AND3    gate20528  (.A(g19933), .B(g17896), .C(g23403), .Z(g24529) ) ;
AND3    gate20529  (.A(g18548), .B(g23089), .C(g23403), .Z(g24540) ) ;
AND3    gate20530  (.A(g23420), .B(g17896), .C(g23052), .Z(g24541) ) ;
AND3    gate20531  (.A(g19950), .B(g18007), .C(g23410), .Z(g24542) ) ;
AND3    gate20532  (.A(g18548), .B(g23420), .C(g19948), .Z(g24550) ) ;
AND3    gate20533  (.A(g18598), .B(g23107), .C(g23410), .Z(g24552) ) ;
AND3    gate20534  (.A(g23429), .B(g18007), .C(g23071), .Z(g24553) ) ;
AND3    gate20535  (.A(g19977), .B(g18124), .C(g23415), .Z(g24554) ) ;
AND2    gate20536  (.A(g79), .B(g23448), .Z(g24559) ) ;
AND3    gate20537  (.A(g18598), .B(g23429), .C(g19975), .Z(g24561) ) ;
AND3    gate20538  (.A(g18630), .B(g23120), .C(g23415), .Z(g24563) ) ;
AND3    gate20539  (.A(g23435), .B(g18124), .C(g23084), .Z(g24564) ) ;
AND3    gate20540  (.A(g20007), .B(g18240), .C(g23424), .Z(g24565) ) ;
AND2    gate20541  (.A(g767), .B(g23455), .Z(g24569) ) ;
AND3    gate20542  (.A(g18630), .B(g23435), .C(g20005), .Z(g24571) ) ;
AND3    gate20543  (.A(g18639), .B(g23129), .C(g23424), .Z(g24573) ) ;
AND3    gate20544  (.A(g23441), .B(g18240), .C(g23100), .Z(g24574) ) ;
AND2    gate20545  (.A(g1453), .B(g23464), .Z(g24578) ) ;
AND3    gate20546  (.A(g18639), .B(g23441), .C(g20043), .Z(g24580) ) ;
AND2    gate20547  (.A(g2147), .B(g23473), .Z(g24585) ) ;
AND2    gate20548  (.A(g23486), .B(g23478), .Z(g24590) ) ;
AND2    gate20549  (.A(g83), .B(g23853), .Z(g24591) ) ;
AND2    gate20550  (.A(g23502), .B(g23489), .Z(g24595) ) ;
AND2    gate20551  (.A(g771), .B(g23887), .Z(g24596) ) ;
AND2    gate20552  (.A(g23518), .B(g23505), .Z(g24603) ) ;
AND2    gate20553  (.A(g1457), .B(g23908), .Z(g24604) ) ;
AND2    gate20554  (.A(g23533), .B(g23521), .Z(g24610) ) ;
AND2    gate20555  (.A(g2151), .B(g23940), .Z(g24611) ) ;
AND2    gate20556  (.A(g17203), .B(g24115), .Z(g24644) ) ;
AND2    gate20557  (.A(g17208), .B(g24134), .Z(g24664) ) ;
AND2    gate20558  (.A(g17214), .B(g24153), .Z(g24683) ) ;
AND2    gate20559  (.A(g17217), .B(g24168), .Z(g24700) ) ;
NAND3   gate20560  (.A(g9232), .B(g9150), .C(g12780), .Z(g15454) ) ;
AND2    gate20561  (.A(g15454), .B(g24096), .Z(g24745) ) ;
AND2    gate20562  (.A(g15454), .B(g24098), .Z(g24746) ) ;
AND2    gate20563  (.A(g9427), .B(g24099), .Z(g24747) ) ;
AND2    gate20564  (.A(g672), .B(g24101), .Z(g24748) ) ;
NAND3   gate20565  (.A(g9310), .B(g9174), .C(g12819), .Z(g15540) ) ;
AND2    gate20566  (.A(g15540), .B(g24102), .Z(g24749) ) ;
AND2    gate20567  (.A(g15454), .B(g24104), .Z(g24750) ) ;
AND2    gate20568  (.A(g9427), .B(g24105), .Z(g24751) ) ;
AND2    gate20569  (.A(g9507), .B(g24106), .Z(g24752) ) ;
AND2    gate20570  (.A(g15540), .B(g24107), .Z(g24754) ) ;
AND2    gate20571  (.A(g9569), .B(g24108), .Z(g24755) ) ;
AND2    gate20572  (.A(g1358), .B(g24110), .Z(g24757) ) ;
NAND3   gate20573  (.A(g9391), .B(g9216), .C(g12857), .Z(g15618) ) ;
AND2    gate20574  (.A(g15618), .B(g24111), .Z(g24758) ) ;
AND2    gate20575  (.A(g21825), .B(g23885), .Z(g24759) ) ;
AND2    gate20576  (.A(g9427), .B(g24112), .Z(g24760) ) ;
AND2    gate20577  (.A(g9507), .B(g24113), .Z(g24761) ) ;
AND2    gate20578  (.A(g12876), .B(g24114), .Z(g24762) ) ;
AND2    gate20579  (.A(g15540), .B(g24121), .Z(g24767) ) ;
AND2    gate20580  (.A(g9569), .B(g24122), .Z(g24768) ) ;
AND2    gate20581  (.A(g9649), .B(g24123), .Z(g24769) ) ;
AND2    gate20582  (.A(g15618), .B(g24124), .Z(g24772) ) ;
AND2    gate20583  (.A(g9711), .B(g24125), .Z(g24773) ) ;
AND2    gate20584  (.A(g2052), .B(g24127), .Z(g24774) ) ;
NAND3   gate20585  (.A(g9488), .B(g9277), .C(g12898), .Z(g15694) ) ;
AND2    gate20586  (.A(g15694), .B(g24128), .Z(g24775) ) ;
AND2    gate20587  (.A(g9507), .B(g24129), .Z(g24776) ) ;
AND2    gate20588  (.A(g12876), .B(g24130), .Z(g24777) ) ;
AND2    gate20589  (.A(g9569), .B(g24131), .Z(g24779) ) ;
AND2    gate20590  (.A(g9649), .B(g24132), .Z(g24780) ) ;
AND2    gate20591  (.A(g12916), .B(g24133), .Z(g24781) ) ;
AND2    gate20592  (.A(g15618), .B(g24140), .Z(g24788) ) ;
AND2    gate20593  (.A(g9711), .B(g24141), .Z(g24789) ) ;
AND2    gate20594  (.A(g9795), .B(g24142), .Z(g24790) ) ;
AND2    gate20595  (.A(g15694), .B(g24143), .Z(g24792) ) ;
AND2    gate20596  (.A(g9857), .B(g24144), .Z(g24793) ) ;
AND2    gate20597  (.A(g2746), .B(g24146), .Z(g24794) ) ;
NOR2    gate20598  (.A(g22637), .B(g22665), .Z(g24232) ) ;
AND2    gate20599  (.A(g12017), .B(g24232), .Z(g24795) ) ;
AND2    gate20600  (.A(g12876), .B(g24147), .Z(g24796) ) ;
AND2    gate20601  (.A(g9649), .B(g24148), .Z(g24798) ) ;
AND2    gate20602  (.A(g12916), .B(g24149), .Z(g24799) ) ;
AND2    gate20603  (.A(g9711), .B(g24150), .Z(g24802) ) ;
AND2    gate20604  (.A(g9795), .B(g24151), .Z(g24803) ) ;
AND2    gate20605  (.A(g12945), .B(g24152), .Z(g24804) ) ;
AND2    gate20606  (.A(g15694), .B(g24159), .Z(g24809) ) ;
AND2    gate20607  (.A(g9857), .B(g24160), .Z(g24810) ) ;
AND2    gate20608  (.A(g9941), .B(g24161), .Z(g24811) ) ;
AND2    gate20609  (.A(g21825), .B(g23905), .Z(g24813) ) ;
AND2    gate20610  (.A(g12916), .B(g24162), .Z(g24818) ) ;
AND2    gate20611  (.A(g9795), .B(g24163), .Z(g24821) ) ;
AND2    gate20612  (.A(g12945), .B(g24164), .Z(g24822) ) ;
AND2    gate20613  (.A(g9857), .B(g24165), .Z(g24824) ) ;
AND2    gate20614  (.A(g9941), .B(g24166), .Z(g24825) ) ;
AND2    gate20615  (.A(g12974), .B(g24167), .Z(g24826) ) ;
NAND2   gate20616  (.A(g20885), .B(g22175), .Z(g24100) ) ;
AND2    gate20617  (.A(g24100), .B(g20401), .Z(g24831) ) ;
AND2    gate20618  (.A(g12945), .B(g24175), .Z(g24838) ) ;
AND2    gate20619  (.A(g9941), .B(g24176), .Z(g24840) ) ;
AND2    gate20620  (.A(g12974), .B(g24177), .Z(g24841) ) ;
AND2    gate20621  (.A(g21825), .B(g23918), .Z(g24843) ) ;
NAND2   gate20622  (.A(g20904), .B(g22190), .Z(g24109) ) ;
AND2    gate20623  (.A(g24109), .B(g20426), .Z(g24846) ) ;
AND2    gate20624  (.A(g12974), .B(g24180), .Z(g24853) ) ;
AND2    gate20625  (.A(g18174), .B(g23731), .Z(g24855) ) ;
AND2    gate20626  (.A(g24047), .B(g18873), .Z(g24858) ) ;
NAND2   gate20627  (.A(g20928), .B(g22199), .Z(g24126) ) ;
AND2    gate20628  (.A(g24126), .B(g20448), .Z(g24861) ) ;
AND2    gate20629  (.A(g666), .B(g23779), .Z(g24867) ) ;
AND2    gate20630  (.A(g24047), .B(g18894), .Z(g24869) ) ;
AND2    gate20631  (.A(g18281), .B(g23786), .Z(g24870) ) ;
AND2    gate20632  (.A(g24060), .B(g18899), .Z(g24874) ) ;
NAND2   gate20633  (.A(g20956), .B(g22205), .Z(g24145) ) ;
AND2    gate20634  (.A(g24145), .B(g20467), .Z(g24876) ) ;
AND2    gate20635  (.A(g19830), .B(g24210), .Z(g24878) ) ;
AND2    gate20636  (.A(g24047), .B(g18912), .Z(g24881) ) ;
AND2    gate20637  (.A(g1352), .B(g23832), .Z(g24882) ) ;
AND2    gate20638  (.A(g24060), .B(g18917), .Z(g24884) ) ;
AND2    gate20639  (.A(g18374), .B(g23839), .Z(g24885) ) ;
AND2    gate20640  (.A(g24073), .B(g18922), .Z(g24888) ) ;
AND2    gate20641  (.A(g24060), .B(g18931), .Z(g24898) ) ;
AND2    gate20642  (.A(g2046), .B(g23867), .Z(g24899) ) ;
AND2    gate20643  (.A(g24073), .B(g18936), .Z(g24901) ) ;
AND2    gate20644  (.A(g18469), .B(g23874), .Z(g24902) ) ;
AND2    gate20645  (.A(g24084), .B(g18941), .Z(g24905) ) ;
AND2    gate20646  (.A(g18886), .B(g23879), .Z(g24906) ) ;
AND2    gate20647  (.A(g7466), .B(g24220), .Z(g24907) ) ;
AND2    gate20648  (.A(g7342), .B(g23882), .Z(g24908) ) ;
AND2    gate20649  (.A(g24073), .B(g18951), .Z(g24921) ) ;
AND2    gate20650  (.A(g2740), .B(g23901), .Z(g24922) ) ;
AND2    gate20651  (.A(g24084), .B(g18956), .Z(g24924) ) ;
AND2    gate20652  (.A(g24084), .B(g18967), .Z(g24938) ) ;
AND2    gate20653  (.A(g7595), .B(g24251), .Z(g24964) ) ;
AND2    gate20654  (.A(g7600), .B(g24030), .Z(g24974) ) ;
AND2    gate20655  (.A(g23444), .B(g10880), .Z(g25086) ) ;
AND2    gate20656  (.A(g23444), .B(g10915), .Z(g25102) ) ;
AND2    gate20657  (.A(g23444), .B(g10974), .Z(g25117) ) ;
AND3    gate20658  (.A(g17051), .B(g24115), .C(g13614), .Z(g25128) ) ;
NOR2    gate20659  (.A(g24183), .B(g529), .Z(g24623) ) ;
AND2    gate20660  (.A(g24623), .B(g20634), .Z(g25178) ) ;
NOR2    gate20661  (.A(g24183), .B(g530), .Z(g24636) ) ;
AND2    gate20662  (.A(g24636), .B(g20673), .Z(g25181) ) ;
NOR2    gate20663  (.A(g24183), .B(g533), .Z(g24681) ) ;
AND2    gate20664  (.A(g24681), .B(g20676), .Z(g25182) ) ;
NOR2    gate20665  (.A(g24183), .B(g534), .Z(g24694) ) ;
AND2    gate20666  (.A(g24694), .B(g20735), .Z(g25184) ) ;
OR2     gate20667  (.A(g24094), .B(g20842), .Z(g24633) ) ;
AND2    gate20668  (.A(g24633), .B(g16608), .Z(g25187) ) ;
NOR2    gate20669  (.A(g24183), .B(g531), .Z(g24652) ) ;
AND2    gate20670  (.A(g24652), .B(g20763), .Z(g25188) ) ;
NOR2    gate20671  (.A(g24183), .B(g536), .Z(g24711) ) ;
AND2    gate20672  (.A(g24711), .B(g20790), .Z(g25192) ) ;
OR2     gate20673  (.A(g24095), .B(g20850), .Z(g24653) ) ;
AND2    gate20674  (.A(g24653), .B(g16626), .Z(g25193) ) ;
OR2     gate20675  (.A(g24097), .B(g20858), .Z(g24672) ) ;
AND2    gate20676  (.A(g24672), .B(g16640), .Z(g25196) ) ;
OR2     gate20677  (.A(g24103), .B(g20866), .Z(g24691) ) ;
AND2    gate20678  (.A(g24691), .B(g16651), .Z(g25198) ) ;
AND2    gate20679  (.A(g24648), .B(g8700), .Z(g25269) ) ;
AND2    gate20680  (.A(g24648), .B(g8714), .Z(g25277) ) ;
AND2    gate20681  (.A(g24668), .B(g8719), .Z(g25278) ) ;
AND2    gate20682  (.A(g5606), .B(g24815), .Z(g25281) ) ;
AND2    gate20683  (.A(g24648), .B(g8748), .Z(g25282) ) ;
AND2    gate20684  (.A(g24668), .B(g8752), .Z(g25286) ) ;
AND2    gate20685  (.A(g24687), .B(g8757), .Z(g25287) ) ;
AND2    gate20686  (.A(g5631), .B(g24834), .Z(g25289) ) ;
AND2    gate20687  (.A(g24668), .B(g8771), .Z(g25290) ) ;
AND2    gate20688  (.A(g24687), .B(g8775), .Z(g25294) ) ;
AND2    gate20689  (.A(g24704), .B(g8780), .Z(g25295) ) ;
AND2    gate20690  (.A(g5659), .B(g24850), .Z(g25299) ) ;
AND2    gate20691  (.A(g24687), .B(g8794), .Z(g25300) ) ;
AND2    gate20692  (.A(g24704), .B(g8798), .Z(g25304) ) ;
AND2    gate20693  (.A(g5697), .B(g24864), .Z(g25309) ) ;
AND2    gate20694  (.A(g24704), .B(g8813), .Z(g25310) ) ;
NOR2    gate20695  (.A(g23688), .B(g24183), .Z(g24682) ) ;
AND3    gate20696  (.A(g24682), .B(g19358), .C(g19335), .Z(g25318) ) ;
NOR2    gate20697  (.A(g13880), .B(g23483), .Z(g25075) ) ;
AND2    gate20698  (.A(g25075), .B(g9669), .Z(g25321) ) ;
AND2    gate20699  (.A(g24644), .B(g17892), .Z(g25328) ) ;
AND2    gate20700  (.A(g24644), .B(g17984), .Z(g25334) ) ;
AND2    gate20701  (.A(g24664), .B(g18003), .Z(g25337) ) ;
AND2    gate20702  (.A(g5851), .B(g24600), .Z(g25342) ) ;
AND2    gate20703  (.A(g24644), .B(g18084), .Z(g25346) ) ;
AND2    gate20704  (.A(g24664), .B(g18101), .Z(g25348) ) ;
AND2    gate20705  (.A(g24683), .B(g18120), .Z(g25351) ) ;
AND2    gate20706  (.A(g5898), .B(g24607), .Z(g25356) ) ;
AND2    gate20707  (.A(g24664), .B(g18200), .Z(g25360) ) ;
AND2    gate20708  (.A(g24683), .B(g18217), .Z(g25362) ) ;
AND2    gate20709  (.A(g24700), .B(g18236), .Z(g25365) ) ;
AND2    gate20710  (.A(g5937), .B(g24619), .Z(g25371) ) ;
AND2    gate20711  (.A(g24683), .B(g18307), .Z(g25375) ) ;
AND2    gate20712  (.A(g24700), .B(g18324), .Z(g25377) ) ;
AND2    gate20713  (.A(g5971), .B(g24630), .Z(g25388) ) ;
AND2    gate20714  (.A(g24700), .B(g18400), .Z(g25392) ) ;
AND2    gate20715  (.A(g6142), .B(g24763), .Z(g25453) ) ;
AND2    gate20716  (.A(g6163), .B(g24784), .Z(g25457) ) ;
AND2    gate20717  (.A(g6190), .B(g24805), .Z(g25461) ) ;
AND2    gate20718  (.A(g6222), .B(g24827), .Z(g25466) ) ;
NOR2    gate20719  (.A(g23593), .B(g22516), .Z(g24479) ) ;
AND2    gate20720  (.A(g24479), .B(g20400), .Z(g25470) ) ;
AND2    gate20721  (.A(g14148), .B(g25087), .Z(g25475) ) ;
NOR2    gate20722  (.A(g23617), .B(g23659), .Z(g24480) ) ;
AND2    gate20723  (.A(g24480), .B(g17567), .Z(g25482) ) ;
NOR2    gate20724  (.A(g23618), .B(g19696), .Z(g24481) ) ;
AND2    gate20725  (.A(g24481), .B(g20421), .Z(g25483) ) ;
NOR2    gate20726  (.A(g23625), .B(g22556), .Z(g24485) ) ;
AND2    gate20727  (.A(g24485), .B(g20425), .Z(g25487) ) ;
AND2    gate20728  (.A(g6707), .B(g25094), .Z(g25505) ) ;
AND2    gate20729  (.A(g14263), .B(g25095), .Z(g25506) ) ;
NOR2    gate20730  (.A(g23666), .B(g23709), .Z(g24487) ) ;
AND2    gate20731  (.A(g24487), .B(g17664), .Z(g25513) ) ;
NOR2    gate20732  (.A(g23667), .B(g19740), .Z(g24488) ) ;
AND2    gate20733  (.A(g24488), .B(g20443), .Z(g25514) ) ;
NOR2    gate20734  (.A(g23674), .B(g22596), .Z(g24489) ) ;
AND2    gate20735  (.A(g24489), .B(g20447), .Z(g25518) ) ;
AND2    gate20736  (.A(g7009), .B(g25104), .Z(g25552) ) ;
AND2    gate20737  (.A(g14385), .B(g25105), .Z(g25553) ) ;
NOR2    gate20738  (.A(g23716), .B(g23763), .Z(g24494) ) ;
AND2    gate20739  (.A(g24494), .B(g17764), .Z(g25560) ) ;
NOR2    gate20740  (.A(g23717), .B(g19783), .Z(g24495) ) ;
AND2    gate20741  (.A(g24495), .B(g20462), .Z(g25561) ) ;
NOR2    gate20742  (.A(g23724), .B(g22633), .Z(g24496) ) ;
AND2    gate20743  (.A(g24496), .B(g20466), .Z(g25565) ) ;
AND2    gate20744  (.A(g7259), .B(g25110), .Z(g25618) ) ;
AND2    gate20745  (.A(g14497), .B(g25111), .Z(g25619) ) ;
NOR2    gate20746  (.A(g23770), .B(g23818), .Z(g24504) ) ;
AND2    gate20747  (.A(g24504), .B(g17865), .Z(g25626) ) ;
NOR2    gate20748  (.A(g23771), .B(g19825), .Z(g24505) ) ;
AND2    gate20749  (.A(g24505), .B(g20477), .Z(g25627) ) ;
NOR2    gate20750  (.A(g19836), .B(g17877), .Z(g21008) ) ;
AND2    gate20751  (.A(g21008), .B(g25115), .Z(g25628) ) ;
AND2    gate20752  (.A(g3024), .B(g25116), .Z(g25629) ) ;
AND2    gate20753  (.A(g7455), .B(g25120), .Z(g25697) ) ;
AND2    gate20754  (.A(g2908), .B(g25126), .Z(g25881) ) ;
NOR2    gate20755  (.A(g16211), .B(g24229), .Z(g24800) ) ;
AND2    gate20756  (.A(g24800), .B(g13670), .Z(g25951) ) ;
NOR2    gate20757  (.A(g16161), .B(g24224), .Z(g24783) ) ;
AND2    gate20758  (.A(g24783), .B(g13699), .Z(g25953) ) ;
NOR2    gate20759  (.A(g16160), .B(g24221), .Z(g24782) ) ;
AND2    gate20760  (.A(g24782), .B(g11869), .Z(g25957) ) ;
NOR2    gate20761  (.A(g16119), .B(g24217), .Z(g24770) ) ;
AND2    gate20762  (.A(g24770), .B(g11901), .Z(g25961) ) ;
NOR2    gate20763  (.A(g16089), .B(g24211), .Z(g24756) ) ;
AND2    gate20764  (.A(g24756), .B(g11944), .Z(g25963) ) ;
NOR2    gate20765  (.A(g16422), .B(g24256), .Z(g24871) ) ;
AND2    gate20766  (.A(g24871), .B(g11986), .Z(g25968) ) ;
NOR2    gate20767  (.A(g16390), .B(g24253), .Z(g24859) ) ;
AND2    gate20768  (.A(g24859), .B(g12042), .Z(g25972) ) ;
NOR2    gate20769  (.A(g16356), .B(g24247), .Z(g24847) ) ;
AND2    gate20770  (.A(g24847), .B(g13838), .Z(g25973) ) ;
NOR2    gate20771  (.A(g24183), .B(g537), .Z(g24606) ) ;
AND2    gate20772  (.A(g24606), .B(g21917), .Z(g25975) ) ;
NOR2    gate20773  (.A(g16350), .B(g24246), .Z(g24845) ) ;
AND2    gate20774  (.A(g24845), .B(g12089), .Z(g25977) ) ;
NOR2    gate20775  (.A(g16309), .B(g24241), .Z(g24836) ) ;
AND2    gate20776  (.A(g24836), .B(g13850), .Z(g25978) ) ;
NOR2    gate20777  (.A(g24183), .B(g532), .Z(g24663) ) ;
AND2    gate20778  (.A(g24663), .B(g21928), .Z(g25980) ) ;
NOR2    gate20779  (.A(g16262), .B(g24236), .Z(g24819) ) ;
AND2    gate20780  (.A(g24819), .B(g13858), .Z(g25981) ) ;
AND2    gate20781  (.A(g25422), .B(g24912), .Z(g26023) ) ;
AND2    gate20782  (.A(g25301), .B(g21102), .Z(g26024) ) ;
AND2    gate20783  (.A(g25431), .B(g24929), .Z(g26026) ) ;
NOR2    gate20784  (.A(g24482), .B(g22319), .Z(g25418) ) ;
AND2    gate20785  (.A(g25418), .B(g22271), .Z(g26027) ) ;
AND2    gate20786  (.A(g25438), .B(g24941), .Z(g26028) ) ;
AND2    gate20787  (.A(g25445), .B(g24952), .Z(g26029) ) ;
NOR2    gate20788  (.A(g24482), .B(g22319), .Z(g25429) ) ;
AND2    gate20789  (.A(g25429), .B(g22304), .Z(g26030) ) ;
AND2    gate20790  (.A(g25379), .B(g19415), .Z(g26032) ) ;
AND2    gate20791  (.A(g25395), .B(g19452), .Z(g26033) ) ;
AND2    gate20792  (.A(g25405), .B(g19479), .Z(g26034) ) ;
NOR2    gate20793  (.A(g20842), .B(g24429), .Z(g25523) ) ;
AND2    gate20794  (.A(g25523), .B(g19483), .Z(g26035) ) ;
AND2    gate20795  (.A(g25413), .B(g19502), .Z(g26036) ) ;
NOR2    gate20796  (.A(g20850), .B(g24433), .Z(g25589) ) ;
AND2    gate20797  (.A(g25589), .B(g19504), .Z(g26038) ) ;
NOR2    gate20798  (.A(g20858), .B(g24437), .Z(g25668) ) ;
AND2    gate20799  (.A(g25668), .B(g19523), .Z(g26039) ) ;
NOR2    gate20800  (.A(g20866), .B(g24440), .Z(g25745) ) ;
AND2    gate20801  (.A(g25745), .B(g19533), .Z(g26040) ) ;
AND2    gate20802  (.A(g70), .B(g25296), .Z(g26051) ) ;
NOR2    gate20803  (.A(g24529), .B(g24540), .Z(g25941) ) ;
AND2    gate20804  (.A(g25941), .B(g21087), .Z(g26052) ) ;
AND2    gate20805  (.A(g758), .B(g25306), .Z(g26053) ) ;
NOR2    gate20806  (.A(g24542), .B(g24552), .Z(g25944) ) ;
AND2    gate20807  (.A(g25944), .B(g21099), .Z(g26054) ) ;
NOR2    gate20808  (.A(g24541), .B(g24550), .Z(g25943) ) ;
AND2    gate20809  (.A(g25943), .B(g21108), .Z(g26060) ) ;
AND2    gate20810  (.A(g1444), .B(g25315), .Z(g26061) ) ;
NOR2    gate20811  (.A(g24554), .B(g24563), .Z(g25947) ) ;
AND2    gate20812  (.A(g25947), .B(g21113), .Z(g26062) ) ;
NOR2    gate20813  (.A(g24553), .B(g24561), .Z(g25946) ) ;
AND2    gate20814  (.A(g25946), .B(g21125), .Z(g26067) ) ;
AND2    gate20815  (.A(g2138), .B(g25324), .Z(g26068) ) ;
NOR2    gate20816  (.A(g24565), .B(g24573), .Z(g25949) ) ;
AND2    gate20817  (.A(g25949), .B(g21130), .Z(g26069) ) ;
NOR2    gate20818  (.A(g24564), .B(g24571), .Z(g25948) ) ;
AND2    gate20819  (.A(g25948), .B(g21144), .Z(g26074) ) ;
AND2    gate20820  (.A(g74), .B(g25698), .Z(g26075) ) ;
NOR2    gate20821  (.A(g24574), .B(g24580), .Z(g25950) ) ;
AND2    gate20822  (.A(g25950), .B(g21164), .Z(g26080) ) ;
AND2    gate20823  (.A(g762), .B(g25771), .Z(g26082) ) ;
AND2    gate20824  (.A(g1448), .B(g25825), .Z(g26085) ) ;
AND2    gate20825  (.A(g2142), .B(g25860), .Z(g26091) ) ;
AND2    gate20826  (.A(g21825), .B(g25630), .Z(g26157) ) ;
AND2    gate20827  (.A(g679), .B(g25937), .Z(g26158) ) ;
AND2    gate20828  (.A(g1365), .B(g25939), .Z(g26163) ) ;
AND2    gate20829  (.A(g686), .B(g25454), .Z(g26166) ) ;
AND2    gate20830  (.A(g2059), .B(g25942), .Z(g26171) ) ;
AND2    gate20831  (.A(g1372), .B(g25458), .Z(g26186) ) ;
AND2    gate20832  (.A(g2753), .B(g25945), .Z(g26188) ) ;
AND2    gate20833  (.A(g2066), .B(g25463), .Z(g26207) ) ;
AND2    gate20834  (.A(g4217), .B(g25467), .Z(g26212) ) ;
AND2    gate20835  (.A(g25895), .B(g9306), .Z(g26213) ) ;
AND2    gate20836  (.A(g2760), .B(g25472), .Z(g26231) ) ;
AND2    gate20837  (.A(g4340), .B(g25476), .Z(g26233) ) ;
AND2    gate20838  (.A(g4343), .B(g25479), .Z(g26234) ) ;
AND2    gate20839  (.A(g25895), .B(g9368), .Z(g26235) ) ;
AND2    gate20840  (.A(g25899), .B(g9371), .Z(g26236) ) ;
AND2    gate20841  (.A(g4372), .B(g25484), .Z(g26243) ) ;
AND2    gate20842  (.A(g25903), .B(g9387), .Z(g26244) ) ;
AND2    gate20843  (.A(g4465), .B(g25493), .Z(g26257) ) ;
AND2    gate20844  (.A(g4468), .B(g25496), .Z(g26258) ) ;
AND2    gate20845  (.A(g4471), .B(g25499), .Z(g26259) ) ;
NOR2    gate20846  (.A(g24831), .B(g23687), .Z(g25254) ) ;
AND2    gate20847  (.A(g25254), .B(g17649), .Z(g26260) ) ;
AND2    gate20848  (.A(g25895), .B(g9443), .Z(g26261) ) ;
AND2    gate20849  (.A(g25899), .B(g9446), .Z(g26262) ) ;
AND2    gate20850  (.A(g4476), .B(g25502), .Z(g26263) ) ;
AND2    gate20851  (.A(g4509), .B(g25507), .Z(g26268) ) ;
AND2    gate20852  (.A(g4512), .B(g25510), .Z(g26269) ) ;
AND2    gate20853  (.A(g25903), .B(g9465), .Z(g26270) ) ;
AND2    gate20854  (.A(g25907), .B(g9468), .Z(g26271) ) ;
AND2    gate20855  (.A(g4541), .B(g25515), .Z(g26278) ) ;
AND2    gate20856  (.A(g25911), .B(g9484), .Z(g26279) ) ;
AND2    gate20857  (.A(g4592), .B(g25524), .Z(g26288) ) ;
AND2    gate20858  (.A(g4595), .B(g25527), .Z(g26289) ) ;
AND2    gate20859  (.A(g4598), .B(g25530), .Z(g26290) ) ;
AND2    gate20860  (.A(g25899), .B(g9524), .Z(g26291) ) ;
AND2    gate20861  (.A(g4603), .B(g25533), .Z(g26292) ) ;
AND2    gate20862  (.A(g4606), .B(g25536), .Z(g26293) ) ;
AND2    gate20863  (.A(g4641), .B(g25540), .Z(g26298) ) ;
AND2    gate20864  (.A(g4644), .B(g25543), .Z(g26299) ) ;
AND2    gate20865  (.A(g4647), .B(g25546), .Z(g26300) ) ;
NOR2    gate20866  (.A(g24846), .B(g23741), .Z(g25258) ) ;
AND2    gate20867  (.A(g25258), .B(g17749), .Z(g26301) ) ;
AND2    gate20868  (.A(g25903), .B(g9585), .Z(g26302) ) ;
AND2    gate20869  (.A(g25907), .B(g9588), .Z(g26303) ) ;
AND2    gate20870  (.A(g4652), .B(g25549), .Z(g26307) ) ;
AND2    gate20871  (.A(g4685), .B(g25554), .Z(g26309) ) ;
AND2    gate20872  (.A(g4688), .B(g25557), .Z(g26310) ) ;
AND2    gate20873  (.A(g25911), .B(g9607), .Z(g26311) ) ;
AND2    gate20874  (.A(g25915), .B(g9610), .Z(g26312) ) ;
AND2    gate20875  (.A(g4717), .B(g25562), .Z(g26316) ) ;
AND2    gate20876  (.A(g25919), .B(g9626), .Z(g26317) ) ;
AND2    gate20877  (.A(g4737), .B(g25573), .Z(g26318) ) ;
AND2    gate20878  (.A(g4740), .B(g25576), .Z(g26319) ) ;
AND2    gate20879  (.A(g4743), .B(g25579), .Z(g26324) ) ;
AND2    gate20880  (.A(g4746), .B(g25582), .Z(g26325) ) ;
AND2    gate20881  (.A(g4749), .B(g25585), .Z(g26326) ) ;
AND2    gate20882  (.A(g4769), .B(g25590), .Z(g26332) ) ;
AND2    gate20883  (.A(g4772), .B(g25593), .Z(g26333) ) ;
AND2    gate20884  (.A(g4775), .B(g25596), .Z(g26334) ) ;
AND2    gate20885  (.A(g25907), .B(g9666), .Z(g26335) ) ;
AND2    gate20886  (.A(g4780), .B(g25599), .Z(g26339) ) ;
AND2    gate20887  (.A(g4783), .B(g25602), .Z(g26340) ) ;
AND2    gate20888  (.A(g4818), .B(g25606), .Z(g26342) ) ;
AND2    gate20889  (.A(g4821), .B(g25609), .Z(g26343) ) ;
AND2    gate20890  (.A(g4824), .B(g25612), .Z(g26344) ) ;
NOR2    gate20891  (.A(g24861), .B(g23796), .Z(g25261) ) ;
AND2    gate20892  (.A(g25261), .B(g17850), .Z(g26345) ) ;
AND2    gate20893  (.A(g25911), .B(g9727), .Z(g26346) ) ;
AND2    gate20894  (.A(g25915), .B(g9730), .Z(g26347) ) ;
AND2    gate20895  (.A(g4829), .B(g25615), .Z(g26348) ) ;
AND2    gate20896  (.A(g4862), .B(g25620), .Z(g26350) ) ;
AND2    gate20897  (.A(g4865), .B(g25623), .Z(g26351) ) ;
AND2    gate20898  (.A(g25919), .B(g9749), .Z(g26352) ) ;
AND2    gate20899  (.A(g25923), .B(g9752), .Z(g26353) ) ;
AND2    gate20900  (.A(g4882), .B(g25634), .Z(g26357) ) ;
AND2    gate20901  (.A(g4888), .B(g25637), .Z(g26361) ) ;
AND2    gate20902  (.A(g4891), .B(g25640), .Z(g26362) ) ;
AND2    gate20903  (.A(g4894), .B(g25643), .Z(g26363) ) ;
AND2    gate20904  (.A(g4913), .B(g25652), .Z(g26365) ) ;
AND2    gate20905  (.A(g4916), .B(g25655), .Z(g26366) ) ;
AND2    gate20906  (.A(g4919), .B(g25658), .Z(g26371) ) ;
AND2    gate20907  (.A(g4922), .B(g25661), .Z(g26372) ) ;
AND2    gate20908  (.A(g4925), .B(g25664), .Z(g26373) ) ;
AND2    gate20909  (.A(g4945), .B(g25669), .Z(g26379) ) ;
AND2    gate20910  (.A(g4948), .B(g25672), .Z(g26380) ) ;
AND2    gate20911  (.A(g4951), .B(g25675), .Z(g26381) ) ;
AND2    gate20912  (.A(g25915), .B(g9812), .Z(g26382) ) ;
AND2    gate20913  (.A(g4956), .B(g25678), .Z(g26383) ) ;
AND2    gate20914  (.A(g4959), .B(g25681), .Z(g26384) ) ;
AND2    gate20915  (.A(g4994), .B(g25685), .Z(g26386) ) ;
AND2    gate20916  (.A(g4997), .B(g25688), .Z(g26387) ) ;
AND2    gate20917  (.A(g5000), .B(g25691), .Z(g26388) ) ;
NOR2    gate20918  (.A(g24876), .B(g23849), .Z(g25264) ) ;
AND2    gate20919  (.A(g25264), .B(g17962), .Z(g26389) ) ;
AND2    gate20920  (.A(g25919), .B(g9873), .Z(g26390) ) ;
AND2    gate20921  (.A(g25923), .B(g9876), .Z(g26391) ) ;
AND2    gate20922  (.A(g5005), .B(g25694), .Z(g26392) ) ;
AND2    gate20923  (.A(g5027), .B(g25700), .Z(g26396) ) ;
AND2    gate20924  (.A(g5030), .B(g25703), .Z(g26397) ) ;
AND2    gate20925  (.A(g5041), .B(g25711), .Z(g26400) ) ;
AND2    gate20926  (.A(g5047), .B(g25714), .Z(g26404) ) ;
AND2    gate20927  (.A(g5050), .B(g25717), .Z(g26405) ) ;
AND2    gate20928  (.A(g5053), .B(g25720), .Z(g26406) ) ;
AND2    gate20929  (.A(g5072), .B(g25729), .Z(g26408) ) ;
AND2    gate20930  (.A(g5075), .B(g25732), .Z(g26409) ) ;
AND2    gate20931  (.A(g5078), .B(g25735), .Z(g26414) ) ;
AND2    gate20932  (.A(g5081), .B(g25738), .Z(g26415) ) ;
AND2    gate20933  (.A(g5084), .B(g25741), .Z(g26416) ) ;
AND2    gate20934  (.A(g5104), .B(g25746), .Z(g26422) ) ;
AND2    gate20935  (.A(g5107), .B(g25749), .Z(g26423) ) ;
AND2    gate20936  (.A(g5110), .B(g25752), .Z(g26424) ) ;
AND2    gate20937  (.A(g25923), .B(g9958), .Z(g26425) ) ;
AND2    gate20938  (.A(g5115), .B(g25755), .Z(g26426) ) ;
AND2    gate20939  (.A(g5118), .B(g25758), .Z(g26427) ) ;
AND2    gate20940  (.A(g5145), .B(g25767), .Z(g26432) ) ;
AND2    gate20941  (.A(g5156), .B(g25773), .Z(g26437) ) ;
AND2    gate20942  (.A(g5159), .B(g25776), .Z(g26438) ) ;
AND2    gate20943  (.A(g5170), .B(g25784), .Z(g26441) ) ;
AND2    gate20944  (.A(g5176), .B(g25787), .Z(g26445) ) ;
AND2    gate20945  (.A(g5179), .B(g25790), .Z(g26446) ) ;
AND2    gate20946  (.A(g5182), .B(g25793), .Z(g26447) ) ;
AND2    gate20947  (.A(g5201), .B(g25802), .Z(g26449) ) ;
AND2    gate20948  (.A(g5204), .B(g25805), .Z(g26450) ) ;
AND2    gate20949  (.A(g5207), .B(g25808), .Z(g26455) ) ;
AND2    gate20950  (.A(g5210), .B(g25811), .Z(g26456) ) ;
AND2    gate20951  (.A(g5213), .B(g25814), .Z(g26457) ) ;
AND2    gate20952  (.A(g5238), .B(g25821), .Z(g26464) ) ;
AND2    gate20953  (.A(g5249), .B(g25827), .Z(g26469) ) ;
AND2    gate20954  (.A(g5252), .B(g25830), .Z(g26470) ) ;
AND2    gate20955  (.A(g5263), .B(g25838), .Z(g26473) ) ;
AND2    gate20956  (.A(g5269), .B(g25841), .Z(g26477) ) ;
AND2    gate20957  (.A(g5272), .B(g25844), .Z(g26478) ) ;
AND2    gate20958  (.A(g5275), .B(g25847), .Z(g26479) ) ;
AND2    gate20959  (.A(g5301), .B(g25856), .Z(g26488) ) ;
AND2    gate20960  (.A(g5312), .B(g25862), .Z(g26493) ) ;
AND2    gate20961  (.A(g5315), .B(g25865), .Z(g26494) ) ;
AND2    gate20962  (.A(g5338), .B(g25877), .Z(g26504) ) ;
AND2    gate20963  (.A(g25274), .B(g21066), .Z(g26663) ) ;
AND2    gate20964  (.A(g25283), .B(g21076), .Z(g26668) ) ;
NOR2    gate20965  (.A(g8580), .B(g10730), .Z(g12431) ) ;
AND2    gate20966  (.A(g12431), .B(g25318), .Z(g26673) ) ;
AND2    gate20967  (.A(g25291), .B(g21090), .Z(g26674) ) ;
AND2    gate20968  (.A(g14657), .B(g26508), .Z(g26754) ) ;
NOR2    gate20969  (.A(g25426), .B(g22319), .Z(g26083) ) ;
AND2    gate20970  (.A(g26083), .B(g22239), .Z(g26755) ) ;
NOR2    gate20971  (.A(g25426), .B(g22319), .Z(g26113) ) ;
AND2    gate20972  (.A(g26113), .B(g22240), .Z(g26756) ) ;
NOR3    gate20973  (.A(g15962), .B(g15942), .C(g14677), .Z(g16614) ) ;
AND3    gate20974  (.A(g16614), .B(g26521), .C(g13637), .Z(g26758) ) ;
NAND2   gate20975  (.A(g16539), .B(g25183), .Z(g26356) ) ;
AND2    gate20976  (.A(g26356), .B(g19251), .Z(g26759) ) ;
NOR3    gate20977  (.A(g6068), .B(g24183), .C(g25355), .Z(g26137) ) ;
AND2    gate20978  (.A(g26137), .B(g22256), .Z(g26760) ) ;
NOR3    gate20979  (.A(g6068), .B(g24183), .C(g25329), .Z(g26154) ) ;
AND2    gate20980  (.A(g26154), .B(g22257), .Z(g26761) ) ;
AND2    gate20981  (.A(g14691), .B(g26516), .Z(g26763) ) ;
NOR3    gate20982  (.A(g15981), .B(g15971), .C(g14711), .Z(g16632) ) ;
AND3    gate20983  (.A(g16632), .B(g26525), .C(g13649), .Z(g26764) ) ;
NAND2   gate20984  (.A(g16571), .B(g25186), .Z(g26399) ) ;
AND2    gate20985  (.A(g26399), .B(g19265), .Z(g26765) ) ;
AND2    gate20986  (.A(g14725), .B(g26521), .Z(g26766) ) ;
NOR3    gate20987  (.A(g6068), .B(g24183), .C(g25319), .Z(g26087) ) ;
AND2    gate20988  (.A(g26087), .B(g22287), .Z(g26767) ) ;
NAND2   gate20989  (.A(g16595), .B(g25190), .Z(g26440) ) ;
AND2    gate20990  (.A(g26440), .B(g19280), .Z(g26768) ) ;
AND2    gate20991  (.A(g14753), .B(g26525), .Z(g26769) ) ;
NAND3   gate20992  (.A(g25422), .B(g25379), .C(g25274), .Z(g26059) ) ;
AND2    gate20993  (.A(g26059), .B(g19287), .Z(g26770) ) ;
AND3    gate20994  (.A(g24912), .B(g26508), .C(g13614), .Z(g26771) ) ;
NOR3    gate20995  (.A(g6068), .B(g24183), .C(g25347), .Z(g26145) ) ;
AND2    gate20996  (.A(g26145), .B(g22303), .Z(g26773) ) ;
NAND2   gate20997  (.A(g16615), .B(g25195), .Z(g26472) ) ;
AND2    gate20998  (.A(g26472), .B(g19299), .Z(g26774) ) ;
NOR3    gate20999  (.A(g6068), .B(g24183), .C(g25313), .Z(g26099) ) ;
AND2    gate21000  (.A(g26099), .B(g22318), .Z(g26775) ) ;
NAND3   gate21001  (.A(g25431), .B(g25395), .C(g25283), .Z(g26066) ) ;
AND2    gate21002  (.A(g26066), .B(g19305), .Z(g26777) ) ;
AND3    gate21003  (.A(g24929), .B(g26516), .C(g13626), .Z(g26778) ) ;
NAND4   gate21004  (.A(g8278), .B(g14657), .C(g25422), .D(g25379), .Z(g26119) ) ;
AND2    gate21005  (.A(g26119), .B(g16622), .Z(g26780) ) ;
NAND3   gate21006  (.A(g25438), .B(g25405), .C(g25291), .Z(g26073) ) ;
AND2    gate21007  (.A(g26073), .B(g19326), .Z(g26783) ) ;
AND3    gate21008  (.A(g24941), .B(g26521), .C(g13637), .Z(g26784) ) ;
NAND4   gate21009  (.A(g8287), .B(g14691), .C(g25431), .D(g25395), .Z(g26129) ) ;
AND2    gate21010  (.A(g26129), .B(g16636), .Z(g26787) ) ;
NAND3   gate21011  (.A(g25445), .B(g25413), .C(g25301), .Z(g26079) ) ;
AND2    gate21012  (.A(g26079), .B(g19353), .Z(g26790) ) ;
AND3    gate21013  (.A(g24952), .B(g26525), .C(g13649), .Z(g26791) ) ;
NAND4   gate21014  (.A(g8296), .B(g14725), .C(g25438), .D(g25405), .Z(g26143) ) ;
AND2    gate21015  (.A(g26143), .B(g16647), .Z(g26794) ) ;
NAND4   gate21016  (.A(g8305), .B(g14753), .C(g25445), .D(g25413), .Z(g26148) ) ;
AND2    gate21017  (.A(g26148), .B(g16659), .Z(g26797) ) ;
AND2    gate21018  (.A(g5623), .B(g26209), .Z(g26829) ) ;
AND2    gate21019  (.A(g5651), .B(g26237), .Z(g26833) ) ;
AND2    gate21020  (.A(g5689), .B(g26275), .Z(g26842) ) ;
AND2    gate21021  (.A(g5664), .B(g26056), .Z(g26845) ) ;
AND2    gate21022  (.A(g5741), .B(g26313), .Z(g26851) ) ;
AND2    gate21023  (.A(g5716), .B(g26063), .Z(g26853) ) ;
AND2    gate21024  (.A(g5774), .B(g26070), .Z(g26860) ) ;
AND2    gate21025  (.A(g5833), .B(g26076), .Z(g26866) ) ;
AND2    gate21026  (.A(g6157), .B(g26533), .Z(g26955) ) ;
AND2    gate21027  (.A(g6184), .B(g26538), .Z(g26958) ) ;
AND2    gate21028  (.A(g13907), .B(g26175), .Z(g26961) ) ;
AND2    gate21029  (.A(g6180), .B(g26178), .Z(g26962) ) ;
AND2    gate21030  (.A(g6216), .B(g26539), .Z(g26963) ) ;
NAND2   gate21031  (.A(g23066), .B(g23051), .Z(g23320) ) ;
AND2    gate21032  (.A(g23320), .B(g26540), .Z(g26965) ) ;
AND2    gate21033  (.A(g13963), .B(g26196), .Z(g26966) ) ;
AND2    gate21034  (.A(g6212), .B(g26202), .Z(g26967) ) ;
AND2    gate21035  (.A(g6305), .B(g26542), .Z(g26968) ) ;
AND2    gate21036  (.A(g23320), .B(g26543), .Z(g26969) ) ;
NAND3   gate21037  (.A(g19242), .B(g21120), .C(g19275), .Z(g21976) ) ;
AND2    gate21038  (.A(g21976), .B(g26544), .Z(g26970) ) ;
NAND2   gate21039  (.A(g23080), .B(g23070), .Z(g23325) ) ;
AND2    gate21040  (.A(g23325), .B(g26546), .Z(g26971) ) ;
AND2    gate21041  (.A(g14033), .B(g26223), .Z(g26972) ) ;
AND2    gate21042  (.A(g6301), .B(g26226), .Z(g26973) ) ;
AND2    gate21043  (.A(g23320), .B(g26550), .Z(g26977) ) ;
AND2    gate21044  (.A(g21976), .B(g26551), .Z(g26978) ) ;
NAND2   gate21045  (.A(g22999), .B(g22174), .Z(g23331) ) ;
AND2    gate21046  (.A(g23331), .B(g26552), .Z(g26979) ) ;
NAND2   gate21047  (.A(g21980), .B(g21975), .Z(g23360) ) ;
AND2    gate21048  (.A(g23360), .B(g26554), .Z(g26980) ) ;
AND2    gate21049  (.A(g23325), .B(g26555), .Z(g26981) ) ;
NAND3   gate21050  (.A(g19255), .B(g21139), .C(g19294), .Z(g21983) ) ;
AND2    gate21051  (.A(g21983), .B(g26556), .Z(g26982) ) ;
NAND2   gate21052  (.A(g23096), .B(g23083), .Z(g23335) ) ;
AND2    gate21053  (.A(g23335), .B(g26558), .Z(g26984) ) ;
AND2    gate21054  (.A(g14124), .B(g26251), .Z(g26985) ) ;
AND2    gate21055  (.A(g6438), .B(g26254), .Z(g26986) ) ;
AND2    gate21056  (.A(g21976), .B(g26561), .Z(g26993) ) ;
AND2    gate21057  (.A(g23331), .B(g26562), .Z(g26994) ) ;
NAND2   gate21058  (.A(g21501), .B(g21536), .Z(g21991) ) ;
AND2    gate21059  (.A(g21991), .B(g26563), .Z(g26995) ) ;
AND2    gate21060  (.A(g23360), .B(g26564), .Z(g26996) ) ;
NAND3   gate21061  (.A(g19450), .B(g21244), .C(g19503), .Z(g22050) ) ;
AND2    gate21062  (.A(g22050), .B(g26565), .Z(g26997) ) ;
AND2    gate21063  (.A(g23325), .B(g26566), .Z(g26998) ) ;
AND2    gate21064  (.A(g21983), .B(g26567), .Z(g26999) ) ;
NAND2   gate21065  (.A(g23013), .B(g22189), .Z(g23340) ) ;
AND2    gate21066  (.A(g23340), .B(g26568), .Z(g27000) ) ;
NAND2   gate21067  (.A(g21987), .B(g21981), .Z(g23364) ) ;
AND2    gate21068  (.A(g23364), .B(g26570), .Z(g27001) ) ;
AND2    gate21069  (.A(g23335), .B(g26571), .Z(g27002) ) ;
NAND3   gate21070  (.A(g19268), .B(g21159), .C(g19312), .Z(g21996) ) ;
AND2    gate21071  (.A(g21996), .B(g26572), .Z(g27003) ) ;
NAND2   gate21072  (.A(g23113), .B(g23099), .Z(g23344) ) ;
AND2    gate21073  (.A(g23344), .B(g26574), .Z(g27004) ) ;
AND2    gate21074  (.A(g23331), .B(g26578), .Z(g27005) ) ;
AND2    gate21075  (.A(g21991), .B(g26579), .Z(g27006) ) ;
AND2    gate21076  (.A(g23360), .B(g26580), .Z(g27007) ) ;
AND2    gate21077  (.A(g22050), .B(g26581), .Z(g27008) ) ;
NAND2   gate21078  (.A(g23135), .B(g22288), .Z(g23368) ) ;
AND2    gate21079  (.A(g23368), .B(g26582), .Z(g27009) ) ;
AND2    gate21080  (.A(g21983), .B(g26584), .Z(g27016) ) ;
AND2    gate21081  (.A(g23340), .B(g26585), .Z(g27017) ) ;
NAND2   gate21082  (.A(g21540), .B(g21572), .Z(g22005) ) ;
AND2    gate21083  (.A(g22005), .B(g26586), .Z(g27018) ) ;
AND2    gate21084  (.A(g23364), .B(g26587), .Z(g27019) ) ;
NAND3   gate21085  (.A(g19477), .B(g21253), .C(g19522), .Z(g22069) ) ;
AND2    gate21086  (.A(g22069), .B(g26588), .Z(g27020) ) ;
AND2    gate21087  (.A(g23335), .B(g26589), .Z(g27021) ) ;
AND2    gate21088  (.A(g21996), .B(g26590), .Z(g27022) ) ;
NAND2   gate21089  (.A(g23029), .B(g22198), .Z(g23349) ) ;
AND2    gate21090  (.A(g23349), .B(g26591), .Z(g27023) ) ;
NAND2   gate21091  (.A(g22000), .B(g21988), .Z(g23372) ) ;
AND2    gate21092  (.A(g23372), .B(g26593), .Z(g27024) ) ;
AND2    gate21093  (.A(g23344), .B(g26594), .Z(g27025) ) ;
NAND3   gate21094  (.A(g19283), .B(g21179), .C(g19333), .Z(g22009) ) ;
AND2    gate21095  (.A(g22009), .B(g26595), .Z(g27026) ) ;
AND2    gate21096  (.A(g21991), .B(g26598), .Z(g27027) ) ;
AND2    gate21097  (.A(g22050), .B(g26599), .Z(g27028) ) ;
AND2    gate21098  (.A(g23368), .B(g26600), .Z(g27029) ) ;
NAND2   gate21099  (.A(g21774), .B(g21787), .Z(g22083) ) ;
AND2    gate21100  (.A(g22083), .B(g26601), .Z(g27030) ) ;
AND2    gate21101  (.A(g23340), .B(g26602), .Z(g27031) ) ;
AND2    gate21102  (.A(g22005), .B(g26603), .Z(g27032) ) ;
AND2    gate21103  (.A(g23364), .B(g26604), .Z(g27033) ) ;
AND2    gate21104  (.A(g22069), .B(g26605), .Z(g27034) ) ;
NAND2   gate21105  (.A(g21968), .B(g22308), .Z(g23377) ) ;
AND2    gate21106  (.A(g23377), .B(g26606), .Z(g27035) ) ;
AND2    gate21107  (.A(g21996), .B(g26608), .Z(g27042) ) ;
AND2    gate21108  (.A(g23349), .B(g26609), .Z(g27043) ) ;
NAND2   gate21109  (.A(g21576), .B(g21605), .Z(g22016) ) ;
AND2    gate21110  (.A(g22016), .B(g26610), .Z(g27044) ) ;
AND2    gate21111  (.A(g23372), .B(g26611), .Z(g27045) ) ;
NAND3   gate21112  (.A(g19500), .B(g21261), .C(g19532), .Z(g22093) ) ;
AND2    gate21113  (.A(g22093), .B(g26612), .Z(g27046) ) ;
AND2    gate21114  (.A(g23344), .B(g26613), .Z(g27047) ) ;
AND2    gate21115  (.A(g22009), .B(g26614), .Z(g27048) ) ;
NAND2   gate21116  (.A(g23046), .B(g22204), .Z(g23353) ) ;
AND2    gate21117  (.A(g23353), .B(g26615), .Z(g27049) ) ;
NAND2   gate21118  (.A(g22013), .B(g22001), .Z(g23381) ) ;
AND2    gate21119  (.A(g23381), .B(g26617), .Z(g27050) ) ;
AND2    gate21120  (.A(g4885), .B(g26358), .Z(g27052) ) ;
AND2    gate21121  (.A(g23368), .B(g26619), .Z(g27053) ) ;
AND2    gate21122  (.A(g22083), .B(g26620), .Z(g27054) ) ;
AND2    gate21123  (.A(g22005), .B(g26621), .Z(g27055) ) ;
AND2    gate21124  (.A(g22069), .B(g26622), .Z(g27056) ) ;
AND2    gate21125  (.A(g23377), .B(g26623), .Z(g27057) ) ;
NAND2   gate21126  (.A(g21789), .B(g21801), .Z(g22108) ) ;
AND2    gate21127  (.A(g22108), .B(g26624), .Z(g27058) ) ;
AND2    gate21128  (.A(g23349), .B(g26625), .Z(g27059) ) ;
AND2    gate21129  (.A(g22016), .B(g26626), .Z(g27060) ) ;
AND2    gate21130  (.A(g23372), .B(g26627), .Z(g27061) ) ;
AND2    gate21131  (.A(g22093), .B(g26628), .Z(g27062) ) ;
NAND2   gate21132  (.A(g21971), .B(g22336), .Z(g23388) ) ;
AND2    gate21133  (.A(g23388), .B(g26629), .Z(g27063) ) ;
AND2    gate21134  (.A(g22009), .B(g26631), .Z(g27070) ) ;
AND2    gate21135  (.A(g23353), .B(g26632), .Z(g27071) ) ;
NAND2   gate21136  (.A(g21609), .B(g21634), .Z(g22021) ) ;
AND2    gate21137  (.A(g22021), .B(g26633), .Z(g27072) ) ;
AND2    gate21138  (.A(g23381), .B(g26634), .Z(g27073) ) ;
NAND3   gate21139  (.A(g19521), .B(g21269), .C(g19542), .Z(g22118) ) ;
AND2    gate21140  (.A(g22118), .B(g26635), .Z(g27074) ) ;
AND2    gate21141  (.A(g5024), .B(g26393), .Z(g27076) ) ;
AND2    gate21142  (.A(g22083), .B(g26636), .Z(g27077) ) ;
AND2    gate21143  (.A(g5044), .B(g26401), .Z(g27079) ) ;
AND2    gate21144  (.A(g23377), .B(g26637), .Z(g27080) ) ;
AND2    gate21145  (.A(g22108), .B(g26638), .Z(g27081) ) ;
AND2    gate21146  (.A(g22016), .B(g26639), .Z(g27082) ) ;
AND2    gate21147  (.A(g22093), .B(g26640), .Z(g27083) ) ;
AND2    gate21148  (.A(g23388), .B(g26641), .Z(g27084) ) ;
NAND2   gate21149  (.A(g21803), .B(g21809), .Z(g22134) ) ;
AND2    gate21150  (.A(g22134), .B(g26642), .Z(g27085) ) ;
AND2    gate21151  (.A(g23353), .B(g26643), .Z(g27086) ) ;
AND2    gate21152  (.A(g22021), .B(g26644), .Z(g27087) ) ;
AND2    gate21153  (.A(g23381), .B(g26645), .Z(g27088) ) ;
AND2    gate21154  (.A(g22118), .B(g26646), .Z(g27089) ) ;
NAND2   gate21155  (.A(g21973), .B(g22361), .Z(g23395) ) ;
AND2    gate21156  (.A(g23395), .B(g26647), .Z(g27090) ) ;
AND2    gate21157  (.A(g5142), .B(g26429), .Z(g27091) ) ;
AND2    gate21158  (.A(g5153), .B(g26434), .Z(g27092) ) ;
AND2    gate21159  (.A(g22108), .B(g26648), .Z(g27093) ) ;
AND2    gate21160  (.A(g5173), .B(g26442), .Z(g27095) ) ;
AND2    gate21161  (.A(g23388), .B(g26649), .Z(g27096) ) ;
AND2    gate21162  (.A(g22134), .B(g26650), .Z(g27097) ) ;
AND2    gate21163  (.A(g22021), .B(g26651), .Z(g27098) ) ;
AND2    gate21164  (.A(g22118), .B(g26652), .Z(g27099) ) ;
AND2    gate21165  (.A(g23395), .B(g26653), .Z(g27100) ) ;
NAND2   gate21166  (.A(g21811), .B(g21816), .Z(g22157) ) ;
AND2    gate21167  (.A(g22157), .B(g26654), .Z(g27101) ) ;
AND2    gate21168  (.A(g5235), .B(g26461), .Z(g27103) ) ;
AND2    gate21169  (.A(g5246), .B(g26466), .Z(g27104) ) ;
AND2    gate21170  (.A(g22134), .B(g26656), .Z(g27105) ) ;
AND2    gate21171  (.A(g5266), .B(g26474), .Z(g27107) ) ;
AND2    gate21172  (.A(g23395), .B(g26657), .Z(g27108) ) ;
AND2    gate21173  (.A(g22157), .B(g26658), .Z(g27109) ) ;
AND2    gate21174  (.A(g5298), .B(g26485), .Z(g27110) ) ;
AND2    gate21175  (.A(g5309), .B(g26490), .Z(g27111) ) ;
AND2    gate21176  (.A(g22157), .B(g26662), .Z(g27112) ) ;
AND2    gate21177  (.A(g5335), .B(g26501), .Z(g27115) ) ;
NOR3    gate21178  (.A(g6068), .B(g24183), .C(g25305), .Z(g26110) ) ;
AND2    gate21179  (.A(g26110), .B(g22213), .Z(g27178) ) ;
NOR3    gate21180  (.A(g15904), .B(g15880), .C(g14630), .Z(g16570) ) ;
AND3    gate21181  (.A(g16570), .B(g26508), .C(g13614), .Z(g27181) ) ;
NOR3    gate21182  (.A(g6068), .B(g24183), .C(g25335), .Z(g26151) ) ;
AND2    gate21183  (.A(g26151), .B(g22217), .Z(g27182) ) ;
NOR3    gate21184  (.A(g6068), .B(g24183), .C(g25368), .Z(g26126) ) ;
AND2    gate21185  (.A(g26126), .B(g22230), .Z(g27185) ) ;
NOR3    gate21186  (.A(g15933), .B(g15913), .C(g14650), .Z(g16594) ) ;
AND3    gate21187  (.A(g16594), .B(g26516), .C(g13626), .Z(g27187) ) ;
NOR2    gate21188  (.A(g26096), .B(g22319), .Z(g26905) ) ;
AND2    gate21189  (.A(g26905), .B(g22241), .Z(g27240) ) ;
NAND2   gate21190  (.A(II35124), .B(II35125), .Z(g26934) ) ;
AND2    gate21191  (.A(g10730), .B(g26934), .Z(g27241) ) ;
AND2    gate21192  (.A(g26793), .B(g8357), .Z(g27242) ) ;
NOR2    gate21193  (.A(g26107), .B(g22319), .Z(g26914) ) ;
AND2    gate21194  (.A(g26914), .B(g22258), .Z(g27244) ) ;
NOR2    gate21195  (.A(g26140), .B(g22319), .Z(g26877) ) ;
AND2    gate21196  (.A(g26877), .B(g22286), .Z(g27245) ) ;
NOR2    gate21197  (.A(g24893), .B(g26023), .Z(g26988) ) ;
AND2    gate21198  (.A(g26988), .B(g16676), .Z(g27246) ) ;
NOR2    gate21199  (.A(g24916), .B(g26026), .Z(g27011) ) ;
AND2    gate21200  (.A(g27011), .B(g16702), .Z(g27247) ) ;
NOR2    gate21201  (.A(g24933), .B(g26028), .Z(g27037) ) ;
AND2    gate21202  (.A(g27037), .B(g16733), .Z(g27248) ) ;
NOR2    gate21203  (.A(g24945), .B(g26029), .Z(g27065) ) ;
AND2    gate21204  (.A(g27065), .B(g16775), .Z(g27249) ) ;
AND2    gate21205  (.A(g61), .B(g26837), .Z(g27355) ) ;
AND2    gate21206  (.A(g65), .B(g26987), .Z(g27356) ) ;
AND2    gate21207  (.A(g749), .B(g26846), .Z(g27358) ) ;
AND2    gate21208  (.A(g753), .B(g27010), .Z(g27359) ) ;
AND2    gate21209  (.A(g1435), .B(g26855), .Z(g27364) ) ;
AND2    gate21210  (.A(g1439), .B(g27036), .Z(g27365) ) ;
AND2    gate21211  (.A(g27126), .B(g8874), .Z(g27370) ) ;
AND2    gate21212  (.A(g2129), .B(g26861), .Z(g27371) ) ;
AND2    gate21213  (.A(g2133), .B(g27064), .Z(g27372) ) ;
AND2    gate21214  (.A(g17802), .B(g27134), .Z(g27394) ) ;
AND2    gate21215  (.A(g692), .B(g27135), .Z(g27396) ) ;
AND2    gate21216  (.A(g17914), .B(g27136), .Z(g27407) ) ;
AND2    gate21217  (.A(g1378), .B(g27137), .Z(g27409) ) ;
AND2    gate21218  (.A(g18025), .B(g27138), .Z(g27425) ) ;
AND2    gate21219  (.A(g2072), .B(g27139), .Z(g27427) ) ;
AND2    gate21220  (.A(g18142), .B(g27141), .Z(g27446) ) ;
AND2    gate21221  (.A(g2766), .B(g27142), .Z(g27448) ) ;
NOR3    gate21222  (.A(g4456), .B(g13565), .C(g23009), .Z(g23945) ) ;
AND2    gate21223  (.A(g23945), .B(g27146), .Z(g27495) ) ;
AND2    gate21224  (.A(g23945), .B(g27148), .Z(g27509) ) ;
NOR3    gate21225  (.A(g4632), .B(g13573), .C(g23025), .Z(g23974) ) ;
AND2    gate21226  (.A(g23974), .B(g27151), .Z(g27516) ) ;
AND2    gate21227  (.A(g23945), .B(g27153), .Z(g27530) ) ;
AND2    gate21228  (.A(g23974), .B(g27155), .Z(g27534) ) ;
NOR3    gate21229  (.A(g4809), .B(g13582), .C(g23042), .Z(g24004) ) ;
AND2    gate21230  (.A(g24004), .B(g27159), .Z(g27541) ) ;
AND2    gate21231  (.A(g23974), .B(g27162), .Z(g27552) ) ;
AND2    gate21232  (.A(g24004), .B(g27164), .Z(g27554) ) ;
NOR3    gate21233  (.A(g4985), .B(g13602), .C(g23061), .Z(g24038) ) ;
AND2    gate21234  (.A(g24038), .B(g27167), .Z(g27561) ) ;
AND2    gate21235  (.A(g24004), .B(g27172), .Z(g27568) ) ;
AND2    gate21236  (.A(g24038), .B(g27173), .Z(g27570) ) ;
AND2    gate21237  (.A(g24038), .B(g27177), .Z(g27578) ) ;
AND2    gate21238  (.A(g26796), .B(g11004), .Z(g27656) ) ;
AND2    gate21239  (.A(g27114), .B(g11051), .Z(g27657) ) ;
AND2    gate21240  (.A(g27132), .B(g11114), .Z(g27659) ) ;
AND2    gate21241  (.A(g26835), .B(g11117), .Z(g27660) ) ;
AND2    gate21242  (.A(g26841), .B(g11173), .Z(g27661) ) ;
AND2    gate21243  (.A(g26849), .B(g11243), .Z(g27666) ) ;
NOR2    gate21244  (.A(g26140), .B(g22319), .Z(g26885) ) ;
AND2    gate21245  (.A(g26885), .B(g22212), .Z(g27671) ) ;
AND2    gate21246  (.A(g26854), .B(g11312), .Z(g27673) ) ;
AND2    gate21247  (.A(g26782), .B(g11386), .Z(g27679) ) ;
AND2    gate21248  (.A(g26983), .B(g11392), .Z(g27680) ) ;
AND2    gate21249  (.A(g26788), .B(g11456), .Z(g27681) ) ;
NOR2    gate21250  (.A(g27185), .B(g25178), .Z(g27496) ) ;
AND2    gate21251  (.A(g27496), .B(g20649), .Z(g27719) ) ;
NOR2    gate21252  (.A(g27182), .B(g25980), .Z(g27481) ) ;
AND2    gate21253  (.A(g27481), .B(g20652), .Z(g27720) ) ;
NOR2    gate21254  (.A(g26775), .B(g25192), .Z(g27579) ) ;
AND2    gate21255  (.A(g27579), .B(g20655), .Z(g27721) ) ;
NOR2    gate21256  (.A(g27178), .B(g25975), .Z(g27464) ) ;
AND2    gate21257  (.A(g27464), .B(g20679), .Z(g27723) ) ;
NOR2    gate21258  (.A(g26761), .B(g25182), .Z(g27532) ) ;
AND2    gate21259  (.A(g27532), .B(g20704), .Z(g27725) ) ;
NOR2    gate21260  (.A(g26760), .B(g25181), .Z(g27531) ) ;
AND2    gate21261  (.A(g27531), .B(g20732), .Z(g27726) ) ;
NOR2    gate21262  (.A(g26770), .B(g25187), .Z(g27414) ) ;
AND2    gate21263  (.A(g27414), .B(g19301), .Z(g27727) ) ;
NOR2    gate21264  (.A(g26767), .B(g25184), .Z(g27564) ) ;
AND2    gate21265  (.A(g27564), .B(g20766), .Z(g27728) ) ;
NOR2    gate21266  (.A(g26777), .B(g25193), .Z(g27435) ) ;
AND2    gate21267  (.A(g27435), .B(g19322), .Z(g27729) ) ;
NOR2    gate21268  (.A(g26783), .B(g25196), .Z(g27454) ) ;
AND2    gate21269  (.A(g27454), .B(g19349), .Z(g27730) ) ;
NOR2    gate21270  (.A(g26790), .B(g25198), .Z(g27470) ) ;
AND2    gate21271  (.A(g27470), .B(g19383), .Z(g27731) ) ;
NOR3    gate21272  (.A(g24958), .B(g24633), .C(g26771), .Z(g27492) ) ;
AND2    gate21273  (.A(g27492), .B(g16758), .Z(g27732) ) ;
NOR3    gate21274  (.A(g24969), .B(g24653), .C(g26778), .Z(g27513) ) ;
AND2    gate21275  (.A(g27513), .B(g16785), .Z(g27733) ) ;
NOR3    gate21276  (.A(g24982), .B(g24672), .C(g26784), .Z(g27538) ) ;
AND2    gate21277  (.A(g27538), .B(g16814), .Z(g27734) ) ;
NOR3    gate21278  (.A(g24993), .B(g24691), .C(g26791), .Z(g27558) ) ;
AND2    gate21279  (.A(g27558), .B(g16832), .Z(g27737) ) ;
AND2    gate21280  (.A(g5642), .B(g27449), .Z(g27770) ) ;
AND2    gate21281  (.A(g5680), .B(g27465), .Z(g27772) ) ;
AND2    gate21282  (.A(g5732), .B(g27484), .Z(g27773) ) ;
AND2    gate21283  (.A(g5702), .B(g27361), .Z(g27774) ) ;
AND2    gate21284  (.A(g5790), .B(g27506), .Z(g27775) ) ;
AND2    gate21285  (.A(g5760), .B(g27367), .Z(g27779) ) ;
AND2    gate21286  (.A(g5819), .B(g27373), .Z(g27783) ) ;
AND2    gate21287  (.A(g5875), .B(g27376), .Z(g27790) ) ;
AND2    gate21288  (.A(g13873), .B(g27387), .Z(g27904) ) ;
AND2    gate21289  (.A(g13886), .B(g27391), .Z(g27908) ) ;
AND2    gate21290  (.A(g13895), .B(g27397), .Z(g27909) ) ;
AND2    gate21291  (.A(g4017), .B(g27401), .Z(g27913) ) ;
AND2    gate21292  (.A(g13927), .B(g27404), .Z(g27914) ) ;
AND2    gate21293  (.A(g13936), .B(g27410), .Z(g27915) ) ;
AND2    gate21294  (.A(g4112), .B(g27416), .Z(g27922) ) ;
AND2    gate21295  (.A(g4144), .B(g27419), .Z(g27923) ) ;
AND2    gate21296  (.A(g13983), .B(g27422), .Z(g27924) ) ;
AND2    gate21297  (.A(g13992), .B(g27428), .Z(g27926) ) ;
AND2    gate21298  (.A(g4221), .B(g27432), .Z(g27931) ) ;
AND2    gate21299  (.A(g4251), .B(g27437), .Z(g27935) ) ;
AND2    gate21300  (.A(g4283), .B(g27440), .Z(g27936) ) ;
AND2    gate21301  (.A(g14053), .B(g27443), .Z(g27938) ) ;
AND2    gate21302  (.A(g4376), .B(g27451), .Z(g27945) ) ;
AND2    gate21303  (.A(g4406), .B(g27456), .Z(g27949) ) ;
AND2    gate21304  (.A(g4438), .B(g27459), .Z(g27951) ) ;
AND2    gate21305  (.A(g4545), .B(g27467), .Z(g27963) ) ;
AND2    gate21306  (.A(g4575), .B(g27472), .Z(g27968) ) ;
AND2    gate21307  (.A(g14238), .B(g27475), .Z(g27970) ) ;
AND2    gate21308  (.A(g4721), .B(g27486), .Z(g27984) ) ;
AND2    gate21309  (.A(g14342), .B(g27489), .Z(g27985) ) ;
AND2    gate21310  (.A(g14360), .B(g27498), .Z(g27991) ) ;
AND2    gate21311  (.A(g27590), .B(g9770), .Z(g28008) ) ;
AND2    gate21312  (.A(g14454), .B(g27510), .Z(g28009) ) ;
AND2    gate21313  (.A(g14472), .B(g27518), .Z(g28015) ) ;
AND2    gate21314  (.A(g27590), .B(g9895), .Z(g28027) ) ;
AND2    gate21315  (.A(g27595), .B(g9898), .Z(g28028) ) ;
AND2    gate21316  (.A(g27599), .B(g9916), .Z(g28035) ) ;
AND2    gate21317  (.A(g14541), .B(g27535), .Z(g28036) ) ;
AND2    gate21318  (.A(g14559), .B(g27543), .Z(g28042) ) ;
AND2    gate21319  (.A(g27590), .B(g10018), .Z(g28050) ) ;
AND2    gate21320  (.A(g27595), .B(g10021), .Z(g28051) ) ;
AND2    gate21321  (.A(g27599), .B(g10049), .Z(g28057) ) ;
AND2    gate21322  (.A(g27604), .B(g10052), .Z(g28058) ) ;
AND2    gate21323  (.A(g27608), .B(g10070), .Z(g28065) ) ;
AND2    gate21324  (.A(g14596), .B(g27555), .Z(g28066) ) ;
AND2    gate21325  (.A(g27595), .B(g10109), .Z(g28073) ) ;
AND2    gate21326  (.A(g27599), .B(g10127), .Z(g28079) ) ;
AND2    gate21327  (.A(g27604), .B(g10130), .Z(g28080) ) ;
AND2    gate21328  (.A(g27608), .B(g10158), .Z(g28086) ) ;
AND2    gate21329  (.A(g27613), .B(g10161), .Z(g28087) ) ;
AND2    gate21330  (.A(g27617), .B(g10179), .Z(g28094) ) ;
AND2    gate21331  (.A(g27604), .B(g10214), .Z(g28098) ) ;
AND2    gate21332  (.A(g27608), .B(g10232), .Z(g28104) ) ;
AND2    gate21333  (.A(g27613), .B(g10235), .Z(g28105) ) ;
AND2    gate21334  (.A(g27617), .B(g10263), .Z(g28111) ) ;
AND2    gate21335  (.A(g27622), .B(g10266), .Z(g28112) ) ;
AND2    gate21336  (.A(g27613), .B(g10316), .Z(g28116) ) ;
AND2    gate21337  (.A(g27617), .B(g10334), .Z(g28122) ) ;
AND2    gate21338  (.A(g27622), .B(g10337), .Z(g28123) ) ;
AND2    gate21339  (.A(g27622), .B(g10409), .Z(g28127) ) ;
AND2    gate21340  (.A(g27349), .B(g10898), .Z(g28171) ) ;
AND2    gate21341  (.A(g27349), .B(g10940), .Z(g28176) ) ;
AND2    gate21342  (.A(g27349), .B(g11008), .Z(g28188) ) ;
NOR2    gate21343  (.A(g26773), .B(g25188), .Z(g27573) ) ;
AND2    gate21344  (.A(g27573), .B(g21914), .Z(g28193) ) ;
NOR3    gate21345  (.A(g6087), .B(g27632), .C(g25385), .Z(g27855) ) ;
AND2    gate21346  (.A(g27855), .B(g22246), .Z(g28319) ) ;
NOR2    gate21347  (.A(g27632), .B(g1218), .Z(g27854) ) ;
AND2    gate21348  (.A(g27854), .B(g20637), .Z(g28320) ) ;
NOR2    gate21349  (.A(g16321), .B(g27666), .Z(g27937) ) ;
AND2    gate21350  (.A(g27937), .B(g13868), .Z(g28322) ) ;
NAND2   gate21351  (.A(II36301), .B(II36302), .Z(g27838) ) ;
AND2    gate21352  (.A(g8580), .B(g27838), .Z(g28323) ) ;
NOR2    gate21353  (.A(g27632), .B(g1215), .Z(g27810) ) ;
AND2    gate21354  (.A(g27810), .B(g20659), .Z(g28324) ) ;
NOR3    gate21355  (.A(g6087), .B(g27632), .C(g25370), .Z(g27865) ) ;
AND2    gate21356  (.A(g27865), .B(g22274), .Z(g28326) ) ;
NOR3    gate21357  (.A(g6087), .B(g27632), .C(g25338), .Z(g27900) ) ;
AND2    gate21358  (.A(g27900), .B(g22275), .Z(g28327) ) ;
NOR2    gate21359  (.A(g27632), .B(g1216), .Z(g27823) ) ;
AND2    gate21360  (.A(g27823), .B(g20708), .Z(g28329) ) ;
NOR2    gate21361  (.A(g27632), .B(g1219), .Z(g27864) ) ;
AND2    gate21362  (.A(g27864), .B(g20711), .Z(g28330) ) ;
NOR3    gate21363  (.A(g6087), .B(g27632), .C(g25330), .Z(g27802) ) ;
AND2    gate21364  (.A(g27802), .B(g22307), .Z(g28331) ) ;
NOR3    gate21365  (.A(g6087), .B(g27632), .C(g25361), .Z(g27883) ) ;
AND2    gate21366  (.A(g27883), .B(g22331), .Z(g28332) ) ;
NOR2    gate21367  (.A(g27632), .B(g1220), .Z(g27882) ) ;
AND2    gate21368  (.A(g27882), .B(g20772), .Z(g28333) ) ;
NOR2    gate21369  (.A(g27632), .B(g1217), .Z(g27842) ) ;
AND2    gate21370  (.A(g27842), .B(g20793), .Z(g28334) ) ;
NOR3    gate21371  (.A(g6087), .B(g27632), .C(g25322), .Z(g27814) ) ;
AND2    gate21372  (.A(g27814), .B(g22343), .Z(g28335) ) ;
NOR2    gate21373  (.A(g27632), .B(g1222), .Z(g27896) ) ;
AND2    gate21374  (.A(g27896), .B(g20810), .Z(g28336) ) ;
NOR2    gate21375  (.A(g26032), .B(g27246), .Z(g28002) ) ;
AND2    gate21376  (.A(g28002), .B(g19448), .Z(g28337) ) ;
NOR2    gate21377  (.A(g26033), .B(g27247), .Z(g28029) ) ;
AND2    gate21378  (.A(g28029), .B(g19475), .Z(g28338) ) ;
NOR2    gate21379  (.A(g26034), .B(g27248), .Z(g28059) ) ;
AND2    gate21380  (.A(g28059), .B(g19498), .Z(g28339) ) ;
NOR2    gate21381  (.A(g26036), .B(g27249), .Z(g28088) ) ;
AND2    gate21382  (.A(g28088), .B(g19519), .Z(g28340) ) ;
AND2    gate21383  (.A(g56), .B(g27969), .Z(g28373) ) ;
AND2    gate21384  (.A(g744), .B(g27990), .Z(g28376) ) ;
AND2    gate21385  (.A(g52), .B(g27776), .Z(g28378) ) ;
NOR2    gate21386  (.A(g23742), .B(g27632), .Z(g27868) ) ;
AND3    gate21387  (.A(g27868), .B(g19390), .C(g19369), .Z(g28379) ) ;
AND2    gate21388  (.A(g1430), .B(g28014), .Z(g28380) ) ;
NOR2    gate21389  (.A(g13902), .B(g27370), .Z(g28157) ) ;
AND2    gate21390  (.A(g28157), .B(g9815), .Z(g28381) ) ;
AND2    gate21391  (.A(g740), .B(g27780), .Z(g28383) ) ;
AND2    gate21392  (.A(g2124), .B(g28041), .Z(g28385) ) ;
AND2    gate21393  (.A(g1426), .B(g27787), .Z(g28387) ) ;
AND2    gate21394  (.A(g2120), .B(g27794), .Z(g28389) ) ;
AND2    gate21395  (.A(g7754), .B(g27806), .Z(g28396) ) ;
AND2    gate21396  (.A(g7769), .B(g27817), .Z(g28398) ) ;
AND2    gate21397  (.A(g7776), .B(g27820), .Z(g28399) ) ;
AND2    gate21398  (.A(g7782), .B(g27831), .Z(g28401) ) ;
AND2    gate21399  (.A(g7785), .B(g27839), .Z(g28402) ) ;
AND2    gate21400  (.A(g7792), .B(g27843), .Z(g28404) ) ;
AND2    gate21401  (.A(g7796), .B(g27847), .Z(g28405) ) ;
AND2    gate21402  (.A(g7799), .B(g27858), .Z(g28407) ) ;
AND2    gate21403  (.A(g7806), .B(g27861), .Z(g28408) ) ;
AND2    gate21404  (.A(g7809), .B(g27872), .Z(g28411) ) ;
AND2    gate21405  (.A(g7812), .B(g27879), .Z(g28412) ) ;
AND2    gate21406  (.A(g7823), .B(g27889), .Z(g28416) ) ;
AND2    gate21407  (.A(g17640), .B(g28150), .Z(g28422) ) ;
AND2    gate21408  (.A(g17724), .B(g28152), .Z(g28423) ) ;
AND2    gate21409  (.A(g17741), .B(g28153), .Z(g28424) ) ;
AND2    gate21410  (.A(g28128), .B(g9170), .Z(g28426) ) ;
AND2    gate21411  (.A(g26092), .B(g28154), .Z(g28427) ) ;
AND2    gate21412  (.A(g17825), .B(g28155), .Z(g28428) ) ;
AND2    gate21413  (.A(g17842), .B(g28156), .Z(g28429) ) ;
AND2    gate21414  (.A(g28128), .B(g9196), .Z(g28430) ) ;
AND2    gate21415  (.A(g26092), .B(g28158), .Z(g28431) ) ;
AND2    gate21416  (.A(g28133), .B(g9212), .Z(g28433) ) ;
AND2    gate21417  (.A(g26114), .B(g28159), .Z(g28434) ) ;
AND2    gate21418  (.A(g17937), .B(g28160), .Z(g28435) ) ;
AND2    gate21419  (.A(g17954), .B(g28161), .Z(g28436) ) ;
AND2    gate21420  (.A(g17882), .B(g27919), .Z(g28438) ) ;
AND2    gate21421  (.A(g28128), .B(g9242), .Z(g28439) ) ;
AND2    gate21422  (.A(g26092), .B(g28162), .Z(g28440) ) ;
AND2    gate21423  (.A(g28133), .B(g9257), .Z(g28441) ) ;
AND2    gate21424  (.A(g26114), .B(g28163), .Z(g28442) ) ;
AND2    gate21425  (.A(g28137), .B(g9273), .Z(g28444) ) ;
AND2    gate21426  (.A(g26121), .B(g28164), .Z(g28445) ) ;
AND2    gate21427  (.A(g18048), .B(g28165), .Z(g28446) ) ;
AND2    gate21428  (.A(g17974), .B(g27928), .Z(g28448) ) ;
AND2    gate21429  (.A(g17993), .B(g27932), .Z(g28450) ) ;
AND2    gate21430  (.A(g28133), .B(g9320), .Z(g28451) ) ;
AND2    gate21431  (.A(g26114), .B(g28166), .Z(g28452) ) ;
AND2    gate21432  (.A(g28137), .B(g9335), .Z(g28453) ) ;
AND2    gate21433  (.A(g26121), .B(g28167), .Z(g28454) ) ;
AND2    gate21434  (.A(g28141), .B(g9351), .Z(g28456) ) ;
AND2    gate21435  (.A(g26131), .B(g28168), .Z(g28457) ) ;
AND2    gate21436  (.A(g18074), .B(g27939), .Z(g28459) ) ;
AND2    gate21437  (.A(g18091), .B(g27942), .Z(g28460) ) ;
AND2    gate21438  (.A(g18110), .B(g27946), .Z(g28462) ) ;
AND2    gate21439  (.A(g28137), .B(g9401), .Z(g28463) ) ;
AND2    gate21440  (.A(g26121), .B(g28169), .Z(g28464) ) ;
AND2    gate21441  (.A(g28141), .B(g9416), .Z(g28465) ) ;
AND2    gate21442  (.A(g26131), .B(g28170), .Z(g28466) ) ;
AND2    gate21443  (.A(g18265), .B(g28172), .Z(g28468) ) ;
AND2    gate21444  (.A(g18179), .B(g27952), .Z(g28469) ) ;
AND2    gate21445  (.A(g18190), .B(g27956), .Z(g28471) ) ;
AND2    gate21446  (.A(g18207), .B(g27959), .Z(g28472) ) ;
AND2    gate21447  (.A(g18226), .B(g27965), .Z(g28474) ) ;
AND2    gate21448  (.A(g28141), .B(g9498), .Z(g28475) ) ;
AND2    gate21449  (.A(g26131), .B(g28173), .Z(g28476) ) ;
AND2    gate21450  (.A(g18341), .B(g28174), .Z(g28477) ) ;
AND2    gate21451  (.A(g18358), .B(g28175), .Z(g28478) ) ;
AND2    gate21452  (.A(g18286), .B(g27973), .Z(g28479) ) ;
AND2    gate21453  (.A(g18297), .B(g27977), .Z(g28480) ) ;
AND2    gate21454  (.A(g18314), .B(g27981), .Z(g28481) ) ;
AND2    gate21455  (.A(g18436), .B(g28177), .Z(g28484) ) ;
AND2    gate21456  (.A(g18453), .B(g28178), .Z(g28485) ) ;
AND2    gate21457  (.A(g18379), .B(g27994), .Z(g28486) ) ;
AND2    gate21458  (.A(g18390), .B(g27999), .Z(g28487) ) ;
AND2    gate21459  (.A(g18509), .B(g28186), .Z(g28492) ) ;
AND2    gate21460  (.A(g18526), .B(g28187), .Z(g28493) ) ;
AND2    gate21461  (.A(g18474), .B(g28018), .Z(g28494) ) ;
AND2    gate21462  (.A(g18573), .B(g28190), .Z(g28497) ) ;
NOR2    gate21463  (.A(g16276), .B(g27661), .Z(g27925) ) ;
AND2    gate21464  (.A(g27925), .B(g13700), .Z(g28657) ) ;
NOR2    gate21465  (.A(g16220), .B(g27660), .Z(g27917) ) ;
AND2    gate21466  (.A(g27917), .B(g13736), .Z(g28659) ) ;
NOR2    gate21467  (.A(g16219), .B(g27659), .Z(g27916) ) ;
AND2    gate21468  (.A(g27916), .B(g11911), .Z(g28660) ) ;
NOR2    gate21469  (.A(g16170), .B(g27657), .Z(g27911) ) ;
AND2    gate21470  (.A(g27911), .B(g11951), .Z(g28662) ) ;
NOR2    gate21471  (.A(g16127), .B(g27656), .Z(g27906) ) ;
AND2    gate21472  (.A(g27906), .B(g11997), .Z(g28663) ) ;
NOR2    gate21473  (.A(g16456), .B(g27242), .Z(g27997) ) ;
AND2    gate21474  (.A(g27997), .B(g12055), .Z(g28664) ) ;
NOR3    gate21475  (.A(g6087), .B(g27632), .C(g25314), .Z(g27827) ) ;
AND2    gate21476  (.A(g27827), .B(g22222), .Z(g28665) ) ;
NOR2    gate21477  (.A(g16428), .B(g27681), .Z(g27980) ) ;
AND2    gate21478  (.A(g27980), .B(g12106), .Z(g28666) ) ;
NOR2    gate21479  (.A(g16400), .B(g27680), .Z(g27964) ) ;
AND2    gate21480  (.A(g27964), .B(g13852), .Z(g28667) ) ;
NOR3    gate21481  (.A(g6087), .B(g27632), .C(g25349), .Z(g27897) ) ;
AND2    gate21482  (.A(g27897), .B(g22233), .Z(g28669) ) ;
NOR2    gate21483  (.A(g27632), .B(g1223), .Z(g27798) ) ;
AND2    gate21484  (.A(g27798), .B(g21935), .Z(g28670) ) ;
NOR2    gate21485  (.A(g16394), .B(g27679), .Z(g27962) ) ;
AND2    gate21486  (.A(g27962), .B(g12161), .Z(g28671) ) ;
NOR2    gate21487  (.A(g16367), .B(g27673), .Z(g27950) ) ;
AND2    gate21488  (.A(g27950), .B(g13859), .Z(g28672) ) ;
NOR2    gate21489  (.A(g8587), .B(g10749), .Z(g12436) ) ;
AND2    gate21490  (.A(g12436), .B(g28379), .Z(g28707) ) ;
NOR2    gate21491  (.A(g27886), .B(g22344), .Z(g28392) ) ;
AND2    gate21492  (.A(g28392), .B(g22260), .Z(g28708) ) ;
NOR2    gate21493  (.A(g27886), .B(g22344), .Z(g28400) ) ;
AND2    gate21494  (.A(g28400), .B(g22261), .Z(g28709) ) ;
NOR2    gate21495  (.A(g27811), .B(g22344), .Z(g28403) ) ;
AND2    gate21496  (.A(g28403), .B(g22262), .Z(g28710) ) ;
NAND2   gate21497  (.A(II37357), .B(II37358), .Z(g28415) ) ;
AND2    gate21498  (.A(g10749), .B(g28415), .Z(g28711) ) ;
NOR2    gate21499  (.A(g27824), .B(g22344), .Z(g28406) ) ;
AND2    gate21500  (.A(g28406), .B(g22276), .Z(g28712) ) ;
NOR2    gate21501  (.A(g27748), .B(g22344), .Z(g28410) ) ;
AND2    gate21502  (.A(g28410), .B(g22290), .Z(g28713) ) ;
NOR2    gate21503  (.A(g27869), .B(g22344), .Z(g28394) ) ;
AND2    gate21504  (.A(g28394), .B(g22306), .Z(g28714) ) ;
NOR2    gate21505  (.A(g27748), .B(g22344), .Z(g28414) ) ;
AND2    gate21506  (.A(g28414), .B(g22332), .Z(g28715) ) ;
NOR2    gate21507  (.A(g27727), .B(g26780), .Z(g28449) ) ;
AND2    gate21508  (.A(g28449), .B(g19319), .Z(g28716) ) ;
NOR2    gate21509  (.A(g27729), .B(g26787), .Z(g28461) ) ;
AND2    gate21510  (.A(g28461), .B(g19346), .Z(g28717) ) ;
NOR2    gate21511  (.A(g27730), .B(g26794), .Z(g28473) ) ;
AND2    gate21512  (.A(g28473), .B(g19380), .Z(g28718) ) ;
NOR2    gate21513  (.A(g27731), .B(g26797), .Z(g28482) ) ;
AND2    gate21514  (.A(g28482), .B(g19412), .Z(g28719) ) ;
NOR2    gate21515  (.A(g26035), .B(g27732), .Z(g28523) ) ;
AND2    gate21516  (.A(g28523), .B(g16694), .Z(g28722) ) ;
NOR2    gate21517  (.A(g26038), .B(g27733), .Z(g28551) ) ;
AND2    gate21518  (.A(g28551), .B(g16725), .Z(g28724) ) ;
NOR2    gate21519  (.A(g26039), .B(g27734), .Z(g28578) ) ;
AND2    gate21520  (.A(g28578), .B(g16767), .Z(g28726) ) ;
NOR2    gate21521  (.A(g26040), .B(g27737), .Z(g28606) ) ;
AND2    gate21522  (.A(g28606), .B(g16794), .Z(g28729) ) ;
AND2    gate21523  (.A(g5751), .B(g28483), .Z(g28834) ) ;
AND2    gate21524  (.A(g5810), .B(g28491), .Z(g28836) ) ;
AND2    gate21525  (.A(g5866), .B(g28496), .Z(g28838) ) ;
AND2    gate21526  (.A(g5913), .B(g28500), .Z(g28840) ) ;
NOR2    gate21527  (.A(g27478), .B(g14630), .Z(g27834) ) ;
AND2    gate21528  (.A(g27834), .B(g28554), .Z(g28841) ) ;
AND2    gate21529  (.A(g27834), .B(g28581), .Z(g28843) ) ;
NOR2    gate21530  (.A(g27501), .B(g14650), .Z(g27850) ) ;
AND2    gate21531  (.A(g27850), .B(g28582), .Z(g28844) ) ;
AND2    gate21532  (.A(g27834), .B(g28608), .Z(g28846) ) ;
AND2    gate21533  (.A(g27850), .B(g28609), .Z(g28847) ) ;
NOR2    gate21534  (.A(g27521), .B(g14677), .Z(g27875) ) ;
AND2    gate21535  (.A(g27875), .B(g28610), .Z(g28848) ) ;
AND2    gate21536  (.A(g27850), .B(g28616), .Z(g28849) ) ;
AND2    gate21537  (.A(g27875), .B(g28617), .Z(g28850) ) ;
NOR2    gate21538  (.A(g27546), .B(g14711), .Z(g27892) ) ;
AND2    gate21539  (.A(g27892), .B(g28618), .Z(g28851) ) ;
AND2    gate21540  (.A(g27875), .B(g28623), .Z(g28852) ) ;
AND2    gate21541  (.A(g27892), .B(g28624), .Z(g28853) ) ;
AND2    gate21542  (.A(g27892), .B(g28629), .Z(g28854) ) ;
AND2    gate21543  (.A(g13946), .B(g28639), .Z(g28880) ) ;
AND2    gate21544  (.A(g28612), .B(g9199), .Z(g28881) ) ;
AND2    gate21545  (.A(g14001), .B(g28640), .Z(g28892) ) ;
AND2    gate21546  (.A(g28612), .B(g9245), .Z(g28893) ) ;
AND2    gate21547  (.A(g14016), .B(g28641), .Z(g28897) ) ;
AND2    gate21548  (.A(g28619), .B(g9260), .Z(g28898) ) ;
AND2    gate21549  (.A(g14062), .B(g28642), .Z(g28909) ) ;
AND2    gate21550  (.A(g28612), .B(g9303), .Z(g28910) ) ;
AND2    gate21551  (.A(g14092), .B(g28643), .Z(g28914) ) ;
AND2    gate21552  (.A(g28619), .B(g9323), .Z(g28915) ) ;
AND2    gate21553  (.A(g14107), .B(g28644), .Z(g28919) ) ;
AND2    gate21554  (.A(g28625), .B(g9338), .Z(g28923) ) ;
AND2    gate21555  (.A(g14153), .B(g28645), .Z(g28931) ) ;
AND2    gate21556  (.A(g14177), .B(g28646), .Z(g28935) ) ;
AND2    gate21557  (.A(g28619), .B(g9384), .Z(g28936) ) ;
AND2    gate21558  (.A(g14207), .B(g28647), .Z(g28940) ) ;
AND2    gate21559  (.A(g28625), .B(g9404), .Z(g28944) ) ;
AND2    gate21560  (.A(g14222), .B(g28648), .Z(g28948) ) ;
AND2    gate21561  (.A(g28630), .B(g9419), .Z(g28949) ) ;
AND2    gate21562  (.A(g14268), .B(g28649), .Z(g28958) ) ;
AND2    gate21563  (.A(g14292), .B(g28650), .Z(g28962) ) ;
AND2    gate21564  (.A(g28625), .B(g9481), .Z(g28966) ) ;
AND2    gate21565  (.A(g14322), .B(g28651), .Z(g28970) ) ;
AND2    gate21566  (.A(g28630), .B(g9501), .Z(g28971) ) ;
AND2    gate21567  (.A(g14390), .B(g28652), .Z(g28986) ) ;
AND2    gate21568  (.A(g14414), .B(g28653), .Z(g28996) ) ;
AND2    gate21569  (.A(g28630), .B(g9623), .Z(g28997) ) ;
AND2    gate21570  (.A(g14502), .B(g28655), .Z(g29022) ) ;
NOR2    gate21571  (.A(g27869), .B(g22344), .Z(g28397) ) ;
AND2    gate21572  (.A(g28397), .B(g22221), .Z(g29130) ) ;
NOR2    gate21573  (.A(g28319), .B(g28324), .Z(g29031) ) ;
AND2    gate21574  (.A(g29031), .B(g20684), .Z(g29174) ) ;
NOR2    gate21575  (.A(g28669), .B(g28320), .Z(g29009) ) ;
AND2    gate21576  (.A(g29009), .B(g20687), .Z(g29175) ) ;
NOR2    gate21577  (.A(g28335), .B(g28336), .Z(g29097) ) ;
AND2    gate21578  (.A(g29097), .B(g20690), .Z(g29176) ) ;
NOR2    gate21579  (.A(g28665), .B(g28670), .Z(g28982) ) ;
AND2    gate21580  (.A(g28982), .B(g20714), .Z(g29180) ) ;
NOR2    gate21581  (.A(g28327), .B(g28330), .Z(g29064) ) ;
AND2    gate21582  (.A(g29064), .B(g20739), .Z(g29183) ) ;
NOR2    gate21583  (.A(g28326), .B(g28329), .Z(g29063) ) ;
AND2    gate21584  (.A(g29063), .B(g20769), .Z(g29186) ) ;
NOR2    gate21585  (.A(g28331), .B(g28333), .Z(g29083) ) ;
AND2    gate21586  (.A(g29083), .B(g20796), .Z(g29188) ) ;
AND2    gate21587  (.A(g15022), .B(g28741), .Z(g29196) ) ;
AND2    gate21588  (.A(g15096), .B(g28751), .Z(g29200) ) ;
AND2    gate21589  (.A(g15118), .B(g28755), .Z(g29203) ) ;
AND2    gate21590  (.A(g15188), .B(g28764), .Z(g29208) ) ;
AND2    gate21591  (.A(g15210), .B(g28768), .Z(g29211) ) ;
AND2    gate21592  (.A(g15274), .B(g28775), .Z(g29217) ) ;
AND2    gate21593  (.A(g15296), .B(g28779), .Z(g29220) ) ;
AND2    gate21594  (.A(g15366), .B(g28785), .Z(g29225) ) ;
AND2    gate21595  (.A(g9293), .B(g28791), .Z(g29229) ) ;
AND2    gate21596  (.A(g9356), .B(g28796), .Z(g29232) ) ;
AND2    gate21597  (.A(g9374), .B(g28799), .Z(g29233) ) ;
AND2    gate21598  (.A(g9427), .B(g28804), .Z(g29234) ) ;
AND2    gate21599  (.A(g9453), .B(g28807), .Z(g29235) ) ;
AND2    gate21600  (.A(g9471), .B(g28810), .Z(g29236) ) ;
AND2    gate21601  (.A(g9569), .B(g28814), .Z(g29238) ) ;
AND2    gate21602  (.A(g9595), .B(g28817), .Z(g29239) ) ;
AND2    gate21603  (.A(g9613), .B(g28820), .Z(g29240) ) ;
AND2    gate21604  (.A(g9711), .B(g28823), .Z(g29241) ) ;
AND2    gate21605  (.A(g9737), .B(g28826), .Z(g29242) ) ;
AND2    gate21606  (.A(g9857), .B(g28829), .Z(g29243) ) ;
AND2    gate21607  (.A(g28855), .B(g8836), .Z(g29248) ) ;
AND2    gate21608  (.A(g28855), .B(g8856), .Z(g29251) ) ;
AND2    gate21609  (.A(g28859), .B(g8863), .Z(g29252) ) ;
AND2    gate21610  (.A(g28855), .B(g8885), .Z(g29255) ) ;
AND2    gate21611  (.A(g28859), .B(g8894), .Z(g29256) ) ;
AND2    gate21612  (.A(g28863), .B(g8901), .Z(g29257) ) ;
AND2    gate21613  (.A(g28859), .B(g8925), .Z(g29259) ) ;
AND2    gate21614  (.A(g28863), .B(g8934), .Z(g29260) ) ;
AND2    gate21615  (.A(g28867), .B(g8941), .Z(g29261) ) ;
AND2    gate21616  (.A(g28863), .B(g8965), .Z(g29262) ) ;
AND2    gate21617  (.A(g28867), .B(g8974), .Z(g29263) ) ;
AND2    gate21618  (.A(g28867), .B(g8997), .Z(g29264) ) ;
NAND2   gate21619  (.A(g9161), .B(g28512), .Z(g29001) ) ;
AND2    gate21620  (.A(g29001), .B(g28871), .Z(g29284) ) ;
NAND2   gate21621  (.A(g9203), .B(g28540), .Z(g29030) ) ;
AND2    gate21622  (.A(g29030), .B(g28883), .Z(g29289) ) ;
NAND2   gate21623  (.A(g9264), .B(g28567), .Z(g29053) ) ;
AND2    gate21624  (.A(g29053), .B(g28900), .Z(g29294) ) ;
NAND2   gate21625  (.A(g9342), .B(g28595), .Z(g29072) ) ;
AND2    gate21626  (.A(g29072), .B(g28925), .Z(g29300) ) ;
NAND2   gate21627  (.A(g9187), .B(g28512), .Z(g29026) ) ;
AND2    gate21628  (.A(g29026), .B(g28928), .Z(g29302) ) ;
NAND2   gate21629  (.A(g9150), .B(g28512), .Z(g28978) ) ;
AND2    gate21630  (.A(g28978), .B(g28951), .Z(g29310) ) ;
NAND2   gate21631  (.A(g9248), .B(g28540), .Z(g29049) ) ;
AND2    gate21632  (.A(g29049), .B(g28955), .Z(g29312) ) ;
NAND2   gate21633  (.A(g9507), .B(g28512), .Z(g29088) ) ;
AND2    gate21634  (.A(g29088), .B(g28972), .Z(g29320) ) ;
NAND2   gate21635  (.A(g9174), .B(g28540), .Z(g29008) ) ;
AND2    gate21636  (.A(g29008), .B(g28979), .Z(g29321) ) ;
NAND2   gate21637  (.A(g9326), .B(g28567), .Z(g29068) ) ;
AND2    gate21638  (.A(g29068), .B(g28983), .Z(g29323) ) ;
NAND2   gate21639  (.A(g9649), .B(g28540), .Z(g29096) ) ;
AND2    gate21640  (.A(g29096), .B(g29002), .Z(g29329) ) ;
NAND2   gate21641  (.A(g9216), .B(g28567), .Z(g29038) ) ;
AND2    gate21642  (.A(g29038), .B(g29010), .Z(g29330) ) ;
NAND2   gate21643  (.A(g9407), .B(g28595), .Z(g29080) ) ;
AND2    gate21644  (.A(g29080), .B(g29019), .Z(g29332) ) ;
NAND2   gate21645  (.A(g9232), .B(g28512), .Z(g29045) ) ;
AND2    gate21646  (.A(g29045), .B(g29023), .Z(g29336) ) ;
NAND2   gate21647  (.A(g9795), .B(g28567), .Z(g29103) ) ;
AND2    gate21648  (.A(g29103), .B(g29032), .Z(g29337) ) ;
NAND2   gate21649  (.A(g9277), .B(g28595), .Z(g29060) ) ;
AND2    gate21650  (.A(g29060), .B(g29042), .Z(g29338) ) ;
NAND2   gate21651  (.A(g9310), .B(g28540), .Z(g29062) ) ;
AND2    gate21652  (.A(g29062), .B(g29046), .Z(g29341) ) ;
NAND2   gate21653  (.A(g9941), .B(g28595), .Z(g29107) ) ;
AND2    gate21654  (.A(g29107), .B(g29054), .Z(g29342) ) ;
NAND2   gate21655  (.A(g9391), .B(g28567), .Z(g29076) ) ;
AND2    gate21656  (.A(g29076), .B(g29065), .Z(g29344) ) ;
NAND2   gate21657  (.A(g9488), .B(g28595), .Z(g29087) ) ;
AND2    gate21658  (.A(g29087), .B(g29077), .Z(g29346) ) ;
NOR2    gate21659  (.A(g28332), .B(g28334), .Z(g29090) ) ;
AND2    gate21660  (.A(g29090), .B(g21932), .Z(g29411) ) ;
AND2    gate21661  (.A(g29190), .B(g8375), .Z(g29464) ) ;
AND2    gate21662  (.A(g29191), .B(g8424), .Z(g29465) ) ;
NAND2   gate21663  (.A(II38379), .B(II38380), .Z(g29265) ) ;
AND2    gate21664  (.A(g8587), .B(g29265), .Z(g29466) ) ;
NOR2    gate21665  (.A(g28337), .B(g28722), .Z(g29340) ) ;
AND2    gate21666  (.A(g29340), .B(g19467), .Z(g29467) ) ;
NOR2    gate21667  (.A(g28338), .B(g28724), .Z(g29343) ) ;
AND2    gate21668  (.A(g29343), .B(g19490), .Z(g29468) ) ;
NOR2    gate21669  (.A(g28339), .B(g28726), .Z(g29345) ) ;
AND2    gate21670  (.A(g29345), .B(g19511), .Z(g29469) ) ;
NOR2    gate21671  (.A(g28340), .B(g28729), .Z(g29347) ) ;
AND2    gate21672  (.A(g29347), .B(g19530), .Z(g29470) ) ;
AND2    gate21673  (.A(g21461), .B(g29266), .Z(g29471) ) ;
AND2    gate21674  (.A(g21461), .B(g29268), .Z(g29472) ) ;
AND2    gate21675  (.A(g21508), .B(g29269), .Z(g29473) ) ;
AND2    gate21676  (.A(g21508), .B(g29271), .Z(g29474) ) ;
AND2    gate21677  (.A(g21544), .B(g29272), .Z(g29475) ) ;
AND2    gate21678  (.A(g21544), .B(g29274), .Z(g29476) ) ;
AND2    gate21679  (.A(g21580), .B(g29275), .Z(g29477) ) ;
AND2    gate21680  (.A(g21580), .B(g29277), .Z(g29478) ) ;
AND2    gate21681  (.A(g21461), .B(g29280), .Z(g29479) ) ;
AND2    gate21682  (.A(g21461), .B(g29282), .Z(g29480) ) ;
AND2    gate21683  (.A(g21508), .B(g29283), .Z(g29481) ) ;
AND2    gate21684  (.A(g21461), .B(g29285), .Z(g29482) ) ;
AND2    gate21685  (.A(g21508), .B(g29286), .Z(g29483) ) ;
AND2    gate21686  (.A(g21544), .B(g29287), .Z(g29484) ) ;
AND2    gate21687  (.A(g21508), .B(g29290), .Z(g29485) ) ;
AND2    gate21688  (.A(g21544), .B(g29291), .Z(g29486) ) ;
AND2    gate21689  (.A(g21580), .B(g29292), .Z(g29487) ) ;
AND2    gate21690  (.A(g21544), .B(g29295), .Z(g29488) ) ;
AND2    gate21691  (.A(g21580), .B(g29296), .Z(g29489) ) ;
AND2    gate21692  (.A(g21580), .B(g29301), .Z(g29490) ) ;
AND2    gate21693  (.A(g29350), .B(g8912), .Z(g29502) ) ;
NOR2    gate21694  (.A(g28422), .B(g27904), .Z(g28728) ) ;
AND2    gate21695  (.A(g28728), .B(g29360), .Z(g29518) ) ;
NOR2    gate21696  (.A(g28423), .B(g27908), .Z(g28731) ) ;
AND2    gate21697  (.A(g28731), .B(g29361), .Z(g29520) ) ;
NOR2    gate21698  (.A(g28424), .B(g27909), .Z(g28733) ) ;
AND2    gate21699  (.A(g28733), .B(g29362), .Z(g29521) ) ;
NOR2    gate21700  (.A(g27394), .B(g26961), .Z(g27735) ) ;
AND2    gate21701  (.A(g27735), .B(g29363), .Z(g29522) ) ;
NOR2    gate21702  (.A(g28428), .B(g27914), .Z(g28737) ) ;
AND2    gate21703  (.A(g28737), .B(g29364), .Z(g29523) ) ;
NOR2    gate21704  (.A(g28429), .B(g27915), .Z(g28739) ) ;
AND2    gate21705  (.A(g28739), .B(g29365), .Z(g29524) ) ;
NOR2    gate21706  (.A(g28880), .B(g28438), .Z(g29195) ) ;
AND2    gate21707  (.A(g29195), .B(g29366), .Z(g29525) ) ;
NOR2    gate21708  (.A(g27407), .B(g26966), .Z(g27741) ) ;
AND2    gate21709  (.A(g27741), .B(g29367), .Z(g29526) ) ;
NOR2    gate21710  (.A(g28435), .B(g27924), .Z(g28748) ) ;
AND2    gate21711  (.A(g28748), .B(g29368), .Z(g29527) ) ;
NOR2    gate21712  (.A(g28436), .B(g27926), .Z(g28750) ) ;
AND2    gate21713  (.A(g28750), .B(g29369), .Z(g29528) ) ;
NOR2    gate21714  (.A(g28892), .B(g28448), .Z(g29199) ) ;
AND2    gate21715  (.A(g29199), .B(g29370), .Z(g29529) ) ;
NOR2    gate21716  (.A(g28897), .B(g28450), .Z(g29202) ) ;
AND2    gate21717  (.A(g29202), .B(g29371), .Z(g29531) ) ;
NOR2    gate21718  (.A(g27425), .B(g26972), .Z(g27746) ) ;
AND2    gate21719  (.A(g27746), .B(g29372), .Z(g29532) ) ;
NOR2    gate21720  (.A(g28446), .B(g27938), .Z(g28762) ) ;
AND2    gate21721  (.A(g28762), .B(g29373), .Z(g29533) ) ;
NOR2    gate21722  (.A(g28909), .B(g28459), .Z(g29206) ) ;
AND2    gate21723  (.A(g29206), .B(g29374), .Z(g29534) ) ;
NOR2    gate21724  (.A(g28914), .B(g28460), .Z(g29207) ) ;
AND2    gate21725  (.A(g29207), .B(g29375), .Z(g29536) ) ;
NOR2    gate21726  (.A(g28919), .B(g28462), .Z(g29210) ) ;
AND2    gate21727  (.A(g29210), .B(g29376), .Z(g29538) ) ;
NOR2    gate21728  (.A(g27446), .B(g26985), .Z(g27754) ) ;
AND2    gate21729  (.A(g27754), .B(g29377), .Z(g29539) ) ;
NOR2    gate21730  (.A(g25475), .B(g24855), .Z(g26041) ) ;
AND2    gate21731  (.A(g26041), .B(g29378), .Z(g29540) ) ;
NOR2    gate21732  (.A(g28931), .B(g28469), .Z(g29214) ) ;
AND2    gate21733  (.A(g29214), .B(g29379), .Z(g29541) ) ;
NOR2    gate21734  (.A(g28935), .B(g28471), .Z(g29215) ) ;
AND2    gate21735  (.A(g29215), .B(g29380), .Z(g29543) ) ;
NOR2    gate21736  (.A(g28940), .B(g28472), .Z(g29216) ) ;
AND2    gate21737  (.A(g29216), .B(g29381), .Z(g29545) ) ;
NOR2    gate21738  (.A(g28948), .B(g28474), .Z(g29219) ) ;
AND2    gate21739  (.A(g29219), .B(g29382), .Z(g29547) ) ;
NOR2    gate21740  (.A(g28468), .B(g27970), .Z(g28784) ) ;
AND2    gate21741  (.A(g28784), .B(g29383), .Z(g29548) ) ;
NOR2    gate21742  (.A(g25506), .B(g24870), .Z(g26043) ) ;
AND2    gate21743  (.A(g26043), .B(g29384), .Z(g29549) ) ;
NOR2    gate21744  (.A(g28958), .B(g28479), .Z(g29222) ) ;
AND2    gate21745  (.A(g29222), .B(g29385), .Z(g29550) ) ;
NOR2    gate21746  (.A(g28962), .B(g28480), .Z(g29223) ) ;
AND2    gate21747  (.A(g29223), .B(g29386), .Z(g29553) ) ;
NOR2    gate21748  (.A(g28970), .B(g28481), .Z(g29224) ) ;
AND2    gate21749  (.A(g29224), .B(g29387), .Z(g29555) ) ;
NOR2    gate21750  (.A(g28477), .B(g27985), .Z(g28789) ) ;
AND2    gate21751  (.A(g28789), .B(g29388), .Z(g29557) ) ;
NOR2    gate21752  (.A(g28478), .B(g27991), .Z(g28790) ) ;
AND2    gate21753  (.A(g28790), .B(g29389), .Z(g29558) ) ;
NOR2    gate21754  (.A(g25553), .B(g24885), .Z(g26045) ) ;
AND2    gate21755  (.A(g26045), .B(g29390), .Z(g29559) ) ;
NOR2    gate21756  (.A(g28986), .B(g28486), .Z(g29227) ) ;
AND2    gate21757  (.A(g29227), .B(g29391), .Z(g29560) ) ;
NOR2    gate21758  (.A(g28996), .B(g28487), .Z(g29228) ) ;
AND2    gate21759  (.A(g29228), .B(g29392), .Z(g29562) ) ;
NOR2    gate21760  (.A(g28484), .B(g28009), .Z(g28794) ) ;
AND2    gate21761  (.A(g28794), .B(g29393), .Z(g29564) ) ;
NOR2    gate21762  (.A(g28485), .B(g28015), .Z(g28795) ) ;
AND2    gate21763  (.A(g28795), .B(g29394), .Z(g29565) ) ;
NOR2    gate21764  (.A(g25619), .B(g24902), .Z(g26047) ) ;
AND2    gate21765  (.A(g26047), .B(g29395), .Z(g29566) ) ;
NOR2    gate21766  (.A(g29022), .B(g28494), .Z(g29231) ) ;
AND2    gate21767  (.A(g29231), .B(g29396), .Z(g29567) ) ;
NOR2    gate21768  (.A(g28492), .B(g28036), .Z(g28802) ) ;
AND2    gate21769  (.A(g28802), .B(g29397), .Z(g29572) ) ;
NOR2    gate21770  (.A(g28493), .B(g28042), .Z(g28803) ) ;
AND2    gate21771  (.A(g28803), .B(g29398), .Z(g29573) ) ;
NOR2    gate21772  (.A(g28497), .B(g28066), .Z(g28813) ) ;
AND2    gate21773  (.A(g28813), .B(g29402), .Z(g29575) ) ;
AND2    gate21774  (.A(g29193), .B(g11056), .Z(g29607) ) ;
AND2    gate21775  (.A(g29349), .B(g11123), .Z(g29610) ) ;
AND2    gate21776  (.A(g29359), .B(g11182), .Z(g29614) ) ;
AND2    gate21777  (.A(g29245), .B(g11185), .Z(g29615) ) ;
AND2    gate21778  (.A(g29247), .B(g11259), .Z(g29619) ) ;
AND2    gate21779  (.A(g29250), .B(g11327), .Z(g29622) ) ;
AND2    gate21780  (.A(g29254), .B(g11407), .Z(g29624) ) ;
AND2    gate21781  (.A(g29189), .B(g11472), .Z(g29625) ) ;
AND2    gate21782  (.A(g29318), .B(g11478), .Z(g29626) ) ;
AND2    gate21783  (.A(g29491), .B(g10918), .Z(g29790) ) ;
AND2    gate21784  (.A(g29491), .B(g10977), .Z(g29792) ) ;
AND2    gate21785  (.A(g29491), .B(g11063), .Z(g29793) ) ;
NOR3    gate21786  (.A(g6104), .B(g29583), .C(g25363), .Z(g29748) ) ;
AND2    gate21787  (.A(g29748), .B(g22248), .Z(g29810) ) ;
NOR2    gate21788  (.A(g29583), .B(g1917), .Z(g29703) ) ;
AND2    gate21789  (.A(g29703), .B(g20644), .Z(g29811) ) ;
NOR2    gate21790  (.A(g16432), .B(g29625), .Z(g29762) ) ;
AND2    gate21791  (.A(g29762), .B(g12223), .Z(g29812) ) ;
NOR2    gate21792  (.A(g16411), .B(g29624), .Z(g29760) ) ;
AND2    gate21793  (.A(g29760), .B(g13869), .Z(g29813) ) ;
NOR3    gate21794  (.A(g6104), .B(g29583), .C(g25401), .Z(g29728) ) ;
AND2    gate21795  (.A(g29728), .B(g22266), .Z(g29814) ) ;
NOR2    gate21796  (.A(g29583), .B(g1912), .Z(g29727) ) ;
AND2    gate21797  (.A(g29727), .B(g20662), .Z(g29815) ) ;
NOR2    gate21798  (.A(g16379), .B(g29622), .Z(g29759) ) ;
AND2    gate21799  (.A(g29759), .B(g13883), .Z(g29816) ) ;
NOR2    gate21800  (.A(g29583), .B(g1909), .Z(g29709) ) ;
AND2    gate21801  (.A(g29709), .B(g20694), .Z(g29817) ) ;
NOR3    gate21802  (.A(g6104), .B(g29583), .C(g25387), .Z(g29732) ) ;
AND2    gate21803  (.A(g29732), .B(g22293), .Z(g29818) ) ;
NOR3    gate21804  (.A(g6104), .B(g29583), .C(g25352), .Z(g29751) ) ;
AND2    gate21805  (.A(g29751), .B(g22294), .Z(g29819) ) ;
NOR2    gate21806  (.A(g29583), .B(g1910), .Z(g29717) ) ;
AND2    gate21807  (.A(g29717), .B(g20743), .Z(g29820) ) ;
NOR2    gate21808  (.A(g29583), .B(g1913), .Z(g29731) ) ;
AND2    gate21809  (.A(g29731), .B(g20746), .Z(g29821) ) ;
NOR3    gate21810  (.A(g6104), .B(g29583), .C(g25339), .Z(g29705) ) ;
AND2    gate21811  (.A(g29705), .B(g22335), .Z(g29822) ) ;
NOR3    gate21812  (.A(g6104), .B(g29583), .C(g25376), .Z(g29741) ) ;
AND2    gate21813  (.A(g29741), .B(g22356), .Z(g29827) ) ;
NOR2    gate21814  (.A(g29583), .B(g1914), .Z(g29740) ) ;
AND2    gate21815  (.A(g29740), .B(g20802), .Z(g29828) ) ;
NOR2    gate21816  (.A(g29583), .B(g1911), .Z(g29725) ) ;
AND2    gate21817  (.A(g29725), .B(g20813), .Z(g29833) ) ;
NOR3    gate21818  (.A(g6104), .B(g29583), .C(g25332), .Z(g29713) ) ;
AND2    gate21819  (.A(g29713), .B(g22366), .Z(g29834) ) ;
NOR2    gate21820  (.A(g29583), .B(g1916), .Z(g29747) ) ;
AND2    gate21821  (.A(g29747), .B(g20827), .Z(g29839) ) ;
NOR2    gate21822  (.A(g23797), .B(g29583), .Z(g29735) ) ;
AND3    gate21823  (.A(g29735), .B(g19420), .C(g19401), .Z(g29909) ) ;
NOR2    gate21824  (.A(g13943), .B(g29502), .Z(g29779) ) ;
AND2    gate21825  (.A(g29779), .B(g9961), .Z(g29910) ) ;
NOR2    gate21826  (.A(g29472), .B(g29200), .Z(g29771) ) ;
AND2    gate21827  (.A(g29771), .B(g28877), .Z(g29942) ) ;
NOR2    gate21828  (.A(g29482), .B(g29234), .Z(g29782) ) ;
AND2    gate21829  (.A(g29782), .B(g28889), .Z(g29944) ) ;
NOR2    gate21830  (.A(g29474), .B(g29208), .Z(g29773) ) ;
AND2    gate21831  (.A(g29773), .B(g28894), .Z(g29945) ) ;
NOR2    gate21832  (.A(g29479), .B(g29229), .Z(g29778) ) ;
AND2    gate21833  (.A(g29778), .B(g28906), .Z(g29946) ) ;
NOR2    gate21834  (.A(g29485), .B(g29238), .Z(g29785) ) ;
AND2    gate21835  (.A(g29785), .B(g28911), .Z(g29947) ) ;
NOR2    gate21836  (.A(g29476), .B(g29217), .Z(g29775) ) ;
AND2    gate21837  (.A(g29775), .B(g28916), .Z(g29948) ) ;
NOR2    gate21838  (.A(g29481), .B(g29233), .Z(g29781) ) ;
AND2    gate21839  (.A(g29781), .B(g28932), .Z(g29949) ) ;
NOR2    gate21840  (.A(g29488), .B(g29241), .Z(g29788) ) ;
AND2    gate21841  (.A(g29788), .B(g28937), .Z(g29950) ) ;
NOR2    gate21842  (.A(g29478), .B(g29225), .Z(g29777) ) ;
AND2    gate21843  (.A(g29777), .B(g28945), .Z(g29951) ) ;
NOR2    gate21844  (.A(g29484), .B(g29236), .Z(g29784) ) ;
AND2    gate21845  (.A(g29784), .B(g28959), .Z(g29952) ) ;
NOR2    gate21846  (.A(g29490), .B(g29243), .Z(g29791) ) ;
AND2    gate21847  (.A(g29791), .B(g28967), .Z(g29953) ) ;
NOR2    gate21848  (.A(g29471), .B(g29196), .Z(g29770) ) ;
AND2    gate21849  (.A(g29770), .B(g28975), .Z(g29954) ) ;
NOR2    gate21850  (.A(g29487), .B(g29240), .Z(g29787) ) ;
AND2    gate21851  (.A(g29787), .B(g28993), .Z(g29955) ) ;
NOR2    gate21852  (.A(g29480), .B(g29232), .Z(g29780) ) ;
AND2    gate21853  (.A(g29780), .B(g28998), .Z(g29956) ) ;
NOR2    gate21854  (.A(g29473), .B(g29203), .Z(g29772) ) ;
AND2    gate21855  (.A(g29772), .B(g29005), .Z(g29957) ) ;
NOR2    gate21856  (.A(g29483), .B(g29235), .Z(g29783) ) ;
AND2    gate21857  (.A(g29783), .B(g29027), .Z(g29958) ) ;
NOR2    gate21858  (.A(g29475), .B(g29211), .Z(g29774) ) ;
AND2    gate21859  (.A(g29774), .B(g29035), .Z(g29959) ) ;
NOR2    gate21860  (.A(g29486), .B(g29239), .Z(g29786) ) ;
AND2    gate21861  (.A(g29786), .B(g29050), .Z(g29960) ) ;
NOR2    gate21862  (.A(g29477), .B(g29220), .Z(g29776) ) ;
AND2    gate21863  (.A(g29776), .B(g29057), .Z(g29961) ) ;
NOR2    gate21864  (.A(g29489), .B(g29242), .Z(g29789) ) ;
AND2    gate21865  (.A(g29789), .B(g29069), .Z(g29962) ) ;
NOR2    gate21866  (.A(g16335), .B(g29619), .Z(g29758) ) ;
AND2    gate21867  (.A(g29758), .B(g13737), .Z(g29963) ) ;
NOR2    gate21868  (.A(g16285), .B(g29615), .Z(g29757) ) ;
AND2    gate21869  (.A(g29757), .B(g13786), .Z(g29964) ) ;
NOR2    gate21870  (.A(g16284), .B(g29614), .Z(g29756) ) ;
AND2    gate21871  (.A(g29756), .B(g11961), .Z(g29965) ) ;
NOR2    gate21872  (.A(g16229), .B(g29610), .Z(g29755) ) ;
AND2    gate21873  (.A(g29755), .B(g12004), .Z(g29966) ) ;
NOR2    gate21874  (.A(g16178), .B(g29607), .Z(g29754) ) ;
AND2    gate21875  (.A(g29754), .B(g12066), .Z(g29967) ) ;
NOR2    gate21876  (.A(g13492), .B(g29465), .Z(g29765) ) ;
AND2    gate21877  (.A(g29765), .B(g12119), .Z(g29968) ) ;
NOR3    gate21878  (.A(g6104), .B(g29583), .C(g25323), .Z(g29721) ) ;
AND2    gate21879  (.A(g29721), .B(g22237), .Z(g29969) ) ;
NOR2    gate21880  (.A(g16462), .B(g29464), .Z(g29764) ) ;
AND2    gate21881  (.A(g29764), .B(g12178), .Z(g29970) ) ;
NOR2    gate21882  (.A(g16438), .B(g29626), .Z(g29763) ) ;
AND2    gate21883  (.A(g29763), .B(g13861), .Z(g29971) ) ;
AND2    gate21884  (.A(g29881), .B(g8324), .Z(g29980) ) ;
AND2    gate21885  (.A(g29869), .B(g8330), .Z(g29981) ) ;
AND2    gate21886  (.A(g29893), .B(g8336), .Z(g29982) ) ;
AND2    gate21887  (.A(g29885), .B(g8344), .Z(g29983) ) ;
AND2    gate21888  (.A(g29873), .B(g8351), .Z(g29984) ) ;
AND2    gate21889  (.A(g29897), .B(g8363), .Z(g29985) ) ;
AND2    gate21890  (.A(g29877), .B(g8366), .Z(g29986) ) ;
AND2    gate21891  (.A(g29889), .B(g8369), .Z(g29987) ) ;
AND2    gate21892  (.A(g29881), .B(g8382), .Z(g29988) ) ;
AND2    gate21893  (.A(g29893), .B(g8391), .Z(g29989) ) ;
AND2    gate21894  (.A(g29885), .B(g8397), .Z(g29990) ) ;
AND2    gate21895  (.A(g29901), .B(g8403), .Z(g29991) ) ;
NOR2    gate21896  (.A(g8594), .B(g10767), .Z(g12441) ) ;
AND2    gate21897  (.A(g12441), .B(g29909), .Z(g29992) ) ;
AND2    gate21898  (.A(g29897), .B(g8411), .Z(g29993) ) ;
AND2    gate21899  (.A(g29889), .B(g8418), .Z(g29994) ) ;
AND2    gate21900  (.A(g29893), .B(g8434), .Z(g29995) ) ;
AND2    gate21901  (.A(g29901), .B(g8443), .Z(g29996) ) ;
NOR2    gate21902  (.A(g29744), .B(g22367), .Z(g29918) ) ;
AND2    gate21903  (.A(g29918), .B(g22277), .Z(g29997) ) ;
NOR2    gate21904  (.A(g29744), .B(g22367), .Z(g29922) ) ;
AND2    gate21905  (.A(g29922), .B(g22278), .Z(g29998) ) ;
NOR2    gate21906  (.A(g29710), .B(g22367), .Z(g29924) ) ;
AND2    gate21907  (.A(g29924), .B(g22279), .Z(g29999) ) ;
NAND2   gate21908  (.A(II39385), .B(II39386), .Z(g29930) ) ;
AND2    gate21909  (.A(g10767), .B(g29930), .Z(g30000) ) ;
AND2    gate21910  (.A(g29897), .B(g8449), .Z(g30001) ) ;
AND2    gate21911  (.A(g29905), .B(g8455), .Z(g30002) ) ;
AND2    gate21912  (.A(g29901), .B(g8469), .Z(g30003) ) ;
NOR2    gate21913  (.A(g29718), .B(g22367), .Z(g29926) ) ;
AND2    gate21914  (.A(g29926), .B(g22295), .Z(g30004) ) ;
AND2    gate21915  (.A(g29905), .B(g8478), .Z(g30005) ) ;
NOR2    gate21916  (.A(g29673), .B(g22367), .Z(g29928) ) ;
AND2    gate21917  (.A(g29928), .B(g22310), .Z(g30006) ) ;
AND2    gate21918  (.A(g29905), .B(g8494), .Z(g30007) ) ;
NOR2    gate21919  (.A(g29736), .B(g22367), .Z(g29919) ) ;
AND2    gate21920  (.A(g29919), .B(g22334), .Z(g30008) ) ;
NOR2    gate21921  (.A(g29673), .B(g22367), .Z(g29929) ) ;
AND2    gate21922  (.A(g29929), .B(g22357), .Z(g30009) ) ;
AND2    gate21923  (.A(g29823), .B(g10963), .Z(g30077) ) ;
AND2    gate21924  (.A(g29823), .B(g10988), .Z(g30079) ) ;
AND2    gate21925  (.A(g29829), .B(g10996), .Z(g30080) ) ;
AND2    gate21926  (.A(g29823), .B(g11022), .Z(g30081) ) ;
AND2    gate21927  (.A(g29829), .B(g11036), .Z(g30082) ) ;
AND2    gate21928  (.A(g29835), .B(g11048), .Z(g30083) ) ;
AND2    gate21929  (.A(g29829), .B(g11092), .Z(g30085) ) ;
AND2    gate21930  (.A(g29835), .B(g11108), .Z(g30086) ) ;
AND2    gate21931  (.A(g29840), .B(g11120), .Z(g30087) ) ;
AND2    gate21932  (.A(g29844), .B(g11138), .Z(g30088) ) ;
AND2    gate21933  (.A(g29835), .B(g11160), .Z(g30089) ) ;
AND2    gate21934  (.A(g29840), .B(g11176), .Z(g30090) ) ;
AND2    gate21935  (.A(g29844), .B(g11202), .Z(g30091) ) ;
AND2    gate21936  (.A(g29849), .B(g11205), .Z(g30092) ) ;
AND2    gate21937  (.A(g29853), .B(g11222), .Z(g30093) ) ;
AND2    gate21938  (.A(g29840), .B(g11246), .Z(g30094) ) ;
AND2    gate21939  (.A(g29857), .B(g11265), .Z(g30095) ) ;
AND2    gate21940  (.A(g29844), .B(g11268), .Z(g30096) ) ;
AND2    gate21941  (.A(g29849), .B(g11271), .Z(g30097) ) ;
AND2    gate21942  (.A(g29853), .B(g11284), .Z(g30098) ) ;
AND2    gate21943  (.A(g29861), .B(g11287), .Z(g30099) ) ;
AND2    gate21944  (.A(g29865), .B(g11306), .Z(g30100) ) ;
AND2    gate21945  (.A(g29857), .B(g11341), .Z(g30101) ) ;
AND2    gate21946  (.A(g29849), .B(g11348), .Z(g30102) ) ;
AND2    gate21947  (.A(g29869), .B(g11358), .Z(g30103) ) ;
AND2    gate21948  (.A(g29853), .B(g11361), .Z(g30104) ) ;
AND2    gate21949  (.A(g29861), .B(g11364), .Z(g30105) ) ;
AND2    gate21950  (.A(g29865), .B(g11379), .Z(g30106) ) ;
AND2    gate21951  (.A(g29873), .B(g11382), .Z(g30107) ) ;
AND2    gate21952  (.A(g29877), .B(g11401), .Z(g30108) ) ;
AND2    gate21953  (.A(g29857), .B(g11411), .Z(g30109) ) ;
AND2    gate21954  (.A(g29881), .B(g11417), .Z(g30110) ) ;
AND2    gate21955  (.A(g29869), .B(g11425), .Z(g30111) ) ;
AND2    gate21956  (.A(g29861), .B(g11432), .Z(g30112) ) ;
AND2    gate21957  (.A(g29885), .B(g11444), .Z(g30113) ) ;
AND2    gate21958  (.A(g29865), .B(g11447), .Z(g30114) ) ;
AND2    gate21959  (.A(g29873), .B(g11450), .Z(g30115) ) ;
NOR2    gate21960  (.A(g29736), .B(g22367), .Z(g29921) ) ;
AND2    gate21961  (.A(g29921), .B(g22236), .Z(g30116) ) ;
AND2    gate21962  (.A(g29877), .B(g11465), .Z(g30117) ) ;
AND2    gate21963  (.A(g29889), .B(g11468), .Z(g30118) ) ;
NOR2    gate21964  (.A(g29827), .B(g29833), .Z(g30070) ) ;
AND2    gate21965  (.A(g30070), .B(g20641), .Z(g30123) ) ;
NOR2    gate21966  (.A(g29814), .B(g29817), .Z(g30065) ) ;
AND2    gate21967  (.A(g30065), .B(g20719), .Z(g30127) ) ;
NOR2    gate21968  (.A(g29810), .B(g29815), .Z(g30062) ) ;
AND2    gate21969  (.A(g30062), .B(g20722), .Z(g30128) ) ;
NOR2    gate21970  (.A(g29834), .B(g29839), .Z(g30071) ) ;
AND2    gate21971  (.A(g30071), .B(g20725), .Z(g30129) ) ;
NOR2    gate21972  (.A(g29969), .B(g29811), .Z(g30059) ) ;
AND2    gate21973  (.A(g30059), .B(g20749), .Z(g30131) ) ;
NOR2    gate21974  (.A(g29819), .B(g29821), .Z(g30068) ) ;
AND2    gate21975  (.A(g30068), .B(g20776), .Z(g30132) ) ;
NOR2    gate21976  (.A(g29818), .B(g29820), .Z(g30067) ) ;
AND2    gate21977  (.A(g30067), .B(g20799), .Z(g30133) ) ;
NOR2    gate21978  (.A(g29822), .B(g29828), .Z(g30069) ) ;
AND2    gate21979  (.A(g30069), .B(g20816), .Z(g30138) ) ;
AND2    gate21980  (.A(g30036), .B(g8921), .Z(g30216) ) ;
AND2    gate21981  (.A(g30036), .B(g8955), .Z(g30217) ) ;
AND2    gate21982  (.A(g30040), .B(g8961), .Z(g30218) ) ;
AND2    gate21983  (.A(g30036), .B(g8980), .Z(g30219) ) ;
AND2    gate21984  (.A(g30040), .B(g8987), .Z(g30220) ) ;
AND2    gate21985  (.A(g30044), .B(g8993), .Z(g30221) ) ;
AND2    gate21986  (.A(g30040), .B(g9010), .Z(g30222) ) ;
AND2    gate21987  (.A(g30044), .B(g9016), .Z(g30223) ) ;
AND2    gate21988  (.A(g30048), .B(g9022), .Z(g30224) ) ;
AND2    gate21989  (.A(g30044), .B(g9035), .Z(g30225) ) ;
AND2    gate21990  (.A(g30048), .B(g9041), .Z(g30226) ) ;
AND2    gate21991  (.A(g30048), .B(g9058), .Z(g30227) ) ;
AND2    gate21992  (.A(g30187), .B(g8321), .Z(g30327) ) ;
AND2    gate21993  (.A(g30195), .B(g8333), .Z(g30330) ) ;
AND2    gate21994  (.A(g30191), .B(g8341), .Z(g30333) ) ;
AND2    gate21995  (.A(g30203), .B(g8347), .Z(g30334) ) ;
AND2    gate21996  (.A(g30199), .B(g8354), .Z(g30337) ) ;
AND2    gate21997  (.A(g30207), .B(g8372), .Z(g30340) ) ;
AND2    gate21998  (.A(g30195), .B(g8388), .Z(g30345) ) ;
AND2    gate21999  (.A(g30203), .B(g8400), .Z(g30348) ) ;
AND2    gate22000  (.A(g30199), .B(g8408), .Z(g30351) ) ;
AND2    gate22001  (.A(g30211), .B(g8414), .Z(g30352) ) ;
AND2    gate22002  (.A(g30207), .B(g8421), .Z(g30355) ) ;
AND2    gate22003  (.A(g30203), .B(g8440), .Z(g30361) ) ;
AND2    gate22004  (.A(g30211), .B(g8452), .Z(g30364) ) ;
AND2    gate22005  (.A(g30207), .B(g8460), .Z(g30367) ) ;
NAND2   gate22006  (.A(II39690), .B(II39691), .Z(g30228) ) ;
AND2    gate22007  (.A(g8594), .B(g30228), .Z(g30372) ) ;
AND2    gate22008  (.A(g30211), .B(g8475), .Z(g30374) ) ;
AND2    gate22009  (.A(g30229), .B(g8888), .Z(g30387) ) ;
AND2    gate22010  (.A(g30229), .B(g8918), .Z(g30388) ) ;
AND2    gate22011  (.A(g30233), .B(g8928), .Z(g30389) ) ;
AND2    gate22012  (.A(g30229), .B(g8952), .Z(g30390) ) ;
AND2    gate22013  (.A(g30233), .B(g8958), .Z(g30391) ) ;
AND2    gate22014  (.A(g30237), .B(g8968), .Z(g30392) ) ;
AND2    gate22015  (.A(g30233), .B(g8984), .Z(g30393) ) ;
AND2    gate22016  (.A(g30237), .B(g8990), .Z(g30394) ) ;
AND2    gate22017  (.A(g30241), .B(g9000), .Z(g30395) ) ;
AND2    gate22018  (.A(g30237), .B(g9013), .Z(g30396) ) ;
AND2    gate22019  (.A(g30241), .B(g9019), .Z(g30397) ) ;
AND2    gate22020  (.A(g30241), .B(g9038), .Z(g30398) ) ;
AND2    gate22021  (.A(g30134), .B(g10991), .Z(g30407) ) ;
AND2    gate22022  (.A(g30134), .B(g11025), .Z(g30409) ) ;
AND2    gate22023  (.A(g30139), .B(g11028), .Z(g30410) ) ;
AND2    gate22024  (.A(g30143), .B(g11039), .Z(g30411) ) ;
AND2    gate22025  (.A(g30134), .B(g11079), .Z(g30436) ) ;
AND2    gate22026  (.A(g30139), .B(g11082), .Z(g30437) ) ;
AND2    gate22027  (.A(g30147), .B(g11085), .Z(g30438) ) ;
AND2    gate22028  (.A(g30143), .B(g11095), .Z(g30440) ) ;
AND2    gate22029  (.A(g30151), .B(g11098), .Z(g30441) ) ;
AND2    gate22030  (.A(g30155), .B(g11111), .Z(g30442) ) ;
AND2    gate22031  (.A(g30139), .B(g11132), .Z(g30444) ) ;
AND2    gate22032  (.A(g30147), .B(g11135), .Z(g30445) ) ;
AND2    gate22033  (.A(g30143), .B(g11145), .Z(g30447) ) ;
AND2    gate22034  (.A(g30151), .B(g11148), .Z(g30448) ) ;
AND2    gate22035  (.A(g30159), .B(g11151), .Z(g30449) ) ;
AND2    gate22036  (.A(g30155), .B(g11163), .Z(g30451) ) ;
AND2    gate22037  (.A(g30163), .B(g11166), .Z(g30452) ) ;
AND2    gate22038  (.A(g30167), .B(g11179), .Z(g30453) ) ;
AND2    gate22039  (.A(g30147), .B(g11199), .Z(g30454) ) ;
AND2    gate22040  (.A(g30151), .B(g11216), .Z(g30457) ) ;
AND2    gate22041  (.A(g30159), .B(g11219), .Z(g30458) ) ;
AND2    gate22042  (.A(g30155), .B(g11231), .Z(g30460) ) ;
AND2    gate22043  (.A(g30163), .B(g11234), .Z(g30461) ) ;
AND2    gate22044  (.A(g30171), .B(g11237), .Z(g30462) ) ;
AND2    gate22045  (.A(g30167), .B(g11249), .Z(g30464) ) ;
AND2    gate22046  (.A(g30175), .B(g11252), .Z(g30465) ) ;
AND2    gate22047  (.A(g30179), .B(g11274), .Z(g30467) ) ;
AND2    gate22048  (.A(g30159), .B(g11281), .Z(g30469) ) ;
AND2    gate22049  (.A(g30163), .B(g11300), .Z(g30472) ) ;
AND2    gate22050  (.A(g30171), .B(g11303), .Z(g30473) ) ;
AND2    gate22051  (.A(g30167), .B(g11315), .Z(g30475) ) ;
AND2    gate22052  (.A(g30175), .B(g11318), .Z(g30476) ) ;
AND2    gate22053  (.A(g30183), .B(g11321), .Z(g30477) ) ;
AND2    gate22054  (.A(g30187), .B(g11344), .Z(g30478) ) ;
AND2    gate22055  (.A(g30179), .B(g11351), .Z(g30481) ) ;
AND2    gate22056  (.A(g30191), .B(g11367), .Z(g30484) ) ;
AND2    gate22057  (.A(g30171), .B(g11376), .Z(g30486) ) ;
AND2    gate22058  (.A(g30175), .B(g11395), .Z(g30489) ) ;
AND2    gate22059  (.A(g30183), .B(g11398), .Z(g30490) ) ;
AND2    gate22060  (.A(g30187), .B(g11414), .Z(g30492) ) ;
AND2    gate22061  (.A(g30179), .B(g11422), .Z(g30495) ) ;
AND2    gate22062  (.A(g30195), .B(g11428), .Z(g30496) ) ;
AND2    gate22063  (.A(g30191), .B(g11435), .Z(g30499) ) ;
AND2    gate22064  (.A(g30199), .B(g11453), .Z(g30502) ) ;
AND2    gate22065  (.A(g30183), .B(g11462), .Z(g30504) ) ;
AND2    gate22066  (.A(g30383), .B(g10943), .Z(g30696) ) ;
AND2    gate22067  (.A(g30383), .B(g11011), .Z(g30697) ) ;
AND2    gate22068  (.A(g30383), .B(g11126), .Z(g30698) ) ;
NOR3    gate22069  (.A(g6119), .B(g30412), .C(g25333), .Z(g30605) ) ;
AND2    gate22070  (.A(g30605), .B(g22252), .Z(g30728) ) ;
NOR3    gate22071  (.A(g6119), .B(g30412), .C(g25378), .Z(g30629) ) ;
AND2    gate22072  (.A(g30629), .B(g22268), .Z(g30735) ) ;
NOR2    gate22073  (.A(g30412), .B(g2611), .Z(g30584) ) ;
AND2    gate22074  (.A(g30584), .B(g20669), .Z(g30736) ) ;
NOR3    gate22075  (.A(g6119), .B(g30412), .C(g25411), .Z(g30610) ) ;
AND2    gate22076  (.A(g30610), .B(g22283), .Z(g30743) ) ;
NOR2    gate22077  (.A(g30412), .B(g2606), .Z(g30609) ) ;
AND2    gate22078  (.A(g30609), .B(g20697), .Z(g30744) ) ;
NOR2    gate22079  (.A(g30412), .B(g2603), .Z(g30593) ) ;
AND2    gate22080  (.A(g30593), .B(g20729), .Z(g30750) ) ;
NOR3    gate22081  (.A(g6119), .B(g30412), .C(g25403), .Z(g30614) ) ;
AND2    gate22082  (.A(g30614), .B(g22313), .Z(g30754) ) ;
NOR3    gate22083  (.A(g6119), .B(g30412), .C(g25366), .Z(g30632) ) ;
AND2    gate22084  (.A(g30632), .B(g22314), .Z(g30755) ) ;
NOR2    gate22085  (.A(g30412), .B(g2604), .Z(g30601) ) ;
AND2    gate22086  (.A(g30601), .B(g20780), .Z(g30757) ) ;
NOR2    gate22087  (.A(g30412), .B(g2607), .Z(g30613) ) ;
AND2    gate22088  (.A(g30613), .B(g20783), .Z(g30758) ) ;
NOR3    gate22089  (.A(g6119), .B(g30412), .C(g25353), .Z(g30588) ) ;
AND2    gate22090  (.A(g30588), .B(g22360), .Z(g30759) ) ;
NOR3    gate22091  (.A(g6119), .B(g30412), .C(g25393), .Z(g30622) ) ;
AND2    gate22092  (.A(g30622), .B(g22379), .Z(g30760) ) ;
NOR2    gate22093  (.A(g30412), .B(g2608), .Z(g30621) ) ;
AND2    gate22094  (.A(g30621), .B(g20822), .Z(g30761) ) ;
NOR2    gate22095  (.A(g30412), .B(g2605), .Z(g30608) ) ;
AND2    gate22096  (.A(g30608), .B(g20830), .Z(g30762) ) ;
NOR3    gate22097  (.A(g6119), .B(g30412), .C(g25341), .Z(g30597) ) ;
AND2    gate22098  (.A(g30597), .B(g22386), .Z(g30763) ) ;
NOR2    gate22099  (.A(g30412), .B(g2610), .Z(g30628) ) ;
AND2    gate22100  (.A(g30628), .B(g20837), .Z(g30764) ) ;
NOR2    gate22101  (.A(g23850), .B(g30412), .Z(g30617) ) ;
AND3    gate22102  (.A(g30617), .B(g19457), .C(g19431), .Z(g30766) ) ;
NOR2    gate22103  (.A(g30618), .B(g22387), .Z(g30785) ) ;
AND2    gate22104  (.A(g30785), .B(g22251), .Z(g30916) ) ;
NOR2    gate22105  (.A(g8605), .B(g10773), .Z(g12446) ) ;
AND2    gate22106  (.A(g12446), .B(g30766), .Z(g30917) ) ;
NOR2    gate22107  (.A(g30625), .B(g22387), .Z(g30780) ) ;
AND2    gate22108  (.A(g30780), .B(g22296), .Z(g30918) ) ;
NOR2    gate22109  (.A(g30625), .B(g22387), .Z(g30786) ) ;
AND2    gate22110  (.A(g30786), .B(g22297), .Z(g30919) ) ;
NOR2    gate22111  (.A(g30594), .B(g22387), .Z(g30787) ) ;
AND2    gate22112  (.A(g30787), .B(g22298), .Z(g30920) ) ;
NAND2   gate22113  (.A(II40628), .B(II40629), .Z(g30791) ) ;
AND2    gate22114  (.A(g10773), .B(g30791), .Z(g30921) ) ;
NOR2    gate22115  (.A(g30602), .B(g22387), .Z(g30788) ) ;
AND2    gate22116  (.A(g30788), .B(g22315), .Z(g30922) ) ;
NOR2    gate22117  (.A(g30575), .B(g22387), .Z(g30789) ) ;
AND2    gate22118  (.A(g30789), .B(g22338), .Z(g30923) ) ;
NOR2    gate22119  (.A(g30618), .B(g22387), .Z(g30783) ) ;
AND2    gate22120  (.A(g30783), .B(g22359), .Z(g30924) ) ;
NOR2    gate22121  (.A(g30575), .B(g22387), .Z(g30790) ) ;
AND2    gate22122  (.A(g30790), .B(g22380), .Z(g30925) ) ;
NOR2    gate22123  (.A(g30760), .B(g30762), .Z(g30935) ) ;
AND2    gate22124  (.A(g30935), .B(g20666), .Z(g30944) ) ;
NOR2    gate22125  (.A(g30743), .B(g30750), .Z(g30931) ) ;
AND2    gate22126  (.A(g30931), .B(g20754), .Z(g30945) ) ;
NOR2    gate22127  (.A(g30735), .B(g30744), .Z(g30930) ) ;
AND2    gate22128  (.A(g30930), .B(g20757), .Z(g30946) ) ;
NOR2    gate22129  (.A(g30763), .B(g30764), .Z(g30936) ) ;
AND2    gate22130  (.A(g30936), .B(g20760), .Z(g30947) ) ;
NOR2    gate22131  (.A(g30728), .B(g30736), .Z(g30929) ) ;
AND2    gate22132  (.A(g30929), .B(g20786), .Z(g30948) ) ;
NOR2    gate22133  (.A(g30755), .B(g30758), .Z(g30933) ) ;
AND2    gate22134  (.A(g30933), .B(g20806), .Z(g30949) ) ;
NOR2    gate22135  (.A(g30754), .B(g30757), .Z(g30932) ) ;
AND2    gate22136  (.A(g30932), .B(g20819), .Z(g30950) ) ;
NOR2    gate22137  (.A(g30759), .B(g30761), .Z(g30934) ) ;
AND2    gate22138  (.A(g30934), .B(g20833), .Z(g30951) ) ;
NAND2   gate22139  (.A(II41065), .B(II41066), .Z(g30952) ) ;
AND2    gate22140  (.A(g8605), .B(g30952), .Z(g30953) ) ;
OR2     gate22141  (.A(g2986), .B(g5389), .Z(g9144) ) ;
OR2     gate22142  (.A(g2929), .B(g8022), .Z(g10778) ) ;
OR2     gate22143  (.A(g7553), .B(g11059), .Z(g12377) ) ;
OR2     gate22144  (.A(g7573), .B(g10779), .Z(g12407) ) ;
OR2     gate22145  (.A(g9534), .B(g3398), .Z(g12886) ) ;
OR2     gate22146  (.A(g9676), .B(g3554), .Z(g12926) ) ;
OR2     gate22147  (.A(g9822), .B(g3710), .Z(g12955) ) ;
OR2     gate22148  (.A(g9968), .B(g3866), .Z(g12984) ) ;
OR2     gate22149  (.A(g15880), .B(g14657), .Z(g16539) ) ;
OR2     gate22150  (.A(g15913), .B(g14691), .Z(g16571) ) ;
OR2     gate22151  (.A(g15942), .B(g14725), .Z(g16595) ) ;
OR2     gate22152  (.A(g15971), .B(g14753), .Z(g16615) ) ;
NAND2   gate22153  (.A(II23807), .B(II23808), .Z(g17729) ) ;
NAND2   gate22154  (.A(II24016), .B(II24017), .Z(g17979) ) ;
OR2     gate22155  (.A(g17729), .B(g17979), .Z(g19181) ) ;
NAND2   gate22156  (.A(II24437), .B(II24438), .Z(g18419) ) ;
NAND2   gate22157  (.A(II23942), .B(II23943), .Z(g17887) ) ;
OR2     gate22158  (.A(g18419), .B(g17887), .Z(g19186) ) ;
OR2     gate22159  (.A(g18419), .B(g17729), .Z(g19187) ) ;
NAND2   gate22160  (.A(II23894), .B(II23895), .Z(g17830) ) ;
NAND2   gate22161  (.A(II24111), .B(II24112), .Z(g18096) ) ;
OR2     gate22162  (.A(g17830), .B(g18096), .Z(g19188) ) ;
NAND2   gate22163  (.A(II23879), .B(II23880), .Z(g17807) ) ;
OR2     gate22164  (.A(g17807), .B(g17887), .Z(g19191) ) ;
NAND2   gate22165  (.A(II24179), .B(II24180), .Z(g18183) ) ;
NAND2   gate22166  (.A(II24264), .B(II24265), .Z(g18270) ) ;
OR2     gate22167  (.A(g18183), .B(g18270), .Z(g19192) ) ;
NAND2   gate22168  (.A(II24538), .B(II24539), .Z(g18492) ) ;
NAND2   gate22169  (.A(II24037), .B(II24038), .Z(g17998) ) ;
OR2     gate22170  (.A(g18492), .B(g17998), .Z(g19193) ) ;
OR2     gate22171  (.A(g18492), .B(g17830), .Z(g19194) ) ;
NAND2   gate22172  (.A(II23982), .B(II23983), .Z(g17942) ) ;
NAND2   gate22173  (.A(II24214), .B(II24215), .Z(g18212) ) ;
OR2     gate22174  (.A(g17942), .B(g18212), .Z(g19195) ) ;
NAND2   gate22175  (.A(II24352), .B(II24353), .Z(g18346) ) ;
NAND2   gate22176  (.A(II24444), .B(II24445), .Z(g18424) ) ;
OR2     gate22177  (.A(g18346), .B(g18424), .Z(g19200) ) ;
OR2     gate22178  (.A(g18183), .B(g18424), .Z(g19201) ) ;
NAND2   gate22179  (.A(II23967), .B(II23968), .Z(g17919) ) ;
OR2     gate22180  (.A(g17919), .B(g17998), .Z(g19202) ) ;
NAND2   gate22181  (.A(II24291), .B(II24292), .Z(g18290) ) ;
NAND2   gate22182  (.A(II24373), .B(II24374), .Z(g18363) ) ;
OR2     gate22183  (.A(g18290), .B(g18363), .Z(g19203) ) ;
NAND2   gate22184  (.A(II24640), .B(II24641), .Z(g18556) ) ;
NAND2   gate22185  (.A(II24132), .B(II24133), .Z(g18115) ) ;
OR2     gate22186  (.A(g18556), .B(g18115), .Z(g19204) ) ;
OR2     gate22187  (.A(g18556), .B(g17942), .Z(g19205) ) ;
NAND2   gate22188  (.A(II24077), .B(II24078), .Z(g18053) ) ;
NAND2   gate22189  (.A(II24326), .B(II24327), .Z(g18319) ) ;
OR2     gate22190  (.A(g18053), .B(g18319), .Z(g19206) ) ;
NAND2   gate22191  (.A(II24092), .B(II24093), .Z(g18079) ) ;
OR2     gate22192  (.A(g18079), .B(g18346), .Z(g19209) ) ;
OR2     gate22193  (.A(g18079), .B(g18183), .Z(g19210) ) ;
NAND2   gate22194  (.A(II24465), .B(II24466), .Z(g18441) ) ;
NAND2   gate22195  (.A(II24545), .B(II24546), .Z(g18497) ) ;
OR2     gate22196  (.A(g18441), .B(g18497), .Z(g19211) ) ;
OR2     gate22197  (.A(g18290), .B(g18497), .Z(g19212) ) ;
NAND2   gate22198  (.A(II24062), .B(II24063), .Z(g18030) ) ;
OR2     gate22199  (.A(g18030), .B(g18115), .Z(g19213) ) ;
NAND2   gate22200  (.A(II24400), .B(II24401), .Z(g18383) ) ;
NAND2   gate22201  (.A(II24486), .B(II24487), .Z(g18458) ) ;
OR2     gate22202  (.A(g18383), .B(g18458), .Z(g19214) ) ;
NAND2   gate22203  (.A(II24710), .B(II24711), .Z(g18606) ) ;
NAND2   gate22204  (.A(II24235), .B(II24236), .Z(g18231) ) ;
OR2     gate22205  (.A(g18606), .B(g18231), .Z(g19215) ) ;
OR2     gate22206  (.A(g18606), .B(g18053), .Z(g19216) ) ;
OR2     gate22207  (.A(g18270), .B(g18346), .Z(g19221) ) ;
NAND2   gate22208  (.A(II24195), .B(II24196), .Z(g18195) ) ;
OR2     gate22209  (.A(g18195), .B(g18441), .Z(g19222) ) ;
OR2     gate22210  (.A(g18195), .B(g18290), .Z(g19223) ) ;
NAND2   gate22211  (.A(II24566), .B(II24567), .Z(g18514) ) ;
NAND2   gate22212  (.A(II24647), .B(II24648), .Z(g18561) ) ;
OR2     gate22213  (.A(g18514), .B(g18561), .Z(g19224) ) ;
OR2     gate22214  (.A(g18383), .B(g18561), .Z(g19225) ) ;
NAND2   gate22215  (.A(II24157), .B(II24158), .Z(g18147) ) ;
OR2     gate22216  (.A(g18147), .B(g18231), .Z(g19226) ) ;
NAND2   gate22217  (.A(II24513), .B(II24514), .Z(g18478) ) ;
NAND2   gate22218  (.A(II24587), .B(II24588), .Z(g18531) ) ;
OR2     gate22219  (.A(g18478), .B(g18531), .Z(g19227) ) ;
NAND2   gate22220  (.A(II22999), .B(II23000), .Z(g17024) ) ;
NAND2   gate22221  (.A(II22963), .B(II22964), .Z(g17000) ) ;
NAND2   gate22222  (.A(II22937), .B(II22938), .Z(g16992) ) ;
OR3     gate22223  (.A(g17024), .B(g17000), .C(g16992), .Z(II25477) ) ;
NAND2   gate22224  (.A(II22918), .B(II22919), .Z(g16985) ) ;
NAND2   gate22225  (.A(II22901), .B(II22902), .Z(g16965) ) ;
OR3     gate22226  (.A(g16985), .B(g16965), .C(II25477), .Z(g19230) ) ;
OR2     gate22227  (.A(g18363), .B(g18441), .Z(g19231) ) ;
NAND2   gate22228  (.A(II24307), .B(II24308), .Z(g18302) ) ;
OR2     gate22229  (.A(g18302), .B(g18514), .Z(g19232) ) ;
OR2     gate22230  (.A(g18302), .B(g18383), .Z(g19233) ) ;
NAND2   gate22231  (.A(II24668), .B(II24669), .Z(g18578) ) ;
NAND2   gate22232  (.A(II24717), .B(II24718), .Z(g18611) ) ;
OR2     gate22233  (.A(g18578), .B(g18611), .Z(g19234) ) ;
OR2     gate22234  (.A(g18478), .B(g18611), .Z(g19235) ) ;
NAND2   gate22235  (.A(II23191), .B(II23192), .Z(g17158) ) ;
NAND2   gate22236  (.A(II23153), .B(II23154), .Z(g17137) ) ;
NAND2   gate22237  (.A(II23114), .B(II23115), .Z(g17115) ) ;
OR3     gate22238  (.A(g17158), .B(g17137), .C(g17115), .Z(II25495) ) ;
NAND2   gate22239  (.A(II23075), .B(II23076), .Z(g17083) ) ;
NAND2   gate22240  (.A(II23035), .B(II23036), .Z(g17050) ) ;
OR3     gate22241  (.A(g17083), .B(g17050), .C(II25495), .Z(g19240) ) ;
OR2     gate22242  (.A(g14244), .B(g16501), .Z(g19242) ) ;
NAND2   gate22243  (.A(II23046), .B(II23047), .Z(g17058) ) ;
NAND2   gate22244  (.A(II23009), .B(II23010), .Z(g17030) ) ;
NAND2   gate22245  (.A(II22973), .B(II22974), .Z(g17016) ) ;
OR3     gate22246  (.A(g17058), .B(g17030), .C(g17016), .Z(II25500) ) ;
NAND2   gate22247  (.A(II22946), .B(II22947), .Z(g16995) ) ;
NAND2   gate22248  (.A(II22925), .B(II22926), .Z(g16986) ) ;
OR3     gate22249  (.A(g16995), .B(g16986), .C(II25500), .Z(g19243) ) ;
OR2     gate22250  (.A(g18458), .B(g18514), .Z(g19244) ) ;
NAND2   gate22251  (.A(II24416), .B(II24417), .Z(g18395) ) ;
OR2     gate22252  (.A(g18395), .B(g18578), .Z(g19245) ) ;
OR2     gate22253  (.A(g18395), .B(g18478), .Z(g19246) ) ;
OR2     gate22254  (.A(g17729), .B(g17807), .Z(g19250) ) ;
NAND2   gate22255  (.A(II23226), .B(II23227), .Z(g17173) ) ;
NAND2   gate22256  (.A(II23199), .B(II23200), .Z(g17160) ) ;
NAND2   gate22257  (.A(II23162), .B(II23163), .Z(g17142) ) ;
OR3     gate22258  (.A(g17173), .B(g17160), .C(g17142), .Z(II25516) ) ;
NAND2   gate22259  (.A(II23124), .B(II23125), .Z(g17121) ) ;
NAND2   gate22260  (.A(II23083), .B(II23084), .Z(g17085) ) ;
OR3     gate22261  (.A(g17121), .B(g17085), .C(II25516), .Z(g19253) ) ;
OR2     gate22262  (.A(g14366), .B(g16523), .Z(g19255) ) ;
NAND2   gate22263  (.A(II23094), .B(II23095), .Z(g17093) ) ;
NAND2   gate22264  (.A(II23056), .B(II23057), .Z(g17064) ) ;
NAND2   gate22265  (.A(II23019), .B(II23020), .Z(g17046) ) ;
OR3     gate22266  (.A(g17093), .B(g17064), .C(g17046), .Z(II25521) ) ;
NAND2   gate22267  (.A(II22982), .B(II22983), .Z(g17019) ) ;
NAND2   gate22268  (.A(II22953), .B(II22954), .Z(g16996) ) ;
OR3     gate22269  (.A(g17019), .B(g16996), .C(II25521), .Z(g19256) ) ;
OR2     gate22270  (.A(g18531), .B(g18578), .Z(g19257) ) ;
OR2     gate22271  (.A(g17887), .B(g17979), .Z(g19263) ) ;
OR2     gate22272  (.A(g17830), .B(g17919), .Z(g19264) ) ;
NAND2   gate22273  (.A(II23257), .B(II23258), .Z(g17190) ) ;
NAND2   gate22274  (.A(II23234), .B(II23235), .Z(g17175) ) ;
NAND2   gate22275  (.A(II23208), .B(II23209), .Z(g17165) ) ;
OR3     gate22276  (.A(g17190), .B(g17175), .C(g17165), .Z(II25549) ) ;
NAND2   gate22277  (.A(II23172), .B(II23173), .Z(g17148) ) ;
NAND2   gate22278  (.A(II23132), .B(II23133), .Z(g17123) ) ;
OR3     gate22279  (.A(g17148), .B(g17123), .C(II25549), .Z(g19266) ) ;
OR2     gate22280  (.A(g14478), .B(g16554), .Z(g19268) ) ;
NAND2   gate22281  (.A(II23143), .B(II23144), .Z(g17131) ) ;
NAND2   gate22282  (.A(II23104), .B(II23105), .Z(g17099) ) ;
NAND2   gate22283  (.A(II23066), .B(II23067), .Z(g17080) ) ;
OR3     gate22284  (.A(g17131), .B(g17099), .C(g17080), .Z(II25554) ) ;
NAND2   gate22285  (.A(II23028), .B(II23029), .Z(g17049) ) ;
NAND2   gate22286  (.A(II22989), .B(II22990), .Z(g17020) ) ;
OR3     gate22287  (.A(g17049), .B(g17020), .C(II25554), .Z(g19269) ) ;
OR3     gate22288  (.A(g16867), .B(g16515), .C(g19001), .Z(g19275) ) ;
OR2     gate22289  (.A(g17998), .B(g18096), .Z(g19278) ) ;
OR2     gate22290  (.A(g17942), .B(g18030), .Z(g19279) ) ;
NAND2   gate22291  (.A(II23278), .B(II23279), .Z(g17201) ) ;
NAND2   gate22292  (.A(II23265), .B(II23266), .Z(g17192) ) ;
NAND2   gate22293  (.A(II23243), .B(II23244), .Z(g17180) ) ;
OR3     gate22294  (.A(g17201), .B(g17192), .C(g17180), .Z(II25588) ) ;
NAND2   gate22295  (.A(II23218), .B(II23219), .Z(g17171) ) ;
NAND2   gate22296  (.A(II23180), .B(II23181), .Z(g17150) ) ;
OR3     gate22297  (.A(g17171), .B(g17150), .C(II25588), .Z(g19281) ) ;
OR2     gate22298  (.A(g14565), .B(g16586), .Z(g19283) ) ;
OR3     gate22299  (.A(g16895), .B(g16546), .C(g16507), .Z(g19294) ) ;
OR2     gate22300  (.A(g18115), .B(g18212), .Z(g19297) ) ;
OR2     gate22301  (.A(g18053), .B(g18147), .Z(g19298) ) ;
OR3     gate22302  (.A(g16924), .B(g16578), .C(g16529), .Z(g19312) ) ;
OR2     gate22303  (.A(g18231), .B(g18319), .Z(g19315) ) ;
OR3     gate22304  (.A(g16954), .B(g16602), .C(g16560), .Z(g19333) ) ;
OR2     gate22305  (.A(g14837), .B(g16682), .Z(g19450) ) ;
OR2     gate22306  (.A(g14910), .B(g16708), .Z(g19477) ) ;
OR2     gate22307  (.A(g14991), .B(g16739), .Z(g19500) ) ;
OR3     gate22308  (.A(g16884), .B(g16697), .C(g16665), .Z(g19503) ) ;
OR2     gate22309  (.A(g15080), .B(g16781), .Z(g19521) ) ;
OR3     gate22310  (.A(g16913), .B(g16728), .C(g16686), .Z(g19522) ) ;
OR3     gate22311  (.A(g16943), .B(g16770), .C(g16712), .Z(g19532) ) ;
OR3     gate22312  (.A(g16974), .B(g16797), .C(g16743), .Z(g19542) ) ;
OR3     gate22313  (.A(g17979), .B(g17887), .C(g17807), .Z(II26429) ) ;
OR3     gate22314  (.A(g17729), .B(g18419), .C(II26429), .Z(g19981) ) ;
OR3     gate22315  (.A(g18424), .B(g18346), .C(g18270), .Z(II26455) ) ;
OR3     gate22316  (.A(g18183), .B(g18079), .C(II26455), .Z(g20015) ) ;
OR3     gate22317  (.A(g18096), .B(g17998), .C(g17919), .Z(II26461) ) ;
OR3     gate22318  (.A(g17830), .B(g18492), .C(II26461), .Z(g20019) ) ;
OR3     gate22319  (.A(g18497), .B(g18441), .C(g18363), .Z(II26491) ) ;
OR3     gate22320  (.A(g18290), .B(g18195), .C(II26491), .Z(g20057) ) ;
OR3     gate22321  (.A(g18212), .B(g18115), .C(g18030), .Z(II26497) ) ;
OR3     gate22322  (.A(g17942), .B(g18556), .C(II26497), .Z(g20061) ) ;
OR3     gate22323  (.A(g18561), .B(g18514), .C(g18458), .Z(II26532) ) ;
OR3     gate22324  (.A(g18383), .B(g18302), .C(II26532), .Z(g20098) ) ;
OR3     gate22325  (.A(g18319), .B(g18231), .C(g18147), .Z(II26538) ) ;
OR3     gate22326  (.A(g18053), .B(g18606), .C(II26538), .Z(g20102) ) ;
OR3     gate22327  (.A(g18611), .B(g18578), .C(g18531), .Z(II26571) ) ;
OR3     gate22328  (.A(g18478), .B(g18395), .C(II26571), .Z(g20123) ) ;
OR3     gate22329  (.A(g19484), .B(g16515), .C(g14071), .Z(g21120) ) ;
OR3     gate22330  (.A(g19505), .B(g16546), .C(g14186), .Z(g21139) ) ;
OR3     gate22331  (.A(g19524), .B(g16578), .C(g14301), .Z(g21159) ) ;
OR3     gate22332  (.A(g19534), .B(g16602), .C(g14423), .Z(g21179) ) ;
OR3     gate22333  (.A(g19578), .B(g16697), .C(g14776), .Z(g21244) ) ;
OR3     gate22334  (.A(g19608), .B(g16728), .C(g14811), .Z(g21253) ) ;
OR3     gate22335  (.A(g19641), .B(g16770), .C(g14863), .Z(g21261) ) ;
OR3     gate22336  (.A(g19681), .B(g16797), .C(g14936), .Z(g21269) ) ;
NAND2   gate22337  (.A(g16501), .B(g16515), .Z(g20522) ) ;
OR3     gate22338  (.A(g20522), .B(g16867), .C(g14071), .Z(g21501) ) ;
OR3     gate22339  (.A(g20522), .B(g19484), .C(g19001), .Z(g21536) ) ;
NAND2   gate22340  (.A(g16523), .B(g16546), .Z(g20542) ) ;
OR3     gate22341  (.A(g20542), .B(g16895), .C(g14186), .Z(g21540) ) ;
OR3     gate22342  (.A(g20542), .B(g19505), .C(g16507), .Z(g21572) ) ;
NAND2   gate22343  (.A(g16554), .B(g16578), .Z(g19067) ) ;
OR3     gate22344  (.A(g19067), .B(g16924), .C(g14301), .Z(g21576) ) ;
OR3     gate22345  (.A(g19067), .B(g19524), .C(g16529), .Z(g21605) ) ;
NAND2   gate22346  (.A(g16586), .B(g16602), .Z(g19084) ) ;
OR3     gate22347  (.A(g19084), .B(g16954), .C(g14423), .Z(g21609) ) ;
OR3     gate22348  (.A(g19084), .B(g19534), .C(g16560), .Z(g21634) ) ;
NAND2   gate22349  (.A(g16682), .B(g16697), .Z(g19121) ) ;
OR3     gate22350  (.A(g19121), .B(g16884), .C(g14776), .Z(g21774) ) ;
OR3     gate22351  (.A(g19121), .B(g19578), .C(g16665), .Z(g21787) ) ;
OR3     gate22352  (.A(g20197), .B(g20177), .C(g20145), .Z(II28305) ) ;
OR3     gate22353  (.A(g20117), .B(g20094), .C(II28305), .Z(g21788) ) ;
NAND2   gate22354  (.A(g16708), .B(g16728), .Z(g19128) ) ;
OR3     gate22355  (.A(g19128), .B(g16913), .C(g14811), .Z(g21789) ) ;
OR3     gate22356  (.A(g19092), .B(g19088), .C(g19079), .Z(II28318) ) ;
OR4     gate22357  (.A(g16505), .B(g20538), .C(g18994), .D(II28318), .Z(g21799) ) ;
OR4     gate22358  (.A(g18665), .B(g20270), .C(g20248), .D(g18647), .Z(g21800) ) ;
OR3     gate22359  (.A(g19128), .B(g19608), .C(g16686), .Z(g21801) ) ;
OR3     gate22360  (.A(g20227), .B(g20211), .C(g20183), .Z(II28323) ) ;
OR3     gate22361  (.A(g20147), .B(g20119), .C(II28323), .Z(g21802) ) ;
NAND2   gate22362  (.A(g16739), .B(g16770), .Z(g19135) ) ;
OR3     gate22363  (.A(g19135), .B(g16943), .C(g14863), .Z(g21803) ) ;
OR4     gate22364  (.A(g20116), .B(g20093), .C(g18547), .D(g19097), .Z(g21806) ) ;
OR3     gate22365  (.A(g19099), .B(g19094), .C(g19089), .Z(II28330) ) ;
OR4     gate22366  (.A(g16527), .B(g19063), .C(g19007), .D(II28330), .Z(g21807) ) ;
OR4     gate22367  (.A(g18688), .B(g20282), .C(g20271), .D(g18650), .Z(g21808) ) ;
OR3     gate22368  (.A(g19135), .B(g19641), .C(g16712), .Z(g21809) ) ;
OR3     gate22369  (.A(g20254), .B(g20241), .C(g20217), .Z(II28335) ) ;
OR3     gate22370  (.A(g20185), .B(g20149), .C(II28335), .Z(g21810) ) ;
NAND2   gate22371  (.A(g16781), .B(g16797), .Z(g19138) ) ;
OR3     gate22372  (.A(g19138), .B(g16974), .C(g14936), .Z(g21811) ) ;
OR4     gate22373  (.A(g20146), .B(g20118), .C(g18597), .D(g19104), .Z(g21813) ) ;
OR3     gate22374  (.A(g19106), .B(g19101), .C(g19095), .Z(II28341) ) ;
OR4     gate22375  (.A(g16558), .B(g19080), .C(g16513), .D(II28341), .Z(g21814) ) ;
OR4     gate22376  (.A(g18717), .B(g20293), .C(g20283), .D(g18654), .Z(g21815) ) ;
OR3     gate22377  (.A(g19138), .B(g19681), .C(g16743), .Z(g21816) ) ;
OR3     gate22378  (.A(g20277), .B(g20268), .C(g20247), .Z(II28346) ) ;
OR3     gate22379  (.A(g20219), .B(g20187), .C(II28346), .Z(g21817) ) ;
OR4     gate22380  (.A(g20184), .B(g20148), .C(g18629), .D(g19109), .Z(g21819) ) ;
OR3     gate22381  (.A(g19111), .B(g19108), .C(g19102), .Z(II28351) ) ;
OR4     gate22382  (.A(g16590), .B(g19090), .C(g16535), .D(II28351), .Z(g21820) ) ;
OR4     gate22383  (.A(g18753), .B(g20309), .C(g20294), .D(g18668), .Z(g21821) ) ;
OR4     gate22384  (.A(g20218), .B(g20186), .C(g18638), .D(g19116), .Z(g21823) ) ;
OR3     gate22385  (.A(g20280), .B(g18652), .C(g18649), .Z(II28365) ) ;
OR3     gate22386  (.A(g20222), .B(g18645), .C(II28365), .Z(g21844) ) ;
OR3     gate22387  (.A(g20291), .B(g18666), .C(g18653), .Z(II28369) ) ;
OR3     gate22388  (.A(g20249), .B(g18648), .C(II28369), .Z(g21846) ) ;
OR3     gate22389  (.A(g20307), .B(g18689), .C(g18667), .Z(II28374) ) ;
OR3     gate22390  (.A(g20272), .B(g18651), .C(II28374), .Z(g21849) ) ;
OR3     gate22391  (.A(g20326), .B(g18718), .C(g18690), .Z(II28380) ) ;
OR3     gate22392  (.A(g20284), .B(g18655), .C(II28380), .Z(g21856) ) ;
OR2     gate22393  (.A(g16075), .B(g20842), .Z(g22175) ) ;
OR2     gate22394  (.A(g16113), .B(g20850), .Z(g22190) ) ;
OR2     gate22395  (.A(g16164), .B(g20858), .Z(g22199) ) ;
OR2     gate22396  (.A(g16223), .B(g20866), .Z(g22205) ) ;
NOR2    gate22397  (.A(g499), .B(g8983), .Z(g12451) ) ;
NAND3   gate22398  (.A(g21207), .B(g21266), .C(g21196), .Z(g22385) ) ;
OR2     gate22399  (.A(g14493), .B(g22385), .Z(g23319) ) ;
OR2     gate22400  (.A(g23106), .B(g21906), .Z(g23688) ) ;
OR2     gate22401  (.A(g23119), .B(g21920), .Z(g23742) ) ;
OR2     gate22402  (.A(g23128), .B(g21938), .Z(g23797) ) ;
OR2     gate22403  (.A(g23139), .B(g20647), .Z(g23850) ) ;
OR2     gate22404  (.A(g19387), .B(g22401), .Z(g24239) ) ;
NAND3   gate22405  (.A(g21152), .B(g21241), .C(g21136), .Z(g22317) ) ;
OR2     gate22406  (.A(g14144), .B(g22317), .Z(g24244) ) ;
OR2     gate22407  (.A(g19417), .B(g22402), .Z(g24245) ) ;
NAND3   gate22408  (.A(g21172), .B(g21249), .C(g21156), .Z(g22342) ) ;
OR2     gate22409  (.A(g14259), .B(g22342), .Z(g24252) ) ;
OR2     gate22410  (.A(g19454), .B(g22403), .Z(g24254) ) ;
NAND3   gate22411  (.A(g21192), .B(g21258), .C(g21176), .Z(g22365) ) ;
OR2     gate22412  (.A(g14381), .B(g22365), .Z(g24257) ) ;
OR2     gate22413  (.A(g19481), .B(g22404), .Z(g24258) ) ;
NOR2    gate22414  (.A(g4456), .B(g22985), .Z(g23922) ) ;
OR2     gate22415  (.A(g23922), .B(g23945), .Z(g24965) ) ;
NOR2    gate22416  (.A(g4632), .B(g22987), .Z(g23954) ) ;
OR2     gate22417  (.A(g23954), .B(g23974), .Z(g24978) ) ;
NOR2    gate22418  (.A(g4809), .B(g22990), .Z(g23983) ) ;
OR2     gate22419  (.A(g23983), .B(g24004), .Z(g24989) ) ;
NOR2    gate22420  (.A(g4985), .B(g22997), .Z(g24013) ) ;
OR2     gate22421  (.A(g24013), .B(g24038), .Z(g25000) ) ;
OR2     gate22422  (.A(g24958), .B(g24893), .Z(g25183) ) ;
OR2     gate22423  (.A(g24969), .B(g24916), .Z(g25186) ) ;
OR2     gate22424  (.A(g24982), .B(g24933), .Z(g25190) ) ;
OR2     gate22425  (.A(g24993), .B(g24945), .Z(g25195) ) ;
NOR3    gate22426  (.A(g4456), .B(g14831), .C(g25078), .Z(g25852) ) ;
OR2     gate22427  (.A(g25852), .B(g25870), .Z(g26320) ) ;
NOR3    gate22428  (.A(g4632), .B(g14904), .C(g25082), .Z(g25873) ) ;
OR2     gate22429  (.A(g25873), .B(g25882), .Z(g26367) ) ;
NOR3    gate22430  (.A(g4809), .B(g14985), .C(g25091), .Z(g25885) ) ;
OR2     gate22431  (.A(g25885), .B(g25887), .Z(g26410) ) ;
NOR3    gate22432  (.A(g4985), .B(g15074), .C(g25099), .Z(g25890) ) ;
OR2     gate22433  (.A(g25890), .B(g25892), .Z(g26451) ) ;
NAND2   gate22434  (.A(g25367), .B(g27415), .Z(g27738) ) ;
NAND2   gate22435  (.A(g25384), .B(g27436), .Z(g27743) ) ;
NAND2   gate22436  (.A(g25400), .B(g27455), .Z(g27751) ) ;
NAND2   gate22437  (.A(g25410), .B(g27471), .Z(g27756) ) ;
NAND2   gate22438  (.A(g2981), .B(g2874), .Z(II15167) ) ;
NAND2   gate22439  (.A(g2981), .B(II15167), .Z(II15168) ) ;
NAND2   gate22440  (.A(g2874), .B(II15167), .Z(II15169) ) ;
NAND2   gate22441  (.A(II15168), .B(II15169), .Z(g7855) ) ;
NAND2   gate22442  (.A(g2975), .B(g2978), .Z(II15183) ) ;
NAND2   gate22443  (.A(g2975), .B(II15183), .Z(II15184) ) ;
NAND2   gate22444  (.A(g2978), .B(II15183), .Z(II15185) ) ;
NAND2   gate22445  (.A(II15184), .B(II15185), .Z(g7875) ) ;
NAND2   gate22446  (.A(g2956), .B(g2959), .Z(II15190) ) ;
NAND2   gate22447  (.A(g2956), .B(II15190), .Z(II15191) ) ;
NAND2   gate22448  (.A(g2959), .B(II15190), .Z(II15192) ) ;
NAND2   gate22449  (.A(II15191), .B(II15192), .Z(g7876) ) ;
NAND2   gate22450  (.A(g2969), .B(g2972), .Z(II15204) ) ;
NAND2   gate22451  (.A(g2969), .B(II15204), .Z(II15205) ) ;
NAND2   gate22452  (.A(g2972), .B(II15204), .Z(II15206) ) ;
NAND2   gate22453  (.A(II15205), .B(II15206), .Z(g7895) ) ;
NAND2   gate22454  (.A(g2947), .B(g2953), .Z(II15211) ) ;
NAND2   gate22455  (.A(g2947), .B(II15211), .Z(II15212) ) ;
NAND2   gate22456  (.A(g2953), .B(II15211), .Z(II15213) ) ;
NAND2   gate22457  (.A(II15212), .B(II15213), .Z(g7896) ) ;
NAND2   gate22458  (.A(g2963), .B(g2966), .Z(II15237) ) ;
NAND2   gate22459  (.A(g2963), .B(II15237), .Z(II15238) ) ;
NAND2   gate22460  (.A(g2966), .B(II15237), .Z(II15239) ) ;
NAND2   gate22461  (.A(II15238), .B(II15239), .Z(g7922) ) ;
NAND2   gate22462  (.A(g2941), .B(g2944), .Z(II15244) ) ;
NAND2   gate22463  (.A(g2941), .B(II15244), .Z(II15245) ) ;
NAND2   gate22464  (.A(g2944), .B(II15244), .Z(II15246) ) ;
NAND2   gate22465  (.A(II15245), .B(II15246), .Z(g7923) ) ;
NAND2   gate22466  (.A(g2935), .B(g2938), .Z(II15276) ) ;
NAND2   gate22467  (.A(g2935), .B(II15276), .Z(II15277) ) ;
NAND2   gate22468  (.A(g2938), .B(II15276), .Z(II15278) ) ;
NAND2   gate22469  (.A(II15277), .B(II15278), .Z(g7970) ) ;
NAND2   gate22470  (.A(g4203), .B(g3998), .Z(II16879) ) ;
NAND2   gate22471  (.A(g4203), .B(II16879), .Z(II16880) ) ;
NAND2   gate22472  (.A(g3998), .B(II16879), .Z(II16881) ) ;
NAND2   gate22473  (.A(II16880), .B(II16881), .Z(g9883) ) ;
NAND2   gate22474  (.A(g4734), .B(g4452), .Z(II16965) ) ;
NAND2   gate22475  (.A(g4734), .B(II16965), .Z(II16966) ) ;
NAND2   gate22476  (.A(g4452), .B(II16965), .Z(II16967) ) ;
NAND2   gate22477  (.A(II16966), .B(II16967), .Z(g10003) ) ;
NAND2   gate22478  (.A(g6637), .B(g6309), .Z(II17059) ) ;
NAND2   gate22479  (.A(g6637), .B(II17059), .Z(II17060) ) ;
NAND2   gate22480  (.A(g6309), .B(II17059), .Z(II17061) ) ;
NAND2   gate22481  (.A(II17060), .B(II17061), .Z(g10095) ) ;
NAND2   gate22482  (.A(g7465), .B(g7142), .Z(II17149) ) ;
NAND2   gate22483  (.A(g7465), .B(II17149), .Z(II17150) ) ;
NAND2   gate22484  (.A(g7142), .B(II17149), .Z(II17151) ) ;
NAND2   gate22485  (.A(II17150), .B(II17151), .Z(g10185) ) ;
NAND2   gate22486  (.A(g7875), .B(g7855), .Z(II18106) ) ;
NAND2   gate22487  (.A(g7875), .B(II18106), .Z(II18107) ) ;
NAND2   gate22488  (.A(g7855), .B(II18106), .Z(II18108) ) ;
NAND2   gate22489  (.A(II18107), .B(II18108), .Z(g11188) ) ;
NAND2   gate22490  (.A(g3997), .B(g8181), .Z(II18113) ) ;
NAND2   gate22491  (.A(g3997), .B(II18113), .Z(II18114) ) ;
NAND2   gate22492  (.A(g8181), .B(II18113), .Z(II18115) ) ;
NAND2   gate22493  (.A(II18114), .B(II18115), .Z(g11189) ) ;
NAND2   gate22494  (.A(g7922), .B(g7895), .Z(II18190) ) ;
NAND2   gate22495  (.A(g7922), .B(II18190), .Z(II18191) ) ;
NAND2   gate22496  (.A(g7895), .B(II18190), .Z(II18192) ) ;
NAND2   gate22497  (.A(II18191), .B(II18192), .Z(g11262) ) ;
NAND2   gate22498  (.A(g7896), .B(g7876), .Z(II18197) ) ;
NAND2   gate22499  (.A(g7896), .B(II18197), .Z(II18198) ) ;
NAND2   gate22500  (.A(g7876), .B(II18197), .Z(II18199) ) ;
NAND2   gate22501  (.A(II18198), .B(II18199), .Z(g11263) ) ;
NAND2   gate22502  (.A(g7975), .B(g4202), .Z(II18204) ) ;
NAND2   gate22503  (.A(g7975), .B(II18204), .Z(II18205) ) ;
NAND2   gate22504  (.A(g4202), .B(II18204), .Z(II18206) ) ;
NAND2   gate22505  (.A(II18205), .B(II18206), .Z(g11264) ) ;
NAND2   gate22506  (.A(g7970), .B(g7923), .Z(II18280) ) ;
NAND2   gate22507  (.A(g7970), .B(II18280), .Z(II18281) ) ;
NAND2   gate22508  (.A(g7923), .B(II18280), .Z(II18282) ) ;
NAND2   gate22509  (.A(II18281), .B(II18282), .Z(g11330) ) ;
NAND2   gate22510  (.A(g8256), .B(g8102), .Z(II18287) ) ;
NAND2   gate22511  (.A(g8256), .B(II18287), .Z(II18288) ) ;
NAND2   gate22512  (.A(g8102), .B(II18287), .Z(II18289) ) ;
NAND2   gate22513  (.A(II18288), .B(II18289), .Z(g11331) ) ;
NAND2   gate22514  (.A(g4325), .B(g4093), .Z(II18368) ) ;
NAND2   gate22515  (.A(g4325), .B(II18368), .Z(II18369) ) ;
NAND2   gate22516  (.A(g4093), .B(II18368), .Z(II18370) ) ;
NAND2   gate22517  (.A(II18369), .B(II18370), .Z(g11410) ) ;
NAND2   gate22518  (.A(g11410), .B(g11331), .Z(II18799) ) ;
NAND2   gate22519  (.A(g11410), .B(II18799), .Z(II18800) ) ;
NAND2   gate22520  (.A(g11331), .B(II18799), .Z(II18801) ) ;
NAND2   gate22521  (.A(II18800), .B(II18801), .Z(g11621) ) ;
NAND2   gate22522  (.A(g10003), .B(g9883), .Z(II20031) ) ;
NAND2   gate22523  (.A(g10003), .B(II20031), .Z(II20032) ) ;
NAND2   gate22524  (.A(g9883), .B(II20031), .Z(II20033) ) ;
NAND2   gate22525  (.A(II20032), .B(II20033), .Z(g12988) ) ;
NAND2   gate22526  (.A(g10185), .B(g10095), .Z(II20048) ) ;
NAND2   gate22527  (.A(g10185), .B(II20048), .Z(II20049) ) ;
NAND2   gate22528  (.A(g10095), .B(II20048), .Z(II20050) ) ;
NAND2   gate22529  (.A(II20049), .B(II20050), .Z(g12999) ) ;
NAND2   gate22530  (.A(g11262), .B(g11188), .Z(II20429) ) ;
NAND2   gate22531  (.A(g11262), .B(II20429), .Z(II20430) ) ;
NAND2   gate22532  (.A(g11188), .B(II20429), .Z(II20431) ) ;
NAND2   gate22533  (.A(II20430), .B(II20431), .Z(g13348) ) ;
NAND2   gate22534  (.A(g11330), .B(g11263), .Z(II20465) ) ;
NAND2   gate22535  (.A(g11330), .B(II20465), .Z(II20466) ) ;
NAND2   gate22536  (.A(g11263), .B(II20465), .Z(II20467) ) ;
NAND2   gate22537  (.A(II20466), .B(II20467), .Z(g13370) ) ;
NAND2   gate22538  (.A(g11264), .B(g11189), .Z(II20504) ) ;
NAND2   gate22539  (.A(g11264), .B(II20504), .Z(II20505) ) ;
NAND2   gate22540  (.A(g11189), .B(II20504), .Z(II20506) ) ;
NAND2   gate22541  (.A(II20505), .B(II20506), .Z(g13399) ) ;
NAND2   gate22542  (.A(g11621), .B(g13399), .Z(II20743) ) ;
NAND2   gate22543  (.A(g11621), .B(II20743), .Z(II20744) ) ;
NAND2   gate22544  (.A(g13399), .B(II20743), .Z(II20745) ) ;
NAND2   gate22545  (.A(II20744), .B(II20745), .Z(g13507) ) ;
NAND2   gate22546  (.A(g8580), .B(g12463), .Z(g13893) ) ;
NAND3   gate22547  (.A(g8822), .B(g12473), .C(g12463), .Z(g13915) ) ;
NAND2   gate22548  (.A(g8587), .B(g12478), .Z(g13934) ) ;
NAND2   gate22549  (.A(g10730), .B(g12473), .Z(g13957) ) ;
NAND3   gate22550  (.A(g8846), .B(g12490), .C(g12478), .Z(g13971) ) ;
NAND2   gate22551  (.A(g8594), .B(g12495), .Z(g13990) ) ;
NAND2   gate22552  (.A(g10749), .B(g12490), .Z(g14027) ) ;
NAND3   gate22553  (.A(g8873), .B(g12510), .C(g12495), .Z(g14041) ) ;
NAND2   gate22554  (.A(g8605), .B(g12515), .Z(g14060) ) ;
NAND2   gate22555  (.A(g10767), .B(g12510), .Z(g14118) ) ;
NAND3   gate22556  (.A(g8911), .B(g12527), .C(g12515), .Z(g14132) ) ;
NAND2   gate22557  (.A(g10773), .B(g12527), .Z(g14233) ) ;
NOR2    gate22558  (.A(g9187), .B(g9161), .Z(g12780) ) ;
NOR2    gate22559  (.A(g9248), .B(g9203), .Z(g12819) ) ;
NOR2    gate22560  (.A(g9326), .B(g9264), .Z(g12857) ) ;
NOR4    gate22561  (.A(g11481), .B(g11332), .C(g7928), .D(g11069), .Z(g13401) ) ;
NOR2    gate22562  (.A(g9407), .B(g9342), .Z(g12898) ) ;
NOR4    gate22563  (.A(g11481), .B(g11332), .C(g11190), .D(g7880), .Z(g13286) ) ;
NOR4    gate22564  (.A(g8183), .B(g11332), .C(g11190), .D(g7880), .Z(g13313) ) ;
NOR4    gate22565  (.A(g8183), .B(g11332), .C(g7928), .D(g11069), .Z(g11622) ) ;
NOR4    gate22566  (.A(g11481), .B(g8045), .C(g11190), .D(g7880), .Z(g13332) ) ;
NOR4    gate22567  (.A(g11481), .B(g8045), .C(g7928), .D(g11069), .Z(g11643) ) ;
NOR4    gate22568  (.A(g11481), .B(g11332), .C(g7928), .D(g7880), .Z(g13375) ) ;
NOR4    gate22569  (.A(g8183), .B(g8045), .C(g7928), .D(g11069), .Z(g11660) ) ;
NAND2   gate22570  (.A(g12999), .B(g12988), .Z(II22062) ) ;
NAND2   gate22571  (.A(g12999), .B(II22062), .Z(II22063) ) ;
NAND2   gate22572  (.A(g12988), .B(II22062), .Z(II22064) ) ;
NAND2   gate22573  (.A(II22063), .B(II22064), .Z(g15814) ) ;
NOR4    gate22574  (.A(g11481), .B(g8045), .C(g7928), .D(g7880), .Z(g13024) ) ;
NOR4    gate22575  (.A(g11481), .B(g11332), .C(g11190), .D(g11069), .Z(g13310) ) ;
NOR4    gate22576  (.A(g8183), .B(g11332), .C(g11190), .D(g11069), .Z(g13331) ) ;
NOR4    gate22577  (.A(g11481), .B(g8045), .C(g11190), .D(g11069), .Z(g13353) ) ;
NOR4    gate22578  (.A(g8183), .B(g8045), .C(g11190), .D(g7880), .Z(g13354) ) ;
NOR4    gate22579  (.A(g8183), .B(g8045), .C(g11190), .D(g11069), .Z(g13374) ) ;
NOR4    gate22580  (.A(g8183), .B(g11332), .C(g7928), .D(g7880), .Z(g13404) ) ;
NAND2   gate22581  (.A(g2962), .B(g13348), .Z(II22282) ) ;
NAND2   gate22582  (.A(g2962), .B(II22282), .Z(II22283) ) ;
NAND2   gate22583  (.A(g13348), .B(II22282), .Z(II22284) ) ;
NAND2   gate22584  (.A(g2934), .B(g13370), .Z(II22316) ) ;
NAND2   gate22585  (.A(g2934), .B(II22316), .Z(II22317) ) ;
NAND2   gate22586  (.A(g13370), .B(II22316), .Z(II22318) ) ;
NOR2    gate22587  (.A(g11737), .B(g7152), .Z(g15978) ) ;
NAND2   gate22588  (.A(g13507), .B(g15978), .Z(II22630) ) ;
NAND2   gate22589  (.A(g13507), .B(II22630), .Z(II22631) ) ;
NAND2   gate22590  (.A(g15978), .B(II22630), .Z(II22632) ) ;
NOR2    gate22591  (.A(g11737), .B(g7345), .Z(g15661) ) ;
NAND2   gate22592  (.A(g13348), .B(g15661), .Z(II22705) ) ;
NAND2   gate22593  (.A(g13348), .B(II22705), .Z(II22706) ) ;
NAND2   gate22594  (.A(g15661), .B(II22705), .Z(II22707) ) ;
NAND2   gate22595  (.A(g13370), .B(g15661), .Z(II22884) ) ;
NAND2   gate22596  (.A(g13370), .B(II22884), .Z(II22885) ) ;
NAND2   gate22597  (.A(g15661), .B(II22884), .Z(II22886) ) ;
NAND2   gate22598  (.A(g15022), .B(g14000), .Z(II22900) ) ;
NAND2   gate22599  (.A(g15022), .B(II22900), .Z(II22901) ) ;
NAND2   gate22600  (.A(g14000), .B(II22900), .Z(II22902) ) ;
NAND2   gate22601  (.A(g15096), .B(g13945), .Z(II22917) ) ;
NAND2   gate22602  (.A(g15096), .B(II22917), .Z(II22918) ) ;
NAND2   gate22603  (.A(g13945), .B(II22917), .Z(II22919) ) ;
NAND2   gate22604  (.A(g15118), .B(g14091), .Z(II22924) ) ;
NAND2   gate22605  (.A(g15118), .B(II22924), .Z(II22925) ) ;
NAND2   gate22606  (.A(g14091), .B(II22924), .Z(II22926) ) ;
NAND2   gate22607  (.A(g9150), .B(g13906), .Z(II22936) ) ;
NAND2   gate22608  (.A(g9150), .B(II22936), .Z(II22937) ) ;
NAND2   gate22609  (.A(g13906), .B(II22936), .Z(II22938) ) ;
NAND2   gate22610  (.A(g15188), .B(g14015), .Z(II22945) ) ;
NAND2   gate22611  (.A(g15188), .B(II22945), .Z(II22946) ) ;
NAND2   gate22612  (.A(g14015), .B(II22945), .Z(II22947) ) ;
NAND2   gate22613  (.A(g15210), .B(g14206), .Z(II22952) ) ;
NAND2   gate22614  (.A(g15210), .B(II22952), .Z(II22953) ) ;
NAND2   gate22615  (.A(g14206), .B(II22952), .Z(II22954) ) ;
NAND2   gate22616  (.A(g9161), .B(g13885), .Z(II22962) ) ;
NAND2   gate22617  (.A(g9161), .B(II22962), .Z(II22963) ) ;
NAND2   gate22618  (.A(g13885), .B(II22962), .Z(II22964) ) ;
NAND2   gate22619  (.A(g9174), .B(g13962), .Z(II22972) ) ;
NAND2   gate22620  (.A(g9174), .B(II22972), .Z(II22973) ) ;
NAND2   gate22621  (.A(g13962), .B(II22972), .Z(II22974) ) ;
NAND2   gate22622  (.A(g15274), .B(g14106), .Z(II22981) ) ;
NAND2   gate22623  (.A(g15274), .B(II22981), .Z(II22982) ) ;
NAND2   gate22624  (.A(g14106), .B(II22981), .Z(II22983) ) ;
NAND2   gate22625  (.A(g15296), .B(g14321), .Z(II22988) ) ;
NAND2   gate22626  (.A(g15296), .B(II22988), .Z(II22989) ) ;
NAND2   gate22627  (.A(g14321), .B(II22988), .Z(II22990) ) ;
NAND2   gate22628  (.A(g9187), .B(g13872), .Z(II22998) ) ;
NAND2   gate22629  (.A(g9187), .B(II22998), .Z(II22999) ) ;
NAND2   gate22630  (.A(g13872), .B(II22998), .Z(II23000) ) ;
NAND2   gate22631  (.A(g9203), .B(g13926), .Z(II23008) ) ;
NAND2   gate22632  (.A(g9203), .B(II23008), .Z(II23009) ) ;
NAND2   gate22633  (.A(g13926), .B(II23008), .Z(II23010) ) ;
NAND2   gate22634  (.A(g9216), .B(g14032), .Z(II23018) ) ;
NAND2   gate22635  (.A(g9216), .B(II23018), .Z(II23019) ) ;
NAND2   gate22636  (.A(g14032), .B(II23018), .Z(II23020) ) ;
NAND2   gate22637  (.A(g15366), .B(g14221), .Z(II23027) ) ;
NAND2   gate22638  (.A(g15366), .B(II23027), .Z(II23028) ) ;
NAND2   gate22639  (.A(g14221), .B(II23027), .Z(II23029) ) ;
NAND2   gate22640  (.A(g9232), .B(g13864), .Z(II23034) ) ;
NAND2   gate22641  (.A(g9232), .B(II23034), .Z(II23035) ) ;
NAND2   gate22642  (.A(g13864), .B(II23034), .Z(II23036) ) ;
NAND2   gate22643  (.A(g9248), .B(g13894), .Z(II23045) ) ;
NAND2   gate22644  (.A(g9248), .B(II23045), .Z(II23046) ) ;
NAND2   gate22645  (.A(g13894), .B(II23045), .Z(II23047) ) ;
NAND2   gate22646  (.A(g9264), .B(g13982), .Z(II23055) ) ;
NAND2   gate22647  (.A(g9264), .B(II23055), .Z(II23056) ) ;
NAND2   gate22648  (.A(g13982), .B(II23055), .Z(II23057) ) ;
NAND2   gate22649  (.A(g9277), .B(g14123), .Z(II23065) ) ;
NAND2   gate22650  (.A(g9277), .B(II23065), .Z(II23066) ) ;
NAND2   gate22651  (.A(g14123), .B(II23065), .Z(II23067) ) ;
NAND2   gate22652  (.A(g9293), .B(g13856), .Z(II23074) ) ;
NAND2   gate22653  (.A(g9293), .B(II23074), .Z(II23075) ) ;
NAND2   gate22654  (.A(g13856), .B(II23074), .Z(II23076) ) ;
NAND2   gate22655  (.A(g9310), .B(g13879), .Z(II23082) ) ;
NAND2   gate22656  (.A(g9310), .B(II23082), .Z(II23083) ) ;
NAND2   gate22657  (.A(g13879), .B(II23082), .Z(II23084) ) ;
NAND2   gate22658  (.A(g9326), .B(g13935), .Z(II23093) ) ;
NAND2   gate22659  (.A(g9326), .B(II23093), .Z(II23094) ) ;
NAND2   gate22660  (.A(g13935), .B(II23093), .Z(II23095) ) ;
NAND2   gate22661  (.A(g9342), .B(g14052), .Z(II23103) ) ;
NAND2   gate22662  (.A(g9342), .B(II23103), .Z(II23104) ) ;
NAND2   gate22663  (.A(g14052), .B(II23103), .Z(II23105) ) ;
NAND2   gate22664  (.A(g9356), .B(g13848), .Z(II23113) ) ;
NAND2   gate22665  (.A(g9356), .B(II23113), .Z(II23114) ) ;
NAND2   gate22666  (.A(g13848), .B(II23113), .Z(II23115) ) ;
NAND2   gate22667  (.A(g9374), .B(g13866), .Z(II23123) ) ;
NAND2   gate22668  (.A(g9374), .B(II23123), .Z(II23124) ) ;
NAND2   gate22669  (.A(g13866), .B(II23123), .Z(II23125) ) ;
NAND2   gate22670  (.A(g9391), .B(g13901), .Z(II23131) ) ;
NAND2   gate22671  (.A(g9391), .B(II23131), .Z(II23132) ) ;
NAND2   gate22672  (.A(g13901), .B(II23131), .Z(II23133) ) ;
NAND2   gate22673  (.A(g9407), .B(g13991), .Z(II23142) ) ;
NAND2   gate22674  (.A(g9407), .B(II23142), .Z(II23143) ) ;
NAND2   gate22675  (.A(g13991), .B(II23142), .Z(II23144) ) ;
NAND2   gate22676  (.A(g9427), .B(g14061), .Z(II23152) ) ;
NAND2   gate22677  (.A(g9427), .B(II23152), .Z(II23153) ) ;
NAND2   gate22678  (.A(g14061), .B(II23152), .Z(II23154) ) ;
NAND2   gate22679  (.A(g9453), .B(g13857), .Z(II23161) ) ;
NAND2   gate22680  (.A(g9453), .B(II23161), .Z(II23162) ) ;
NAND2   gate22681  (.A(g13857), .B(II23161), .Z(II23163) ) ;
NAND2   gate22682  (.A(g9471), .B(g13881), .Z(II23171) ) ;
NAND2   gate22683  (.A(g9471), .B(II23171), .Z(II23172) ) ;
NAND2   gate22684  (.A(g13881), .B(II23171), .Z(II23173) ) ;
NAND2   gate22685  (.A(g9488), .B(g13942), .Z(II23179) ) ;
NAND2   gate22686  (.A(g9488), .B(II23179), .Z(II23180) ) ;
NAND2   gate22687  (.A(g13942), .B(II23179), .Z(II23181) ) ;
NAND2   gate22688  (.A(g9507), .B(g13999), .Z(II23190) ) ;
NAND2   gate22689  (.A(g9507), .B(II23190), .Z(II23191) ) ;
NAND2   gate22690  (.A(g13999), .B(II23190), .Z(II23192) ) ;
NAND2   gate22691  (.A(g9569), .B(g14176), .Z(II23198) ) ;
NAND2   gate22692  (.A(g9569), .B(II23198), .Z(II23199) ) ;
NAND2   gate22693  (.A(g14176), .B(II23198), .Z(II23200) ) ;
NAND2   gate22694  (.A(g9595), .B(g13867), .Z(II23207) ) ;
NAND2   gate22695  (.A(g9595), .B(II23207), .Z(II23208) ) ;
NAND2   gate22696  (.A(g13867), .B(II23207), .Z(II23209) ) ;
NAND2   gate22697  (.A(g9613), .B(g13903), .Z(II23217) ) ;
NAND2   gate22698  (.A(g9613), .B(II23217), .Z(II23218) ) ;
NAND2   gate22699  (.A(g13903), .B(II23217), .Z(II23219) ) ;
NAND2   gate22700  (.A(g9649), .B(g14090), .Z(II23225) ) ;
NAND2   gate22701  (.A(g9649), .B(II23225), .Z(II23226) ) ;
NAND2   gate22702  (.A(g14090), .B(II23225), .Z(II23227) ) ;
NAND2   gate22703  (.A(g9711), .B(g14291), .Z(II23233) ) ;
NAND2   gate22704  (.A(g9711), .B(II23233), .Z(II23234) ) ;
NAND2   gate22705  (.A(g14291), .B(II23233), .Z(II23235) ) ;
NAND2   gate22706  (.A(g9737), .B(g13882), .Z(II23242) ) ;
NAND2   gate22707  (.A(g9737), .B(II23242), .Z(II23243) ) ;
NAND2   gate22708  (.A(g13882), .B(II23242), .Z(II23244) ) ;
NAND2   gate22709  (.A(g9795), .B(g14205), .Z(II23256) ) ;
NAND2   gate22710  (.A(g9795), .B(II23256), .Z(II23257) ) ;
NAND2   gate22711  (.A(g14205), .B(II23256), .Z(II23258) ) ;
NAND2   gate22712  (.A(g9857), .B(g14413), .Z(II23264) ) ;
NAND2   gate22713  (.A(g9857), .B(II23264), .Z(II23265) ) ;
NAND2   gate22714  (.A(g14413), .B(II23264), .Z(II23266) ) ;
NAND2   gate22715  (.A(g9941), .B(g14320), .Z(II23277) ) ;
NAND2   gate22716  (.A(g9941), .B(II23277), .Z(II23278) ) ;
NAND2   gate22717  (.A(g14320), .B(II23277), .Z(II23279) ) ;
NAND2   gate22718  (.A(g14062), .B(g9150), .Z(II23806) ) ;
NAND2   gate22719  (.A(g14062), .B(II23806), .Z(II23807) ) ;
NAND2   gate22720  (.A(g9150), .B(II23806), .Z(II23808) ) ;
NAND2   gate22721  (.A(g14001), .B(g9187), .Z(II23878) ) ;
NAND2   gate22722  (.A(g14001), .B(II23878), .Z(II23879) ) ;
NAND2   gate22723  (.A(g9187), .B(II23878), .Z(II23880) ) ;
NAND2   gate22724  (.A(g14177), .B(g9174), .Z(II23893) ) ;
NAND2   gate22725  (.A(g14177), .B(II23893), .Z(II23894) ) ;
NAND2   gate22726  (.A(g9174), .B(II23893), .Z(II23895) ) ;
NAND2   gate22727  (.A(g13946), .B(g9293), .Z(II23941) ) ;
NAND2   gate22728  (.A(g13946), .B(II23941), .Z(II23942) ) ;
NAND2   gate22729  (.A(g9293), .B(II23941), .Z(II23943) ) ;
NAND2   gate22730  (.A(g6513), .B(g14171), .Z(II23958) ) ;
NAND2   gate22731  (.A(g6513), .B(II23958), .Z(II23959) ) ;
NAND2   gate22732  (.A(g14171), .B(II23958), .Z(II23960) ) ;
NAND2   gate22733  (.A(g14092), .B(g9248), .Z(II23966) ) ;
NAND2   gate22734  (.A(g14092), .B(II23966), .Z(II23967) ) ;
NAND2   gate22735  (.A(g9248), .B(II23966), .Z(II23968) ) ;
NAND2   gate22736  (.A(g14292), .B(g9216), .Z(II23981) ) ;
NAND2   gate22737  (.A(g14292), .B(II23981), .Z(II23982) ) ;
NAND2   gate22738  (.A(g9216), .B(II23981), .Z(II23983) ) ;
NAND2   gate22739  (.A(g7548), .B(g15814), .Z(II24005) ) ;
NAND2   gate22740  (.A(g7548), .B(II24005), .Z(II24006) ) ;
NAND2   gate22741  (.A(g15814), .B(II24005), .Z(II24007) ) ;
NAND2   gate22742  (.A(g13907), .B(g9427), .Z(II24015) ) ;
NAND2   gate22743  (.A(g13907), .B(II24015), .Z(II24016) ) ;
NAND2   gate22744  (.A(g9427), .B(II24015), .Z(II24017) ) ;
NAND2   gate22745  (.A(g6201), .B(g14086), .Z(II24028) ) ;
NAND2   gate22746  (.A(g6201), .B(II24028), .Z(II24029) ) ;
NAND2   gate22747  (.A(g14086), .B(II24028), .Z(II24030) ) ;
NAND2   gate22748  (.A(g14016), .B(g9374), .Z(II24036) ) ;
NAND2   gate22749  (.A(g14016), .B(II24036), .Z(II24037) ) ;
NAND2   gate22750  (.A(g9374), .B(II24036), .Z(II24038) ) ;
NAND2   gate22751  (.A(g6777), .B(g14286), .Z(II24053) ) ;
NAND2   gate22752  (.A(g6777), .B(II24053), .Z(II24054) ) ;
NAND2   gate22753  (.A(g14286), .B(II24053), .Z(II24055) ) ;
NAND2   gate22754  (.A(g14207), .B(g9326), .Z(II24061) ) ;
NAND2   gate22755  (.A(g14207), .B(II24061), .Z(II24062) ) ;
NAND2   gate22756  (.A(g9326), .B(II24061), .Z(II24063) ) ;
NAND2   gate22757  (.A(g14414), .B(g9277), .Z(II24076) ) ;
NAND2   gate22758  (.A(g14414), .B(II24076), .Z(II24077) ) ;
NAND2   gate22759  (.A(g9277), .B(II24076), .Z(II24078) ) ;
NAND2   gate22760  (.A(g13886), .B(g15096), .Z(II24091) ) ;
NAND2   gate22761  (.A(g13886), .B(II24091), .Z(II24092) ) ;
NAND2   gate22762  (.A(g15096), .B(II24091), .Z(II24093) ) ;
NAND2   gate22763  (.A(g6363), .B(g14011), .Z(II24102) ) ;
NAND2   gate22764  (.A(g6363), .B(II24102), .Z(II24103) ) ;
NAND2   gate22765  (.A(g14011), .B(II24102), .Z(II24104) ) ;
NAND2   gate22766  (.A(g13963), .B(g9569), .Z(II24110) ) ;
NAND2   gate22767  (.A(g13963), .B(II24110), .Z(II24111) ) ;
NAND2   gate22768  (.A(g9569), .B(II24110), .Z(II24112) ) ;
NAND2   gate22769  (.A(g6290), .B(g14201), .Z(II24123) ) ;
NAND2   gate22770  (.A(g6290), .B(II24123), .Z(II24124) ) ;
NAND2   gate22771  (.A(g14201), .B(II24123), .Z(II24125) ) ;
NAND2   gate22772  (.A(g14107), .B(g9471), .Z(II24131) ) ;
NAND2   gate22773  (.A(g14107), .B(II24131), .Z(II24132) ) ;
NAND2   gate22774  (.A(g9471), .B(II24131), .Z(II24133) ) ;
NAND2   gate22775  (.A(g7079), .B(g14408), .Z(II24148) ) ;
NAND2   gate22776  (.A(g7079), .B(II24148), .Z(II24149) ) ;
NAND2   gate22777  (.A(g14408), .B(II24148), .Z(II24150) ) ;
NAND2   gate22778  (.A(g14322), .B(g9407), .Z(II24156) ) ;
NAND2   gate22779  (.A(g14322), .B(II24156), .Z(II24157) ) ;
NAND2   gate22780  (.A(g9407), .B(II24156), .Z(II24158) ) ;
NAND2   gate22781  (.A(g13873), .B(g9161), .Z(II24178) ) ;
NAND2   gate22782  (.A(g13873), .B(II24178), .Z(II24179) ) ;
NAND2   gate22783  (.A(g9161), .B(II24178), .Z(II24180) ) ;
NAND2   gate22784  (.A(g6177), .B(g13958), .Z(II24186) ) ;
NAND2   gate22785  (.A(g6177), .B(II24186), .Z(II24187) ) ;
NAND2   gate22786  (.A(g13958), .B(II24186), .Z(II24188) ) ;
NAND2   gate22787  (.A(g13927), .B(g15188), .Z(II24194) ) ;
NAND2   gate22788  (.A(g13927), .B(II24194), .Z(II24195) ) ;
NAND2   gate22789  (.A(g15188), .B(II24194), .Z(II24196) ) ;
NAND2   gate22790  (.A(g6568), .B(g14102), .Z(II24205) ) ;
NAND2   gate22791  (.A(g6568), .B(II24205), .Z(II24206) ) ;
NAND2   gate22792  (.A(g14102), .B(II24205), .Z(II24207) ) ;
NAND2   gate22793  (.A(g14033), .B(g9711), .Z(II24213) ) ;
NAND2   gate22794  (.A(g14033), .B(II24213), .Z(II24214) ) ;
NAND2   gate22795  (.A(g9711), .B(II24213), .Z(II24215) ) ;
NAND2   gate22796  (.A(g6427), .B(g14316), .Z(II24226) ) ;
NAND2   gate22797  (.A(g6427), .B(II24226), .Z(II24227) ) ;
NAND2   gate22798  (.A(g14316), .B(II24226), .Z(II24228) ) ;
NAND2   gate22799  (.A(g14222), .B(g9613), .Z(II24234) ) ;
NAND2   gate22800  (.A(g14222), .B(II24234), .Z(II24235) ) ;
NAND2   gate22801  (.A(g9613), .B(II24234), .Z(II24236) ) ;
NAND2   gate22802  (.A(g7329), .B(g14520), .Z(II24251) ) ;
NAND2   gate22803  (.A(g7329), .B(II24251), .Z(II24252) ) ;
NAND2   gate22804  (.A(g14520), .B(II24251), .Z(II24253) ) ;
NAND2   gate22805  (.A(g14342), .B(g9232), .Z(II24263) ) ;
NAND2   gate22806  (.A(g14342), .B(II24263), .Z(II24264) ) ;
NAND2   gate22807  (.A(g9232), .B(II24263), .Z(II24265) ) ;
NAND2   gate22808  (.A(g6180), .B(g13922), .Z(II24271) ) ;
NAND2   gate22809  (.A(g6180), .B(II24271), .Z(II24272) ) ;
NAND2   gate22810  (.A(g13922), .B(II24271), .Z(II24273) ) ;
NAND2   gate22811  (.A(g6284), .B(g13918), .Z(II24278) ) ;
NAND2   gate22812  (.A(g6284), .B(II24278), .Z(II24279) ) ;
NAND2   gate22813  (.A(g13918), .B(II24278), .Z(II24280) ) ;
NAND2   gate22814  (.A(g13895), .B(g9203), .Z(II24290) ) ;
NAND2   gate22815  (.A(g13895), .B(II24290), .Z(II24291) ) ;
NAND2   gate22816  (.A(g9203), .B(II24290), .Z(II24292) ) ;
NAND2   gate22817  (.A(g6209), .B(g14028), .Z(II24298) ) ;
NAND2   gate22818  (.A(g6209), .B(II24298), .Z(II24299) ) ;
NAND2   gate22819  (.A(g14028), .B(II24298), .Z(II24300) ) ;
NAND2   gate22820  (.A(g13983), .B(g15274), .Z(II24306) ) ;
NAND2   gate22821  (.A(g13983), .B(II24306), .Z(II24307) ) ;
NAND2   gate22822  (.A(g15274), .B(II24306), .Z(II24308) ) ;
NAND2   gate22823  (.A(g6832), .B(g14217), .Z(II24317) ) ;
NAND2   gate22824  (.A(g6832), .B(II24317), .Z(II24318) ) ;
NAND2   gate22825  (.A(g14217), .B(II24317), .Z(II24319) ) ;
NAND2   gate22826  (.A(g14124), .B(g9857), .Z(II24325) ) ;
NAND2   gate22827  (.A(g14124), .B(II24325), .Z(II24326) ) ;
NAND2   gate22828  (.A(g9857), .B(II24325), .Z(II24327) ) ;
NAND2   gate22829  (.A(g6632), .B(g14438), .Z(II24338) ) ;
NAND2   gate22830  (.A(g6632), .B(II24338), .Z(II24339) ) ;
NAND2   gate22831  (.A(g14438), .B(II24338), .Z(II24340) ) ;
NAND2   gate22832  (.A(g14238), .B(g9356), .Z(II24351) ) ;
NAND2   gate22833  (.A(g14238), .B(II24351), .Z(II24352) ) ;
NAND2   gate22834  (.A(g9356), .B(II24351), .Z(II24353) ) ;
NAND2   gate22835  (.A(g6157), .B(g14525), .Z(II24361) ) ;
NAND2   gate22836  (.A(g6157), .B(II24361), .Z(II24362) ) ;
NAND2   gate22837  (.A(g14525), .B(II24361), .Z(II24363) ) ;
NAND2   gate22838  (.A(g14454), .B(g9310), .Z(II24372) ) ;
NAND2   gate22839  (.A(g14454), .B(II24372), .Z(II24373) ) ;
NAND2   gate22840  (.A(g9310), .B(II24372), .Z(II24374) ) ;
NAND2   gate22841  (.A(g6212), .B(g13978), .Z(II24380) ) ;
NAND2   gate22842  (.A(g6212), .B(II24380), .Z(II24381) ) ;
NAND2   gate22843  (.A(g13978), .B(II24380), .Z(II24382) ) ;
NAND2   gate22844  (.A(g6421), .B(g13974), .Z(II24387) ) ;
NAND2   gate22845  (.A(g6421), .B(II24387), .Z(II24388) ) ;
NAND2   gate22846  (.A(g13974), .B(II24387), .Z(II24389) ) ;
NAND2   gate22847  (.A(g13936), .B(g9264), .Z(II24399) ) ;
NAND2   gate22848  (.A(g13936), .B(II24399), .Z(II24400) ) ;
NAND2   gate22849  (.A(g9264), .B(II24399), .Z(II24401) ) ;
NAND2   gate22850  (.A(g6298), .B(g14119), .Z(II24407) ) ;
NAND2   gate22851  (.A(g6298), .B(II24407), .Z(II24408) ) ;
NAND2   gate22852  (.A(g14119), .B(II24407), .Z(II24409) ) ;
NAND2   gate22853  (.A(g14053), .B(g15366), .Z(II24415) ) ;
NAND2   gate22854  (.A(g14053), .B(II24415), .Z(II24416) ) ;
NAND2   gate22855  (.A(g15366), .B(II24415), .Z(II24417) ) ;
NAND2   gate22856  (.A(g7134), .B(g14332), .Z(II24426) ) ;
NAND2   gate22857  (.A(g7134), .B(II24426), .Z(II24427) ) ;
NAND2   gate22858  (.A(g14332), .B(II24426), .Z(II24428) ) ;
NAND2   gate22859  (.A(g14153), .B(g15022), .Z(II24436) ) ;
NAND2   gate22860  (.A(g14153), .B(II24436), .Z(II24437) ) ;
NAND2   gate22861  (.A(g15022), .B(II24436), .Z(II24438) ) ;
NAND2   gate22862  (.A(g14148), .B(g9507), .Z(II24443) ) ;
NAND2   gate22863  (.A(g14148), .B(II24443), .Z(II24444) ) ;
NAND2   gate22864  (.A(g9507), .B(II24443), .Z(II24445) ) ;
NAND2   gate22865  (.A(g6142), .B(g14450), .Z(II24452) ) ;
NAND2   gate22866  (.A(g6142), .B(II24452), .Z(II24453) ) ;
NAND2   gate22867  (.A(g14450), .B(II24452), .Z(II24454) ) ;
NAND2   gate22868  (.A(g14360), .B(g9453), .Z(II24464) ) ;
NAND2   gate22869  (.A(g14360), .B(II24464), .Z(II24465) ) ;
NAND2   gate22870  (.A(g9453), .B(II24464), .Z(II24466) ) ;
NAND2   gate22871  (.A(g6184), .B(g14580), .Z(II24474) ) ;
NAND2   gate22872  (.A(g6184), .B(II24474), .Z(II24475) ) ;
NAND2   gate22873  (.A(g14580), .B(II24474), .Z(II24476) ) ;
NAND2   gate22874  (.A(g14541), .B(g9391), .Z(II24485) ) ;
NAND2   gate22875  (.A(g14541), .B(II24485), .Z(II24486) ) ;
NAND2   gate22876  (.A(g9391), .B(II24485), .Z(II24487) ) ;
NAND2   gate22877  (.A(g6301), .B(g14048), .Z(II24493) ) ;
NAND2   gate22878  (.A(g6301), .B(II24493), .Z(II24494) ) ;
NAND2   gate22879  (.A(g14048), .B(II24493), .Z(II24495) ) ;
NAND2   gate22880  (.A(g6626), .B(g14044), .Z(II24500) ) ;
NAND2   gate22881  (.A(g6626), .B(II24500), .Z(II24501) ) ;
NAND2   gate22882  (.A(g14044), .B(II24500), .Z(II24502) ) ;
NAND2   gate22883  (.A(g13992), .B(g9342), .Z(II24512) ) ;
NAND2   gate22884  (.A(g13992), .B(II24512), .Z(II24513) ) ;
NAND2   gate22885  (.A(g9342), .B(II24512), .Z(II24514) ) ;
NAND2   gate22886  (.A(g6435), .B(g14234), .Z(II24520) ) ;
NAND2   gate22887  (.A(g6435), .B(II24520), .Z(II24521) ) ;
NAND2   gate22888  (.A(g14234), .B(II24520), .Z(II24522) ) ;
NAND2   gate22889  (.A(g6707), .B(g14355), .Z(II24530) ) ;
NAND2   gate22890  (.A(g6707), .B(II24530), .Z(II24531) ) ;
NAND2   gate22891  (.A(g14355), .B(II24530), .Z(II24532) ) ;
NAND2   gate22892  (.A(g14268), .B(g15118), .Z(II24537) ) ;
NAND2   gate22893  (.A(g14268), .B(II24537), .Z(II24538) ) ;
NAND2   gate22894  (.A(g15118), .B(II24537), .Z(II24539) ) ;
NAND2   gate22895  (.A(g14263), .B(g9649), .Z(II24544) ) ;
NAND2   gate22896  (.A(g14263), .B(II24544), .Z(II24545) ) ;
NAND2   gate22897  (.A(g9649), .B(II24544), .Z(II24546) ) ;
NAND2   gate22898  (.A(g6163), .B(g14537), .Z(II24553) ) ;
NAND2   gate22899  (.A(g6163), .B(II24553), .Z(II24554) ) ;
NAND2   gate22900  (.A(g14537), .B(II24553), .Z(II24555) ) ;
NAND2   gate22901  (.A(g14472), .B(g9595), .Z(II24565) ) ;
NAND2   gate22902  (.A(g14472), .B(II24565), .Z(II24566) ) ;
NAND2   gate22903  (.A(g9595), .B(II24565), .Z(II24567) ) ;
NAND2   gate22904  (.A(g6216), .B(g14614), .Z(II24575) ) ;
NAND2   gate22905  (.A(g6216), .B(II24575), .Z(II24576) ) ;
NAND2   gate22906  (.A(g14614), .B(II24575), .Z(II24577) ) ;
NAND2   gate22907  (.A(g14596), .B(g9488), .Z(II24586) ) ;
NAND2   gate22908  (.A(g14596), .B(II24586), .Z(II24587) ) ;
NAND2   gate22909  (.A(g9488), .B(II24586), .Z(II24588) ) ;
NAND2   gate22910  (.A(g6438), .B(g14139), .Z(II24594) ) ;
NAND2   gate22911  (.A(g6438), .B(II24594), .Z(II24595) ) ;
NAND2   gate22912  (.A(g14139), .B(II24594), .Z(II24596) ) ;
NAND2   gate22913  (.A(g6890), .B(g14135), .Z(II24601) ) ;
NAND2   gate22914  (.A(g6890), .B(II24601), .Z(II24602) ) ;
NAND2   gate22915  (.A(g14135), .B(II24601), .Z(II24603) ) ;
NAND2   gate22916  (.A(g15814), .B(g15978), .Z(II24611) ) ;
NAND2   gate22917  (.A(g15814), .B(II24611), .Z(II24612) ) ;
NAND2   gate22918  (.A(g15978), .B(II24611), .Z(II24613) ) ;
NAND2   gate22919  (.A(g6136), .B(g14252), .Z(II24624) ) ;
NAND2   gate22920  (.A(g6136), .B(II24624), .Z(II24625) ) ;
NAND2   gate22921  (.A(g14252), .B(II24624), .Z(II24626) ) ;
NAND2   gate22922  (.A(g7009), .B(g14467), .Z(II24632) ) ;
NAND2   gate22923  (.A(g7009), .B(II24632), .Z(II24633) ) ;
NAND2   gate22924  (.A(g14467), .B(II24632), .Z(II24634) ) ;
NAND2   gate22925  (.A(g14390), .B(g15210), .Z(II24639) ) ;
NAND2   gate22926  (.A(g14390), .B(II24639), .Z(II24640) ) ;
NAND2   gate22927  (.A(g15210), .B(II24639), .Z(II24641) ) ;
NAND2   gate22928  (.A(g14385), .B(g9795), .Z(II24646) ) ;
NAND2   gate22929  (.A(g14385), .B(II24646), .Z(II24647) ) ;
NAND2   gate22930  (.A(g9795), .B(II24646), .Z(II24648) ) ;
NAND2   gate22931  (.A(g6190), .B(g14592), .Z(II24655) ) ;
NAND2   gate22932  (.A(g6190), .B(II24655), .Z(II24656) ) ;
NAND2   gate22933  (.A(g14592), .B(II24655), .Z(II24657) ) ;
NAND2   gate22934  (.A(g14559), .B(g9737), .Z(II24667) ) ;
NAND2   gate22935  (.A(g14559), .B(II24667), .Z(II24668) ) ;
NAND2   gate22936  (.A(g9737), .B(II24667), .Z(II24669) ) ;
NAND2   gate22937  (.A(g6305), .B(g14637), .Z(II24677) ) ;
NAND2   gate22938  (.A(g6305), .B(II24677), .Z(II24678) ) ;
NAND2   gate22939  (.A(g14637), .B(II24677), .Z(II24679) ) ;
NAND2   gate22940  (.A(g6146), .B(g14374), .Z(II24694) ) ;
NAND2   gate22941  (.A(g6146), .B(II24694), .Z(II24695) ) ;
NAND2   gate22942  (.A(g14374), .B(II24694), .Z(II24696) ) ;
NAND2   gate22943  (.A(g7259), .B(g14554), .Z(II24702) ) ;
NAND2   gate22944  (.A(g7259), .B(II24702), .Z(II24703) ) ;
NAND2   gate22945  (.A(g14554), .B(II24702), .Z(II24704) ) ;
NAND2   gate22946  (.A(g14502), .B(g15296), .Z(II24709) ) ;
NAND2   gate22947  (.A(g14502), .B(II24709), .Z(II24710) ) ;
NAND2   gate22948  (.A(g15296), .B(II24709), .Z(II24711) ) ;
NAND2   gate22949  (.A(g14497), .B(g9941), .Z(II24716) ) ;
NAND2   gate22950  (.A(g14497), .B(II24716), .Z(II24717) ) ;
NAND2   gate22951  (.A(g9941), .B(II24716), .Z(II24718) ) ;
NAND2   gate22952  (.A(g6222), .B(g14626), .Z(II24725) ) ;
NAND2   gate22953  (.A(g6222), .B(II24725), .Z(II24726) ) ;
NAND2   gate22954  (.A(g14626), .B(II24725), .Z(II24727) ) ;
NAND2   gate22955  (.A(g6167), .B(g14486), .Z(II24743) ) ;
NAND2   gate22956  (.A(g6167), .B(II24743), .Z(II24744) ) ;
NAND2   gate22957  (.A(g14486), .B(II24743), .Z(II24745) ) ;
NAND2   gate22958  (.A(g7455), .B(g14609), .Z(II24751) ) ;
NAND2   gate22959  (.A(g7455), .B(II24751), .Z(II24752) ) ;
NAND2   gate22960  (.A(g14609), .B(II24751), .Z(II24753) ) ;
NAND2   gate22961  (.A(g6194), .B(g14573), .Z(II24763) ) ;
NAND2   gate22962  (.A(g6194), .B(II24763), .Z(II24764) ) ;
NAND2   gate22963  (.A(g14573), .B(II24763), .Z(II24765) ) ;
NAND2   gate22964  (.A(g8029), .B(g13507), .Z(II25030) ) ;
NAND2   gate22965  (.A(g8029), .B(II25030), .Z(II25031) ) ;
NAND2   gate22966  (.A(g13507), .B(II25030), .Z(II25032) ) ;
NAND2   gate22967  (.A(g52), .B(g18179), .Z(II25532) ) ;
NAND2   gate22968  (.A(g52), .B(II25532), .Z(II25533) ) ;
NAND2   gate22969  (.A(g18179), .B(II25532), .Z(II25534) ) ;
NAND2   gate22970  (.A(g92), .B(g18174), .Z(II25539) ) ;
NAND2   gate22971  (.A(g92), .B(II25539), .Z(II25540) ) ;
NAND2   gate22972  (.A(g18174), .B(II25539), .Z(II25541) ) ;
NAND2   gate22973  (.A(g56), .B(g17724), .Z(II25560) ) ;
NAND2   gate22974  (.A(g56), .B(II25560), .Z(II25561) ) ;
NAND2   gate22975  (.A(g17724), .B(II25560), .Z(II25562) ) ;
NAND2   gate22976  (.A(g740), .B(g18286), .Z(II25571) ) ;
NAND2   gate22977  (.A(g740), .B(II25571), .Z(II25572) ) ;
NAND2   gate22978  (.A(g18286), .B(II25571), .Z(II25573) ) ;
NAND2   gate22979  (.A(g780), .B(g18281), .Z(II25578) ) ;
NAND2   gate22980  (.A(g780), .B(II25578), .Z(II25579) ) ;
NAND2   gate22981  (.A(g18281), .B(II25578), .Z(II25580) ) ;
NAND2   gate22982  (.A(g61), .B(g18074), .Z(II25595) ) ;
NAND2   gate22983  (.A(g61), .B(II25595), .Z(II25596) ) ;
NAND2   gate22984  (.A(g18074), .B(II25595), .Z(II25597) ) ;
NAND2   gate22985  (.A(g744), .B(g17825), .Z(II25605) ) ;
NAND2   gate22986  (.A(g744), .B(II25605), .Z(II25606) ) ;
NAND2   gate22987  (.A(g17825), .B(II25605), .Z(II25607) ) ;
NAND2   gate22988  (.A(g1426), .B(g18379), .Z(II25616) ) ;
NAND2   gate22989  (.A(g1426), .B(II25616), .Z(II25617) ) ;
NAND2   gate22990  (.A(g18379), .B(II25616), .Z(II25618) ) ;
NAND2   gate22991  (.A(g1466), .B(g18374), .Z(II25623) ) ;
NAND2   gate22992  (.A(g1466), .B(II25623), .Z(II25624) ) ;
NAND2   gate22993  (.A(g18374), .B(II25623), .Z(II25625) ) ;
NAND2   gate22994  (.A(g65), .B(g17640), .Z(II25633) ) ;
NAND2   gate22995  (.A(g65), .B(II25633), .Z(II25634) ) ;
NAND2   gate22996  (.A(g17640), .B(II25633), .Z(II25635) ) ;
NAND2   gate22997  (.A(g749), .B(g18190), .Z(II25643) ) ;
NAND2   gate22998  (.A(g749), .B(II25643), .Z(II25644) ) ;
NAND2   gate22999  (.A(g18190), .B(II25643), .Z(II25645) ) ;
NAND2   gate23000  (.A(g1430), .B(g17937), .Z(II25653) ) ;
NAND2   gate23001  (.A(g1430), .B(II25653), .Z(II25654) ) ;
NAND2   gate23002  (.A(g17937), .B(II25653), .Z(II25655) ) ;
NAND2   gate23003  (.A(g2120), .B(g18474), .Z(II25664) ) ;
NAND2   gate23004  (.A(g2120), .B(II25664), .Z(II25665) ) ;
NAND2   gate23005  (.A(g18474), .B(II25664), .Z(II25666) ) ;
NAND2   gate23006  (.A(g2160), .B(g18469), .Z(II25671) ) ;
NAND2   gate23007  (.A(g2160), .B(II25671), .Z(II25672) ) ;
NAND2   gate23008  (.A(g18469), .B(II25671), .Z(II25673) ) ;
NAND2   gate23009  (.A(g70), .B(g17974), .Z(II25681) ) ;
NAND2   gate23010  (.A(g70), .B(II25681), .Z(II25682) ) ;
NAND2   gate23011  (.A(g17974), .B(II25681), .Z(II25683) ) ;
NAND2   gate23012  (.A(g753), .B(g17741), .Z(II25690) ) ;
NAND2   gate23013  (.A(g753), .B(II25690), .Z(II25691) ) ;
NAND2   gate23014  (.A(g17741), .B(II25690), .Z(II25692) ) ;
NAND2   gate23015  (.A(g1435), .B(g18297), .Z(II25700) ) ;
NAND2   gate23016  (.A(g1435), .B(II25700), .Z(II25701) ) ;
NAND2   gate23017  (.A(g18297), .B(II25700), .Z(II25702) ) ;
NAND2   gate23018  (.A(g2124), .B(g18048), .Z(II25710) ) ;
NAND2   gate23019  (.A(g2124), .B(II25710), .Z(II25711) ) ;
NAND2   gate23020  (.A(g18048), .B(II25710), .Z(II25712) ) ;
NAND2   gate23021  (.A(g74), .B(g18341), .Z(II25721) ) ;
NAND2   gate23022  (.A(g74), .B(II25721), .Z(II25722) ) ;
NAND2   gate23023  (.A(g18341), .B(II25721), .Z(II25723) ) ;
NAND2   gate23024  (.A(g758), .B(g18091), .Z(II25731) ) ;
NAND2   gate23025  (.A(g758), .B(II25731), .Z(II25732) ) ;
NAND2   gate23026  (.A(g18091), .B(II25731), .Z(II25733) ) ;
NAND2   gate23027  (.A(g1439), .B(g17842), .Z(II25740) ) ;
NAND2   gate23028  (.A(g1439), .B(II25740), .Z(II25741) ) ;
NAND2   gate23029  (.A(g17842), .B(II25740), .Z(II25742) ) ;
NAND2   gate23030  (.A(g2129), .B(g18390), .Z(II25750) ) ;
NAND2   gate23031  (.A(g2129), .B(II25750), .Z(II25751) ) ;
NAND2   gate23032  (.A(g18390), .B(II25750), .Z(II25752) ) ;
NAND2   gate23033  (.A(g79), .B(g17882), .Z(II25761) ) ;
NAND2   gate23034  (.A(g79), .B(II25761), .Z(II25762) ) ;
NAND2   gate23035  (.A(g17882), .B(II25761), .Z(II25763) ) ;
NAND2   gate23036  (.A(g762), .B(g18436), .Z(II25771) ) ;
NAND2   gate23037  (.A(g762), .B(II25771), .Z(II25772) ) ;
NAND2   gate23038  (.A(g18436), .B(II25771), .Z(II25773) ) ;
NAND2   gate23039  (.A(g1444), .B(g18207), .Z(II25781) ) ;
NAND2   gate23040  (.A(g1444), .B(II25781), .Z(II25782) ) ;
NAND2   gate23041  (.A(g18207), .B(II25781), .Z(II25783) ) ;
NAND2   gate23042  (.A(g2133), .B(g17954), .Z(II25790) ) ;
NAND2   gate23043  (.A(g2133), .B(II25790), .Z(II25791) ) ;
NAND2   gate23044  (.A(g17954), .B(II25790), .Z(II25792) ) ;
NAND2   gate23045  (.A(g83), .B(g18265), .Z(II25800) ) ;
NAND2   gate23046  (.A(g83), .B(II25800), .Z(II25801) ) ;
NAND2   gate23047  (.A(g18265), .B(II25800), .Z(II25802) ) ;
NAND2   gate23048  (.A(g767), .B(g17993), .Z(II25809) ) ;
NAND2   gate23049  (.A(g767), .B(II25809), .Z(II25810) ) ;
NAND2   gate23050  (.A(g17993), .B(II25809), .Z(II25811) ) ;
NAND2   gate23051  (.A(g1448), .B(g18509), .Z(II25819) ) ;
NAND2   gate23052  (.A(g1448), .B(II25819), .Z(II25820) ) ;
NAND2   gate23053  (.A(g18509), .B(II25819), .Z(II25821) ) ;
NAND2   gate23054  (.A(g2138), .B(g18314), .Z(II25829) ) ;
NAND2   gate23055  (.A(g2138), .B(II25829), .Z(II25830) ) ;
NAND2   gate23056  (.A(g18314), .B(II25829), .Z(II25831) ) ;
NAND2   gate23057  (.A(g88), .B(g17802), .Z(II25838) ) ;
NAND2   gate23058  (.A(g88), .B(II25838), .Z(II25839) ) ;
NAND2   gate23059  (.A(g17802), .B(II25838), .Z(II25840) ) ;
NAND2   gate23060  (.A(g771), .B(g18358), .Z(II25846) ) ;
NAND2   gate23061  (.A(g771), .B(II25846), .Z(II25847) ) ;
NAND2   gate23062  (.A(g18358), .B(II25846), .Z(II25848) ) ;
NAND2   gate23063  (.A(g1453), .B(g18110), .Z(II25855) ) ;
NAND2   gate23064  (.A(g1453), .B(II25855), .Z(II25856) ) ;
NAND2   gate23065  (.A(g18110), .B(II25855), .Z(II25857) ) ;
NAND2   gate23066  (.A(g2142), .B(g18573), .Z(II25865) ) ;
NAND2   gate23067  (.A(g2142), .B(II25865), .Z(II25866) ) ;
NAND2   gate23068  (.A(g18573), .B(II25865), .Z(II25867) ) ;
NAND2   gate23069  (.A(g776), .B(g17914), .Z(II25880) ) ;
NAND2   gate23070  (.A(g776), .B(II25880), .Z(II25881) ) ;
NAND2   gate23071  (.A(g17914), .B(II25880), .Z(II25882) ) ;
NAND2   gate23072  (.A(g1457), .B(g18453), .Z(II25888) ) ;
NAND2   gate23073  (.A(g1457), .B(II25888), .Z(II25889) ) ;
NAND2   gate23074  (.A(g18453), .B(II25888), .Z(II25890) ) ;
NAND2   gate23075  (.A(g2147), .B(g18226), .Z(II25897) ) ;
NAND2   gate23076  (.A(g2147), .B(II25897), .Z(II25898) ) ;
NAND2   gate23077  (.A(g18226), .B(II25897), .Z(II25899) ) ;
NAND2   gate23078  (.A(g1462), .B(g18025), .Z(II25913) ) ;
NAND2   gate23079  (.A(g1462), .B(II25913), .Z(II25914) ) ;
NAND2   gate23080  (.A(g18025), .B(II25913), .Z(II25915) ) ;
NAND2   gate23081  (.A(g2151), .B(g18526), .Z(II25921) ) ;
NAND2   gate23082  (.A(g2151), .B(II25921), .Z(II25922) ) ;
NAND2   gate23083  (.A(g18526), .B(II25921), .Z(II25923) ) ;
NAND2   gate23084  (.A(g2156), .B(g18142), .Z(II25938) ) ;
NAND2   gate23085  (.A(g2156), .B(II25938), .Z(II25939) ) ;
NAND2   gate23086  (.A(g18142), .B(II25938), .Z(II25940) ) ;
NOR2    gate23087  (.A(g18165), .B(g15753), .Z(g19219) ) ;
NAND2   gate23088  (.A(g14079), .B(g19444), .Z(II28189) ) ;
NAND2   gate23089  (.A(g14079), .B(II28189), .Z(II28190) ) ;
NAND2   gate23090  (.A(g19444), .B(II28189), .Z(II28191) ) ;
NAND2   gate23091  (.A(II28190), .B(II28191), .Z(g21660) ) ;
NAND2   gate23092  (.A(g14194), .B(g19471), .Z(II28217) ) ;
NAND2   gate23093  (.A(g14194), .B(II28217), .Z(II28218) ) ;
NAND2   gate23094  (.A(g19471), .B(II28217), .Z(II28219) ) ;
NAND2   gate23095  (.A(II28218), .B(II28219), .Z(g21689) ) ;
NAND2   gate23096  (.A(g14309), .B(g19494), .Z(II28247) ) ;
NAND2   gate23097  (.A(g14309), .B(II28247), .Z(II28248) ) ;
NAND2   gate23098  (.A(g19494), .B(II28247), .Z(II28249) ) ;
NAND2   gate23099  (.A(II28248), .B(II28249), .Z(g21725) ) ;
NAND2   gate23100  (.A(g14431), .B(g19515), .Z(II28271) ) ;
NAND2   gate23101  (.A(g14431), .B(II28271), .Z(II28272) ) ;
NAND2   gate23102  (.A(g19515), .B(II28271), .Z(II28273) ) ;
NAND2   gate23103  (.A(II28272), .B(II28273), .Z(g21751) ) ;
NAND3   gate23104  (.A(g17807), .B(g19181), .C(g19186), .Z(g21848) ) ;
NAND3   gate23105  (.A(g17979), .B(g19187), .C(g19191), .Z(g21850) ) ;
NAND3   gate23106  (.A(g17919), .B(g19188), .C(g19193), .Z(g21855) ) ;
NAND3   gate23107  (.A(g18079), .B(g19192), .C(g19200), .Z(g21857) ) ;
NAND3   gate23108  (.A(g18096), .B(g19194), .C(g19202), .Z(g21858) ) ;
NAND3   gate23109  (.A(g18030), .B(g19195), .C(g19204), .Z(g21859) ) ;
NAND3   gate23110  (.A(g18270), .B(g19201), .C(g19209), .Z(g21860) ) ;
NAND3   gate23111  (.A(g18195), .B(g19203), .C(g19211), .Z(g21862) ) ;
NAND3   gate23112  (.A(g18212), .B(g19205), .C(g19213), .Z(g21863) ) ;
NAND3   gate23113  (.A(g18147), .B(g19206), .C(g19215), .Z(g21864) ) ;
NAND3   gate23114  (.A(g18424), .B(g19210), .C(g19221), .Z(g21865) ) ;
NAND3   gate23115  (.A(g18363), .B(g19212), .C(g19222), .Z(g21866) ) ;
NAND3   gate23116  (.A(g18302), .B(g19214), .C(g19224), .Z(g21868) ) ;
NAND3   gate23117  (.A(g18319), .B(g19216), .C(g19226), .Z(g21869) ) ;
NAND3   gate23118  (.A(g18497), .B(g19223), .C(g19231), .Z(g21870) ) ;
NAND3   gate23119  (.A(g18458), .B(g19225), .C(g19232), .Z(g21871) ) ;
NAND3   gate23120  (.A(g18395), .B(g19227), .C(g19234), .Z(g21873) ) ;
NAND3   gate23121  (.A(g18561), .B(g19233), .C(g19244), .Z(g21874) ) ;
NAND3   gate23122  (.A(g18531), .B(g19235), .C(g19245), .Z(g21875) ) ;
NAND3   gate23123  (.A(g18611), .B(g19246), .C(g19257), .Z(g21877) ) ;
NAND3   gate23124  (.A(g18419), .B(g19250), .C(g19263), .Z(g21879) ) ;
NAND3   gate23125  (.A(g18492), .B(g19264), .C(g19278), .Z(g21881) ) ;
NAND3   gate23126  (.A(g18556), .B(g19279), .C(g19297), .Z(g21885) ) ;
NAND3   gate23127  (.A(g18606), .B(g19298), .C(g19315), .Z(g21888) ) ;
NOR2    gate23128  (.A(g19889), .B(g18062), .Z(g21048) ) ;
NOR2    gate23129  (.A(g19914), .B(g18169), .Z(g21065) ) ;
NOR2    gate23130  (.A(g13519), .B(g19289), .Z(g21887) ) ;
NAND2   gate23131  (.A(g21887), .B(g13519), .Z(II28726) ) ;
NAND2   gate23132  (.A(g21887), .B(II28726), .Z(II28727) ) ;
NAND2   gate23133  (.A(g13519), .B(II28726), .Z(II28728) ) ;
NOR2    gate23134  (.A(g13530), .B(g19307), .Z(g21890) ) ;
NAND2   gate23135  (.A(g21890), .B(g13530), .Z(II28741) ) ;
NAND2   gate23136  (.A(g21890), .B(II28741), .Z(II28742) ) ;
NAND2   gate23137  (.A(g13530), .B(II28741), .Z(II28743) ) ;
NOR2    gate23138  (.A(g13541), .B(g19328), .Z(g21893) ) ;
NAND2   gate23139  (.A(g21893), .B(g13541), .Z(II28753) ) ;
NAND2   gate23140  (.A(g21893), .B(II28753), .Z(II28754) ) ;
NAND2   gate23141  (.A(g13541), .B(II28753), .Z(II28755) ) ;
NOR2    gate23142  (.A(g13552), .B(g19355), .Z(g21901) ) ;
NAND2   gate23143  (.A(g21901), .B(g13552), .Z(II28765) ) ;
NAND2   gate23144  (.A(g21901), .B(II28765), .Z(II28766) ) ;
NAND2   gate23145  (.A(g13552), .B(II28765), .Z(II28767) ) ;
NOR2    gate23146  (.A(g19240), .B(g19230), .Z(g21211) ) ;
NOR2    gate23147  (.A(g19253), .B(g19243), .Z(g21219) ) ;
NOR2    gate23148  (.A(g19266), .B(g19256), .Z(g21230) ) ;
NOR2    gate23149  (.A(g19281), .B(g19269), .Z(g21235) ) ;
NAND3   gate23150  (.A(g21850), .B(g21848), .C(g21879), .Z(g22809) ) ;
NAND3   gate23151  (.A(g21865), .B(g21860), .C(g21857), .Z(g22844) ) ;
NAND2   gate23152  (.A(g8278), .B(g21660), .Z(g22846) ) ;
NAND3   gate23153  (.A(g21858), .B(g21855), .C(g21881), .Z(g22850) ) ;
NAND3   gate23154  (.A(g21870), .B(g21866), .C(g21862), .Z(g22879) ) ;
NAND2   gate23155  (.A(g8287), .B(g21689), .Z(g22881) ) ;
NAND3   gate23156  (.A(g21863), .B(g21859), .C(g21885), .Z(g22885) ) ;
NAND3   gate23157  (.A(g21874), .B(g21871), .C(g21868), .Z(g22914) ) ;
NAND2   gate23158  (.A(g8296), .B(g21725), .Z(g22916) ) ;
NAND3   gate23159  (.A(g21869), .B(g21864), .C(g21888), .Z(g22920) ) ;
NAND3   gate23160  (.A(g21877), .B(g21875), .C(g21873), .Z(g22939) ) ;
NAND2   gate23161  (.A(g8305), .B(g21751), .Z(g22941) ) ;
NOR3    gate23162  (.A(g21138), .B(g19303), .C(g19320), .Z(g23066) ) ;
NOR2    gate23163  (.A(g21121), .B(g21153), .Z(g23051) ) ;
NOR3    gate23164  (.A(g21158), .B(g19324), .C(g19347), .Z(g23080) ) ;
NOR2    gate23165  (.A(g21140), .B(g21173), .Z(g23070) ) ;
NOR2    gate23166  (.A(g21085), .B(g19241), .Z(g22999) ) ;
NOR2    gate23167  (.A(g19868), .B(g21593), .Z(g22174) ) ;
NOR3    gate23168  (.A(g21178), .B(g19351), .C(g19381), .Z(g23096) ) ;
NOR2    gate23169  (.A(g21160), .B(g21193), .Z(g23083) ) ;
NOR2    gate23170  (.A(g21097), .B(g19254), .Z(g23013) ) ;
NOR2    gate23171  (.A(g19899), .B(g21622), .Z(g22189) ) ;
NOR3    gate23172  (.A(g21198), .B(g19385), .C(g19413), .Z(g23113) ) ;
NOR2    gate23173  (.A(g21180), .B(g21208), .Z(g23099) ) ;
NOR2    gate23174  (.A(g21111), .B(g19267), .Z(g23029) ) ;
NOR2    gate23175  (.A(g19924), .B(g21650), .Z(g22198) ) ;
NOR2    gate23176  (.A(g21128), .B(g19282), .Z(g23046) ) ;
NOR2    gate23177  (.A(g19939), .B(g21681), .Z(g22204) ) ;
NOR3    gate23178  (.A(g21252), .B(g19531), .C(g19540), .Z(g21980) ) ;
NOR2    gate23179  (.A(g21245), .B(g21259), .Z(g21975) ) ;
NOR3    gate23180  (.A(g21260), .B(g19541), .C(g19544), .Z(g21987) ) ;
NOR2    gate23181  (.A(g21254), .B(g21267), .Z(g21981) ) ;
NOR2    gate23182  (.A(g21229), .B(g19449), .Z(g23135) ) ;
NOR2    gate23183  (.A(g20144), .B(g21805), .Z(g22288) ) ;
NOR3    gate23184  (.A(g21268), .B(g19545), .C(g19547), .Z(g22000) ) ;
NOR2    gate23185  (.A(g21262), .B(g21276), .Z(g21988) ) ;
NAND2   gate23186  (.A(g18435), .B(g22812), .Z(g23376) ) ;
NOR2    gate23187  (.A(g21234), .B(g19476), .Z(g21968) ) ;
NOR2    gate23188  (.A(g20182), .B(g21812), .Z(g22308) ) ;
NOR3    gate23189  (.A(g21277), .B(g19548), .C(g19551), .Z(g22013) ) ;
NOR2    gate23190  (.A(g21270), .B(g21283), .Z(g22001) ) ;
NAND2   gate23191  (.A(g18508), .B(g22852), .Z(g23387) ) ;
NOR2    gate23192  (.A(g21243), .B(g19499), .Z(g21971) ) ;
NOR2    gate23193  (.A(g20216), .B(g21818), .Z(g22336) ) ;
NAND2   gate23194  (.A(g18572), .B(g22887), .Z(g23394) ) ;
NOR2    gate23195  (.A(g21251), .B(g19520), .Z(g21973) ) ;
NOR2    gate23196  (.A(g20246), .B(g21822), .Z(g22361) ) ;
NAND2   gate23197  (.A(g18622), .B(g22922), .Z(g23402) ) ;
NAND2   gate23198  (.A(g22846), .B(g14079), .Z(II30790) ) ;
NAND2   gate23199  (.A(g22846), .B(II30790), .Z(II30791) ) ;
NAND2   gate23200  (.A(g14079), .B(II30790), .Z(II30792) ) ;
NAND2   gate23201  (.A(g22881), .B(g14194), .Z(II30868) ) ;
NAND2   gate23202  (.A(g22881), .B(II30868), .Z(II30869) ) ;
NAND2   gate23203  (.A(g14194), .B(II30868), .Z(II30870) ) ;
NAND2   gate23204  (.A(g22916), .B(g14309), .Z(II30952) ) ;
NAND2   gate23205  (.A(g22916), .B(II30952), .Z(II30953) ) ;
NAND2   gate23206  (.A(g14309), .B(II30952), .Z(II30954) ) ;
NAND2   gate23207  (.A(g22941), .B(g14431), .Z(II31035) ) ;
NAND2   gate23208  (.A(g22941), .B(II31035), .Z(II31036) ) ;
NAND2   gate23209  (.A(g14431), .B(II31035), .Z(II31037) ) ;
NAND2   gate23210  (.A(g22812), .B(g13958), .Z(g23906) ) ;
NAND2   gate23211  (.A(g22812), .B(g13922), .Z(g23936) ) ;
NAND2   gate23212  (.A(g22812), .B(g13918), .Z(g23937) ) ;
NAND2   gate23213  (.A(g22852), .B(g14028), .Z(g23938) ) ;
NAND2   gate23214  (.A(g22812), .B(g14525), .Z(g23953) ) ;
NAND2   gate23215  (.A(g22852), .B(g13978), .Z(g23968) ) ;
NAND2   gate23216  (.A(g22852), .B(g13974), .Z(g23969) ) ;
NAND2   gate23217  (.A(g22887), .B(g14119), .Z(g23970) ) ;
NAND2   gate23218  (.A(g22812), .B(g14450), .Z(g23973) ) ;
NAND2   gate23219  (.A(g22852), .B(g14580), .Z(g23982) ) ;
NAND2   gate23220  (.A(g22887), .B(g14048), .Z(g23997) ) ;
NAND2   gate23221  (.A(g22887), .B(g14044), .Z(g23998) ) ;
NAND2   gate23222  (.A(g22922), .B(g14234), .Z(g23999) ) ;
NAND2   gate23223  (.A(g22812), .B(g14355), .Z(g24002) ) ;
NAND2   gate23224  (.A(g22852), .B(g14537), .Z(g24003) ) ;
NAND2   gate23225  (.A(g22887), .B(g14614), .Z(g24012) ) ;
NAND2   gate23226  (.A(g22922), .B(g14139), .Z(g24027) ) ;
NAND2   gate23227  (.A(g22922), .B(g14135), .Z(g24028) ) ;
NAND2   gate23228  (.A(g22812), .B(g14252), .Z(g24034) ) ;
NAND2   gate23229  (.A(g22852), .B(g14467), .Z(g24036) ) ;
NAND2   gate23230  (.A(g22887), .B(g14592), .Z(g24037) ) ;
NAND2   gate23231  (.A(g22922), .B(g14637), .Z(g24046) ) ;
NAND2   gate23232  (.A(g22812), .B(g14171), .Z(g24052) ) ;
NAND2   gate23233  (.A(g22852), .B(g14374), .Z(g24054) ) ;
NAND2   gate23234  (.A(g22887), .B(g14554), .Z(g24056) ) ;
NAND2   gate23235  (.A(g22922), .B(g14626), .Z(g24057) ) ;
NAND2   gate23236  (.A(g22812), .B(g14086), .Z(g24058) ) ;
NAND2   gate23237  (.A(g22852), .B(g14286), .Z(g24065) ) ;
NAND2   gate23238  (.A(g22887), .B(g14486), .Z(g24067) ) ;
NAND2   gate23239  (.A(g22922), .B(g14609), .Z(g24069) ) ;
NAND2   gate23240  (.A(g22812), .B(g14011), .Z(g24070) ) ;
NAND2   gate23241  (.A(g22852), .B(g14201), .Z(g24071) ) ;
NAND2   gate23242  (.A(g22887), .B(g14408), .Z(g24078) ) ;
NAND2   gate23243  (.A(g22922), .B(g14573), .Z(g24080) ) ;
NAND2   gate23244  (.A(g22852), .B(g14102), .Z(g24081) ) ;
NAND2   gate23245  (.A(g22887), .B(g14316), .Z(g24082) ) ;
NAND2   gate23246  (.A(g22922), .B(g14520), .Z(g24089) ) ;
NAND2   gate23247  (.A(g22887), .B(g14217), .Z(g24090) ) ;
NAND2   gate23248  (.A(g22922), .B(g14438), .Z(g24091) ) ;
NAND2   gate23249  (.A(g22922), .B(g14332), .Z(g24093) ) ;
NAND2   gate23250  (.A(g17903), .B(g23936), .Z(II32265) ) ;
NAND2   gate23251  (.A(g17903), .B(II32265), .Z(II32266) ) ;
NAND2   gate23252  (.A(g23936), .B(II32265), .Z(II32267) ) ;
NAND2   gate23253  (.A(g17815), .B(g23953), .Z(II32284) ) ;
NAND2   gate23254  (.A(g17815), .B(II32284), .Z(II32285) ) ;
NAND2   gate23255  (.A(g23953), .B(II32284), .Z(II32286) ) ;
NAND2   gate23256  (.A(g18014), .B(g23968), .Z(II32295) ) ;
NAND2   gate23257  (.A(g18014), .B(II32295), .Z(II32296) ) ;
NAND2   gate23258  (.A(g23968), .B(II32295), .Z(II32297) ) ;
NAND2   gate23259  (.A(g17903), .B(g23973), .Z(II32308) ) ;
NAND2   gate23260  (.A(g17903), .B(II32308), .Z(II32309) ) ;
NAND2   gate23261  (.A(g23973), .B(II32308), .Z(II32310) ) ;
NAND2   gate23262  (.A(g17927), .B(g23982), .Z(II32323) ) ;
NAND2   gate23263  (.A(g17927), .B(II32323), .Z(II32324) ) ;
NAND2   gate23264  (.A(g23982), .B(II32323), .Z(II32325) ) ;
NAND2   gate23265  (.A(g18131), .B(g23997), .Z(II32333) ) ;
NAND2   gate23266  (.A(g18131), .B(II32333), .Z(II32334) ) ;
NAND2   gate23267  (.A(g23997), .B(II32333), .Z(II32335) ) ;
NAND2   gate23268  (.A(g17815), .B(g24002), .Z(II32345) ) ;
NAND2   gate23269  (.A(g17815), .B(II32345), .Z(II32346) ) ;
NAND2   gate23270  (.A(g24002), .B(II32345), .Z(II32347) ) ;
NAND2   gate23271  (.A(g18014), .B(g24003), .Z(II32355) ) ;
NAND2   gate23272  (.A(g18014), .B(II32355), .Z(II32356) ) ;
NAND2   gate23273  (.A(g24003), .B(II32355), .Z(II32357) ) ;
NAND2   gate23274  (.A(g18038), .B(g24012), .Z(II32368) ) ;
NAND2   gate23275  (.A(g18038), .B(II32368), .Z(II32369) ) ;
NAND2   gate23276  (.A(g24012), .B(II32368), .Z(II32370) ) ;
NAND2   gate23277  (.A(g18247), .B(g24027), .Z(II32378) ) ;
NAND2   gate23278  (.A(g18247), .B(II32378), .Z(II32379) ) ;
NAND2   gate23279  (.A(g24027), .B(II32378), .Z(II32380) ) ;
NAND2   gate23280  (.A(g17903), .B(g24034), .Z(II32391) ) ;
NAND2   gate23281  (.A(g17903), .B(II32391), .Z(II32392) ) ;
NAND2   gate23282  (.A(g24034), .B(II32391), .Z(II32393) ) ;
NAND2   gate23283  (.A(g17927), .B(g24036), .Z(II32400) ) ;
NAND2   gate23284  (.A(g17927), .B(II32400), .Z(II32401) ) ;
NAND2   gate23285  (.A(g24036), .B(II32400), .Z(II32402) ) ;
NAND2   gate23286  (.A(g18131), .B(g24037), .Z(II32409) ) ;
NAND2   gate23287  (.A(g18131), .B(II32409), .Z(II32410) ) ;
NAND2   gate23288  (.A(g24037), .B(II32409), .Z(II32411) ) ;
NAND2   gate23289  (.A(g18155), .B(g24046), .Z(II32422) ) ;
NAND2   gate23290  (.A(g18155), .B(II32422), .Z(II32423) ) ;
NAND2   gate23291  (.A(g24046), .B(II32422), .Z(II32424) ) ;
NAND2   gate23292  (.A(g17815), .B(g24052), .Z(II32430) ) ;
NAND2   gate23293  (.A(g17815), .B(II32430), .Z(II32431) ) ;
NAND2   gate23294  (.A(g24052), .B(II32430), .Z(II32432) ) ;
NAND2   gate23295  (.A(g18014), .B(g24054), .Z(II32443) ) ;
NAND2   gate23296  (.A(g18014), .B(II32443), .Z(II32444) ) ;
NAND2   gate23297  (.A(g24054), .B(II32443), .Z(II32445) ) ;
NAND2   gate23298  (.A(g18038), .B(g24056), .Z(II32451) ) ;
NAND2   gate23299  (.A(g18038), .B(II32451), .Z(II32452) ) ;
NAND2   gate23300  (.A(g24056), .B(II32451), .Z(II32453) ) ;
NAND2   gate23301  (.A(g18247), .B(g24057), .Z(II32460) ) ;
NAND2   gate23302  (.A(g18247), .B(II32460), .Z(II32461) ) ;
NAND2   gate23303  (.A(g24057), .B(II32460), .Z(II32462) ) ;
NAND2   gate23304  (.A(g17903), .B(g24058), .Z(II32468) ) ;
NAND2   gate23305  (.A(g17903), .B(II32468), .Z(II32469) ) ;
NAND2   gate23306  (.A(g24058), .B(II32468), .Z(II32470) ) ;
NAND2   gate23307  (.A(g17927), .B(g24065), .Z(II32478) ) ;
NAND2   gate23308  (.A(g17927), .B(II32478), .Z(II32479) ) ;
NAND2   gate23309  (.A(g24065), .B(II32478), .Z(II32480) ) ;
NAND2   gate23310  (.A(g18131), .B(g24067), .Z(II32490) ) ;
NAND2   gate23311  (.A(g18131), .B(II32490), .Z(II32491) ) ;
NAND2   gate23312  (.A(g24067), .B(II32490), .Z(II32492) ) ;
NAND2   gate23313  (.A(g18155), .B(g24069), .Z(II32498) ) ;
NAND2   gate23314  (.A(g18155), .B(II32498), .Z(II32499) ) ;
NAND2   gate23315  (.A(g24069), .B(II32498), .Z(II32500) ) ;
NAND2   gate23316  (.A(g17815), .B(g24070), .Z(II32509) ) ;
NAND2   gate23317  (.A(g17815), .B(II32509), .Z(II32510) ) ;
NAND2   gate23318  (.A(g24070), .B(II32509), .Z(II32511) ) ;
NAND2   gate23319  (.A(g18014), .B(g24071), .Z(II32518) ) ;
NAND2   gate23320  (.A(g18014), .B(II32518), .Z(II32519) ) ;
NAND2   gate23321  (.A(g24071), .B(II32518), .Z(II32520) ) ;
NAND2   gate23322  (.A(g18038), .B(g24078), .Z(II32526) ) ;
NAND2   gate23323  (.A(g18038), .B(II32526), .Z(II32527) ) ;
NAND2   gate23324  (.A(g24078), .B(II32526), .Z(II32528) ) ;
NAND2   gate23325  (.A(g18247), .B(g24080), .Z(II32538) ) ;
NAND2   gate23326  (.A(g18247), .B(II32538), .Z(II32539) ) ;
NAND2   gate23327  (.A(g24080), .B(II32538), .Z(II32540) ) ;
NAND2   gate23328  (.A(g17903), .B(g23906), .Z(II32546) ) ;
NAND2   gate23329  (.A(g17903), .B(II32546), .Z(II32547) ) ;
NAND2   gate23330  (.A(g23906), .B(II32546), .Z(II32548) ) ;
NAND2   gate23331  (.A(g17927), .B(g24081), .Z(II32559) ) ;
NAND2   gate23332  (.A(g17927), .B(II32559), .Z(II32560) ) ;
NAND2   gate23333  (.A(g24081), .B(II32559), .Z(II32561) ) ;
NAND2   gate23334  (.A(g18131), .B(g24082), .Z(II32567) ) ;
NAND2   gate23335  (.A(g18131), .B(II32567), .Z(II32568) ) ;
NAND2   gate23336  (.A(g24082), .B(II32567), .Z(II32569) ) ;
NAND2   gate23337  (.A(g18155), .B(g24089), .Z(II32575) ) ;
NAND2   gate23338  (.A(g18155), .B(II32575), .Z(II32576) ) ;
NAND2   gate23339  (.A(g24089), .B(II32575), .Z(II32577) ) ;
NAND2   gate23340  (.A(g17815), .B(g23937), .Z(II32586) ) ;
NAND2   gate23341  (.A(g17815), .B(II32586), .Z(II32587) ) ;
NAND2   gate23342  (.A(g23937), .B(II32586), .Z(II32588) ) ;
NAND2   gate23343  (.A(g18014), .B(g23938), .Z(II32595) ) ;
NAND2   gate23344  (.A(g18014), .B(II32595), .Z(II32596) ) ;
NAND2   gate23345  (.A(g23938), .B(II32595), .Z(II32597) ) ;
NAND2   gate23346  (.A(g18038), .B(g24090), .Z(II32607) ) ;
NAND2   gate23347  (.A(g18038), .B(II32607), .Z(II32608) ) ;
NAND2   gate23348  (.A(g24090), .B(II32607), .Z(II32609) ) ;
NAND2   gate23349  (.A(g18247), .B(g24091), .Z(II32615) ) ;
NAND2   gate23350  (.A(g18247), .B(II32615), .Z(II32616) ) ;
NAND2   gate23351  (.A(g24091), .B(II32615), .Z(II32617) ) ;
NAND2   gate23352  (.A(g17927), .B(g23969), .Z(II32624) ) ;
NAND2   gate23353  (.A(g17927), .B(II32624), .Z(II32625) ) ;
NAND2   gate23354  (.A(g23969), .B(II32624), .Z(II32626) ) ;
NAND2   gate23355  (.A(g18131), .B(g23970), .Z(II32633) ) ;
NAND2   gate23356  (.A(g18131), .B(II32633), .Z(II32634) ) ;
NAND2   gate23357  (.A(g23970), .B(II32633), .Z(II32635) ) ;
NAND2   gate23358  (.A(g18155), .B(g24093), .Z(II32645) ) ;
NAND2   gate23359  (.A(g18155), .B(II32645), .Z(II32646) ) ;
NAND2   gate23360  (.A(g24093), .B(II32645), .Z(II32647) ) ;
NAND2   gate23361  (.A(g18038), .B(g23998), .Z(II32659) ) ;
NAND2   gate23362  (.A(g18038), .B(II32659), .Z(II32660) ) ;
NAND2   gate23363  (.A(g23998), .B(II32659), .Z(II32661) ) ;
NAND2   gate23364  (.A(g18247), .B(g23999), .Z(II32668) ) ;
NAND2   gate23365  (.A(g18247), .B(II32668), .Z(II32669) ) ;
NAND2   gate23366  (.A(g23999), .B(II32668), .Z(II32670) ) ;
NOR3    gate23367  (.A(g23009), .B(g18490), .C(g4456), .Z(g23823) ) ;
NAND2   gate23368  (.A(g23823), .B(g14165), .Z(II32677) ) ;
NAND2   gate23369  (.A(g23823), .B(II32677), .Z(II32678) ) ;
NAND2   gate23370  (.A(g14165), .B(II32677), .Z(II32679) ) ;
NAND2   gate23371  (.A(g18155), .B(g24028), .Z(II32686) ) ;
NAND2   gate23372  (.A(g18155), .B(II32686), .Z(II32687) ) ;
NAND2   gate23373  (.A(g24028), .B(II32686), .Z(II32688) ) ;
NOR3    gate23374  (.A(g23025), .B(g18554), .C(g4632), .Z(g23858) ) ;
NAND2   gate23375  (.A(g23858), .B(g14280), .Z(II32695) ) ;
NAND2   gate23376  (.A(g23858), .B(II32695), .Z(II32696) ) ;
NAND2   gate23377  (.A(g14280), .B(II32695), .Z(II32697) ) ;
NOR3    gate23378  (.A(g23042), .B(g18604), .C(g4809), .Z(g23892) ) ;
NAND2   gate23379  (.A(g23892), .B(g14402), .Z(II32708) ) ;
NAND2   gate23380  (.A(g23892), .B(II32708), .Z(II32709) ) ;
NAND2   gate23381  (.A(g14402), .B(II32708), .Z(II32710) ) ;
NOR3    gate23382  (.A(g23061), .B(g18636), .C(g4985), .Z(g23913) ) ;
NAND2   gate23383  (.A(g23913), .B(g14514), .Z(II32724) ) ;
NAND2   gate23384  (.A(g23913), .B(II32724), .Z(II32725) ) ;
NAND2   gate23385  (.A(g14514), .B(II32724), .Z(II32726) ) ;
NOR2    gate23386  (.A(g23822), .B(g22701), .Z(g24517) ) ;
NOR2    gate23387  (.A(g23857), .B(g22732), .Z(g24530) ) ;
NOR2    gate23388  (.A(g23891), .B(g22764), .Z(g24543) ) ;
NOR2    gate23389  (.A(g23912), .B(g22798), .Z(g24555) ) ;
NAND2   gate23390  (.A(g26110), .B(g26099), .Z(II35020) ) ;
NAND2   gate23391  (.A(g26110), .B(II35020), .Z(II35021) ) ;
NAND2   gate23392  (.A(g26099), .B(II35020), .Z(II35022) ) ;
NAND2   gate23393  (.A(II35021), .B(II35022), .Z(g26859) ) ;
NAND2   gate23394  (.A(g26087), .B(g26154), .Z(II35034) ) ;
NAND2   gate23395  (.A(g26087), .B(II35034), .Z(II35035) ) ;
NAND2   gate23396  (.A(g26154), .B(II35034), .Z(II35036) ) ;
NAND2   gate23397  (.A(II35035), .B(II35036), .Z(g26865) ) ;
NAND2   gate23398  (.A(g26151), .B(g26145), .Z(II35042) ) ;
NAND2   gate23399  (.A(g26151), .B(II35042), .Z(II35043) ) ;
NAND2   gate23400  (.A(g26145), .B(II35042), .Z(II35044) ) ;
NAND2   gate23401  (.A(II35043), .B(II35044), .Z(g26867) ) ;
NAND2   gate23402  (.A(g26137), .B(g26126), .Z(II35057) ) ;
NAND2   gate23403  (.A(g26137), .B(II35057), .Z(II35058) ) ;
NAND2   gate23404  (.A(g26126), .B(II35057), .Z(II35059) ) ;
NAND2   gate23405  (.A(II35058), .B(II35059), .Z(g26874) ) ;
NOR2    gate23406  (.A(g24613), .B(g24506), .Z(g25699) ) ;
NOR2    gate23407  (.A(g24708), .B(g24490), .Z(g25569) ) ;
NOR2    gate23408  (.A(g24717), .B(g24497), .Z(g25631) ) ;
NOR2    gate23409  (.A(g24624), .B(g24520), .Z(g25772) ) ;
NOR2    gate23410  (.A(g24720), .B(g24500), .Z(g25648) ) ;
NOR2    gate23411  (.A(g24728), .B(g24509), .Z(g25708) ) ;
NOR2    gate23412  (.A(g24638), .B(g24533), .Z(g25826) ) ;
NOR2    gate23413  (.A(g24731), .B(g24512), .Z(g25725) ) ;
NOR2    gate23414  (.A(g24736), .B(g24523), .Z(g25781) ) ;
NOR2    gate23415  (.A(g24657), .B(g24546), .Z(g25861) ) ;
NOR2    gate23416  (.A(g24739), .B(g24526), .Z(g25798) ) ;
NOR2    gate23417  (.A(g24742), .B(g24536), .Z(g25835) ) ;
NOR3    gate23418  (.A(g6068), .B(g24183), .C(g25383), .Z(g26107) ) ;
NOR3    gate23419  (.A(g6068), .B(g24183), .C(g25394), .Z(g26096) ) ;
NAND2   gate23420  (.A(g26107), .B(g26096), .Z(II35123) ) ;
NAND2   gate23421  (.A(g26107), .B(II35123), .Z(II35124) ) ;
NAND2   gate23422  (.A(g26096), .B(II35123), .Z(II35125) ) ;
NAND2   gate23423  (.A(g26867), .B(g26874), .Z(II35701) ) ;
NAND2   gate23424  (.A(g26867), .B(II35701), .Z(II35702) ) ;
NAND2   gate23425  (.A(g26874), .B(II35701), .Z(II35703) ) ;
NAND2   gate23426  (.A(II35702), .B(II35703), .Z(g27379) ) ;
NAND2   gate23427  (.A(g26859), .B(g26865), .Z(II35714) ) ;
NAND2   gate23428  (.A(g26859), .B(II35714), .Z(II35715) ) ;
NAND2   gate23429  (.A(g26865), .B(II35714), .Z(II35716) ) ;
NAND2   gate23430  (.A(II35715), .B(II35716), .Z(g27382) ) ;
NOR2    gate23431  (.A(g26663), .B(g21913), .Z(g26989) ) ;
NOR2    gate23432  (.A(g26668), .B(g21931), .Z(g27012) ) ;
NOR2    gate23433  (.A(g26674), .B(g20640), .Z(g27038) ) ;
NOR2    gate23434  (.A(g26024), .B(g20665), .Z(g27066) ) ;
NOR2    gate23435  (.A(g4456), .B(g26081), .Z(g27051) ) ;
NAND2   gate23436  (.A(g27051), .B(g14831), .Z(II35904) ) ;
NAND2   gate23437  (.A(g27051), .B(II35904), .Z(II35905) ) ;
NAND2   gate23438  (.A(g14831), .B(II35904), .Z(II35906) ) ;
NOR2    gate23439  (.A(g4632), .B(g26084), .Z(g27078) ) ;
NAND2   gate23440  (.A(g27078), .B(g14904), .Z(II35944) ) ;
NAND2   gate23441  (.A(g27078), .B(II35944), .Z(II35945) ) ;
NAND2   gate23442  (.A(g14904), .B(II35944), .Z(II35946) ) ;
NOR2    gate23443  (.A(g4809), .B(g26090), .Z(g27094) ) ;
NAND2   gate23444  (.A(g27094), .B(g14985), .Z(II35974) ) ;
NAND2   gate23445  (.A(g27094), .B(II35974), .Z(II35975) ) ;
NAND2   gate23446  (.A(g14985), .B(II35974), .Z(II35976) ) ;
NOR2    gate23447  (.A(g4985), .B(g26103), .Z(g27106) ) ;
NAND2   gate23448  (.A(g27106), .B(g15074), .Z(II35992) ) ;
NAND2   gate23449  (.A(g27106), .B(II35992), .Z(II35993) ) ;
NAND2   gate23450  (.A(g15074), .B(II35992), .Z(II35994) ) ;
NOR3    gate23451  (.A(g23104), .B(g27181), .C(g25128), .Z(g27415) ) ;
NOR3    gate23452  (.A(g23118), .B(g27187), .C(g24427), .Z(g27436) ) ;
NOR3    gate23453  (.A(g23127), .B(g26758), .C(g24431), .Z(g27455) ) ;
NOR3    gate23454  (.A(g23138), .B(g26764), .C(g24435), .Z(g27471) ) ;
NOR2    gate23455  (.A(g26759), .B(g19087), .Z(g27527) ) ;
NAND2   gate23456  (.A(g27527), .B(g15859), .Z(II36256) ) ;
NAND2   gate23457  (.A(g27527), .B(II36256), .Z(II36257) ) ;
NAND2   gate23458  (.A(g15859), .B(II36256), .Z(II36258) ) ;
NAND2   gate23459  (.A(II36257), .B(II36258), .Z(g27801) ) ;
NOR2    gate23460  (.A(g26765), .B(g19093), .Z(g27549) ) ;
NAND2   gate23461  (.A(g27549), .B(g15890), .Z(II36270) ) ;
NAND2   gate23462  (.A(g27549), .B(II36270), .Z(II36271) ) ;
NAND2   gate23463  (.A(g15890), .B(II36270), .Z(II36272) ) ;
NAND2   gate23464  (.A(II36271), .B(II36272), .Z(g27809) ) ;
NOR2    gate23465  (.A(g26768), .B(g19100), .Z(g27565) ) ;
NAND2   gate23466  (.A(g27565), .B(g15923), .Z(II36289) ) ;
NAND2   gate23467  (.A(g27565), .B(II36289), .Z(II36290) ) ;
NAND2   gate23468  (.A(g15923), .B(II36289), .Z(II36291) ) ;
NAND2   gate23469  (.A(II36290), .B(II36291), .Z(g27830) ) ;
NAND2   gate23470  (.A(g27382), .B(g27379), .Z(II36300) ) ;
NAND2   gate23471  (.A(g27382), .B(II36300), .Z(II36301) ) ;
NAND2   gate23472  (.A(g27379), .B(II36300), .Z(II36302) ) ;
NOR2    gate23473  (.A(g26774), .B(g19107), .Z(g27575) ) ;
NAND2   gate23474  (.A(g27575), .B(g15952), .Z(II36314) ) ;
NAND2   gate23475  (.A(g27575), .B(II36314), .Z(II36315) ) ;
NAND2   gate23476  (.A(g15952), .B(II36314), .Z(II36316) ) ;
NAND2   gate23477  (.A(II36315), .B(II36316), .Z(g27846) ) ;
NOR2    gate23478  (.A(g4456), .B(g26873), .Z(g27529) ) ;
NAND2   gate23479  (.A(g27529), .B(g14885), .Z(II36591) ) ;
NAND2   gate23480  (.A(g27529), .B(II36591), .Z(II36592) ) ;
NAND2   gate23481  (.A(g14885), .B(II36591), .Z(II36593) ) ;
NOR2    gate23482  (.A(g4632), .B(g26882), .Z(g27551) ) ;
NAND2   gate23483  (.A(g27551), .B(g14966), .Z(II36666) ) ;
NAND2   gate23484  (.A(g27551), .B(II36666), .Z(II36667) ) ;
NAND2   gate23485  (.A(g14966), .B(II36666), .Z(II36668) ) ;
NOR2    gate23486  (.A(g4809), .B(g26891), .Z(g27567) ) ;
NAND2   gate23487  (.A(g27567), .B(g15055), .Z(II36731) ) ;
NAND2   gate23488  (.A(g27567), .B(II36731), .Z(II36732) ) ;
NAND2   gate23489  (.A(g15055), .B(II36731), .Z(II36733) ) ;
NOR2    gate23490  (.A(g4985), .B(g26901), .Z(g27577) ) ;
NAND2   gate23491  (.A(g27577), .B(g15151), .Z(II36779) ) ;
NAND2   gate23492  (.A(g27577), .B(II36779), .Z(II36780) ) ;
NAND2   gate23493  (.A(g15151), .B(II36779), .Z(II36781) ) ;
NAND2   gate23494  (.A(g27827), .B(g27814), .Z(II37295) ) ;
NAND2   gate23495  (.A(g27827), .B(II37295), .Z(II37296) ) ;
NAND2   gate23496  (.A(g27814), .B(II37295), .Z(II37297) ) ;
NAND2   gate23497  (.A(II37296), .B(II37297), .Z(g28384) ) ;
NAND2   gate23498  (.A(g27802), .B(g27900), .Z(II37303) ) ;
NAND2   gate23499  (.A(g27802), .B(II37303), .Z(II37304) ) ;
NAND2   gate23500  (.A(g27900), .B(II37303), .Z(II37305) ) ;
NAND2   gate23501  (.A(II37304), .B(II37305), .Z(g28386) ) ;
NAND2   gate23502  (.A(g27897), .B(g27883), .Z(II37311) ) ;
NAND2   gate23503  (.A(g27897), .B(II37311), .Z(II37312) ) ;
NAND2   gate23504  (.A(g27883), .B(II37311), .Z(II37313) ) ;
NAND2   gate23505  (.A(II37312), .B(II37313), .Z(g28388) ) ;
NAND2   gate23506  (.A(g27865), .B(g27855), .Z(II37322) ) ;
NAND2   gate23507  (.A(g27865), .B(II37322), .Z(II37323) ) ;
NAND2   gate23508  (.A(g27855), .B(II37322), .Z(II37324) ) ;
NAND2   gate23509  (.A(II37323), .B(II37324), .Z(g28391) ) ;
NOR3    gate23510  (.A(g6087), .B(g27632), .C(g25399), .Z(g27824) ) ;
NOR3    gate23511  (.A(g6087), .B(g27632), .C(g25404), .Z(g27811) ) ;
NAND2   gate23512  (.A(g27824), .B(g27811), .Z(II37356) ) ;
NAND2   gate23513  (.A(g27824), .B(II37356), .Z(II37357) ) ;
NAND2   gate23514  (.A(g27811), .B(II37356), .Z(II37358) ) ;
NAND2   gate23515  (.A(g28388), .B(g28391), .Z(II37813) ) ;
NAND2   gate23516  (.A(g28388), .B(II37813), .Z(II37814) ) ;
NAND2   gate23517  (.A(g28391), .B(II37813), .Z(II37815) ) ;
NAND2   gate23518  (.A(II37814), .B(II37815), .Z(g28842) ) ;
NAND2   gate23519  (.A(g28384), .B(g28386), .Z(II37822) ) ;
NAND2   gate23520  (.A(g28384), .B(II37822), .Z(II37823) ) ;
NAND2   gate23521  (.A(g28386), .B(II37822), .Z(II37824) ) ;
NAND2   gate23522  (.A(II37823), .B(II37824), .Z(g28845) ) ;
NAND2   gate23523  (.A(g28845), .B(g28842), .Z(II38378) ) ;
NAND2   gate23524  (.A(g28845), .B(II38378), .Z(II38379) ) ;
NAND2   gate23525  (.A(g28842), .B(II38378), .Z(II38380) ) ;
NOR2    gate23526  (.A(g28716), .B(g19112), .Z(g29303) ) ;
NAND2   gate23527  (.A(g29303), .B(g15904), .Z(II38810) ) ;
NAND2   gate23528  (.A(g29303), .B(II38810), .Z(II38811) ) ;
NAND2   gate23529  (.A(g15904), .B(II38810), .Z(II38812) ) ;
NOR2    gate23530  (.A(g28717), .B(g19117), .Z(g29313) ) ;
NAND2   gate23531  (.A(g29313), .B(g15933), .Z(II38820) ) ;
NAND2   gate23532  (.A(g29313), .B(II38820), .Z(II38821) ) ;
NAND2   gate23533  (.A(g15933), .B(II38820), .Z(II38822) ) ;
NOR2    gate23534  (.A(g28718), .B(g19124), .Z(g29324) ) ;
NAND2   gate23535  (.A(g29324), .B(g15962), .Z(II38831) ) ;
NAND2   gate23536  (.A(g29324), .B(II38831), .Z(II38832) ) ;
NAND2   gate23537  (.A(g15962), .B(II38831), .Z(II38833) ) ;
NOR2    gate23538  (.A(g28719), .B(g19131), .Z(g29333) ) ;
NAND2   gate23539  (.A(g29333), .B(g15981), .Z(II38841) ) ;
NAND2   gate23540  (.A(g29333), .B(II38841), .Z(II38842) ) ;
NAND2   gate23541  (.A(g15981), .B(II38841), .Z(II38843) ) ;
NAND2   gate23542  (.A(g29721), .B(g29713), .Z(II39323) ) ;
NAND2   gate23543  (.A(g29721), .B(II39323), .Z(II39324) ) ;
NAND2   gate23544  (.A(g29713), .B(II39323), .Z(II39325) ) ;
NAND2   gate23545  (.A(II39324), .B(II39325), .Z(g29911) ) ;
NAND2   gate23546  (.A(g29705), .B(g29751), .Z(II39331) ) ;
NAND2   gate23547  (.A(g29705), .B(II39331), .Z(II39332) ) ;
NAND2   gate23548  (.A(g29751), .B(II39331), .Z(II39333) ) ;
NAND2   gate23549  (.A(II39332), .B(II39333), .Z(g29913) ) ;
NAND2   gate23550  (.A(g29748), .B(g29741), .Z(II39339) ) ;
NAND2   gate23551  (.A(g29748), .B(II39339), .Z(II39340) ) ;
NAND2   gate23552  (.A(g29741), .B(II39339), .Z(II39341) ) ;
NAND2   gate23553  (.A(II39340), .B(II39341), .Z(g29915) ) ;
NAND2   gate23554  (.A(g29732), .B(g29728), .Z(II39347) ) ;
NAND2   gate23555  (.A(g29732), .B(II39347), .Z(II39348) ) ;
NAND2   gate23556  (.A(g29728), .B(II39347), .Z(II39349) ) ;
NAND2   gate23557  (.A(II39348), .B(II39349), .Z(g29917) ) ;
NOR2    gate23558  (.A(g29467), .B(g19142), .Z(g29766) ) ;
NAND2   gate23559  (.A(g29766), .B(g15880), .Z(II39359) ) ;
NAND2   gate23560  (.A(g29766), .B(II39359), .Z(II39360) ) ;
NAND2   gate23561  (.A(g15880), .B(II39359), .Z(II39361) ) ;
NAND2   gate23562  (.A(II39360), .B(II39361), .Z(g29923) ) ;
NOR2    gate23563  (.A(g29468), .B(g19143), .Z(g29767) ) ;
NAND2   gate23564  (.A(g29767), .B(g15913), .Z(II39367) ) ;
NAND2   gate23565  (.A(g29767), .B(II39367), .Z(II39368) ) ;
NAND2   gate23566  (.A(g15913), .B(II39367), .Z(II39369) ) ;
NAND2   gate23567  (.A(II39368), .B(II39369), .Z(g29925) ) ;
NOR2    gate23568  (.A(g29469), .B(g19146), .Z(g29768) ) ;
NAND2   gate23569  (.A(g29768), .B(g15942), .Z(II39375) ) ;
NAND2   gate23570  (.A(g29768), .B(II39375), .Z(II39376) ) ;
NAND2   gate23571  (.A(g15942), .B(II39375), .Z(II39377) ) ;
NAND2   gate23572  (.A(II39376), .B(II39377), .Z(g29927) ) ;
NOR3    gate23573  (.A(g6104), .B(g29583), .C(g25409), .Z(g29718) ) ;
NOR3    gate23574  (.A(g6104), .B(g29583), .C(g25412), .Z(g29710) ) ;
NAND2   gate23575  (.A(g29718), .B(g29710), .Z(II39384) ) ;
NAND2   gate23576  (.A(g29718), .B(II39384), .Z(II39385) ) ;
NAND2   gate23577  (.A(g29710), .B(II39384), .Z(II39386) ) ;
NOR2    gate23578  (.A(g29470), .B(g19148), .Z(g29769) ) ;
NAND2   gate23579  (.A(g29769), .B(g15971), .Z(II39391) ) ;
NAND2   gate23580  (.A(g29769), .B(II39391), .Z(II39392) ) ;
NAND2   gate23581  (.A(g15971), .B(II39391), .Z(II39393) ) ;
NAND2   gate23582  (.A(II39392), .B(II39393), .Z(g29931) ) ;
NAND2   gate23583  (.A(g29915), .B(g29917), .Z(II39532) ) ;
NAND2   gate23584  (.A(g29915), .B(II39532), .Z(II39533) ) ;
NAND2   gate23585  (.A(g29917), .B(II39532), .Z(II39534) ) ;
NAND2   gate23586  (.A(II39533), .B(II39534), .Z(g30034) ) ;
NAND2   gate23587  (.A(g29911), .B(g29913), .Z(II39539) ) ;
NAND2   gate23588  (.A(g29911), .B(II39539), .Z(II39540) ) ;
NAND2   gate23589  (.A(g29913), .B(II39539), .Z(II39541) ) ;
NAND2   gate23590  (.A(II39540), .B(II39541), .Z(g30035) ) ;
NAND2   gate23591  (.A(g30035), .B(g30034), .Z(II39689) ) ;
NAND2   gate23592  (.A(g30035), .B(II39689), .Z(II39690) ) ;
NAND2   gate23593  (.A(g30034), .B(II39689), .Z(II39691) ) ;
NAND2   gate23594  (.A(g30605), .B(g30597), .Z(II40558) ) ;
NAND2   gate23595  (.A(g30605), .B(II40558), .Z(II40559) ) ;
NAND2   gate23596  (.A(g30597), .B(II40558), .Z(II40560) ) ;
NAND2   gate23597  (.A(II40559), .B(II40560), .Z(g30768) ) ;
NAND2   gate23598  (.A(g30588), .B(g30632), .Z(II40571) ) ;
NAND2   gate23599  (.A(g30588), .B(II40571), .Z(II40572) ) ;
NAND2   gate23600  (.A(g30632), .B(II40571), .Z(II40573) ) ;
NAND2   gate23601  (.A(II40572), .B(II40573), .Z(g30771) ) ;
NAND2   gate23602  (.A(g30629), .B(g30622), .Z(II40587) ) ;
NAND2   gate23603  (.A(g30629), .B(II40587), .Z(II40588) ) ;
NAND2   gate23604  (.A(g30622), .B(II40587), .Z(II40589) ) ;
NAND2   gate23605  (.A(II40588), .B(II40589), .Z(g30775) ) ;
NAND2   gate23606  (.A(g30614), .B(g30610), .Z(II40603) ) ;
NAND2   gate23607  (.A(g30614), .B(II40603), .Z(II40604) ) ;
NAND2   gate23608  (.A(g30610), .B(II40603), .Z(II40605) ) ;
NAND2   gate23609  (.A(II40604), .B(II40605), .Z(g30779) ) ;
NOR3    gate23610  (.A(g6119), .B(g30412), .C(g25417), .Z(g30602) ) ;
NOR3    gate23611  (.A(g6119), .B(g30412), .C(g25419), .Z(g30594) ) ;
NAND2   gate23612  (.A(g30602), .B(g30594), .Z(II40627) ) ;
NAND2   gate23613  (.A(g30602), .B(II40627), .Z(II40628) ) ;
NAND2   gate23614  (.A(g30594), .B(II40627), .Z(II40629) ) ;
NAND2   gate23615  (.A(g30775), .B(g30779), .Z(II41010) ) ;
NAND2   gate23616  (.A(g30775), .B(II41010), .Z(II41011) ) ;
NAND2   gate23617  (.A(g30779), .B(II41010), .Z(II41012) ) ;
NAND2   gate23618  (.A(II41011), .B(II41012), .Z(g30926) ) ;
NAND2   gate23619  (.A(g30768), .B(g30771), .Z(II41017) ) ;
NAND2   gate23620  (.A(g30768), .B(II41017), .Z(II41018) ) ;
NAND2   gate23621  (.A(g30771), .B(II41017), .Z(II41019) ) ;
NAND2   gate23622  (.A(II41018), .B(II41019), .Z(g30927) ) ;
NAND2   gate23623  (.A(g30927), .B(g30926), .Z(II41064) ) ;
NAND2   gate23624  (.A(g30927), .B(II41064), .Z(II41065) ) ;
NAND2   gate23625  (.A(g30926), .B(II41064), .Z(II41066) ) ;
NOR3    gate23626  (.A(g6200), .B(g12457), .C(g10952), .Z(g16020) ) ;
NOR3    gate23627  (.A(g6289), .B(g12467), .C(g10952), .Z(g16036) ) ;
NOR3    gate23628  (.A(g6426), .B(g12482), .C(g10952), .Z(g16058) ) ;
NOR3    gate23629  (.A(g10952), .B(g6140), .C(g12487), .Z(g16082) ) ;
NOR3    gate23630  (.A(g6631), .B(g12499), .C(g10952), .Z(g16094) ) ;
NOR3    gate23631  (.A(g10952), .B(g6161), .C(g12507), .Z(g16120) ) ;
NOR3    gate23632  (.A(g10952), .B(g6188), .C(g12524), .Z(g16171) ) ;
NOR3    gate23633  (.A(g10952), .B(g6220), .C(g12539), .Z(g16230) ) ;
NOR2    gate23634  (.A(g16082), .B(g14249), .Z(g18352) ) ;
NOR2    gate23635  (.A(g16020), .B(g14352), .Z(g18430) ) ;
NOR2    gate23636  (.A(g16120), .B(g14371), .Z(g18447) ) ;
NOR2    gate23637  (.A(g16036), .B(g14464), .Z(g18503) ) ;
NOR2    gate23638  (.A(g16171), .B(g14483), .Z(g18520) ) ;
NOR2    gate23639  (.A(g16058), .B(g14551), .Z(g18567) ) ;
NOR2    gate23640  (.A(g16230), .B(g14570), .Z(g18584) ) ;
NOR2    gate23641  (.A(g16094), .B(g14606), .Z(g18617) ) ;
NOR2    gate23642  (.A(g17446), .B(g15178), .Z(g19160) ) ;
NOR2    gate23643  (.A(g17526), .B(g15264), .Z(g19165) ) ;
NOR2    gate23644  (.A(g17616), .B(g15356), .Z(g19171) ) ;
NOR2    gate23645  (.A(g17713), .B(g15442), .Z(g19177) ) ;
NOR2    gate23646  (.A(g19600), .B(g17395), .Z(g20878) ) ;
NOR2    gate23647  (.A(g19633), .B(g17461), .Z(g20895) ) ;
NOR2    gate23648  (.A(g19673), .B(g17541), .Z(g20914) ) ;
NOR2    gate23649  (.A(g19721), .B(g17631), .Z(g20938) ) ;
NOR2    gate23650  (.A(g19943), .B(g18333), .Z(g21083) ) ;
NOR3    gate23651  (.A(g20016), .B(g14079), .C(g14165), .Z(g21618) ) ;
NOR3    gate23652  (.A(g20058), .B(g14194), .C(g14280), .Z(g21646) ) ;
NOR3    gate23653  (.A(g20099), .B(g14309), .C(g14402), .Z(g21677) ) ;
NOR3    gate23654  (.A(g20124), .B(g14431), .C(g14514), .Z(g21706) ) ;
NOR3    gate23655  (.A(g19444), .B(g17893), .C(g14079), .Z(g21738) ) ;
NOR3    gate23656  (.A(g19471), .B(g18004), .C(g14194), .Z(g21762) ) ;
NOR3    gate23657  (.A(g19494), .B(g18121), .C(g14309), .Z(g21778) ) ;
NOR3    gate23658  (.A(g19515), .B(g18237), .C(g14431), .Z(g21793) ) ;
NOR2    gate23659  (.A(g21410), .B(g19730), .Z(g22144) ) ;
NOR2    gate23660  (.A(g21444), .B(g19773), .Z(g22165) ) ;
NOR2    gate23661  (.A(g21486), .B(g19815), .Z(g22181) ) ;
NOR2    gate23662  (.A(g21497), .B(g19837), .Z(g22186) ) ;
NOR2    gate23663  (.A(g21527), .B(g19859), .Z(g22195) ) ;
NOR2    gate23664  (.A(g21610), .B(g19932), .Z(g22210) ) ;
NOR2    gate23665  (.A(g21635), .B(g19944), .Z(g22216) ) ;
NOR2    gate23666  (.A(g21658), .B(g19953), .Z(g22227) ) ;
NOR2    gate23667  (.A(g21618), .B(g21049), .Z(g22985) ) ;
NOR2    gate23668  (.A(g21646), .B(g21068), .Z(g22987) ) ;
NOR2    gate23669  (.A(g21677), .B(g21078), .Z(g22990) ) ;
NOR2    gate23670  (.A(g21706), .B(g21092), .Z(g22997) ) ;
NOR2    gate23671  (.A(g21738), .B(g21107), .Z(g23009) ) ;
NOR2    gate23672  (.A(g21762), .B(g21124), .Z(g23025) ) ;
NOR2    gate23673  (.A(g21778), .B(g21143), .Z(g23042) ) ;
NOR2    gate23674  (.A(g21793), .B(g21163), .Z(g23061) ) ;
NOR2    gate23675  (.A(g22483), .B(g21388), .Z(g23386) ) ;
NOR2    gate23676  (.A(g22526), .B(g21418), .Z(g23393) ) ;
NOR2    gate23677  (.A(g22566), .B(g21452), .Z(g23401) ) ;
NOR2    gate23678  (.A(g22606), .B(g21494), .Z(g23408) ) ;
NOR2    gate23679  (.A(g22699), .B(g21589), .Z(g23427) ) ;
NOR2    gate23680  (.A(g22726), .B(g21611), .Z(g23433) ) ;
NOR2    gate23681  (.A(g22841), .B(g21707), .Z(g23461) ) ;
NOR2    gate23682  (.A(g22906), .B(g21758), .Z(g23477) ) ;
NOR2    gate23683  (.A(g22270), .B(g21137), .Z(g24227) ) ;
NOR2    gate23684  (.A(g22289), .B(g21157), .Z(g24234) ) ;
NOR2    gate23685  (.A(g22309), .B(g21177), .Z(g24242) ) ;
NOR2    gate23686  (.A(g22337), .B(g21197), .Z(g24249) ) ;
NOR2    gate23687  (.A(g23544), .B(g22398), .Z(g24428) ) ;
NOR2    gate23688  (.A(g23643), .B(g22577), .Z(g24486) ) ;
NOR2    gate23689  (.A(g23686), .B(g22607), .Z(g24490) ) ;
NOR2    gate23690  (.A(g23689), .B(g22610), .Z(g24492) ) ;
NOR2    gate23691  (.A(g23693), .B(g22614), .Z(g24493) ) ;
NOR2    gate23692  (.A(g23734), .B(g22638), .Z(g24497) ) ;
NOR2    gate23693  (.A(g23740), .B(g22643), .Z(g24500) ) ;
NOR2    gate23694  (.A(g23743), .B(g22646), .Z(g24502) ) ;
NOR2    gate23695  (.A(g23747), .B(g22650), .Z(g24503) ) ;
NOR2    gate23696  (.A(g23776), .B(g22667), .Z(g24506) ) ;
NOR2    gate23697  (.A(g23789), .B(g22674), .Z(g24509) ) ;
NOR2    gate23698  (.A(g23795), .B(g22679), .Z(g24512) ) ;
NOR2    gate23699  (.A(g23798), .B(g22682), .Z(g24514) ) ;
NOR2    gate23700  (.A(g23802), .B(g22686), .Z(g24515) ) ;
NOR2    gate23701  (.A(g23820), .B(g22700), .Z(g24516) ) ;
NOR2    gate23702  (.A(g23829), .B(g22707), .Z(g24520) ) ;
NOR2    gate23703  (.A(g23842), .B(g22714), .Z(g24523) ) ;
NOR2    gate23704  (.A(g23848), .B(g22719), .Z(g24526) ) ;
NOR2    gate23705  (.A(g23851), .B(g22722), .Z(g24528) ) ;
NOR2    gate23706  (.A(g23864), .B(g22738), .Z(g24533) ) ;
NOR2    gate23707  (.A(g23877), .B(g22745), .Z(g24536) ) ;
NOR2    gate23708  (.A(g23898), .B(g22770), .Z(g24546) ) ;
NOR2    gate23709  (.A(g23917), .B(g22804), .Z(g24558) ) ;
NOR2    gate23710  (.A(g23944), .B(g22842), .Z(g24566) ) ;
NOR2    gate23711  (.A(g23972), .B(g22874), .Z(g24575) ) ;
NOR2    gate23712  (.A(g23592), .B(g22515), .Z(g24613) ) ;
NOR2    gate23713  (.A(g23616), .B(g22546), .Z(g24622) ) ;
NOR2    gate23714  (.A(g23624), .B(g22555), .Z(g24624) ) ;
NOR2    gate23715  (.A(g23665), .B(g22587), .Z(g24637) ) ;
NOR2    gate23716  (.A(g23673), .B(g22595), .Z(g24638) ) ;
NOR2    gate23717  (.A(g23715), .B(g22624), .Z(g24656) ) ;
NOR2    gate23718  (.A(g23723), .B(g22632), .Z(g24657) ) ;
NOR2    gate23719  (.A(g23769), .B(g22660), .Z(g24675) ) ;
NOR2    gate23720  (.A(g23854), .B(g22727), .Z(g24708) ) ;
NOR2    gate23721  (.A(g23886), .B(g22754), .Z(g24717) ) ;
NOR2    gate23722  (.A(g23888), .B(g22759), .Z(g24720) ) ;
NOR2    gate23723  (.A(g23907), .B(g22788), .Z(g24728) ) ;
NOR2    gate23724  (.A(g23909), .B(g22793), .Z(g24731) ) ;
NOR2    gate23725  (.A(g23939), .B(g22830), .Z(g24736) ) ;
NOR2    gate23726  (.A(g23941), .B(g22835), .Z(g24739) ) ;
NOR2    gate23727  (.A(g23971), .B(g22869), .Z(g24742) ) ;
NOR2    gate23728  (.A(g23409), .B(g22187), .Z(g25076) ) ;
NOR2    gate23729  (.A(g23414), .B(g22196), .Z(g25077) ) ;
NOR2    gate23730  (.A(g23419), .B(g22201), .Z(g25078) ) ;
NOR2    gate23731  (.A(g23423), .B(g22202), .Z(g25081) ) ;
NOR2    gate23732  (.A(g23428), .B(g22207), .Z(g25082) ) ;
NOR2    gate23733  (.A(g23432), .B(g22208), .Z(g25085) ) ;
NOR2    gate23734  (.A(g23434), .B(g22215), .Z(g25091) ) ;
NOR2    gate23735  (.A(g23440), .B(g22224), .Z(g25099) ) ;
NOR2    gate23736  (.A(g23510), .B(g22340), .Z(g25125) ) ;
NOR2    gate23737  (.A(g23525), .B(g22363), .Z(g25127) ) ;
NOR2    gate23738  (.A(g23536), .B(g22383), .Z(g25129) ) ;
NOR2    gate23739  (.A(g24748), .B(g23552), .Z(g25208) ) ;
NOR2    gate23740  (.A(g24757), .B(g23565), .Z(g25216) ) ;
NOR2    gate23741  (.A(g24774), .B(g23584), .Z(g25226) ) ;
NOR2    gate23742  (.A(g24794), .B(g23611), .Z(g25238) ) ;
NOR2    gate23743  (.A(g24907), .B(g23904), .Z(g25273) ) ;
NOR2    gate23744  (.A(g24964), .B(g24029), .Z(g25311) ) ;
NOR2    gate23745  (.A(g24183), .B(g24616), .Z(g25426) ) ;
NOR2    gate23746  (.A(g24591), .B(g23496), .Z(g25962) ) ;
NOR2    gate23747  (.A(g24596), .B(g23512), .Z(g25967) ) ;
NOR2    gate23748  (.A(g24604), .B(g23527), .Z(g25974) ) ;
NOR2    gate23749  (.A(g24611), .B(g23538), .Z(g25979) ) ;
NOR2    gate23750  (.A(g25505), .B(g24867), .Z(g26042) ) ;
NOR2    gate23751  (.A(g25552), .B(g24882), .Z(g26044) ) ;
NOR2    gate23752  (.A(g25618), .B(g24899), .Z(g26046) ) ;
NOR2    gate23753  (.A(g25629), .B(g24908), .Z(g26049) ) ;
NOR2    gate23754  (.A(g25697), .B(g24922), .Z(g26050) ) ;
NOR2    gate23755  (.A(g25881), .B(g24974), .Z(g26055) ) ;
NOR2    gate23756  (.A(g25470), .B(g25482), .Z(g26081) ) ;
NOR2    gate23757  (.A(g25487), .B(g25513), .Z(g26084) ) ;
NOR2    gate23758  (.A(g25518), .B(g25560), .Z(g26090) ) ;
NOR2    gate23759  (.A(g25565), .B(g25626), .Z(g26103) ) ;
NOR2    gate23760  (.A(g24183), .B(g25430), .Z(g26140) ) ;
NOR2    gate23761  (.A(g25281), .B(g24559), .Z(g26560) ) ;
NOR2    gate23762  (.A(g25289), .B(g24569), .Z(g26583) ) ;
NOR2    gate23763  (.A(g25299), .B(g24578), .Z(g26607) ) ;
NOR2    gate23764  (.A(g25309), .B(g24585), .Z(g26630) ) ;
NOR2    gate23765  (.A(g26158), .B(g25453), .Z(g26799) ) ;
NOR2    gate23766  (.A(g26163), .B(g25457), .Z(g26800) ) ;
NOR2    gate23767  (.A(g26171), .B(g25461), .Z(g26801) ) ;
NOR2    gate23768  (.A(g26188), .B(g25466), .Z(g26802) ) ;
NOR2    gate23769  (.A(g25483), .B(g26260), .Z(g26873) ) ;
NOR2    gate23770  (.A(g25514), .B(g26301), .Z(g26882) ) ;
NOR2    gate23771  (.A(g25561), .B(g26345), .Z(g26891) ) ;
NOR2    gate23772  (.A(g25627), .B(g26389), .Z(g26901) ) ;
NOR2    gate23773  (.A(g26075), .B(g25342), .Z(g27175) ) ;
NOR2    gate23774  (.A(g26082), .B(g25356), .Z(g27179) ) ;
NOR2    gate23775  (.A(g26085), .B(g25371), .Z(g27184) ) ;
NOR2    gate23776  (.A(g26091), .B(g25388), .Z(g27188) ) ;
NOR2    gate23777  (.A(g26955), .B(g26166), .Z(g27250) ) ;
NOR2    gate23778  (.A(g26958), .B(g26186), .Z(g27251) ) ;
NOR2    gate23779  (.A(g26963), .B(g26207), .Z(g27252) ) ;
NOR2    gate23780  (.A(g26968), .B(g26231), .Z(g27254) ) ;
NOR2    gate23781  (.A(g26754), .B(g24432), .Z(g27478) ) ;
NOR2    gate23782  (.A(g26763), .B(g24436), .Z(g27501) ) ;
NOR2    gate23783  (.A(g26766), .B(g24439), .Z(g27521) ) ;
NOR2    gate23784  (.A(g26769), .B(g24441), .Z(g27546) ) ;
NOR2    gate23785  (.A(g26829), .B(g26051), .Z(g27629) ) ;
NOR2    gate23786  (.A(g26833), .B(g26053), .Z(g27631) ) ;
NOR2    gate23787  (.A(g26842), .B(g26061), .Z(g27655) ) ;
NOR2    gate23788  (.A(g26851), .B(g26068), .Z(g27658) ) ;
NOR2    gate23789  (.A(g27396), .B(g26962), .Z(g27736) ) ;
NOR2    gate23790  (.A(g27409), .B(g26967), .Z(g27742) ) ;
NOR2    gate23791  (.A(g27427), .B(g26973), .Z(g27747) ) ;
NOR2    gate23792  (.A(g27448), .B(g26986), .Z(g27755) ) ;
NOR2    gate23793  (.A(g27632), .B(g25437), .Z(g27869) ) ;
NOR2    gate23794  (.A(g27632), .B(g24627), .Z(g27886) ) ;
NOR2    gate23795  (.A(g27356), .B(g26845), .Z(g28185) ) ;
NOR2    gate23796  (.A(g27359), .B(g26853), .Z(g28189) ) ;
NOR2    gate23797  (.A(g27365), .B(g26860), .Z(g28191) ) ;
NOR2    gate23798  (.A(g27372), .B(g26866), .Z(g28192) ) ;
NOR2    gate23799  (.A(g27770), .B(g27355), .Z(g28654) ) ;
NOR2    gate23800  (.A(g27772), .B(g27358), .Z(g28656) ) ;
NOR2    gate23801  (.A(g27773), .B(g27364), .Z(g28658) ) ;
NOR2    gate23802  (.A(g27775), .B(g27371), .Z(g28661) ) ;
NOR2    gate23803  (.A(g28373), .B(g27774), .Z(g29126) ) ;
NOR2    gate23804  (.A(g28376), .B(g27779), .Z(g29127) ) ;
NOR2    gate23805  (.A(g28380), .B(g27783), .Z(g29128) ) ;
NOR2    gate23806  (.A(g28385), .B(g27790), .Z(g29129) ) ;
NOR2    gate23807  (.A(g28834), .B(g28378), .Z(g29399) ) ;
NOR2    gate23808  (.A(g28836), .B(g28383), .Z(g29403) ) ;
NOR2    gate23809  (.A(g28838), .B(g28387), .Z(g29406) ) ;
NOR2    gate23810  (.A(g28840), .B(g28389), .Z(g29409) ) ;
NOR2    gate23811  (.A(g29583), .B(g25444), .Z(g29736) ) ;
NOR2    gate23812  (.A(g29583), .B(g24641), .Z(g29744) ) ;
NOR2    gate23813  (.A(g30412), .B(g25449), .Z(g30618) ) ;
NOR2    gate23814  (.A(g30412), .B(g24660), .Z(g30625) ) ;

endmodule
