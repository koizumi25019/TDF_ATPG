module s15850 (g18, g27, g109, g741, g742
    , g743, g744, g872, g873, g877
    , g881, g1712, g1960, g1961, CLK
    , g2355, g2601, g2602, g2603, g2604
    , g2605, g2606, g2607, g2608, g2609
    , g2610, g2611, g2612, g2648, g2986
    , g3007, g3069, g4172, g4173, g4174
    , g4175, g4176, g4177, g4178, g4179
    , g4180, g4181, g4887, g4888, g5101
    , g5105, g5658, g5659, g5816, g6920
    , g6926, g6932, g6942, g6949, g6955
    , g7744, g8061, g8062, g8271, g8313
    , g8316, g8318, g8323, g8328, g8331
    , g8335, g8340, g8347, g8349, g8352
    , g8561, g8562, g8563, g8564, g8565
    , g8566, g8976, g8977, g8978, g8979
    , g8980, g8981, g8982, g8983, g8984
    , g8985, g8986, g9451, g9961, g10377
    , g10379, g10455, g10457, g10459, g10461
    , g10463, g10465, g10628, g10801, g11163
    , g11206, g11489) ;

input   g18, g27, g109, g741, g742
    , g743, g744, g872, g873, g877
    , g881, g1712, g1960, g1961, CLK ;

output  g2355, g2601, g2602, g2603, g2604
    , g2605, g2606, g2607, g2608, g2609
    , g2610, g2611, g2612, g2648, g2986
    , g3007, g3069, g4172, g4173, g4174
    , g4175, g4176, g4177, g4178, g4179
    , g4180, g4181, g4887, g4888, g5101
    , g5105, g5658, g5659, g5816, g6920
    , g6926, g6932, g6942, g6949, g6955
    , g7744, g8061, g8062, g8271, g8313
    , g8316, g8318, g8323, g8328, g8331
    , g8335, g8340, g8347, g8349, g8352
    , g8561, g8562, g8563, g8564, g8565
    , g8566, g8976, g8977, g8978, g8979
    , g8980, g8981, g8982, g8983, g8984
    , g8985, g8986, g9451, g9961, g10377
    , g10379, g10455, g10457, g10459, g10461
    , g10463, g10465, g10628, g10801, g11163
    , g11206, g11489 ;

INV     gate0  (.A(II5435), .Z(g2355) ) ;
INV     gate1  (.A(II5704), .Z(g2601) ) ;
INV     gate2  (.A(II5707), .Z(g2602) ) ;
INV     gate3  (.A(II5710), .Z(g2603) ) ;
INV     gate4  (.A(II5713), .Z(g2604) ) ;
INV     gate5  (.A(II5716), .Z(g2605) ) ;
INV     gate6  (.A(II5719), .Z(g2606) ) ;
INV     gate7  (.A(II5722), .Z(g2607) ) ;
INV     gate8  (.A(II5725), .Z(g2608) ) ;
INV     gate9  (.A(II5728), .Z(g2609) ) ;
INV     gate10  (.A(II5731), .Z(g2610) ) ;
INV     gate11  (.A(II5734), .Z(g2611) ) ;
INV     gate12  (.A(II5737), .Z(g2612) ) ;
INV     gate13  (.A(II5765), .Z(g2648) ) ;
INV     gate14  (.A(II6220), .Z(g2986) ) ;
INV     gate15  (.A(II6240), .Z(g3007) ) ;
INV     gate16  (.A(II6277), .Z(g3069) ) ;
INV     gate17  (.A(II7333), .Z(g4172) ) ;
INV     gate18  (.A(II7336), .Z(g4173) ) ;
INV     gate19  (.A(II7339), .Z(g4174) ) ;
INV     gate20  (.A(II7342), .Z(g4175) ) ;
INV     gate21  (.A(II7345), .Z(g4176) ) ;
INV     gate22  (.A(II7348), .Z(g4177) ) ;
INV     gate23  (.A(II7351), .Z(g4178) ) ;
INV     gate24  (.A(II7354), .Z(g4179) ) ;
INV     gate25  (.A(II7357), .Z(g4180) ) ;
INV     gate26  (.A(II7360), .Z(g4181) ) ;
INV     gate27  (.A(II8234), .Z(g4887) ) ;
INV     gate28  (.A(II8237), .Z(g4888) ) ;
INV     gate29  (.A(II8473), .Z(g5101) ) ;
INV     gate30  (.A(II8487), .Z(g5105) ) ;
INV     gate31  (.A(II9135), .Z(g5658) ) ;
INV     gate32  (.A(II9138), .Z(g5659) ) ;
INV     gate33  (.A(II9424), .Z(g5816) ) ;
INV     gate34  (.A(II11034), .Z(g6920) ) ;
INV     gate35  (.A(II11046), .Z(g6926) ) ;
INV     gate36  (.A(II11058), .Z(g6932) ) ;
INV     gate37  (.A(II11076), .Z(g6942) ) ;
INV     gate38  (.A(II11091), .Z(g6949) ) ;
INV     gate39  (.A(II11103), .Z(g6955) ) ;
INV     gate40  (.A(II12397), .Z(g7744) ) ;
INV     gate41  (.A(II12901), .Z(g8061) ) ;
INV     gate42  (.A(II12904), .Z(g8062) ) ;
INV     gate43  (.A(II13185), .Z(g8271) ) ;
INV     gate44  (.A(II13323), .Z(g8313) ) ;
INV     gate45  (.A(II13332), .Z(g8316) ) ;
INV     gate46  (.A(II13338), .Z(g8318) ) ;
INV     gate47  (.A(II13351), .Z(g8323) ) ;
INV     gate48  (.A(II13364), .Z(g8328) ) ;
INV     gate49  (.A(II13373), .Z(g8331) ) ;
INV     gate50  (.A(II13385), .Z(g8335) ) ;
INV     gate51  (.A(II13400), .Z(g8340) ) ;
INV     gate52  (.A(II13421), .Z(g8347) ) ;
INV     gate53  (.A(II13427), .Z(g8349) ) ;
INV     gate54  (.A(II13436), .Z(g8352) ) ;
INV     gate55  (.A(II13776), .Z(g8561) ) ;
INV     gate56  (.A(II13779), .Z(g8562) ) ;
INV     gate57  (.A(II13782), .Z(g8563) ) ;
INV     gate58  (.A(II13785), .Z(g8564) ) ;
INV     gate59  (.A(II13788), .Z(g8565) ) ;
INV     gate60  (.A(II13791), .Z(g8566) ) ;
INV     gate61  (.A(II14349), .Z(g8976) ) ;
INV     gate62  (.A(II14352), .Z(g8977) ) ;
INV     gate63  (.A(II14355), .Z(g8978) ) ;
INV     gate64  (.A(II14358), .Z(g8979) ) ;
INV     gate65  (.A(II14361), .Z(g8980) ) ;
INV     gate66  (.A(II14364), .Z(g8981) ) ;
INV     gate67  (.A(II14367), .Z(g8982) ) ;
INV     gate68  (.A(II14370), .Z(g8983) ) ;
INV     gate69  (.A(II14373), .Z(g8984) ) ;
INV     gate70  (.A(II14376), .Z(g8985) ) ;
INV     gate71  (.A(II14379), .Z(g8986) ) ;
INV     gate72  (.A(II14642), .Z(g9451) ) ;
INV     gate73  (.A(II15162), .Z(g9961) ) ;
INV     gate74  (.A(II15855), .Z(g10377) ) ;
INV     gate75  (.A(II15861), .Z(g10379) ) ;
INV     gate76  (.A(II15956), .Z(g10455) ) ;
INV     gate77  (.A(II15962), .Z(g10457) ) ;
INV     gate78  (.A(II15968), .Z(g10459) ) ;
INV     gate79  (.A(II15974), .Z(g10461) ) ;
INV     gate80  (.A(II15980), .Z(g10463) ) ;
INV     gate81  (.A(II15986), .Z(g10465) ) ;
INV     gate82  (.A(II16307), .Z(g10628) ) ;
INV     gate83  (.A(II16507), .Z(g10801) ) ;
INV     gate84  (.A(II16920), .Z(g11163) ) ;
INV     gate85  (.A(II16979), .Z(g11206) ) ;
INV     gate86  (.A(II17482), .Z(g11489) ) ;
INV     gate87  (.A(II10021), .Z(g6254) ) ;
DFF     gate88  (.D(g6254), .CP(CLK), .Q(g30) ) ;
INV     gate89  (.A(II10024), .Z(g6255) ) ;
DFF     gate90  (.D(g6255), .CP(CLK), .Q(g31) ) ;
INV     gate91  (.A(II17234), .Z(g11397) ) ;
DFF     gate92  (.D(g11397), .CP(CLK), .Q(g32) ) ;
INV     gate93  (.A(II16571), .Z(g10867) ) ;
DFF     gate94  (.D(g10867), .CP(CLK), .Q(g33) ) ;
INV     gate95  (.A(II16574), .Z(g10868) ) ;
DFF     gate96  (.D(g10868), .CP(CLK), .Q(g34) ) ;
INV     gate97  (.A(II16577), .Z(g10869) ) ;
DFF     gate98  (.D(g10869), .CP(CLK), .Q(g35) ) ;
INV     gate99  (.A(II16580), .Z(g10870) ) ;
DFF     gate100  (.D(g10870), .CP(CLK), .Q(g36) ) ;
INV     gate101  (.A(II16583), .Z(g10871) ) ;
DFF     gate102  (.D(g10871), .CP(CLK), .Q(g37) ) ;
INV     gate103  (.A(II16586), .Z(g10872) ) ;
DFF     gate104  (.D(g10872), .CP(CLK), .Q(g38) ) ;
INV     gate105  (.A(II16458), .Z(g10774) ) ;
DFF     gate106  (.D(g10774), .CP(CLK), .Q(g39) ) ;
INV     gate107  (.A(II16461), .Z(g10775) ) ;
DFF     gate108  (.D(g10775), .CP(CLK), .Q(g40) ) ;
INV     gate109  (.A(II10027), .Z(g6256) ) ;
DFF     gate110  (.D(g6256), .CP(CLK), .Q(g41) ) ;
INV     gate111  (.A(II10030), .Z(g6257) ) ;
DFF     gate112  (.D(g6257), .CP(CLK), .Q(g42) ) ;
INV     gate113  (.A(II10033), .Z(g6258) ) ;
DFF     gate114  (.D(g6258), .CP(CLK), .Q(g43) ) ;
INV     gate115  (.A(II10036), .Z(g6259) ) ;
DFF     gate116  (.D(g6259), .CP(CLK), .Q(g44) ) ;
INV     gate117  (.A(II10039), .Z(g6260) ) ;
DFF     gate118  (.D(g6260), .CP(CLK), .Q(g45) ) ;
INV     gate119  (.A(II10042), .Z(g6261) ) ;
DFF     gate120  (.D(g6261), .CP(CLK), .Q(g46) ) ;
INV     gate121  (.A(II10045), .Z(g6262) ) ;
DFF     gate122  (.D(g6262), .CP(CLK), .Q(g47) ) ;
INV     gate123  (.A(II10048), .Z(g6263) ) ;
DFF     gate124  (.D(g6263), .CP(CLK), .Q(g48) ) ;
INV     gate125  (.A(II10051), .Z(g6264) ) ;
DFF     gate126  (.D(g6264), .CP(CLK), .Q(g82) ) ;
INV     gate127  (.A(II10054), .Z(g6265) ) ;
DFF     gate128  (.D(g6265), .CP(CLK), .Q(g83) ) ;
INV     gate129  (.A(II10057), .Z(g6266) ) ;
DFF     gate130  (.D(g6266), .CP(CLK), .Q(g84) ) ;
INV     gate131  (.A(II10060), .Z(g6267) ) ;
DFF     gate132  (.D(g6267), .CP(CLK), .Q(g85) ) ;
INV     gate133  (.A(II10063), .Z(g6268) ) ;
DFF     gate134  (.D(g6268), .CP(CLK), .Q(g86) ) ;
INV     gate135  (.A(II10066), .Z(g6269) ) ;
DFF     gate136  (.D(g6269), .CP(CLK), .Q(g87) ) ;
INV     gate137  (.A(II10069), .Z(g6270) ) ;
DFF     gate138  (.D(g6270), .CP(CLK), .Q(g88) ) ;
INV     gate139  (.A(II10072), .Z(g6271) ) ;
DFF     gate140  (.D(g6271), .CP(CLK), .Q(g89) ) ;
INV     gate141  (.A(II10075), .Z(g6272) ) ;
DFF     gate142  (.D(g6272), .CP(CLK), .Q(g90) ) ;
INV     gate143  (.A(II10078), .Z(g6273) ) ;
DFF     gate144  (.D(g6273), .CP(CLK), .Q(g91) ) ;
INV     gate145  (.A(II10081), .Z(g6274) ) ;
DFF     gate146  (.D(g6274), .CP(CLK), .Q(g92) ) ;
INV     gate147  (.A(II10084), .Z(g6275) ) ;
DFF     gate148  (.D(g6275), .CP(CLK), .Q(g93) ) ;
INV     gate149  (.A(II10087), .Z(g6276) ) ;
DFF     gate150  (.D(g6276), .CP(CLK), .Q(g94) ) ;
INV     gate151  (.A(II10090), .Z(g6277) ) ;
DFF     gate152  (.D(g6277), .CP(CLK), .Q(g95) ) ;
INV     gate153  (.A(II10093), .Z(g6278) ) ;
DFF     gate154  (.D(g6278), .CP(CLK), .Q(g96) ) ;
INV     gate155  (.A(II10096), .Z(g6279) ) ;
DFF     gate156  (.D(g6279), .CP(CLK), .Q(g99) ) ;
INV     gate157  (.A(II10099), .Z(g6280) ) ;
DFF     gate158  (.D(g6280), .CP(CLK), .Q(g100) ) ;
INV     gate159  (.A(II10102), .Z(g6281) ) ;
DFF     gate160  (.D(g6281), .CP(CLK), .Q(g101) ) ;
INV     gate161  (.A(II10105), .Z(g6282) ) ;
DFF     gate162  (.D(g6282), .CP(CLK), .Q(g102) ) ;
INV     gate163  (.A(II10108), .Z(g6283) ) ;
DFF     gate164  (.D(g6283), .CP(CLK), .Q(g103) ) ;
INV     gate165  (.A(II10111), .Z(g6284) ) ;
DFF     gate166  (.D(g6284), .CP(CLK), .Q(g104) ) ;
INV     gate167  (.A(II10114), .Z(g6285) ) ;
DFF     gate168  (.D(g6285), .CP(CLK), .Q(g28) ) ;
INV     gate169  (.A(II10018), .Z(g6253) ) ;
DFF     gate170  (.D(g6253), .CP(CLK), .Q(g29) ) ;
INV     gate171  (.A(II7402), .Z(g4195) ) ;
DFF     gate172  (.D(g4195), .CP(CLK), .Q(g898) ) ;
INV     gate173  (.A(II7408), .Z(g4197) ) ;
DFF     gate174  (.D(g4197), .CP(CLK), .Q(g901) ) ;
INV     gate175  (.A(II7411), .Z(g4198) ) ;
DFF     gate176  (.D(g4198), .CP(CLK), .Q(g904) ) ;
INV     gate177  (.A(II7414), .Z(g4199) ) ;
DFF     gate178  (.D(g4199), .CP(CLK), .Q(g907) ) ;
INV     gate179  (.A(II7417), .Z(g4200) ) ;
DFF     gate180  (.D(g4200), .CP(CLK), .Q(g910) ) ;
INV     gate181  (.A(II7420), .Z(g4201) ) ;
DFF     gate182  (.D(g4201), .CP(CLK), .Q(g913) ) ;
INV     gate183  (.A(II7423), .Z(g4202) ) ;
DFF     gate184  (.D(g4202), .CP(CLK), .Q(g916) ) ;
INV     gate185  (.A(II7426), .Z(g4203) ) ;
DFF     gate186  (.D(g4203), .CP(CLK), .Q(g919) ) ;
INV     gate187  (.A(II7429), .Z(g4204) ) ;
DFF     gate188  (.D(g4204), .CP(CLK), .Q(g922) ) ;
INV     gate189  (.A(II7405), .Z(g4196) ) ;
DFF     gate190  (.D(g4196), .CP(CLK), .Q(g925) ) ;
INV     gate191  (.A(II17447), .Z(g11470) ) ;
DFF     gate192  (.D(g11470), .CP(CLK), .Q(g971) ) ;
INV     gate193  (.A(II17450), .Z(g11471) ) ;
DFF     gate194  (.D(g11471), .CP(CLK), .Q(g976) ) ;
INV     gate195  (.A(II17453), .Z(g11472) ) ;
DFF     gate196  (.D(g11472), .CP(CLK), .Q(g981) ) ;
INV     gate197  (.A(II17456), .Z(g11473) ) ;
DFF     gate198  (.D(g11473), .CP(CLK), .Q(g986) ) ;
INV     gate199  (.A(II17237), .Z(g11398) ) ;
DFF     gate200  (.D(g11398), .CP(CLK), .Q(g944) ) ;
INV     gate201  (.A(II17240), .Z(g11399) ) ;
DFF     gate202  (.D(g11399), .CP(CLK), .Q(g947) ) ;
INV     gate203  (.A(II17243), .Z(g11400) ) ;
DFF     gate204  (.D(g11400), .CP(CLK), .Q(g950) ) ;
INV     gate205  (.A(II17246), .Z(g11401) ) ;
DFF     gate206  (.D(g11401), .CP(CLK), .Q(g953) ) ;
INV     gate207  (.A(II17249), .Z(g11402) ) ;
DFF     gate208  (.D(g11402), .CP(CLK), .Q(g956) ) ;
INV     gate209  (.A(II17252), .Z(g11403) ) ;
DFF     gate210  (.D(g11403), .CP(CLK), .Q(g959) ) ;
INV     gate211  (.A(II17255), .Z(g11404) ) ;
DFF     gate212  (.D(g11404), .CP(CLK), .Q(g962) ) ;
INV     gate213  (.A(II17258), .Z(g11405) ) ;
DFF     gate214  (.D(g11405), .CP(CLK), .Q(g965) ) ;
INV     gate215  (.A(II17261), .Z(g11406) ) ;
DFF     gate216  (.D(g11406), .CP(CLK), .Q(g968) ) ;
INV     gate217  (.A(II7390), .Z(g4191) ) ;
DFF     gate218  (.D(g4191), .CP(CLK), .Q(g886) ) ;
INV     gate219  (.A(II7393), .Z(g4192) ) ;
DFF     gate220  (.D(g4192), .CP(CLK), .Q(g889) ) ;
INV     gate221  (.A(II7396), .Z(g4193) ) ;
DFF     gate222  (.D(g4193), .CP(CLK), .Q(g892) ) ;
INV     gate223  (.A(II7399), .Z(g4194) ) ;
DFF     gate224  (.D(g4194), .CP(CLK), .Q(g895) ) ;
INV     gate225  (.A(II13800), .Z(g8569) ) ;
DFF     gate226  (.D(g8569), .CP(CLK), .Q(g928) ) ;
INV     gate227  (.A(II13803), .Z(g8570) ) ;
DFF     gate228  (.D(g8570), .CP(CLK), .Q(g932) ) ;
INV     gate229  (.A(II13806), .Z(g8571) ) ;
DFF     gate230  (.D(g8571), .CP(CLK), .Q(g936) ) ;
INV     gate231  (.A(II13809), .Z(g8572) ) ;
DFF     gate232  (.D(g8572), .CP(CLK), .Q(g940) ) ;
INV     gate233  (.A(II8256), .Z(g4897) ) ;
DFF     gate234  (.D(g4897), .CP(CLK), .Q(g883) ) ;
DFF     gate235  (.D(g883), .CP(CLK), .Q(g882) ) ;
INV     gate236  (.A(II8253), .Z(g4896) ) ;
DFF     gate237  (.D(g4896), .CP(CLK), .Q(g878) ) ;
DFF     gate238  (.D(g878), .CP(CLK), .Q(g876) ) ;
INV     gate239  (.A(II16938), .Z(g11179) ) ;
DFF     gate240  (.D(g11179), .CP(CLK), .Q(g757) ) ;
INV     gate241  (.A(II10153), .Z(g6298) ) ;
DFF     gate242  (.D(g6298), .CP(CLK), .Q(g755) ) ;
DFF     gate243  (.D(g755), .CP(CLK), .Q(g756) ) ;
INV     gate244  (.A(II5754), .Z(g2639) ) ;
DFF     gate245  (.D(g2639), .CP(CLK), .Q(g745) ) ;
INV     gate246  (.A(II5751), .Z(g2638) ) ;
DFF     gate247  (.D(g2638), .CP(CLK), .Q(g746) ) ;
INV     gate248  (.A(II7330), .Z(g4171) ) ;
DFF     gate249  (.D(g4171), .CP(CLK), .Q(g750) ) ;
INV     gate250  (.A(II8250), .Z(g4895) ) ;
DFF     gate251  (.D(g4895), .CP(CLK), .Q(g754) ) ;
INV     gate252  (.A(II10801), .Z(g6797) ) ;
DFF     gate253  (.D(g6797), .CP(CLK), .Q(g758) ) ;
INV     gate254  (.A(II10804), .Z(g6798) ) ;
DFF     gate255  (.D(g6798), .CP(CLK), .Q(g762) ) ;
INV     gate256  (.A(II10807), .Z(g6799) ) ;
DFF     gate257  (.D(g6799), .CP(CLK), .Q(g766) ) ;
INV     gate258  (.A(II11540), .Z(g7288) ) ;
DFF     gate259  (.D(g7288), .CP(CLK), .Q(g770) ) ;
INV     gate260  (.A(II12520), .Z(g7785) ) ;
DFF     gate261  (.D(g7785), .CP(CLK), .Q(g774) ) ;
INV     gate262  (.A(II12930), .Z(g8076) ) ;
DFF     gate263  (.D(g8076), .CP(CLK), .Q(g778) ) ;
INV     gate264  (.A(II13191), .Z(g8273) ) ;
DFF     gate265  (.D(g8273), .CP(CLK), .Q(g782) ) ;
INV     gate266  (.A(II13606), .Z(g8436) ) ;
DFF     gate267  (.D(g8436), .CP(CLK), .Q(g786) ) ;
INV     gate268  (.A(II13794), .Z(g8567) ) ;
DFF     gate269  (.D(g8567), .CP(CLK), .Q(g790) ) ;
INV     gate270  (.A(II13197), .Z(g8275) ) ;
DFF     gate271  (.D(g8275), .CP(CLK), .Q(g865) ) ;
INV     gate272  (.A(II10810), .Z(g6800) ) ;
DFF     gate273  (.D(g6800), .CP(CLK), .Q(g794) ) ;
INV     gate274  (.A(II10813), .Z(g6801) ) ;
DFF     gate275  (.D(g6801), .CP(CLK), .Q(g798) ) ;
INV     gate276  (.A(II10816), .Z(g6802) ) ;
DFF     gate277  (.D(g6802), .CP(CLK), .Q(g802) ) ;
INV     gate278  (.A(II11543), .Z(g7289) ) ;
DFF     gate279  (.D(g7289), .CP(CLK), .Q(g806) ) ;
INV     gate280  (.A(II12523), .Z(g7786) ) ;
DFF     gate281  (.D(g7786), .CP(CLK), .Q(g810) ) ;
INV     gate282  (.A(II12933), .Z(g8077) ) ;
DFF     gate283  (.D(g8077), .CP(CLK), .Q(g814) ) ;
INV     gate284  (.A(II13194), .Z(g8274) ) ;
DFF     gate285  (.D(g8274), .CP(CLK), .Q(g818) ) ;
INV     gate286  (.A(II13609), .Z(g8437) ) ;
DFF     gate287  (.D(g8437), .CP(CLK), .Q(g822) ) ;
INV     gate288  (.A(II13797), .Z(g8568) ) ;
DFF     gate289  (.D(g8568), .CP(CLK), .Q(g826) ) ;
INV     gate290  (.A(II7363), .Z(g4182) ) ;
DFF     gate291  (.D(g4182), .CP(CLK), .Q(g829) ) ;
INV     gate292  (.A(II7366), .Z(g4183) ) ;
DFF     gate293  (.D(g4183), .CP(CLK), .Q(g833) ) ;
INV     gate294  (.A(II7369), .Z(g4184) ) ;
DFF     gate295  (.D(g4184), .CP(CLK), .Q(g837) ) ;
INV     gate296  (.A(II7372), .Z(g4185) ) ;
DFF     gate297  (.D(g4185), .CP(CLK), .Q(g841) ) ;
INV     gate298  (.A(II7375), .Z(g4186) ) ;
DFF     gate299  (.D(g4186), .CP(CLK), .Q(g845) ) ;
INV     gate300  (.A(II7378), .Z(g4187) ) ;
DFF     gate301  (.D(g4187), .CP(CLK), .Q(g849) ) ;
INV     gate302  (.A(II7381), .Z(g4188) ) ;
DFF     gate303  (.D(g4188), .CP(CLK), .Q(g853) ) ;
INV     gate304  (.A(II7384), .Z(g4189) ) ;
DFF     gate305  (.D(g4189), .CP(CLK), .Q(g857) ) ;
INV     gate306  (.A(II7387), .Z(g4190) ) ;
DFF     gate307  (.D(g4190), .CP(CLK), .Q(g861) ) ;
INV     gate308  (.A(II14964), .Z(g9821) ) ;
DFF     gate309  (.D(g9821), .CP(CLK), .Q(g874) ) ;
DFF     gate310  (.D(g874), .CP(CLK), .Q(g868) ) ;
INV     gate311  (.A(II14967), .Z(g9822) ) ;
DFF     gate312  (.D(g9822), .CP(CLK), .Q(g875) ) ;
DFF     gate313  (.D(g875), .CP(CLK), .Q(g869) ) ;
INV     gate314  (.A(II9120), .Z(g5653) ) ;
DFF     gate315  (.D(g5653), .CP(CLK), .Q(g590) ) ;
INV     gate316  (.A(II10135), .Z(g6292) ) ;
DFF     gate317  (.D(g6292), .CP(CLK), .Q(g584) ) ;
INV     gate318  (.A(II10138), .Z(g6293) ) ;
DFF     gate319  (.D(g6293), .CP(CLK), .Q(g585) ) ;
INV     gate320  (.A(II10141), .Z(g6294) ) ;
DFF     gate321  (.D(g6294), .CP(CLK), .Q(g586) ) ;
INV     gate322  (.A(II10144), .Z(g6295) ) ;
DFF     gate323  (.D(g6295), .CP(CLK), .Q(g587) ) ;
INV     gate324  (.A(II10147), .Z(g6296) ) ;
DFF     gate325  (.D(g6296), .CP(CLK), .Q(g588) ) ;
INV     gate326  (.A(II10150), .Z(g6297) ) ;
DFF     gate327  (.D(g6297), .CP(CLK), .Q(g589) ) ;
INV     gate328  (.A(II10117), .Z(g6286) ) ;
DFF     gate329  (.D(g6286), .CP(CLK), .Q(g578) ) ;
INV     gate330  (.A(II10120), .Z(g6287) ) ;
DFF     gate331  (.D(g6287), .CP(CLK), .Q(g579) ) ;
INV     gate332  (.A(II10123), .Z(g6288) ) ;
DFF     gate333  (.D(g6288), .CP(CLK), .Q(g580) ) ;
INV     gate334  (.A(II10126), .Z(g6289) ) ;
DFF     gate335  (.D(g6289), .CP(CLK), .Q(g581) ) ;
INV     gate336  (.A(II10129), .Z(g6290) ) ;
DFF     gate337  (.D(g6290), .CP(CLK), .Q(g582) ) ;
INV     gate338  (.A(II10132), .Z(g6291) ) ;
DFF     gate339  (.D(g6291), .CP(CLK), .Q(g583) ) ;
INV     gate340  (.A(II12415), .Z(g7750) ) ;
DFF     gate341  (.D(g7750), .CP(CLK), .Q(g253) ) ;
INV     gate342  (.A(II12421), .Z(g7752) ) ;
DFF     gate343  (.D(g7752), .CP(CLK), .Q(g256) ) ;
INV     gate344  (.A(II12424), .Z(g7753) ) ;
DFF     gate345  (.D(g7753), .CP(CLK), .Q(g257) ) ;
INV     gate346  (.A(II12427), .Z(g7754) ) ;
DFF     gate347  (.D(g7754), .CP(CLK), .Q(g258) ) ;
INV     gate348  (.A(II12430), .Z(g7755) ) ;
DFF     gate349  (.D(g7755), .CP(CLK), .Q(g259) ) ;
INV     gate350  (.A(II12433), .Z(g7756) ) ;
DFF     gate351  (.D(g7756), .CP(CLK), .Q(g260) ) ;
INV     gate352  (.A(II12436), .Z(g7757) ) ;
DFF     gate353  (.D(g7757), .CP(CLK), .Q(g261) ) ;
INV     gate354  (.A(II12439), .Z(g7758) ) ;
DFF     gate355  (.D(g7758), .CP(CLK), .Q(g262) ) ;
INV     gate356  (.A(II12442), .Z(g7759) ) ;
DFF     gate357  (.D(g7759), .CP(CLK), .Q(g254) ) ;
INV     gate358  (.A(II12418), .Z(g7751) ) ;
DFF     gate359  (.D(g7751), .CP(CLK), .Q(g255) ) ;
INV     gate360  (.A(II12403), .Z(g7746) ) ;
DFF     gate361  (.D(g7746), .CP(CLK), .Q(g143) ) ;
INV     gate362  (.A(II12406), .Z(g7747) ) ;
DFF     gate363  (.D(g7747), .CP(CLK), .Q(g166) ) ;
INV     gate364  (.A(II13568), .Z(g8418) ) ;
DFF     gate365  (.D(g8418), .CP(CLK), .Q(g139) ) ;
INV     gate366  (.A(II13571), .Z(g8419) ) ;
DFF     gate367  (.D(g8419), .CP(CLK), .Q(g135) ) ;
INV     gate368  (.A(II13574), .Z(g8420) ) ;
DFF     gate369  (.D(g8420), .CP(CLK), .Q(g131) ) ;
INV     gate370  (.A(II13577), .Z(g8421) ) ;
DFF     gate371  (.D(g8421), .CP(CLK), .Q(g127) ) ;
INV     gate372  (.A(II13580), .Z(g8422) ) ;
DFF     gate373  (.D(g8422), .CP(CLK), .Q(g170) ) ;
INV     gate374  (.A(II13583), .Z(g8423) ) ;
DFF     gate375  (.D(g8423), .CP(CLK), .Q(g174) ) ;
INV     gate376  (.A(II13586), .Z(g8424) ) ;
DFF     gate377  (.D(g8424), .CP(CLK), .Q(g162) ) ;
INV     gate378  (.A(II13589), .Z(g8425) ) ;
DFF     gate379  (.D(g8425), .CP(CLK), .Q(g158) ) ;
INV     gate380  (.A(II13592), .Z(g8426) ) ;
DFF     gate381  (.D(g8426), .CP(CLK), .Q(g153) ) ;
INV     gate382  (.A(II13595), .Z(g8427) ) ;
DFF     gate383  (.D(g8427), .CP(CLK), .Q(g148) ) ;
INV     gate384  (.A(II12409), .Z(g7748) ) ;
DFF     gate385  (.D(g7748), .CP(CLK), .Q(g178) ) ;
INV     gate386  (.A(II12412), .Z(g7749) ) ;
DFF     gate387  (.D(g7749), .CP(CLK), .Q(g182) ) ;
INV     gate388  (.A(II9087), .Z(g5642) ) ;
DFF     gate389  (.D(g5642), .CP(CLK), .Q(g126) ) ;
INV     gate390  (.A(II12445), .Z(g7760) ) ;
DFF     gate391  (.D(g7760), .CP(CLK), .Q(g263) ) ;
INV     gate392  (.A(II12448), .Z(g7761) ) ;
DFF     gate393  (.D(g7761), .CP(CLK), .Q(g266) ) ;
INV     gate394  (.A(II12451), .Z(g7762) ) ;
DFF     gate395  (.D(g7762), .CP(CLK), .Q(g269) ) ;
INV     gate396  (.A(II12454), .Z(g7763) ) ;
DFF     gate397  (.D(g7763), .CP(CLK), .Q(g272) ) ;
INV     gate398  (.A(II12457), .Z(g7764) ) ;
DFF     gate399  (.D(g7764), .CP(CLK), .Q(g275) ) ;
INV     gate400  (.A(II12460), .Z(g7765) ) ;
DFF     gate401  (.D(g7765), .CP(CLK), .Q(g278) ) ;
INV     gate402  (.A(II12463), .Z(g7766) ) ;
DFF     gate403  (.D(g7766), .CP(CLK), .Q(g281) ) ;
INV     gate404  (.A(II12466), .Z(g7767) ) ;
DFF     gate405  (.D(g7767), .CP(CLK), .Q(g284) ) ;
INV     gate406  (.A(II12469), .Z(g7768) ) ;
DFF     gate407  (.D(g7768), .CP(CLK), .Q(g287) ) ;
INV     gate408  (.A(II12472), .Z(g7769) ) ;
DFF     gate409  (.D(g7769), .CP(CLK), .Q(g290) ) ;
INV     gate410  (.A(II12475), .Z(g7770) ) ;
DFF     gate411  (.D(g7770), .CP(CLK), .Q(g293) ) ;
INV     gate412  (.A(II12478), .Z(g7771) ) ;
DFF     gate413  (.D(g7771), .CP(CLK), .Q(g296) ) ;
INV     gate414  (.A(II12481), .Z(g7772) ) ;
DFF     gate415  (.D(g7772), .CP(CLK), .Q(g299) ) ;
INV     gate416  (.A(II12484), .Z(g7773) ) ;
DFF     gate417  (.D(g7773), .CP(CLK), .Q(g302) ) ;
INV     gate418  (.A(II13188), .Z(g8272) ) ;
DFF     gate419  (.D(g8272), .CP(CLK), .Q(g123) ) ;
INV     gate420  (.A(II12400), .Z(g7745) ) ;
DFF     gate421  (.D(g7745), .CP(CLK), .Q(g119) ) ;
INV     gate422  (.A(II15127), .Z(g9930) ) ;
DFF     gate423  (.D(g9930), .CP(CLK), .Q(g611) ) ;
INV     gate424  (.A(II14077), .Z(g8780) ) ;
DFF     gate425  (.D(g8780), .CP(CLK), .Q(g617) ) ;
INV     gate426  (.A(II14955), .Z(g9818) ) ;
DFF     gate427  (.D(g9818), .CP(CLK), .Q(g591) ) ;
INV     gate428  (.A(II14958), .Z(g9819) ) ;
DFF     gate429  (.D(g9819), .CP(CLK), .Q(g599) ) ;
INV     gate430  (.A(II14961), .Z(g9820) ) ;
DFF     gate431  (.D(g9820), .CP(CLK), .Q(g605) ) ;
INV     gate432  (.A(II11537), .Z(g7287) ) ;
DFF     gate433  (.D(g7287), .CP(CLK), .Q(g630) ) ;
INV     gate434  (.A(II9123), .Z(g5654) ) ;
DFF     gate435  (.D(g5654), .CP(CLK), .Q(g631) ) ;
INV     gate436  (.A(II9126), .Z(g5655) ) ;
DFF     gate437  (.D(g5655), .CP(CLK), .Q(g632) ) ;
INV     gate438  (.A(II9129), .Z(g5656) ) ;
DFF     gate439  (.D(g5656), .CP(CLK), .Q(g635) ) ;
INV     gate440  (.A(II9132), .Z(g5657) ) ;
DFF     gate441  (.D(g5657), .CP(CLK), .Q(g627) ) ;
INV     gate442  (.A(II14080), .Z(g8781) ) ;
DFF     gate443  (.D(g8781), .CP(CLK), .Q(g636) ) ;
INV     gate444  (.A(II12907), .Z(g8063) ) ;
DFF     gate445  (.D(g8063), .CP(CLK), .Q(g639) ) ;
INV     gate446  (.A(II14519), .Z(g9338) ) ;
DFF     gate447  (.D(g9338), .CP(CLK), .Q(g622) ) ;
INV     gate448  (.A(II12910), .Z(g8064) ) ;
DFF     gate449  (.D(g8064), .CP(CLK), .Q(g643) ) ;
INV     gate450  (.A(II12913), .Z(g8065) ) ;
DFF     gate451  (.D(g8065), .CP(CLK), .Q(g646) ) ;
INV     gate452  (.A(II12916), .Z(g8066) ) ;
DFF     gate453  (.D(g8066), .CP(CLK), .Q(g650) ) ;
INV     gate454  (.A(II12919), .Z(g8067) ) ;
DFF     gate455  (.D(g8067), .CP(CLK), .Q(g654) ) ;
INV     gate456  (.A(II14522), .Z(g9339) ) ;
DFF     gate457  (.D(g9339), .CP(CLK), .Q(g658) ) ;
INV     gate458  (.A(II14525), .Z(g9340) ) ;
DFF     gate459  (.D(g9340), .CP(CLK), .Q(g668) ) ;
INV     gate460  (.A(II14528), .Z(g9341) ) ;
DFF     gate461  (.D(g9341), .CP(CLK), .Q(g677) ) ;
INV     gate462  (.A(II14531), .Z(g9342) ) ;
DFF     gate463  (.D(g9342), .CP(CLK), .Q(g686) ) ;
INV     gate464  (.A(II14534), .Z(g9343) ) ;
DFF     gate465  (.D(g9343), .CP(CLK), .Q(g695) ) ;
INV     gate466  (.A(II14537), .Z(g9344) ) ;
DFF     gate467  (.D(g9344), .CP(CLK), .Q(g704) ) ;
INV     gate468  (.A(II14540), .Z(g9345) ) ;
DFF     gate469  (.D(g9345), .CP(CLK), .Q(g713) ) ;
INV     gate470  (.A(II14543), .Z(g9346) ) ;
DFF     gate471  (.D(g9346), .CP(CLK), .Q(g722) ) ;
INV     gate472  (.A(II14546), .Z(g9347) ) ;
DFF     gate473  (.D(g9347), .CP(CLK), .Q(g731) ) ;
INV     gate474  (.A(II14083), .Z(g8782) ) ;
DFF     gate475  (.D(g8782), .CP(CLK), .Q(g664) ) ;
OR2     gate476  (.A(g8382), .B(g8068), .Z(g8428) ) ;
DFF     gate477  (.D(g8428), .CP(CLK), .Q(g673) ) ;
OR2     gate478  (.A(g8385), .B(g8069), .Z(g8429) ) ;
DFF     gate479  (.D(g8429), .CP(CLK), .Q(g682) ) ;
OR2     gate480  (.A(g8386), .B(g8070), .Z(g8430) ) ;
DFF     gate481  (.D(g8430), .CP(CLK), .Q(g691) ) ;
OR2     gate482  (.A(g8387), .B(g8071), .Z(g8431) ) ;
DFF     gate483  (.D(g8431), .CP(CLK), .Q(g700) ) ;
OR2     gate484  (.A(g8389), .B(g8072), .Z(g8432) ) ;
DFF     gate485  (.D(g8432), .CP(CLK), .Q(g709) ) ;
OR2     gate486  (.A(g8399), .B(g8073), .Z(g8433) ) ;
DFF     gate487  (.D(g8433), .CP(CLK), .Q(g718) ) ;
OR2     gate488  (.A(g8400), .B(g8074), .Z(g8434) ) ;
DFF     gate489  (.D(g8434), .CP(CLK), .Q(g727) ) ;
OR2     gate490  (.A(g8403), .B(g8075), .Z(g8435) ) ;
DFF     gate491  (.D(g8435), .CP(CLK), .Q(g736) ) ;
INV     gate492  (.A(II5740), .Z(g2613) ) ;
DFF     gate493  (.D(g2613), .CP(CLK), .Q(g8) ) ;
INV     gate494  (.A(II8247), .Z(g4894) ) ;
DFF     gate495  (.D(g4894), .CP(CLK), .Q(g17) ) ;
OR2     gate496  (.A(g11271), .B(g11164), .Z(g11324) ) ;
DFF     gate497  (.D(g11324), .CP(CLK), .Q(g481) ) ;
OR2     gate498  (.A(g11272), .B(g11171), .Z(g11331) ) ;
DFF     gate499  (.D(g11331), .CP(CLK), .Q(g486) ) ;
OR2     gate500  (.A(g11273), .B(g11172), .Z(g11332) ) ;
DFF     gate501  (.D(g11332), .CP(CLK), .Q(g491) ) ;
OR2     gate502  (.A(g11274), .B(g11173), .Z(g11333) ) ;
DFF     gate503  (.D(g11333), .CP(CLK), .Q(g496) ) ;
OR2     gate504  (.A(g11277), .B(g11174), .Z(g11334) ) ;
DFF     gate505  (.D(g11334), .CP(CLK), .Q(g501) ) ;
OR2     gate506  (.A(g11279), .B(g11175), .Z(g11335) ) ;
DFF     gate507  (.D(g11335), .CP(CLK), .Q(g506) ) ;
OR2     gate508  (.A(g11281), .B(g11176), .Z(g11336) ) ;
DFF     gate509  (.D(g11336), .CP(CLK), .Q(g511) ) ;
OR2     gate510  (.A(g11282), .B(g11177), .Z(g11337) ) ;
DFF     gate511  (.D(g11337), .CP(CLK), .Q(g516) ) ;
OR2     gate512  (.A(g11283), .B(g11178), .Z(g11338) ) ;
DFF     gate513  (.D(g11338), .CP(CLK), .Q(g476) ) ;
OR2     gate514  (.A(g11295), .B(g11165), .Z(g11325) ) ;
DFF     gate515  (.D(g11325), .CP(CLK), .Q(g542) ) ;
OR2     gate516  (.A(g11296), .B(g11166), .Z(g11326) ) ;
DFF     gate517  (.D(g11326), .CP(CLK), .Q(g538) ) ;
OR2     gate518  (.A(g11297), .B(g11167), .Z(g11327) ) ;
DFF     gate519  (.D(g11327), .CP(CLK), .Q(g534) ) ;
OR2     gate520  (.A(g11299), .B(g11168), .Z(g11328) ) ;
DFF     gate521  (.D(g11328), .CP(CLK), .Q(g530) ) ;
OR2     gate522  (.A(g11302), .B(g11169), .Z(g11329) ) ;
DFF     gate523  (.D(g11329), .CP(CLK), .Q(g525) ) ;
OR2     gate524  (.A(g11304), .B(g11170), .Z(g11330) ) ;
DFF     gate525  (.D(g11330), .CP(CLK), .Q(g521) ) ;
INV     gate526  (.A(II17435), .Z(g11466) ) ;
DFF     gate527  (.D(g11466), .CP(CLK), .Q(g456) ) ;
INV     gate528  (.A(II17438), .Z(g11467) ) ;
DFF     gate529  (.D(g11467), .CP(CLK), .Q(g461) ) ;
INV     gate530  (.A(II17441), .Z(g11468) ) ;
DFF     gate531  (.D(g11468), .CP(CLK), .Q(g466) ) ;
INV     gate532  (.A(II17444), .Z(g11469) ) ;
DFF     gate533  (.D(g11469), .CP(CLK), .Q(g471) ) ;
INV     gate534  (.A(II9090), .Z(g5643) ) ;
DFF     gate535  (.D(g5643), .CP(CLK), .Q(g305) ) ;
INV     gate536  (.A(II9096), .Z(g5645) ) ;
DFF     gate537  (.D(g5645), .CP(CLK), .Q(g315) ) ;
INV     gate538  (.A(II9099), .Z(g5646) ) ;
DFF     gate539  (.D(g5646), .CP(CLK), .Q(g318) ) ;
INV     gate540  (.A(II9102), .Z(g5647) ) ;
DFF     gate541  (.D(g5647), .CP(CLK), .Q(g321) ) ;
INV     gate542  (.A(II9105), .Z(g5648) ) ;
DFF     gate543  (.D(g5648), .CP(CLK), .Q(g324) ) ;
INV     gate544  (.A(II9108), .Z(g5649) ) ;
DFF     gate545  (.D(g5649), .CP(CLK), .Q(g327) ) ;
INV     gate546  (.A(II9111), .Z(g5650) ) ;
DFF     gate547  (.D(g5650), .CP(CLK), .Q(g330) ) ;
INV     gate548  (.A(II9114), .Z(g5651) ) ;
DFF     gate549  (.D(g5651), .CP(CLK), .Q(g333) ) ;
INV     gate550  (.A(II9117), .Z(g5652) ) ;
DFF     gate551  (.D(g5652), .CP(CLK), .Q(g309) ) ;
INV     gate552  (.A(II9093), .Z(g5644) ) ;
DFF     gate553  (.D(g5644), .CP(CLK), .Q(g312) ) ;
OR2     gate554  (.A(g11186), .B(g11018), .Z(g11256) ) ;
DFF     gate555  (.D(g11256), .CP(CLK), .Q(g426) ) ;
OR2     gate556  (.A(g11187), .B(g11025), .Z(g11263) ) ;
DFF     gate557  (.D(g11263), .CP(CLK), .Q(g386) ) ;
OR2     gate558  (.A(g11188), .B(g11026), .Z(g11264) ) ;
DFF     gate559  (.D(g11264), .CP(CLK), .Q(g391) ) ;
OR2     gate560  (.A(g11189), .B(g11027), .Z(g11265) ) ;
DFF     gate561  (.D(g11265), .CP(CLK), .Q(g396) ) ;
OR2     gate562  (.A(g11190), .B(g11028), .Z(g11266) ) ;
DFF     gate563  (.D(g11266), .CP(CLK), .Q(g401) ) ;
OR2     gate564  (.A(g11192), .B(g11029), .Z(g11267) ) ;
DFF     gate565  (.D(g11267), .CP(CLK), .Q(g406) ) ;
OR2     gate566  (.A(g11194), .B(g11030), .Z(g11268) ) ;
DFF     gate567  (.D(g11268), .CP(CLK), .Q(g411) ) ;
OR2     gate568  (.A(g11196), .B(g11031), .Z(g11269) ) ;
DFF     gate569  (.D(g11269), .CP(CLK), .Q(g416) ) ;
OR2     gate570  (.A(g11198), .B(g11032), .Z(g11270) ) ;
DFF     gate571  (.D(g11270), .CP(CLK), .Q(g421) ) ;
OR2     gate572  (.A(g11234), .B(g11019), .Z(g11257) ) ;
DFF     gate573  (.D(g11257), .CP(CLK), .Q(g452) ) ;
OR2     gate574  (.A(g11235), .B(g11020), .Z(g11258) ) ;
DFF     gate575  (.D(g11258), .CP(CLK), .Q(g448) ) ;
OR2     gate576  (.A(g11236), .B(g11021), .Z(g11259) ) ;
DFF     gate577  (.D(g11259), .CP(CLK), .Q(g444) ) ;
OR2     gate578  (.A(g11237), .B(g11022), .Z(g11260) ) ;
DFF     gate579  (.D(g11260), .CP(CLK), .Q(g440) ) ;
OR2     gate580  (.A(g11238), .B(g11023), .Z(g11261) ) ;
DFF     gate581  (.D(g11261), .CP(CLK), .Q(g435) ) ;
OR2     gate582  (.A(g11240), .B(g11024), .Z(g11262) ) ;
DFF     gate583  (.D(g11262), .CP(CLK), .Q(g431) ) ;
INV     gate584  (.A(II17368), .Z(g11439) ) ;
DFF     gate585  (.D(g11439), .CP(CLK), .Q(g369) ) ;
INV     gate586  (.A(II17371), .Z(g11440) ) ;
DFF     gate587  (.D(g11440), .CP(CLK), .Q(g374) ) ;
INV     gate588  (.A(II17374), .Z(g11441) ) ;
DFF     gate589  (.D(g11441), .CP(CLK), .Q(g378) ) ;
INV     gate590  (.A(II17377), .Z(g11442) ) ;
DFF     gate591  (.D(g11442), .CP(CLK), .Q(g382) ) ;
INV     gate592  (.A(II17761), .Z(g11653) ) ;
DFF     gate593  (.D(g11653), .CP(CLK), .Q(g336) ) ;
INV     gate594  (.A(II17537), .Z(g11506) ) ;
DFF     gate595  (.D(g11506), .CP(CLK), .Q(g348) ) ;
INV     gate596  (.A(II17540), .Z(g11507) ) ;
DFF     gate597  (.D(g11507), .CP(CLK), .Q(g351) ) ;
INV     gate598  (.A(II17543), .Z(g11508) ) ;
DFF     gate599  (.D(g11508), .CP(CLK), .Q(g354) ) ;
INV     gate600  (.A(II17546), .Z(g11509) ) ;
DFF     gate601  (.D(g11509), .CP(CLK), .Q(g357) ) ;
INV     gate602  (.A(II17549), .Z(g11510) ) ;
DFF     gate603  (.D(g11510), .CP(CLK), .Q(g360) ) ;
INV     gate604  (.A(II17552), .Z(g11511) ) ;
DFF     gate605  (.D(g11511), .CP(CLK), .Q(g363) ) ;
INV     gate606  (.A(II17555), .Z(g11512) ) ;
DFF     gate607  (.D(g11512), .CP(CLK), .Q(g366) ) ;
INV     gate608  (.A(II17558), .Z(g11513) ) ;
DFF     gate609  (.D(g11513), .CP(CLK), .Q(g342) ) ;
INV     gate610  (.A(II17534), .Z(g11505) ) ;
DFF     gate611  (.D(g11505), .CP(CLK), .Q(g339) ) ;
INV     gate612  (.A(II17730), .Z(g11642) ) ;
DFF     gate613  (.D(g11642), .CP(CLK), .Q(g345) ) ;
INV     gate614  (.A(II12487), .Z(g7774) ) ;
DFF     gate615  (.D(g7774), .CP(CLK), .Q(g49) ) ;
INV     gate616  (.A(II12496), .Z(g7777) ) ;
DFF     gate617  (.D(g7777), .CP(CLK), .Q(g52) ) ;
INV     gate618  (.A(II12499), .Z(g7778) ) ;
DFF     gate619  (.D(g7778), .CP(CLK), .Q(g55) ) ;
INV     gate620  (.A(II12502), .Z(g7779) ) ;
DFF     gate621  (.D(g7779), .CP(CLK), .Q(g58) ) ;
INV     gate622  (.A(II12505), .Z(g7780) ) ;
DFF     gate623  (.D(g7780), .CP(CLK), .Q(g61) ) ;
INV     gate624  (.A(II12508), .Z(g7781) ) ;
DFF     gate625  (.D(g7781), .CP(CLK), .Q(g64) ) ;
INV     gate626  (.A(II12511), .Z(g7782) ) ;
DFF     gate627  (.D(g7782), .CP(CLK), .Q(g67) ) ;
INV     gate628  (.A(II12514), .Z(g7783) ) ;
DFF     gate629  (.D(g7783), .CP(CLK), .Q(g70) ) ;
INV     gate630  (.A(II12517), .Z(g7784) ) ;
DFF     gate631  (.D(g7784), .CP(CLK), .Q(g73) ) ;
INV     gate632  (.A(II12490), .Z(g7775) ) ;
DFF     gate633  (.D(g7775), .CP(CLK), .Q(g76) ) ;
INV     gate634  (.A(II12493), .Z(g7776) ) ;
DFF     gate635  (.D(g7776), .CP(CLK), .Q(g79) ) ;
INV     gate636  (.A(II11531), .Z(g7285) ) ;
DFF     gate637  (.D(g7285), .CP(CLK), .Q(g113) ) ;
DFF     gate638  (.D(g113), .CP(CLK), .Q(g114) ) ;
INV     gate639  (.A(II10237), .Z(g6338) ) ;
DFF     gate640  (.D(g6338), .CP(CLK), .Q(g1955) ) ;
DFF     gate641  (.D(g1955), .CP(CLK), .Q(g1956) ) ;
DFF     gate642  (.D(g1956), .CP(CLK), .Q(g1957) ) ;
DFF     gate643  (.D(g1957), .CP(CLK), .Q(g1700) ) ;
INV     gate644  (.A(II10898), .Z(g6842) ) ;
DFF     gate645  (.D(g6842), .CP(CLK), .Q(g1696) ) ;
INV     gate646  (.A(II10901), .Z(g6843) ) ;
DFF     gate647  (.D(g6843), .CP(CLK), .Q(g1703) ) ;
INV     gate648  (.A(II8268), .Z(g4901) ) ;
DFF     gate649  (.D(g4901), .CP(CLK), .Q(g1710) ) ;
INV     gate650  (.A(II10231), .Z(g6336) ) ;
DFF     gate651  (.D(g6336), .CP(CLK), .Q(g1713) ) ;
INV     gate652  (.A(II10234), .Z(g6337) ) ;
DFF     gate653  (.D(g6337), .CP(CLK), .Q(g1718) ) ;
INV     gate654  (.A(II12595), .Z(g7810) ) ;
DFF     gate655  (.D(g7810), .CP(CLK), .Q(g1766) ) ;
INV     gate656  (.A(II12598), .Z(g7811) ) ;
DFF     gate657  (.D(g7811), .CP(CLK), .Q(g1771) ) ;
INV     gate658  (.A(II12601), .Z(g7812) ) ;
DFF     gate659  (.D(g7812), .CP(CLK), .Q(g1776) ) ;
INV     gate660  (.A(II12604), .Z(g7813) ) ;
DFF     gate661  (.D(g7813), .CP(CLK), .Q(g1781) ) ;
INV     gate662  (.A(II12607), .Z(g7814) ) ;
DFF     gate663  (.D(g7814), .CP(CLK), .Q(g1786) ) ;
INV     gate664  (.A(II12942), .Z(g8080) ) ;
DFF     gate665  (.D(g8080), .CP(CLK), .Q(g1791) ) ;
INV     gate666  (.A(II13212), .Z(g8280) ) ;
DFF     gate667  (.D(g8280), .CP(CLK), .Q(g1796) ) ;
INV     gate668  (.A(II13648), .Z(g8450) ) ;
DFF     gate669  (.D(g8450), .CP(CLK), .Q(g1801) ) ;
INV     gate670  (.A(II13812), .Z(g8573) ) ;
DFF     gate671  (.D(g8573), .CP(CLK), .Q(g1806) ) ;
INV     gate672  (.A(II10228), .Z(g6335) ) ;
DFF     gate673  (.D(g6335), .CP(CLK), .Q(g1711) ) ;
INV     gate674  (.A(II15088), .Z(g9895) ) ;
DFF     gate675  (.D(g9895), .CP(CLK), .Q(g1834) ) ;
INV     gate676  (.A(II13975), .Z(g8694) ) ;
DFF     gate677  (.D(g8694), .CP(CLK), .Q(g1840) ) ;
INV     gate678  (.A(II14976), .Z(g9825) ) ;
DFF     gate679  (.D(g9825), .CP(CLK), .Q(g1814) ) ;
INV     gate680  (.A(II14979), .Z(g9826) ) ;
DFF     gate681  (.D(g9826), .CP(CLK), .Q(g1822) ) ;
INV     gate682  (.A(II14982), .Z(g9827) ) ;
DFF     gate683  (.D(g9827), .CP(CLK), .Q(g1828) ) ;
INV     gate684  (.A(II11746), .Z(g7366) ) ;
DFF     gate685  (.D(g7366), .CP(CLK), .Q(g1848) ) ;
INV     gate686  (.A(II9171), .Z(g5670) ) ;
DFF     gate687  (.D(g5670), .CP(CLK), .Q(g1849) ) ;
INV     gate688  (.A(II9174), .Z(g5671) ) ;
DFF     gate689  (.D(g5671), .CP(CLK), .Q(g1850) ) ;
INV     gate690  (.A(II9177), .Z(g5672) ) ;
DFF     gate691  (.D(g5672), .CP(CLK), .Q(g1853) ) ;
INV     gate692  (.A(II9180), .Z(g5673) ) ;
DFF     gate693  (.D(g5673), .CP(CLK), .Q(g1845) ) ;
INV     gate694  (.A(II17265), .Z(g11408) ) ;
DFF     gate695  (.D(g11408), .CP(CLK), .Q(g1854) ) ;
INV     gate696  (.A(II17268), .Z(g11409) ) ;
DFF     gate697  (.D(g11409), .CP(CLK), .Q(g1857) ) ;
INV     gate698  (.A(II12610), .Z(g7815) ) ;
DFF     gate699  (.D(g7815), .CP(CLK), .Q(g1861) ) ;
INV     gate700  (.A(II12613), .Z(g7816) ) ;
DFF     gate701  (.D(g7816), .CP(CLK), .Q(g1864) ) ;
INV     gate702  (.A(II12616), .Z(g7817) ) ;
DFF     gate703  (.D(g7817), .CP(CLK), .Q(g1868) ) ;
INV     gate704  (.A(II14549), .Z(g9348) ) ;
DFF     gate705  (.D(g9348), .CP(CLK), .Q(g1872) ) ;
INV     gate706  (.A(II14552), .Z(g9349) ) ;
DFF     gate707  (.D(g9349), .CP(CLK), .Q(g1882) ) ;
INV     gate708  (.A(II14555), .Z(g9350) ) ;
DFF     gate709  (.D(g9350), .CP(CLK), .Q(g1891) ) ;
INV     gate710  (.A(II14558), .Z(g9351) ) ;
DFF     gate711  (.D(g9351), .CP(CLK), .Q(g1900) ) ;
INV     gate712  (.A(II14561), .Z(g9352) ) ;
DFF     gate713  (.D(g9352), .CP(CLK), .Q(g1909) ) ;
INV     gate714  (.A(II14564), .Z(g9353) ) ;
DFF     gate715  (.D(g9353), .CP(CLK), .Q(g1918) ) ;
INV     gate716  (.A(II14567), .Z(g9354) ) ;
DFF     gate717  (.D(g9354), .CP(CLK), .Q(g1927) ) ;
INV     gate718  (.A(II14570), .Z(g9355) ) ;
DFF     gate719  (.D(g9355), .CP(CLK), .Q(g1936) ) ;
INV     gate720  (.A(II14573), .Z(g9356) ) ;
DFF     gate721  (.D(g9356), .CP(CLK), .Q(g1945) ) ;
INV     gate722  (.A(II13978), .Z(g8695) ) ;
DFF     gate723  (.D(g8695), .CP(CLK), .Q(g1878) ) ;
OR2     gate724  (.A(g8097), .B(g7818), .Z(g8281) ) ;
DFF     gate725  (.D(g8281), .CP(CLK), .Q(g1887) ) ;
OR2     gate726  (.A(g8101), .B(g7819), .Z(g8282) ) ;
DFF     gate727  (.D(g8282), .CP(CLK), .Q(g1896) ) ;
OR2     gate728  (.A(g8098), .B(g7820), .Z(g8283) ) ;
DFF     gate729  (.D(g8283), .CP(CLK), .Q(g1905) ) ;
OR2     gate730  (.A(g8102), .B(g7821), .Z(g8284) ) ;
DFF     gate731  (.D(g8284), .CP(CLK), .Q(g1914) ) ;
OR2     gate732  (.A(g8104), .B(g7822), .Z(g8285) ) ;
DFF     gate733  (.D(g8285), .CP(CLK), .Q(g1923) ) ;
OR2     gate734  (.A(g8107), .B(g7823), .Z(g8286) ) ;
DFF     gate735  (.D(g8286), .CP(CLK), .Q(g1932) ) ;
OR2     gate736  (.A(g8117), .B(g7824), .Z(g8287) ) ;
DFF     gate737  (.D(g8287), .CP(CLK), .Q(g1941) ) ;
OR2     gate738  (.A(g8119), .B(g7825), .Z(g8288) ) ;
DFF     gate739  (.D(g8288), .CP(CLK), .Q(g1950) ) ;
INV     gate740  (.A(II8275), .Z(g4906) ) ;
DFF     gate741  (.D(g4906), .CP(CLK), .Q(g16) ) ;
INV     gate742  (.A(II5789), .Z(g2731) ) ;
DFF     gate743  (.D(g2731), .CP(CLK), .Q(g7) ) ;
INV     gate744  (.A(II10910), .Z(g6846) ) ;
DFF     gate745  (.D(g6846), .CP(CLK), .Q(g1736) ) ;
DFF     gate746  (.D(g1736), .CP(CLK), .Q(g1737) ) ;
INV     gate747  (.A(II16944), .Z(g11181) ) ;
DFF     gate748  (.D(g11181), .CP(CLK), .Q(g1648) ) ;
INV     gate749  (.A(II16947), .Z(g11182) ) ;
DFF     gate750  (.D(g11182), .CP(CLK), .Q(g1651) ) ;
INV     gate751  (.A(II16950), .Z(g11183) ) ;
DFF     gate752  (.D(g11183), .CP(CLK), .Q(g1642) ) ;
INV     gate753  (.A(II16953), .Z(g11184) ) ;
DFF     gate754  (.D(g11184), .CP(CLK), .Q(g1645) ) ;
INV     gate755  (.A(II10907), .Z(g6845) ) ;
DFF     gate756  (.D(g6845), .CP(CLK), .Q(g1610) ) ;
INV     gate757  (.A(II6504), .Z(g3329) ) ;
DFF     gate758  (.D(g3329), .CP(CLK), .Q(g1765) ) ;
INV     gate759  (.A(II16956), .Z(g11185) ) ;
DFF     gate760  (.D(g11185), .CP(CLK), .Q(g1811) ) ;
INV     gate761  (.A(II16604), .Z(g10878) ) ;
DFF     gate762  (.D(g10878), .CP(CLK), .Q(g1721) ) ;
INV     gate763  (.A(II16607), .Z(g10879) ) ;
DFF     gate764  (.D(g10879), .CP(CLK), .Q(g1724) ) ;
INV     gate765  (.A(II16610), .Z(g10880) ) ;
DFF     gate766  (.D(g10880), .CP(CLK), .Q(g1727) ) ;
INV     gate767  (.A(II16613), .Z(g10881) ) ;
DFF     gate768  (.D(g10881), .CP(CLK), .Q(g1730) ) ;
INV     gate769  (.A(II16616), .Z(g10882) ) ;
DFF     gate770  (.D(g10882), .CP(CLK), .Q(g1733) ) ;
INV     gate771  (.A(II9144), .Z(g5661) ) ;
DFF     gate772  (.D(g5661), .CP(CLK), .Q(g1738) ) ;
INV     gate773  (.A(II9147), .Z(g5662) ) ;
DFF     gate774  (.D(g5662), .CP(CLK), .Q(g1741) ) ;
INV     gate775  (.A(II9150), .Z(g5663) ) ;
DFF     gate776  (.D(g5663), .CP(CLK), .Q(g1744) ) ;
INV     gate777  (.A(II9153), .Z(g5664) ) ;
DFF     gate778  (.D(g5664), .CP(CLK), .Q(g1747) ) ;
INV     gate779  (.A(II9156), .Z(g5665) ) ;
DFF     gate780  (.D(g5665), .CP(CLK), .Q(g1750) ) ;
INV     gate781  (.A(II9159), .Z(g5666) ) ;
DFF     gate782  (.D(g5666), .CP(CLK), .Q(g1753) ) ;
INV     gate783  (.A(II9162), .Z(g5667) ) ;
DFF     gate784  (.D(g5667), .CP(CLK), .Q(g1756) ) ;
INV     gate785  (.A(II9165), .Z(g5668) ) ;
DFF     gate786  (.D(g5668), .CP(CLK), .Q(g1759) ) ;
INV     gate787  (.A(II9168), .Z(g5669) ) ;
DFF     gate788  (.D(g5669), .CP(CLK), .Q(g1762) ) ;
INV     gate789  (.A(II10240), .Z(g6339) ) ;
DFF     gate790  (.D(g6339), .CP(CLK), .Q(g1958) ) ;
INV     gate791  (.A(II4850), .Z(g2044) ) ;
DFF     gate792  (.D(g2044), .CP(CLK), .Q(g1810) ) ;
INV     gate793  (.A(II7468), .Z(g4217) ) ;
DFF     gate794  (.D(g4217), .CP(CLK), .Q(g1959) ) ;
INV     gate795  (.A(II8278), .Z(g4907) ) ;
DFF     gate796  (.D(g4907), .CP(CLK), .Q(g1707) ) ;
INV     gate797  (.A(II10904), .Z(g6844) ) ;
DFF     gate798  (.D(g6844), .CP(CLK), .Q(g1690) ) ;
INV     gate799  (.A(II7432), .Z(g4205) ) ;
DFF     gate800  (.D(g4205), .CP(CLK), .Q(g1170) ) ;
INV     gate801  (.A(II7444), .Z(g4209) ) ;
DFF     gate802  (.D(g4209), .CP(CLK), .Q(g1173) ) ;
INV     gate803  (.A(II7447), .Z(g4210) ) ;
DFF     gate804  (.D(g4210), .CP(CLK), .Q(g1176) ) ;
INV     gate805  (.A(II7450), .Z(g4211) ) ;
DFF     gate806  (.D(g4211), .CP(CLK), .Q(g1179) ) ;
INV     gate807  (.A(II7453), .Z(g4212) ) ;
DFF     gate808  (.D(g4212), .CP(CLK), .Q(g1182) ) ;
INV     gate809  (.A(II7456), .Z(g4213) ) ;
DFF     gate810  (.D(g4213), .CP(CLK), .Q(g1185) ) ;
INV     gate811  (.A(II7459), .Z(g4214) ) ;
DFF     gate812  (.D(g4214), .CP(CLK), .Q(g1188) ) ;
INV     gate813  (.A(II7462), .Z(g4215) ) ;
DFF     gate814  (.D(g4215), .CP(CLK), .Q(g1191) ) ;
INV     gate815  (.A(II7465), .Z(g4216) ) ;
DFF     gate816  (.D(g4216), .CP(CLK), .Q(g1194) ) ;
INV     gate817  (.A(II7435), .Z(g4206) ) ;
DFF     gate818  (.D(g4206), .CP(CLK), .Q(g1197) ) ;
INV     gate819  (.A(II7438), .Z(g4207) ) ;
DFF     gate820  (.D(g4207), .CP(CLK), .Q(g1200) ) ;
INV     gate821  (.A(II7441), .Z(g4208) ) ;
DFF     gate822  (.D(g4208), .CP(CLK), .Q(g1203) ) ;
INV     gate823  (.A(II10201), .Z(g6314) ) ;
DFF     gate824  (.D(g6314), .CP(CLK), .Q(g1169) ) ;
INV     gate825  (.A(II17633), .Z(g11593) ) ;
DFF     gate826  (.D(g11593), .CP(CLK), .Q(g108) ) ;
INV     gate827  (.A(II17764), .Z(g11654) ) ;
DFF     gate828  (.D(g11654), .CP(CLK), .Q(g1336) ) ;
INV     gate829  (.A(II17767), .Z(g11655) ) ;
DFF     gate830  (.D(g11655), .CP(CLK), .Q(g1341) ) ;
INV     gate831  (.A(II17770), .Z(g11656) ) ;
DFF     gate832  (.D(g11656), .CP(CLK), .Q(g1346) ) ;
INV     gate833  (.A(II17773), .Z(g11657) ) ;
DFF     gate834  (.D(g11657), .CP(CLK), .Q(g1351) ) ;
INV     gate835  (.A(II8259), .Z(g4898) ) ;
DFF     gate836  (.D(g4898), .CP(CLK), .Q(g1206) ) ;
DFF     gate837  (.D(g1206), .CP(CLK), .Q(g1361) ) ;
INV     gate838  (.A(II14973), .Z(g9824) ) ;
DFF     gate839  (.D(g9824), .CP(CLK), .Q(g1360) ) ;
DFF     gate840  (.D(g1360), .CP(CLK), .Q(g1216) ) ;
INV     gate841  (.A(II14970), .Z(g9823) ) ;
DFF     gate842  (.D(g9823), .CP(CLK), .Q(g1217) ) ;
DFF     gate843  (.D(g1217), .CP(CLK), .Q(g1212) ) ;
INV     gate844  (.A(II16589), .Z(g10873) ) ;
DFF     gate845  (.D(g10873), .CP(CLK), .Q(g1209) ) ;
INV     gate846  (.A(II10204), .Z(g6315) ) ;
DFF     gate847  (.D(g6315), .CP(CLK), .Q(g1215) ) ;
INV     gate848  (.A(II10221), .Z(g6330) ) ;
DFF     gate849  (.D(g6330), .CP(CLK), .Q(g1357) ) ;
INV     gate850  (.A(II9141), .Z(g5660) ) ;
DFF     gate851  (.D(g5660), .CP(CLK), .Q(g1289) ) ;
OR2     gate852  (.A(g7130), .B(g11407), .Z(g11443) ) ;
DFF     gate853  (.D(g11443), .CP(CLK), .Q(g1275) ) ;
OR2     gate854  (.A(g7131), .B(g6322), .Z(g7296) ) ;
DFF     gate855  (.D(g7296), .CP(CLK), .Q(g1235) ) ;
OR2     gate856  (.A(g7132), .B(g6323), .Z(g7297) ) ;
DFF     gate857  (.D(g7297), .CP(CLK), .Q(g1240) ) ;
OR2     gate858  (.A(g7136), .B(g6324), .Z(g7298) ) ;
DFF     gate859  (.D(g7298), .CP(CLK), .Q(g1245) ) ;
OR2     gate860  (.A(g7138), .B(g6325), .Z(g7299) ) ;
DFF     gate861  (.D(g7299), .CP(CLK), .Q(g1250) ) ;
OR2     gate862  (.A(g7139), .B(g6326), .Z(g7300) ) ;
DFF     gate863  (.D(g7300), .CP(CLK), .Q(g1255) ) ;
OR2     gate864  (.A(g7140), .B(g6327), .Z(g7301) ) ;
DFF     gate865  (.D(g7301), .CP(CLK), .Q(g1260) ) ;
OR2     gate866  (.A(g7141), .B(g6328), .Z(g7302) ) ;
DFF     gate867  (.D(g7302), .CP(CLK), .Q(g1265) ) ;
OR2     gate868  (.A(g7145), .B(g6329), .Z(g7303) ) ;
DFF     gate869  (.D(g7303), .CP(CLK), .Q(g1270) ) ;
OR2     gate870  (.A(g7046), .B(g6316), .Z(g7290) ) ;
DFF     gate871  (.D(g7290), .CP(CLK), .Q(g1304) ) ;
OR2     gate872  (.A(g7050), .B(g6317), .Z(g7291) ) ;
DFF     gate873  (.D(g7291), .CP(CLK), .Q(g1300) ) ;
OR2     gate874  (.A(g7055), .B(g6318), .Z(g7292) ) ;
DFF     gate875  (.D(g7292), .CP(CLK), .Q(g1296) ) ;
OR2     gate876  (.A(g7063), .B(g6319), .Z(g7293) ) ;
DFF     gate877  (.D(g7293), .CP(CLK), .Q(g1292) ) ;
OR2     gate878  (.A(g7068), .B(g6320), .Z(g7294) ) ;
DFF     gate879  (.D(g7294), .CP(CLK), .Q(g1284) ) ;
OR2     gate880  (.A(g7071), .B(g6321), .Z(g7295) ) ;
DFF     gate881  (.D(g7295), .CP(CLK), .Q(g1280) ) ;
INV     gate882  (.A(II13200), .Z(g8276) ) ;
DFF     gate883  (.D(g8276), .CP(CLK), .Q(g1218) ) ;
INV     gate884  (.A(II13203), .Z(g8277) ) ;
DFF     gate885  (.D(g8277), .CP(CLK), .Q(g1223) ) ;
INV     gate886  (.A(II13206), .Z(g8278) ) ;
DFF     gate887  (.D(g8278), .CP(CLK), .Q(g1227) ) ;
INV     gate888  (.A(II13209), .Z(g8279) ) ;
DFF     gate889  (.D(g8279), .CP(CLK), .Q(g1231) ) ;
INV     gate890  (.A(II10864), .Z(g6818) ) ;
DFF     gate891  (.D(g6818), .CP(CLK), .Q(g1356) ) ;
DFF     gate892  (.D(g1356), .CP(CLK), .Q(g1317) ) ;
INV     gate893  (.A(II17701), .Z(g11629) ) ;
DFF     gate894  (.D(g11629), .CP(CLK), .Q(g1314) ) ;
INV     gate895  (.A(II17704), .Z(g11630) ) ;
DFF     gate896  (.D(g11630), .CP(CLK), .Q(g1318) ) ;
INV     gate897  (.A(II17707), .Z(g11631) ) ;
DFF     gate898  (.D(g11631), .CP(CLK), .Q(g1321) ) ;
INV     gate899  (.A(II17710), .Z(g11632) ) ;
DFF     gate900  (.D(g11632), .CP(CLK), .Q(g1324) ) ;
INV     gate901  (.A(II17713), .Z(g11633) ) ;
DFF     gate902  (.D(g11633), .CP(CLK), .Q(g1327) ) ;
INV     gate903  (.A(II17716), .Z(g11634) ) ;
DFF     gate904  (.D(g11634), .CP(CLK), .Q(g1330) ) ;
INV     gate905  (.A(II17719), .Z(g11635) ) ;
DFF     gate906  (.D(g11635), .CP(CLK), .Q(g1333) ) ;
INV     gate907  (.A(II17695), .Z(g11627) ) ;
DFF     gate908  (.D(g11627), .CP(CLK), .Q(g1308) ) ;
INV     gate909  (.A(II17698), .Z(g11628) ) ;
DFF     gate910  (.D(g11628), .CP(CLK), .Q(g1311) ) ;
INV     gate911  (.A(II12526), .Z(g7787) ) ;
DFF     gate912  (.D(g7787), .CP(CLK), .Q(g1035) ) ;
INV     gate913  (.A(II12535), .Z(g7790) ) ;
DFF     gate914  (.D(g7790), .CP(CLK), .Q(g1047) ) ;
INV     gate915  (.A(II12538), .Z(g7791) ) ;
DFF     gate916  (.D(g7791), .CP(CLK), .Q(g1050) ) ;
INV     gate917  (.A(II12541), .Z(g7792) ) ;
DFF     gate918  (.D(g7792), .CP(CLK), .Q(g1053) ) ;
INV     gate919  (.A(II12544), .Z(g7793) ) ;
DFF     gate920  (.D(g7793), .CP(CLK), .Q(g1056) ) ;
INV     gate921  (.A(II12547), .Z(g7794) ) ;
DFF     gate922  (.D(g7794), .CP(CLK), .Q(g1059) ) ;
INV     gate923  (.A(II12550), .Z(g7795) ) ;
DFF     gate924  (.D(g7795), .CP(CLK), .Q(g1062) ) ;
INV     gate925  (.A(II12553), .Z(g7796) ) ;
DFF     gate926  (.D(g7796), .CP(CLK), .Q(g1065) ) ;
INV     gate927  (.A(II12556), .Z(g7797) ) ;
DFF     gate928  (.D(g7797), .CP(CLK), .Q(g1038) ) ;
INV     gate929  (.A(II12529), .Z(g7788) ) ;
DFF     gate930  (.D(g7788), .CP(CLK), .Q(g1041) ) ;
INV     gate931  (.A(II12532), .Z(g7789) ) ;
DFF     gate932  (.D(g7789), .CP(CLK), .Q(g1044) ) ;
INV     gate933  (.A(II10819), .Z(g6803) ) ;
DFF     gate934  (.D(g6803), .CP(CLK), .Q(g1068) ) ;
INV     gate935  (.A(II10828), .Z(g6806) ) ;
DFF     gate936  (.D(g6806), .CP(CLK), .Q(g1080) ) ;
INV     gate937  (.A(II10831), .Z(g6807) ) ;
DFF     gate938  (.D(g6807), .CP(CLK), .Q(g1083) ) ;
INV     gate939  (.A(II10834), .Z(g6808) ) ;
DFF     gate940  (.D(g6808), .CP(CLK), .Q(g1086) ) ;
INV     gate941  (.A(II10837), .Z(g6809) ) ;
DFF     gate942  (.D(g6809), .CP(CLK), .Q(g1089) ) ;
INV     gate943  (.A(II10840), .Z(g6810) ) ;
DFF     gate944  (.D(g6810), .CP(CLK), .Q(g1092) ) ;
INV     gate945  (.A(II10843), .Z(g6811) ) ;
DFF     gate946  (.D(g6811), .CP(CLK), .Q(g1095) ) ;
INV     gate947  (.A(II10846), .Z(g6812) ) ;
DFF     gate948  (.D(g6812), .CP(CLK), .Q(g1098) ) ;
INV     gate949  (.A(II10849), .Z(g6813) ) ;
DFF     gate950  (.D(g6813), .CP(CLK), .Q(g1074) ) ;
INV     gate951  (.A(II10822), .Z(g6804) ) ;
DFF     gate952  (.D(g6804), .CP(CLK), .Q(g1071) ) ;
INV     gate953  (.A(II10825), .Z(g6805) ) ;
DFF     gate954  (.D(g6805), .CP(CLK), .Q(g1077) ) ;
INV     gate955  (.A(II12559), .Z(g7798) ) ;
DFF     gate956  (.D(g7798), .CP(CLK), .Q(g1027) ) ;
INV     gate957  (.A(II12568), .Z(g7801) ) ;
DFF     gate958  (.D(g7801), .CP(CLK), .Q(g995) ) ;
INV     gate959  (.A(II12571), .Z(g7802) ) ;
DFF     gate960  (.D(g7802), .CP(CLK), .Q(g991) ) ;
INV     gate961  (.A(II12574), .Z(g7803) ) ;
DFF     gate962  (.D(g7803), .CP(CLK), .Q(g1003) ) ;
INV     gate963  (.A(II12577), .Z(g7804) ) ;
DFF     gate964  (.D(g7804), .CP(CLK), .Q(g999) ) ;
INV     gate965  (.A(II12580), .Z(g7805) ) ;
DFF     gate966  (.D(g7805), .CP(CLK), .Q(g1011) ) ;
INV     gate967  (.A(II12583), .Z(g7806) ) ;
DFF     gate968  (.D(g7806), .CP(CLK), .Q(g1007) ) ;
INV     gate969  (.A(II12586), .Z(g7807) ) ;
DFF     gate970  (.D(g7807), .CP(CLK), .Q(g1019) ) ;
INV     gate971  (.A(II12589), .Z(g7808) ) ;
DFF     gate972  (.D(g7808), .CP(CLK), .Q(g1015) ) ;
INV     gate973  (.A(II12562), .Z(g7799) ) ;
DFF     gate974  (.D(g7799), .CP(CLK), .Q(g1023) ) ;
INV     gate975  (.A(II12565), .Z(g7800) ) ;
DFF     gate976  (.D(g7800), .CP(CLK), .Q(g1032) ) ;
INV     gate977  (.A(II16941), .Z(g11180) ) ;
DFF     gate978  (.D(g11180), .CP(CLK), .Q(g105) ) ;
INV     gate979  (.A(II10156), .Z(g6299) ) ;
DFF     gate980  (.D(g6299), .CP(CLK), .Q(g1117) ) ;
INV     gate981  (.A(II10177), .Z(g6306) ) ;
DFF     gate982  (.D(g6306), .CP(CLK), .Q(g1121) ) ;
INV     gate983  (.A(II10180), .Z(g6307) ) ;
DFF     gate984  (.D(g6307), .CP(CLK), .Q(g1125) ) ;
INV     gate985  (.A(II10183), .Z(g6308) ) ;
DFF     gate986  (.D(g6308), .CP(CLK), .Q(g1129) ) ;
INV     gate987  (.A(II10186), .Z(g6309) ) ;
DFF     gate988  (.D(g6309), .CP(CLK), .Q(g1133) ) ;
INV     gate989  (.A(II10189), .Z(g6310) ) ;
DFF     gate990  (.D(g6310), .CP(CLK), .Q(g1137) ) ;
INV     gate991  (.A(II10192), .Z(g6311) ) ;
DFF     gate992  (.D(g6311), .CP(CLK), .Q(g1141) ) ;
INV     gate993  (.A(II10195), .Z(g6312) ) ;
DFF     gate994  (.D(g6312), .CP(CLK), .Q(g1145) ) ;
INV     gate995  (.A(II10198), .Z(g6313) ) ;
DFF     gate996  (.D(g6313), .CP(CLK), .Q(g1113) ) ;
INV     gate997  (.A(II10159), .Z(g6300) ) ;
DFF     gate998  (.D(g6300), .CP(CLK), .Q(g1166) ) ;
INV     gate999  (.A(II10162), .Z(g6301) ) ;
DFF     gate1000  (.D(g6301), .CP(CLK), .Q(g1163) ) ;
INV     gate1001  (.A(II10165), .Z(g6302) ) ;
DFF     gate1002  (.D(g6302), .CP(CLK), .Q(g1160) ) ;
INV     gate1003  (.A(II10168), .Z(g6303) ) ;
DFF     gate1004  (.D(g6303), .CP(CLK), .Q(g1157) ) ;
INV     gate1005  (.A(II10171), .Z(g6304) ) ;
DFF     gate1006  (.D(g6304), .CP(CLK), .Q(g1153) ) ;
INV     gate1007  (.A(II10174), .Z(g6305) ) ;
DFF     gate1008  (.D(g6305), .CP(CLK), .Q(g1149) ) ;
INV     gate1009  (.A(II10852), .Z(g6814) ) ;
DFF     gate1010  (.D(g6814), .CP(CLK), .Q(g1101) ) ;
INV     gate1011  (.A(II10855), .Z(g6815) ) ;
DFF     gate1012  (.D(g6815), .CP(CLK), .Q(g1104) ) ;
INV     gate1013  (.A(II10858), .Z(g6816) ) ;
DFF     gate1014  (.D(g6816), .CP(CLK), .Q(g1107) ) ;
INV     gate1015  (.A(II10861), .Z(g6817) ) ;
DFF     gate1016  (.D(g6817), .CP(CLK), .Q(g1110) ) ;
INV     gate1017  (.A(II17657), .Z(g11611) ) ;
DFF     gate1018  (.D(g11611), .CP(CLK), .Q(g1618) ) ;
INV     gate1019  (.A(II14176), .Z(g8868) ) ;
DFF     gate1020  (.D(g8868), .CP(CLK), .Q(g1615) ) ;
INV     gate1021  (.A(II14179), .Z(g8869) ) ;
DFF     gate1022  (.D(g8869), .CP(CLK), .Q(g1621) ) ;
INV     gate1023  (.A(II14182), .Z(g8870) ) ;
DFF     gate1024  (.D(g8870), .CP(CLK), .Q(g1624) ) ;
INV     gate1025  (.A(II14185), .Z(g8871) ) ;
DFF     gate1026  (.D(g8871), .CP(CLK), .Q(g1627) ) ;
INV     gate1027  (.A(II14188), .Z(g8872) ) ;
DFF     gate1028  (.D(g8872), .CP(CLK), .Q(g1630) ) ;
INV     gate1029  (.A(II14191), .Z(g8873) ) ;
DFF     gate1030  (.D(g8873), .CP(CLK), .Q(g1633) ) ;
INV     gate1031  (.A(II14194), .Z(g8874) ) ;
DFF     gate1032  (.D(g8874), .CP(CLK), .Q(g1636) ) ;
INV     gate1033  (.A(II13642), .Z(g8448) ) ;
DFF     gate1034  (.D(g8448), .CP(CLK), .Q(g1639) ) ;
INV     gate1035  (.A(II13645), .Z(g8449) ) ;
DFF     gate1036  (.D(g8449), .CP(CLK), .Q(g1512) ) ;
INV     gate1037  (.A(II17636), .Z(g11594) ) ;
DFF     gate1038  (.D(g11594), .CP(CLK), .Q(g1448) ) ;
INV     gate1039  (.A(II14382), .Z(g8987) ) ;
DFF     gate1040  (.D(g8987), .CP(CLK), .Q(g1444) ) ;
INV     gate1041  (.A(II14385), .Z(g8988) ) ;
DFF     gate1042  (.D(g8988), .CP(CLK), .Q(g1440) ) ;
INV     gate1043  (.A(II14388), .Z(g8989) ) ;
DFF     gate1044  (.D(g8989), .CP(CLK), .Q(g1436) ) ;
INV     gate1045  (.A(II14391), .Z(g8990) ) ;
DFF     gate1046  (.D(g8990), .CP(CLK), .Q(g1432) ) ;
INV     gate1047  (.A(II14394), .Z(g8991) ) ;
DFF     gate1048  (.D(g8991), .CP(CLK), .Q(g1403) ) ;
INV     gate1049  (.A(II14397), .Z(g8992) ) ;
DFF     gate1050  (.D(g8992), .CP(CLK), .Q(g1428) ) ;
INV     gate1051  (.A(II14400), .Z(g8993) ) ;
DFF     gate1052  (.D(g8993), .CP(CLK), .Q(g1407) ) ;
INV     gate1053  (.A(II11638), .Z(g7330) ) ;
DFF     gate1054  (.D(g7330), .CP(CLK), .Q(g1424) ) ;
INV     gate1055  (.A(II11641), .Z(g7331) ) ;
DFF     gate1056  (.D(g7331), .CP(CLK), .Q(g1411) ) ;
INV     gate1057  (.A(II11644), .Z(g7332) ) ;
DFF     gate1058  (.D(g7332), .CP(CLK), .Q(g1419) ) ;
INV     gate1059  (.A(II11647), .Z(g7333) ) ;
DFF     gate1060  (.D(g7333), .CP(CLK), .Q(g1515) ) ;
INV     gate1061  (.A(II11650), .Z(g7334) ) ;
DFF     gate1062  (.D(g7334), .CP(CLK), .Q(g1520) ) ;
INV     gate1063  (.A(II11653), .Z(g7335) ) ;
DFF     gate1064  (.D(g7335), .CP(CLK), .Q(g1415) ) ;
INV     gate1065  (.A(II11626), .Z(g7326) ) ;
DFF     gate1066  (.D(g7326), .CP(CLK), .Q(g1453) ) ;
INV     gate1067  (.A(II11629), .Z(g7327) ) ;
DFF     gate1068  (.D(g7327), .CP(CLK), .Q(g1458) ) ;
INV     gate1069  (.A(II13612), .Z(g8438) ) ;
DFF     gate1070  (.D(g8438), .CP(CLK), .Q(g1462) ) ;
INV     gate1071  (.A(II13615), .Z(g8439) ) ;
DFF     gate1072  (.D(g8439), .CP(CLK), .Q(g1466) ) ;
INV     gate1073  (.A(II13618), .Z(g8440) ) ;
DFF     gate1074  (.D(g8440), .CP(CLK), .Q(g1470) ) ;
INV     gate1075  (.A(II13621), .Z(g8441) ) ;
DFF     gate1076  (.D(g8441), .CP(CLK), .Q(g1474) ) ;
INV     gate1077  (.A(II13624), .Z(g8442) ) ;
DFF     gate1078  (.D(g8442), .CP(CLK), .Q(g1478) ) ;
INV     gate1079  (.A(II13627), .Z(g8443) ) ;
DFF     gate1080  (.D(g8443), .CP(CLK), .Q(g1482) ) ;
INV     gate1081  (.A(II13630), .Z(g8444) ) ;
DFF     gate1082  (.D(g8444), .CP(CLK), .Q(g1486) ) ;
INV     gate1083  (.A(II13633), .Z(g8445) ) ;
DFF     gate1084  (.D(g8445), .CP(CLK), .Q(g1490) ) ;
INV     gate1085  (.A(II13636), .Z(g8446) ) ;
DFF     gate1086  (.D(g8446), .CP(CLK), .Q(g1494) ) ;
INV     gate1087  (.A(II13639), .Z(g8447) ) ;
DFF     gate1088  (.D(g8447), .CP(CLK), .Q(g1499) ) ;
INV     gate1089  (.A(II11632), .Z(g7328) ) ;
DFF     gate1090  (.D(g7328), .CP(CLK), .Q(g1504) ) ;
INV     gate1091  (.A(II11635), .Z(g7329) ) ;
DFF     gate1092  (.D(g7329), .CP(CLK), .Q(g1508) ) ;
INV     gate1093  (.A(II11608), .Z(g7320) ) ;
DFF     gate1094  (.D(g7320), .CP(CLK), .Q(g1393) ) ;
INV     gate1095  (.A(II12592), .Z(g7809) ) ;
DFF     gate1096  (.D(g7809), .CP(CLK), .Q(g1394) ) ;
INV     gate1097  (.A(II11611), .Z(g7321) ) ;
DFF     gate1098  (.D(g7321), .CP(CLK), .Q(g115) ) ;
INV     gate1099  (.A(II11560), .Z(g7304) ) ;
DFF     gate1100  (.D(g7304), .CP(CLK), .Q(g201) ) ;
INV     gate1101  (.A(II10873), .Z(g6825) ) ;
DFF     gate1102  (.D(g6825), .CP(CLK), .Q(g1374) ) ;
INV     gate1103  (.A(II10885), .Z(g6835) ) ;
DFF     gate1104  (.D(g6835), .CP(CLK), .Q(g197) ) ;
INV     gate1105  (.A(II10888), .Z(g6836) ) ;
DFF     gate1106  (.D(g6836), .CP(CLK), .Q(g1389) ) ;
INV     gate1107  (.A(II10891), .Z(g6837) ) ;
DFF     gate1108  (.D(g6837), .CP(CLK), .Q(g192) ) ;
INV     gate1109  (.A(II11614), .Z(g7322) ) ;
DFF     gate1110  (.D(g7322), .CP(CLK), .Q(g1397) ) ;
INV     gate1111  (.A(II11617), .Z(g7323) ) ;
DFF     gate1112  (.D(g7323), .CP(CLK), .Q(g248) ) ;
INV     gate1113  (.A(II11620), .Z(g7324) ) ;
DFF     gate1114  (.D(g7324), .CP(CLK), .Q(g1400) ) ;
INV     gate1115  (.A(II11623), .Z(g7325) ) ;
DFF     gate1116  (.D(g7325), .CP(CLK), .Q(g243) ) ;
INV     gate1117  (.A(II11563), .Z(g7305) ) ;
DFF     gate1118  (.D(g7305), .CP(CLK), .Q(g1362) ) ;
INV     gate1119  (.A(II11566), .Z(g7306) ) ;
DFF     gate1120  (.D(g7306), .CP(CLK), .Q(g237) ) ;
INV     gate1121  (.A(II11569), .Z(g7307) ) ;
DFF     gate1122  (.D(g7307), .CP(CLK), .Q(g1365) ) ;
INV     gate1123  (.A(II11605), .Z(g7319) ) ;
DFF     gate1124  (.D(g7319), .CP(CLK), .Q(g231) ) ;
INV     gate1125  (.A(II11572), .Z(g7308) ) ;
DFF     gate1126  (.D(g7308), .CP(CLK), .Q(g1368) ) ;
INV     gate1127  (.A(II11575), .Z(g7309) ) ;
DFF     gate1128  (.D(g7309), .CP(CLK), .Q(g225) ) ;
INV     gate1129  (.A(II11581), .Z(g7311) ) ;
DFF     gate1130  (.D(g7311), .CP(CLK), .Q(g1371) ) ;
INV     gate1131  (.A(II11578), .Z(g7310) ) ;
DFF     gate1132  (.D(g7310), .CP(CLK), .Q(g219) ) ;
INV     gate1133  (.A(II11584), .Z(g7312) ) ;
DFF     gate1134  (.D(g7312), .CP(CLK), .Q(g1377) ) ;
INV     gate1135  (.A(II11587), .Z(g7313) ) ;
DFF     gate1136  (.D(g7313), .CP(CLK), .Q(g213) ) ;
INV     gate1137  (.A(II11590), .Z(g7314) ) ;
DFF     gate1138  (.D(g7314), .CP(CLK), .Q(g1380) ) ;
INV     gate1139  (.A(II11593), .Z(g7315) ) ;
DFF     gate1140  (.D(g7315), .CP(CLK), .Q(g207) ) ;
INV     gate1141  (.A(II11596), .Z(g7316) ) ;
DFF     gate1142  (.D(g7316), .CP(CLK), .Q(g1383) ) ;
INV     gate1143  (.A(II11599), .Z(g7317) ) ;
DFF     gate1144  (.D(g7317), .CP(CLK), .Q(g186) ) ;
INV     gate1145  (.A(II11602), .Z(g7318) ) ;
DFF     gate1146  (.D(g7318), .CP(CLK), .Q(g1386) ) ;
INV     gate1147  (.A(II12939), .Z(g8079) ) ;
DFF     gate1148  (.D(g8079), .CP(CLK), .Q(g4) ) ;
INV     gate1149  (.A(II11659), .Z(g7337) ) ;
DFF     gate1150  (.D(g7337), .CP(CLK), .Q(g12) ) ;
INV     gate1151  (.A(II12936), .Z(g8078) ) ;
DFF     gate1152  (.D(g8078), .CP(CLK), .Q(g1) ) ;
INV     gate1153  (.A(II11656), .Z(g7336) ) ;
DFF     gate1154  (.D(g7336), .CP(CLK), .Q(g9) ) ;
INV     gate1155  (.A(II8262), .Z(g4899) ) ;
DFF     gate1156  (.D(g4899), .CP(CLK), .Q(g1527) ) ;
INV     gate1157  (.A(II11662), .Z(g7338) ) ;
DFF     gate1158  (.D(g7338), .CP(CLK), .Q(g1524) ) ;
INV     gate1159  (.A(II11665), .Z(g7339) ) ;
DFF     gate1160  (.D(g7339), .CP(CLK), .Q(g1528) ) ;
INV     gate1161  (.A(II11668), .Z(g7340) ) ;
DFF     gate1162  (.D(g7340), .CP(CLK), .Q(g1531) ) ;
INV     gate1163  (.A(II11671), .Z(g7341) ) ;
DFF     gate1164  (.D(g7341), .CP(CLK), .Q(g1534) ) ;
INV     gate1165  (.A(II11674), .Z(g7342) ) ;
DFF     gate1166  (.D(g7342), .CP(CLK), .Q(g1537) ) ;
INV     gate1167  (.A(II11677), .Z(g7343) ) ;
DFF     gate1168  (.D(g7343), .CP(CLK), .Q(g1540) ) ;
INV     gate1169  (.A(II11680), .Z(g7344) ) ;
DFF     gate1170  (.D(g7344), .CP(CLK), .Q(g1543) ) ;
INV     gate1171  (.A(II11683), .Z(g7345) ) ;
DFF     gate1172  (.D(g7345), .CP(CLK), .Q(g1546) ) ;
INV     gate1173  (.A(II11686), .Z(g7346) ) ;
DFF     gate1174  (.D(g7346), .CP(CLK), .Q(g1549) ) ;
INV     gate1175  (.A(II11689), .Z(g7347) ) ;
DFF     gate1176  (.D(g7347), .CP(CLK), .Q(g1552) ) ;
INV     gate1177  (.A(II11692), .Z(g7348) ) ;
DFF     gate1178  (.D(g7348), .CP(CLK), .Q(g1555) ) ;
INV     gate1179  (.A(II11695), .Z(g7349) ) ;
DFF     gate1180  (.D(g7349), .CP(CLK), .Q(g1558) ) ;
INV     gate1181  (.A(II11698), .Z(g7350) ) ;
DFF     gate1182  (.D(g7350), .CP(CLK), .Q(g1561) ) ;
INV     gate1183  (.A(II11701), .Z(g7351) ) ;
DFF     gate1184  (.D(g7351), .CP(CLK), .Q(g1564) ) ;
INV     gate1185  (.A(II8265), .Z(g4900) ) ;
DFF     gate1186  (.D(g4900), .CP(CLK), .Q(g1570) ) ;
INV     gate1187  (.A(II11704), .Z(g7352) ) ;
DFF     gate1188  (.D(g7352), .CP(CLK), .Q(g1567) ) ;
INV     gate1189  (.A(II11707), .Z(g7353) ) ;
DFF     gate1190  (.D(g7353), .CP(CLK), .Q(g1571) ) ;
INV     gate1191  (.A(II11710), .Z(g7354) ) ;
DFF     gate1192  (.D(g7354), .CP(CLK), .Q(g1574) ) ;
INV     gate1193  (.A(II11713), .Z(g7355) ) ;
DFF     gate1194  (.D(g7355), .CP(CLK), .Q(g1577) ) ;
INV     gate1195  (.A(II11716), .Z(g7356) ) ;
DFF     gate1196  (.D(g7356), .CP(CLK), .Q(g1580) ) ;
INV     gate1197  (.A(II11719), .Z(g7357) ) ;
DFF     gate1198  (.D(g7357), .CP(CLK), .Q(g1583) ) ;
INV     gate1199  (.A(II11722), .Z(g7358) ) ;
DFF     gate1200  (.D(g7358), .CP(CLK), .Q(g1586) ) ;
INV     gate1201  (.A(II11725), .Z(g7359) ) ;
DFF     gate1202  (.D(g7359), .CP(CLK), .Q(g1589) ) ;
INV     gate1203  (.A(II11728), .Z(g7360) ) ;
DFF     gate1204  (.D(g7360), .CP(CLK), .Q(g1592) ) ;
INV     gate1205  (.A(II11731), .Z(g7361) ) ;
DFF     gate1206  (.D(g7361), .CP(CLK), .Q(g1595) ) ;
INV     gate1207  (.A(II11734), .Z(g7362) ) ;
DFF     gate1208  (.D(g7362), .CP(CLK), .Q(g1598) ) ;
INV     gate1209  (.A(II11737), .Z(g7363) ) ;
DFF     gate1210  (.D(g7363), .CP(CLK), .Q(g1601) ) ;
INV     gate1211  (.A(II11740), .Z(g7364) ) ;
DFF     gate1212  (.D(g7364), .CP(CLK), .Q(g1604) ) ;
INV     gate1213  (.A(II11743), .Z(g7365) ) ;
DFF     gate1214  (.D(g7365), .CP(CLK), .Q(g1607) ) ;
INV     gate1215  (.A(II16592), .Z(g10874) ) ;
DFF     gate1216  (.D(g10874), .CP(CLK), .Q(g1654) ) ;
INV     gate1217  (.A(II16595), .Z(g10875) ) ;
DFF     gate1218  (.D(g10875), .CP(CLK), .Q(g1657) ) ;
INV     gate1219  (.A(II16760), .Z(g11033) ) ;
DFF     gate1220  (.D(g11033), .CP(CLK), .Q(g1660) ) ;
INV     gate1221  (.A(II16763), .Z(g11034) ) ;
DFF     gate1222  (.D(g11034), .CP(CLK), .Q(g1663) ) ;
INV     gate1223  (.A(II16766), .Z(g11035) ) ;
DFF     gate1224  (.D(g11035), .CP(CLK), .Q(g1666) ) ;
INV     gate1225  (.A(II16769), .Z(g11036) ) ;
DFF     gate1226  (.D(g11036), .CP(CLK), .Q(g1669) ) ;
INV     gate1227  (.A(II16772), .Z(g11037) ) ;
DFF     gate1228  (.D(g11037), .CP(CLK), .Q(g1672) ) ;
INV     gate1229  (.A(II16775), .Z(g11038) ) ;
DFF     gate1230  (.D(g11038), .CP(CLK), .Q(g1675) ) ;
INV     gate1231  (.A(II16778), .Z(g11039) ) ;
DFF     gate1232  (.D(g11039), .CP(CLK), .Q(g1678) ) ;
INV     gate1233  (.A(II16781), .Z(g11040) ) ;
DFF     gate1234  (.D(g11040), .CP(CLK), .Q(g1681) ) ;
INV     gate1235  (.A(II16784), .Z(g11041) ) ;
DFF     gate1236  (.D(g11041), .CP(CLK), .Q(g1684) ) ;
INV     gate1237  (.A(II16787), .Z(g11042) ) ;
DFF     gate1238  (.D(g11042), .CP(CLK), .Q(g1687) ) ;
INV     gate1239  (.A(II16790), .Z(g11043) ) ;
DFF     gate1240  (.D(g11043), .CP(CLK), .Q(g546) ) ;
INV     gate1241  (.A(II16802), .Z(g11047) ) ;
DFF     gate1242  (.D(g11047), .CP(CLK), .Q(g554) ) ;
INV     gate1243  (.A(II16805), .Z(g11048) ) ;
DFF     gate1244  (.D(g11048), .CP(CLK), .Q(g557) ) ;
INV     gate1245  (.A(II16808), .Z(g11049) ) ;
DFF     gate1246  (.D(g11049), .CP(CLK), .Q(g560) ) ;
INV     gate1247  (.A(II16811), .Z(g11050) ) ;
DFF     gate1248  (.D(g11050), .CP(CLK), .Q(g563) ) ;
INV     gate1249  (.A(II16814), .Z(g11051) ) ;
DFF     gate1250  (.D(g11051), .CP(CLK), .Q(g566) ) ;
INV     gate1251  (.A(II16598), .Z(g10876) ) ;
DFF     gate1252  (.D(g10876), .CP(CLK), .Q(g569) ) ;
INV     gate1253  (.A(II16601), .Z(g10877) ) ;
DFF     gate1254  (.D(g10877), .CP(CLK), .Q(g572) ) ;
INV     gate1255  (.A(II16817), .Z(g11052) ) ;
DFF     gate1256  (.D(g11052), .CP(CLK), .Q(g575) ) ;
INV     gate1257  (.A(II16793), .Z(g11044) ) ;
DFF     gate1258  (.D(g11044), .CP(CLK), .Q(g549) ) ;
INV     gate1259  (.A(II16796), .Z(g11045) ) ;
DFF     gate1260  (.D(g11045), .CP(CLK), .Q(g552) ) ;
INV     gate1261  (.A(II16799), .Z(g11046) ) ;
DFF     gate1262  (.D(g11046), .CP(CLK), .Q(g553) ) ;
INV     gate1263  (.A(II6498), .Z(g3327) ) ;
DFF     gate1264  (.D(g3327), .CP(CLK), .Q(g23) ) ;
INV     gate1265  (.A(II8228), .Z(g4885) ) ;
DFF     gate1266  (.D(g4885), .CP(CLK), .Q(g26) ) ;
INV     gate1267  (.A(g18), .Z(II4777) ) ;
INV     gate1268  (.A(II4777), .Z(g22) ) ;
INV     gate1269  (.A(g872), .Z(II4780) ) ;
INV     gate1270  (.A(II4780), .Z(g97) ) ;
INV     gate1271  (.A(g873), .Z(II4783) ) ;
INV     gate1272  (.A(II4783), .Z(g98) ) ;
INV     gate1273  (.A(g109), .Z(II4786) ) ;
INV     gate1274  (.A(II4786), .Z(g110) ) ;
INV     gate1275  (.A(g27), .Z(g1962) ) ;
INV     gate1276  (.A(g110), .Z(g1963) ) ;
INV     gate1277  (.A(g114), .Z(g1964) ) ;
INV     gate1278  (.A(g119), .Z(g1965) ) ;
INV     gate1279  (.A(g369), .Z(g1968) ) ;
INV     gate1280  (.A(g456), .Z(g1969) ) ;
INV     gate1281  (.A(g461), .Z(g1972) ) ;
INV     gate1282  (.A(g466), .Z(g1973) ) ;
INV     gate1283  (.A(g627), .Z(g1974) ) ;
INV     gate1284  (.A(g622), .Z(g1975) ) ;
INV     gate1285  (.A(g643), .Z(g1976) ) ;
INV     gate1286  (.A(g646), .Z(g1980) ) ;
INV     gate1287  (.A(g650), .Z(g1981) ) ;
INV     gate1288  (.A(g736), .Z(g1982) ) ;
INV     gate1289  (.A(g750), .Z(g1983) ) ;
INV     gate1290  (.A(g758), .Z(g1984) ) ;
INV     gate1291  (.A(g762), .Z(g1987) ) ;
INV     gate1292  (.A(g766), .Z(g1988) ) ;
INV     gate1293  (.A(g770), .Z(g1989) ) ;
INV     gate1294  (.A(g774), .Z(g1990) ) ;
INV     gate1295  (.A(g778), .Z(g1991) ) ;
INV     gate1296  (.A(g782), .Z(g1992) ) ;
INV     gate1297  (.A(g786), .Z(g1993) ) ;
INV     gate1298  (.A(g794), .Z(g1994) ) ;
INV     gate1299  (.A(g798), .Z(g1997) ) ;
INV     gate1300  (.A(g802), .Z(g1998) ) ;
INV     gate1301  (.A(g806), .Z(g1999) ) ;
INV     gate1302  (.A(g810), .Z(g2000) ) ;
INV     gate1303  (.A(g814), .Z(g2001) ) ;
INV     gate1304  (.A(g818), .Z(g2002) ) ;
INV     gate1305  (.A(g822), .Z(g2003) ) ;
INV     gate1306  (.A(g865), .Z(II4820) ) ;
INV     gate1307  (.A(II4820), .Z(g2004) ) ;
INV     gate1308  (.A(g928), .Z(g2005) ) ;
INV     gate1309  (.A(g932), .Z(g2006) ) ;
INV     gate1310  (.A(g936), .Z(g2007) ) ;
INV     gate1311  (.A(g971), .Z(g2008) ) ;
INV     gate1312  (.A(g976), .Z(g2011) ) ;
INV     gate1313  (.A(g981), .Z(g2012) ) ;
INV     gate1314  (.A(g1101), .Z(g2013) ) ;
INV     gate1315  (.A(g1104), .Z(g2014) ) ;
INV     gate1316  (.A(g1107), .Z(g2015) ) ;
INV     gate1317  (.A(g1361), .Z(g2016) ) ;
INV     gate1318  (.A(g1218), .Z(g2017) ) ;
INV     gate1319  (.A(g1336), .Z(g2018) ) ;
INV     gate1320  (.A(g1341), .Z(g2021) ) ;
INV     gate1321  (.A(g1346), .Z(g2022) ) ;
INV     gate1322  (.A(g1357), .Z(g2023) ) ;
INV     gate1323  (.A(g1718), .Z(g2024) ) ;
INV     gate1324  (.A(g1696), .Z(g2025) ) ;
INV     gate1325  (.A(g1703), .Z(g2028) ) ;
INV     gate1326  (.A(g1690), .Z(g2031) ) ;
INV     gate1327  (.A(g1766), .Z(g2034) ) ;
INV     gate1328  (.A(g1771), .Z(g2037) ) ;
INV     gate1329  (.A(g1776), .Z(g2038) ) ;
INV     gate1330  (.A(g1781), .Z(g2039) ) ;
INV     gate1331  (.A(g1786), .Z(g2040) ) ;
INV     gate1332  (.A(g1791), .Z(g2041) ) ;
INV     gate1333  (.A(g1796), .Z(g2042) ) ;
INV     gate1334  (.A(g1801), .Z(g2043) ) ;
INV     gate1335  (.A(g1958), .Z(II4850) ) ;
INV     gate1336  (.A(g1811), .Z(g2045) ) ;
INV     gate1337  (.A(g1845), .Z(g2046) ) ;
INV     gate1338  (.A(g1857), .Z(g2047) ) ;
INV     gate1339  (.A(g1861), .Z(g2050) ) ;
INV     gate1340  (.A(g1864), .Z(g2054) ) ;
INV     gate1341  (.A(g1950), .Z(g2055) ) ;
INV     gate1342  (.A(g578), .Z(II4859) ) ;
INV     gate1343  (.A(II4859), .Z(g2056) ) ;
INV     gate1344  (.A(g754), .Z(g2057) ) ;
INV     gate1345  (.A(g1380), .Z(g2060) ) ;
INV     gate1346  (.A(g1828), .Z(g2061) ) ;
INV     gate1347  (.A(g108), .Z(g2067) ) ;
INV     gate1348  (.A(g579), .Z(II4866) ) ;
INV     gate1349  (.A(II4866), .Z(g2068) ) ;
INV     gate1350  (.A(g253), .Z(II4869) ) ;
INV     gate1351  (.A(II4869), .Z(g2069) ) ;
INV     gate1352  (.A(g213), .Z(g2070) ) ;
INV     gate1353  (.A(g105), .Z(II4873) ) ;
INV     gate1354  (.A(II4873), .Z(g2071) ) ;
INV     gate1355  (.A(g580), .Z(II4876) ) ;
INV     gate1356  (.A(II4876), .Z(g2072) ) ;
INV     gate1357  (.A(g256), .Z(II4879) ) ;
INV     gate1358  (.A(II4879), .Z(g2073) ) ;
INV     gate1359  (.A(g1377), .Z(g2074) ) ;
INV     gate1360  (.A(g581), .Z(II4883) ) ;
INV     gate1361  (.A(II4883), .Z(g2075) ) ;
INV     gate1362  (.A(g257), .Z(II4886) ) ;
INV     gate1363  (.A(II4886), .Z(g2076) ) ;
INV     gate1364  (.A(g219), .Z(g2077) ) ;
INV     gate1365  (.A(g135), .Z(g2078) ) ;
INV     gate1366  (.A(g582), .Z(II4891) ) ;
INV     gate1367  (.A(II4891), .Z(g2079) ) ;
INV     gate1368  (.A(g258), .Z(II4894) ) ;
INV     gate1369  (.A(II4894), .Z(g2080) ) ;
INV     gate1370  (.A(g1371), .Z(g2082) ) ;
INV     gate1371  (.A(g139), .Z(g2083) ) ;
INV     gate1372  (.A(g583), .Z(II4900) ) ;
INV     gate1373  (.A(II4900), .Z(g2084) ) ;
INV     gate1374  (.A(g259), .Z(II4903) ) ;
INV     gate1375  (.A(II4903), .Z(g2085) ) ;
INV     gate1376  (.A(g119), .Z(II4906) ) ;
INV     gate1377  (.A(II4906), .Z(g2086) ) ;
INV     gate1378  (.A(g225), .Z(g2087) ) ;
INV     gate1379  (.A(g584), .Z(II4917) ) ;
INV     gate1380  (.A(II4917), .Z(g2089) ) ;
INV     gate1381  (.A(g260), .Z(II4920) ) ;
INV     gate1382  (.A(II4920), .Z(g2090) ) ;
INV     gate1383  (.A(g123), .Z(II4924) ) ;
INV     gate1384  (.A(II4924), .Z(g2094) ) ;
INV     gate1385  (.A(g143), .Z(g2095) ) ;
INV     gate1386  (.A(g585), .Z(II4935) ) ;
INV     gate1387  (.A(II4935), .Z(g2097) ) ;
INV     gate1388  (.A(g261), .Z(II4938) ) ;
INV     gate1389  (.A(II4938), .Z(g2098) ) ;
INV     gate1390  (.A(g586), .Z(II4948) ) ;
INV     gate1391  (.A(II4948), .Z(g2100) ) ;
INV     gate1392  (.A(g262), .Z(II4951) ) ;
INV     gate1393  (.A(II4951), .Z(g2101) ) ;
INV     gate1394  (.A(g254), .Z(II4961) ) ;
INV     gate1395  (.A(II4961), .Z(g2103) ) ;
INV     gate1396  (.A(g1170), .Z(II4992) ) ;
INV     gate1397  (.A(II4992), .Z(g2108) ) ;
INV     gate1398  (.A(g1173), .Z(II5002) ) ;
INV     gate1399  (.A(II5002), .Z(g2110) ) ;
INV     gate1400  (.A(g639), .Z(g2112) ) ;
INV     gate1401  (.A(g1176), .Z(II5020) ) ;
INV     gate1402  (.A(II5020), .Z(g2116) ) ;
INV     gate1403  (.A(g1854), .Z(g2118) ) ;
INV     gate1404  (.A(g928), .Z(II5031) ) ;
INV     gate1405  (.A(II5031), .Z(g2119) ) ;
INV     gate1406  (.A(g1179), .Z(II5041) ) ;
INV     gate1407  (.A(II5041), .Z(g2121) ) ;
INV     gate1408  (.A(g1182), .Z(II5044) ) ;
INV     gate1409  (.A(II5044), .Z(g2122) ) ;
INV     gate1410  (.A(g1185), .Z(II5047) ) ;
INV     gate1411  (.A(II5047), .Z(g2123) ) ;
INV     gate1412  (.A(g1216), .Z(II5050) ) ;
INV     gate1413  (.A(II5050), .Z(g2124) ) ;
INV     gate1414  (.A(g1188), .Z(II5053) ) ;
INV     gate1415  (.A(II5053), .Z(g2125) ) ;
INV     gate1416  (.A(g12), .Z(g2126) ) ;
INV     gate1417  (.A(g1961), .Z(II5057) ) ;
INV     gate1418  (.A(II5057), .Z(g2130) ) ;
INV     gate1419  (.A(g1191), .Z(II5060) ) ;
INV     gate1420  (.A(II5060), .Z(g2131) ) ;
INV     gate1421  (.A(g1690), .Z(II5064) ) ;
INV     gate1422  (.A(II5064), .Z(g2135) ) ;
INV     gate1423  (.A(g33), .Z(II5067) ) ;
INV     gate1424  (.A(II5067), .Z(g2154) ) ;
INV     gate1425  (.A(g1194), .Z(II5070) ) ;
INV     gate1426  (.A(II5070), .Z(g2155) ) ;
INV     gate1427  (.A(g34), .Z(II5073) ) ;
INV     gate1428  (.A(II5073), .Z(g2156) ) ;
INV     gate1429  (.A(g1703), .Z(g2157) ) ;
INV     gate1430  (.A(g35), .Z(II5077) ) ;
INV     gate1431  (.A(II5077), .Z(g2158) ) ;
INV     gate1432  (.A(g36), .Z(II5080) ) ;
INV     gate1433  (.A(II5080), .Z(g2159) ) ;
INV     gate1434  (.A(g1854), .Z(II5089) ) ;
INV     gate1435  (.A(II5089), .Z(g2162) ) ;
INV     gate1436  (.A(g32), .Z(II5092) ) ;
INV     gate1437  (.A(II5092), .Z(g2163) ) ;
INV     gate1438  (.A(g37), .Z(II5095) ) ;
INV     gate1439  (.A(II5095), .Z(g2164) ) ;
INV     gate1440  (.A(g38), .Z(II5098) ) ;
INV     gate1441  (.A(II5098), .Z(g2165) ) ;
INV     gate1442  (.A(g1960), .Z(II5101) ) ;
INV     gate1443  (.A(II5101), .Z(g2166) ) ;
INV     gate1444  (.A(g39), .Z(II5111) ) ;
INV     gate1445  (.A(II5111), .Z(g2168) ) ;
INV     gate1446  (.A(g42), .Z(g2169) ) ;
INV     gate1447  (.A(g30), .Z(g2170) ) ;
INV     gate1448  (.A(g40), .Z(II5116) ) ;
INV     gate1449  (.A(II5116), .Z(g2171) ) ;
INV     gate1450  (.A(g43), .Z(g2172) ) ;
INV     gate1451  (.A(g622), .Z(II5120) ) ;
INV     gate1452  (.A(II5120), .Z(g2173) ) ;
INV     gate1453  (.A(g31), .Z(g2174) ) ;
INV     gate1454  (.A(g44), .Z(g2175) ) ;
INV     gate1455  (.A(g82), .Z(g2176) ) ;
INV     gate1456  (.A(g45), .Z(g2178) ) ;
INV     gate1457  (.A(g89), .Z(g2179) ) ;
INV     gate1458  (.A(g639), .Z(II5142) ) ;
INV     gate1459  (.A(II5142), .Z(g2181) ) ;
INV     gate1460  (.A(g1806), .Z(g2184) ) ;
INV     gate1461  (.A(g46), .Z(g2185) ) ;
INV     gate1462  (.A(g90), .Z(g2186) ) ;
INV     gate1463  (.A(g746), .Z(g2187) ) ;
INV     gate1464  (.A(g1453), .Z(II5149) ) ;
INV     gate1465  (.A(II5149), .Z(g2190) ) ;
INV     gate1466  (.A(g1696), .Z(g2191) ) ;
INV     gate1467  (.A(g47), .Z(g2194) ) ;
INV     gate1468  (.A(g83), .Z(g2195) ) ;
INV     gate1469  (.A(g91), .Z(g2196) ) ;
INV     gate1470  (.A(g101), .Z(g2197) ) ;
INV     gate1471  (.A(g668), .Z(g2198) ) ;
INV     gate1472  (.A(g48), .Z(g2199) ) ;
INV     gate1473  (.A(g92), .Z(g2200) ) ;
INV     gate1474  (.A(g102), .Z(g2201) ) ;
INV     gate1475  (.A(g148), .Z(g2202) ) ;
INV     gate1476  (.A(g677), .Z(g2203) ) ;
INV     gate1477  (.A(g1419), .Z(II5171) ) ;
INV     gate1478  (.A(II5171), .Z(g2206) ) ;
INV     gate1479  (.A(g52), .Z(II5174) ) ;
INV     gate1480  (.A(II5174), .Z(g2207) ) ;
INV     gate1481  (.A(g84), .Z(g2208) ) ;
INV     gate1482  (.A(g93), .Z(g2209) ) ;
INV     gate1483  (.A(g103), .Z(g2210) ) ;
INV     gate1484  (.A(g153), .Z(g2211) ) ;
INV     gate1485  (.A(g686), .Z(g2212) ) ;
INV     gate1486  (.A(g1110), .Z(g2213) ) ;
INV     gate1487  (.A(g115), .Z(g2214) ) ;
INV     gate1488  (.A(g41), .Z(g2216) ) ;
INV     gate1489  (.A(g55), .Z(II5192) ) ;
INV     gate1490  (.A(II5192), .Z(g2217) ) ;
INV     gate1491  (.A(g85), .Z(g2218) ) ;
INV     gate1492  (.A(g94), .Z(g2219) ) ;
INV     gate1493  (.A(g104), .Z(g2220) ) ;
INV     gate1494  (.A(g143), .Z(II5198) ) ;
INV     gate1495  (.A(II5198), .Z(g2221) ) ;
INV     gate1496  (.A(g158), .Z(g2222) ) ;
INV     gate1497  (.A(g695), .Z(g2224) ) ;
INV     gate1498  (.A(g58), .Z(II5210) ) ;
INV     gate1499  (.A(II5210), .Z(g2225) ) ;
INV     gate1500  (.A(g86), .Z(g2226) ) ;
INV     gate1501  (.A(g95), .Z(g2227) ) ;
INV     gate1502  (.A(g28), .Z(g2228) ) ;
INV     gate1503  (.A(g162), .Z(g2229) ) ;
INV     gate1504  (.A(g704), .Z(g2230) ) ;
INV     gate1505  (.A(g1104), .Z(II5218) ) ;
INV     gate1506  (.A(II5218), .Z(g2231) ) ;
INV     gate1507  (.A(g1407), .Z(II5221) ) ;
INV     gate1508  (.A(II5221), .Z(g2232) ) ;
INV     gate1509  (.A(g61), .Z(II5224) ) ;
INV     gate1510  (.A(II5224), .Z(g2233) ) ;
INV     gate1511  (.A(g87), .Z(g2234) ) ;
INV     gate1512  (.A(g96), .Z(g2235) ) ;
INV     gate1513  (.A(g713), .Z(g2237) ) ;
INV     gate1514  (.A(g1107), .Z(II5237) ) ;
INV     gate1515  (.A(II5237), .Z(g2238) ) ;
INV     gate1516  (.A(g64), .Z(II5240) ) ;
INV     gate1517  (.A(II5240), .Z(g2239) ) ;
INV     gate1518  (.A(g88), .Z(g2240) ) ;
INV     gate1519  (.A(g722), .Z(g2241) ) ;
INV     gate1520  (.A(g925), .Z(II5245) ) ;
INV     gate1521  (.A(II5245), .Z(g2242) ) ;
INV     gate1522  (.A(g1110), .Z(II5248) ) ;
INV     gate1523  (.A(II5248), .Z(g2243) ) ;
INV     gate1524  (.A(g1424), .Z(II5251) ) ;
INV     gate1525  (.A(II5251), .Z(g2244) ) ;
INV     gate1526  (.A(g1700), .Z(II5254) ) ;
INV     gate1527  (.A(II5254), .Z(g2245) ) ;
INV     gate1528  (.A(g1810), .Z(g2246) ) ;
INV     gate1529  (.A(g67), .Z(II5258) ) ;
INV     gate1530  (.A(II5258), .Z(g2247) ) ;
INV     gate1531  (.A(g99), .Z(g2248) ) ;
INV     gate1532  (.A(g127), .Z(g2249) ) ;
INV     gate1533  (.A(g731), .Z(g2251) ) ;
INV     gate1534  (.A(g70), .Z(II5271) ) ;
INV     gate1535  (.A(II5271), .Z(g2252) ) ;
INV     gate1536  (.A(g100), .Z(g2253) ) ;
INV     gate1537  (.A(g131), .Z(g2254) ) ;
INV     gate1538  (.A(g1411), .Z(II5276) ) ;
INV     gate1539  (.A(II5276), .Z(g2255) ) ;
INV     gate1540  (.A(g73), .Z(II5279) ) ;
INV     gate1541  (.A(II5279), .Z(g2256) ) ;
INV     gate1542  (.A(g49), .Z(II5289) ) ;
INV     gate1543  (.A(II5289), .Z(g2258) ) ;
INV     gate1544  (.A(g76), .Z(II5292) ) ;
INV     gate1545  (.A(II5292), .Z(g2259) ) ;
INV     gate1546  (.A(g1713), .Z(g2261) ) ;
INV     gate1547  (.A(g79), .Z(II5304) ) ;
INV     gate1548  (.A(II5304), .Z(g2267) ) ;
INV     gate1549  (.A(g654), .Z(g2268) ) ;
INV     gate1550  (.A(g97), .Z(II5308) ) ;
INV     gate1551  (.A(II5308), .Z(g2269) ) ;
INV     gate1552  (.A(g98), .Z(II5311) ) ;
INV     gate1553  (.A(II5311), .Z(g2270) ) ;
INV     gate1554  (.A(g877), .Z(g2271) ) ;
INV     gate1555  (.A(g881), .Z(g2273) ) ;
INV     gate1556  (.A(g757), .Z(g2275) ) ;
INV     gate1557  (.A(g756), .Z(II5332) ) ;
INV     gate1558  (.A(II5332), .Z(g2296) ) ;
INV     gate1559  (.A(g865), .Z(g2297) ) ;
INV     gate1560  (.A(g1700), .Z(II5336) ) ;
INV     gate1561  (.A(II5336), .Z(g2298) ) ;
INV     gate1562  (.A(g1707), .Z(g2299) ) ;
INV     gate1563  (.A(g29), .Z(g2302) ) ;
INV     gate1564  (.A(g746), .Z(II5348) ) ;
INV     gate1565  (.A(II5348), .Z(g2304) ) ;
INV     gate1566  (.A(g622), .Z(g2317) ) ;
INV     gate1567  (.A(g18), .Z(g2320) ) ;
INV     gate1568  (.A(g1857), .Z(II5378) ) ;
INV     gate1569  (.A(II5378), .Z(g2322) ) ;
INV     gate1570  (.A(g1882), .Z(g2328) ) ;
INV     gate1571  (.A(g886), .Z(II5383) ) ;
INV     gate1572  (.A(II5383), .Z(g2329) ) ;
INV     gate1573  (.A(g1891), .Z(g2330) ) ;
INV     gate1574  (.A(g658), .Z(g2331) ) ;
INV     gate1575  (.A(g889), .Z(II5388) ) ;
INV     gate1576  (.A(II5388), .Z(g2334) ) ;
INV     gate1577  (.A(g1101), .Z(II5391) ) ;
INV     gate1578  (.A(II5391), .Z(g2335) ) ;
INV     gate1579  (.A(g1900), .Z(g2336) ) ;
INV     gate1580  (.A(g892), .Z(II5395) ) ;
INV     gate1581  (.A(II5395), .Z(g2337) ) ;
INV     gate1582  (.A(g1909), .Z(g2338) ) ;
INV     gate1583  (.A(g895), .Z(II5399) ) ;
INV     gate1584  (.A(II5399), .Z(g2339) ) ;
INV     gate1585  (.A(g1918), .Z(g2340) ) ;
INV     gate1586  (.A(g636), .Z(II5403) ) ;
INV     gate1587  (.A(II5403), .Z(g2341) ) ;
INV     gate1588  (.A(g898), .Z(II5406) ) ;
INV     gate1589  (.A(II5406), .Z(g2342) ) ;
INV     gate1590  (.A(g1927), .Z(g2343) ) ;
INV     gate1591  (.A(g901), .Z(II5410) ) ;
INV     gate1592  (.A(II5410), .Z(g2344) ) ;
INV     gate1593  (.A(g1936), .Z(g2345) ) ;
INV     gate1594  (.A(g904), .Z(II5414) ) ;
INV     gate1595  (.A(II5414), .Z(g2346) ) ;
INV     gate1596  (.A(g1945), .Z(g2347) ) ;
INV     gate1597  (.A(g907), .Z(II5418) ) ;
INV     gate1598  (.A(II5418), .Z(g2348) ) ;
INV     gate1599  (.A(g549), .Z(II5421) ) ;
INV     gate1600  (.A(II5421), .Z(g2349) ) ;
INV     gate1601  (.A(g910), .Z(II5424) ) ;
INV     gate1602  (.A(II5424), .Z(g2350) ) ;
INV     gate1603  (.A(g913), .Z(II5427) ) ;
INV     gate1604  (.A(II5427), .Z(g2351) ) ;
INV     gate1605  (.A(g916), .Z(II5430) ) ;
INV     gate1606  (.A(II5430), .Z(g2352) ) ;
INV     gate1607  (.A(g18), .Z(II5435) ) ;
INV     gate1608  (.A(g18), .Z(II5438) ) ;
INV     gate1609  (.A(II5438), .Z(g2356) ) ;
INV     gate1610  (.A(g919), .Z(II5441) ) ;
INV     gate1611  (.A(II5441), .Z(g2363) ) ;
INV     gate1612  (.A(g611), .Z(g2364) ) ;
INV     gate1613  (.A(g922), .Z(II5445) ) ;
INV     gate1614  (.A(II5445), .Z(g2368) ) ;
INV     gate1615  (.A(g617), .Z(g2369) ) ;
INV     gate1616  (.A(g471), .Z(g2373) ) ;
INV     gate1617  (.A(g591), .Z(g2374) ) ;
INV     gate1618  (.A(g1368), .Z(g2381) ) ;
INV     gate1619  (.A(g599), .Z(g2382) ) ;
INV     gate1620  (.A(g1289), .Z(II5475) ) ;
INV     gate1621  (.A(II5475), .Z(g2390) ) ;
INV     gate1622  (.A(g1212), .Z(II5478) ) ;
INV     gate1623  (.A(II5478), .Z(g2391) ) ;
INV     gate1624  (.A(g231), .Z(g2395) ) ;
INV     gate1625  (.A(g1389), .Z(g2396) ) ;
INV     gate1626  (.A(g605), .Z(g2399) ) ;
INV     gate1627  (.A(g1365), .Z(g2406) ) ;
INV     gate1628  (.A(g197), .Z(g2407) ) ;
INV     gate1629  (.A(g1453), .Z(g2410) ) ;
INV     gate1630  (.A(g1690), .Z(II5494) ) ;
INV     gate1631  (.A(II5494), .Z(g2411) ) ;
INV     gate1632  (.A(g587), .Z(II5497) ) ;
INV     gate1633  (.A(II5497), .Z(g2418) ) ;
INV     gate1634  (.A(g237), .Z(g2420) ) ;
INV     gate1635  (.A(g1374), .Z(g2421) ) ;
INV     gate1636  (.A(g1690), .Z(g2424) ) ;
INV     gate1637  (.A(g588), .Z(II5510) ) ;
INV     gate1638  (.A(II5510), .Z(g2431) ) ;
INV     gate1639  (.A(g255), .Z(II5513) ) ;
INV     gate1640  (.A(II5513), .Z(g2432) ) ;
INV     gate1641  (.A(g1362), .Z(g2434) ) ;
INV     gate1642  (.A(g201), .Z(g2435) ) ;
INV     gate1643  (.A(g589), .Z(II5525) ) ;
INV     gate1644  (.A(II5525), .Z(g2436) ) ;
INV     gate1645  (.A(g243), .Z(g2438) ) ;
INV     gate1646  (.A(g876), .Z(g2444) ) ;
INV     gate1647  (.A(g1400), .Z(g2446) ) ;
INV     gate1648  (.A(g790), .Z(g2449) ) ;
INV     gate1649  (.A(g1351), .Z(g2450) ) ;
INV     gate1650  (.A(g248), .Z(g2451) ) ;
INV     gate1651  (.A(g868), .Z(II5549) ) ;
INV     gate1652  (.A(II5549), .Z(g2454) ) ;
INV     gate1653  (.A(g826), .Z(g2455) ) ;
INV     gate1654  (.A(g1397), .Z(g2456) ) ;
INV     gate1655  (.A(g110), .Z(II5555) ) ;
INV     gate1656  (.A(II5555), .Z(g2462) ) ;
INV     gate1657  (.A(g192), .Z(g2475) ) ;
INV     gate1658  (.A(g26), .Z(g2479) ) ;
INV     gate1659  (.A(g869), .Z(II5561) ) ;
INV     gate1660  (.A(II5561), .Z(g2480) ) ;
INV     gate1661  (.A(g882), .Z(g2481) ) ;
INV     gate1662  (.A(g1713), .Z(II5565) ) ;
INV     gate1663  (.A(II5565), .Z(g2482) ) ;
INV     gate1664  (.A(g1197), .Z(II5579) ) ;
INV     gate1665  (.A(II5579), .Z(g2502) ) ;
INV     gate1666  (.A(g1872), .Z(g2503) ) ;
INV     gate1667  (.A(g636), .Z(g2506) ) ;
INV     gate1668  (.A(g1200), .Z(II5584) ) ;
INV     gate1669  (.A(II5584), .Z(g2507) ) ;
INV     gate1670  (.A(g940), .Z(g2508) ) ;
INV     gate1671  (.A(g1203), .Z(II5588) ) ;
INV     gate1672  (.A(II5588), .Z(g2509) ) ;
INV     gate1673  (.A(g590), .Z(g2518) ) ;
INV     gate1674  (.A(g932), .Z(II5632) ) ;
INV     gate1675  (.A(II5632), .Z(g2523) ) ;
INV     gate1676  (.A(g986), .Z(g2524) ) ;
INV     gate1677  (.A(g936), .Z(II5638) ) ;
INV     gate1678  (.A(II5638), .Z(g2529) ) ;
INV     gate1679  (.A(g546), .Z(II5641) ) ;
INV     gate1680  (.A(II5641), .Z(g2530) ) ;
INV     gate1681  (.A(g940), .Z(II5646) ) ;
INV     gate1682  (.A(II5646), .Z(g2537) ) ;
INV     gate1683  (.A(g554), .Z(II5652) ) ;
INV     gate1684  (.A(II5652), .Z(g2539) ) ;
INV     gate1685  (.A(g557), .Z(II5655) ) ;
INV     gate1686  (.A(II5655), .Z(g2540) ) ;
INV     gate1687  (.A(g560), .Z(II5658) ) ;
INV     gate1688  (.A(II5658), .Z(g2541) ) ;
INV     gate1689  (.A(g1868), .Z(g2542) ) ;
INV     gate1690  (.A(g563), .Z(II5662) ) ;
INV     gate1691  (.A(II5662), .Z(g2543) ) ;
INV     gate1692  (.A(g23), .Z(g2547) ) ;
INV     gate1693  (.A(g566), .Z(II5667) ) ;
INV     gate1694  (.A(II5667), .Z(g2548) ) ;
INV     gate1695  (.A(g1386), .Z(g2549) ) ;
INV     gate1696  (.A(g1834), .Z(g2550) ) ;
INV     gate1697  (.A(g569), .Z(II5672) ) ;
INV     gate1698  (.A(II5672), .Z(g2554) ) ;
INV     gate1699  (.A(g186), .Z(g2556) ) ;
INV     gate1700  (.A(g1840), .Z(g2557) ) ;
INV     gate1701  (.A(g572), .Z(II5684) ) ;
INV     gate1702  (.A(II5684), .Z(g2560) ) ;
INV     gate1703  (.A(g1383), .Z(g2562) ) ;
INV     gate1704  (.A(g1814), .Z(g2564) ) ;
INV     gate1705  (.A(g575), .Z(II5695) ) ;
INV     gate1706  (.A(II5695), .Z(g2569) ) ;
INV     gate1707  (.A(g207), .Z(g2570) ) ;
INV     gate1708  (.A(g1822), .Z(g2571) ) ;
INV     gate1709  (.A(g1962), .Z(g2578) ) ;
INV     gate1710  (.A(g1969), .Z(g2579) ) ;
INV     gate1711  (.A(g1972), .Z(g2586) ) ;
INV     gate1712  (.A(g1973), .Z(g2593) ) ;
INV     gate1713  (.A(g2056), .Z(II5704) ) ;
INV     gate1714  (.A(g2418), .Z(II5707) ) ;
INV     gate1715  (.A(g2431), .Z(II5710) ) ;
INV     gate1716  (.A(g2436), .Z(II5713) ) ;
INV     gate1717  (.A(g2068), .Z(II5716) ) ;
INV     gate1718  (.A(g2072), .Z(II5719) ) ;
INV     gate1719  (.A(g2075), .Z(II5722) ) ;
INV     gate1720  (.A(g2079), .Z(II5725) ) ;
INV     gate1721  (.A(g2084), .Z(II5728) ) ;
INV     gate1722  (.A(g2089), .Z(II5731) ) ;
INV     gate1723  (.A(g2097), .Z(II5734) ) ;
INV     gate1724  (.A(g2100), .Z(II5737) ) ;
INV     gate1725  (.A(g2341), .Z(II5740) ) ;
INV     gate1726  (.A(g1994), .Z(g2614) ) ;
INV     gate1727  (.A(g1997), .Z(g2617) ) ;
INV     gate1728  (.A(g1998), .Z(g2620) ) ;
INV     gate1729  (.A(g1999), .Z(g2623) ) ;
INV     gate1730  (.A(g2000), .Z(g2626) ) ;
INV     gate1731  (.A(g2001), .Z(g2629) ) ;
INV     gate1732  (.A(g2002), .Z(g2632) ) ;
INV     gate1733  (.A(g2003), .Z(g2635) ) ;
INV     gate1734  (.A(g2296), .Z(II5751) ) ;
INV     gate1735  (.A(g2304), .Z(II5754) ) ;
INV     gate1736  (.A(g1984), .Z(g2640) ) ;
INV     gate1737  (.A(g1987), .Z(g2641) ) ;
INV     gate1738  (.A(g1988), .Z(g2642) ) ;
INV     gate1739  (.A(g1989), .Z(g2643) ) ;
INV     gate1740  (.A(g1990), .Z(g2644) ) ;
INV     gate1741  (.A(g1991), .Z(g2645) ) ;
INV     gate1742  (.A(g1992), .Z(g2646) ) ;
INV     gate1743  (.A(g1993), .Z(g2647) ) ;
INV     gate1744  (.A(g2004), .Z(II5765) ) ;
INV     gate1745  (.A(g2005), .Z(g2649) ) ;
INV     gate1746  (.A(g2006), .Z(g2650) ) ;
INV     gate1747  (.A(g2007), .Z(g2651) ) ;
INV     gate1748  (.A(g2008), .Z(g2652) ) ;
INV     gate1749  (.A(g2011), .Z(g2653) ) ;
INV     gate1750  (.A(g2012), .Z(g2654) ) ;
INV     gate1751  (.A(g2013), .Z(g2655) ) ;
INV     gate1752  (.A(g2014), .Z(g2662) ) ;
INV     gate1753  (.A(g2015), .Z(g2669) ) ;
INV     gate1754  (.A(g2034), .Z(g2677) ) ;
INV     gate1755  (.A(g2037), .Z(g2683) ) ;
INV     gate1756  (.A(g2038), .Z(g2689) ) ;
INV     gate1757  (.A(g2039), .Z(g2695) ) ;
INV     gate1758  (.A(g2040), .Z(g2701) ) ;
INV     gate1759  (.A(g2041), .Z(g2707) ) ;
INV     gate1760  (.A(g2042), .Z(g2713) ) ;
INV     gate1761  (.A(g2043), .Z(g2719) ) ;
INV     gate1762  (.A(g2018), .Z(g2725) ) ;
INV     gate1763  (.A(g2021), .Z(g2726) ) ;
INV     gate1764  (.A(g2022), .Z(g2727) ) ;
INV     gate1765  (.A(g2025), .Z(g2728) ) ;
INV     gate1766  (.A(g2162), .Z(II5789) ) ;
INV     gate1767  (.A(g2080), .Z(II5792) ) ;
INV     gate1768  (.A(II5792), .Z(g2732) ) ;
INV     gate1769  (.A(g2462), .Z(II5795) ) ;
INV     gate1770  (.A(II5795), .Z(g2733) ) ;
INV     gate1771  (.A(g2085), .Z(II5798) ) ;
INV     gate1772  (.A(II5798), .Z(g2742) ) ;
INV     gate1773  (.A(g1984), .Z(II5801) ) ;
INV     gate1774  (.A(II5801), .Z(g2743) ) ;
INV     gate1775  (.A(g2356), .Z(II5809) ) ;
INV     gate1776  (.A(II5809), .Z(g2745) ) ;
INV     gate1777  (.A(g2090), .Z(II5812) ) ;
INV     gate1778  (.A(II5812), .Z(g2748) ) ;
INV     gate1779  (.A(g1994), .Z(II5815) ) ;
INV     gate1780  (.A(II5815), .Z(g2749) ) ;
INV     gate1781  (.A(g2098), .Z(II5818) ) ;
INV     gate1782  (.A(II5818), .Z(g2750) ) ;
INV     gate1783  (.A(g2101), .Z(II5821) ) ;
INV     gate1784  (.A(II5821), .Z(g2751) ) ;
INV     gate1785  (.A(g2502), .Z(II5824) ) ;
INV     gate1786  (.A(II5824), .Z(g2752) ) ;
INV     gate1787  (.A(g2271), .Z(II5827) ) ;
INV     gate1788  (.A(II5827), .Z(g2753) ) ;
INV     gate1789  (.A(g2067), .Z(II5830) ) ;
INV     gate1790  (.A(II5830), .Z(g2754) ) ;
INV     gate1791  (.A(g2103), .Z(II5833) ) ;
INV     gate1792  (.A(II5833), .Z(g2755) ) ;
INV     gate1793  (.A(g2507), .Z(II5837) ) ;
INV     gate1794  (.A(II5837), .Z(g2757) ) ;
INV     gate1795  (.A(g2432), .Z(II5840) ) ;
INV     gate1796  (.A(II5840), .Z(g2758) ) ;
INV     gate1797  (.A(g2509), .Z(II5843) ) ;
INV     gate1798  (.A(II5843), .Z(g2759) ) ;
INV     gate1799  (.A(g2275), .Z(II5847) ) ;
INV     gate1800  (.A(II5847), .Z(g2763) ) ;
INV     gate1801  (.A(g2273), .Z(II5850) ) ;
INV     gate1802  (.A(II5850), .Z(g2764) ) ;
INV     gate1803  (.A(g2184), .Z(g2765) ) ;
INV     gate1804  (.A(g2523), .Z(II5854) ) ;
INV     gate1805  (.A(II5854), .Z(g2771) ) ;
INV     gate1806  (.A(g2508), .Z(g2772) ) ;
INV     gate1807  (.A(g2529), .Z(II5858) ) ;
INV     gate1808  (.A(II5858), .Z(g2773) ) ;
AND2    gate1809  (.A(g1765), .B(g1610), .Z(g2276) ) ;
INV     gate1810  (.A(g2276), .Z(g2774) ) ;
INV     gate1811  (.A(g2537), .Z(II5862) ) ;
INV     gate1812  (.A(II5862), .Z(g2775) ) ;
INV     gate1813  (.A(g2276), .Z(g2777) ) ;
INV     gate1814  (.A(g2276), .Z(g2778) ) ;
INV     gate1815  (.A(g1974), .Z(g2779) ) ;
INV     gate1816  (.A(g2276), .Z(g2789) ) ;
INV     gate1817  (.A(g2276), .Z(g2790) ) ;
INV     gate1818  (.A(g2276), .Z(g2793) ) ;
INV     gate1819  (.A(g2276), .Z(g2796) ) ;
INV     gate1820  (.A(g2524), .Z(g2797) ) ;
INV     gate1821  (.A(g2449), .Z(g2798) ) ;
INV     gate1822  (.A(g2276), .Z(g2799) ) ;
NAND2   gate1823  (.A(II5024), .B(II5025), .Z(g2117) ) ;
INV     gate1824  (.A(g2117), .Z(g2801) ) ;
INV     gate1825  (.A(g2276), .Z(g2802) ) ;
INV     gate1826  (.A(g2154), .Z(g2803) ) ;
INV     gate1827  (.A(g2156), .Z(g2808) ) ;
INV     gate1828  (.A(g2207), .Z(II5909) ) ;
INV     gate1829  (.A(II5909), .Z(g2809) ) ;
INV     gate1830  (.A(g2158), .Z(g2812) ) ;
INV     gate1831  (.A(g2169), .Z(II5913) ) ;
INV     gate1832  (.A(II5913), .Z(g2813) ) ;
INV     gate1833  (.A(g2217), .Z(II5916) ) ;
INV     gate1834  (.A(II5916), .Z(g2814) ) ;
INV     gate1835  (.A(g2530), .Z(II5919) ) ;
INV     gate1836  (.A(II5919), .Z(g2817) ) ;
INV     gate1837  (.A(g2170), .Z(II5922) ) ;
INV     gate1838  (.A(II5922), .Z(g2818) ) ;
INV     gate1839  (.A(g2159), .Z(g2819) ) ;
INV     gate1840  (.A(g2172), .Z(II5926) ) ;
INV     gate1841  (.A(II5926), .Z(g2820) ) ;
INV     gate1842  (.A(g2225), .Z(II5929) ) ;
INV     gate1843  (.A(II5929), .Z(g2821) ) ;
INV     gate1844  (.A(g2539), .Z(II5932) ) ;
INV     gate1845  (.A(II5932), .Z(g2824) ) ;
INV     gate1846  (.A(g2174), .Z(II5935) ) ;
INV     gate1847  (.A(II5935), .Z(g2825) ) ;
INV     gate1848  (.A(g2163), .Z(g2826) ) ;
INV     gate1849  (.A(g2164), .Z(g2827) ) ;
INV     gate1850  (.A(g2175), .Z(II5940) ) ;
INV     gate1851  (.A(II5940), .Z(g2828) ) ;
INV     gate1852  (.A(g2233), .Z(II5943) ) ;
INV     gate1853  (.A(II5943), .Z(g2829) ) ;
INV     gate1854  (.A(g2176), .Z(II5946) ) ;
INV     gate1855  (.A(II5946), .Z(g2832) ) ;
INV     gate1856  (.A(g2540), .Z(II5949) ) ;
INV     gate1857  (.A(II5949), .Z(g2833) ) ;
INV     gate1858  (.A(g2506), .Z(II5952) ) ;
INV     gate1859  (.A(II5952), .Z(g2834) ) ;
INV     gate1860  (.A(g2130), .Z(g2837) ) ;
INV     gate1861  (.A(g2165), .Z(g2838) ) ;
INV     gate1862  (.A(g2178), .Z(II5957) ) ;
INV     gate1863  (.A(II5957), .Z(g2839) ) ;
INV     gate1864  (.A(g2239), .Z(II5960) ) ;
INV     gate1865  (.A(II5960), .Z(g2840) ) ;
INV     gate1866  (.A(g2179), .Z(II5963) ) ;
INV     gate1867  (.A(II5963), .Z(g2843) ) ;
INV     gate1868  (.A(g2541), .Z(II5966) ) ;
INV     gate1869  (.A(II5966), .Z(g2844) ) ;
INV     gate1870  (.A(g2168), .Z(g2845) ) ;
INV     gate1871  (.A(g2185), .Z(II5970) ) ;
INV     gate1872  (.A(II5970), .Z(g2846) ) ;
INV     gate1873  (.A(g2247), .Z(II5973) ) ;
INV     gate1874  (.A(II5973), .Z(g2847) ) ;
INV     gate1875  (.A(g2186), .Z(II5976) ) ;
INV     gate1876  (.A(II5976), .Z(g2850) ) ;
INV     gate1877  (.A(g2543), .Z(II5979) ) ;
INV     gate1878  (.A(II5979), .Z(g2851) ) ;
NAND2   gate1879  (.A(II5592), .B(II5593), .Z(g2510) ) ;
INV     gate1880  (.A(g2510), .Z(II5982) ) ;
INV     gate1881  (.A(II5982), .Z(g2852) ) ;
INV     gate1882  (.A(g2171), .Z(g2853) ) ;
INV     gate1883  (.A(g2194), .Z(II5986) ) ;
INV     gate1884  (.A(II5986), .Z(g2854) ) ;
INV     gate1885  (.A(g2252), .Z(II5989) ) ;
INV     gate1886  (.A(II5989), .Z(g2855) ) ;
INV     gate1887  (.A(g2195), .Z(II5992) ) ;
INV     gate1888  (.A(II5992), .Z(g2858) ) ;
INV     gate1889  (.A(g2196), .Z(II5995) ) ;
INV     gate1890  (.A(II5995), .Z(g2859) ) ;
INV     gate1891  (.A(g2197), .Z(II5998) ) ;
INV     gate1892  (.A(II5998), .Z(g2860) ) ;
INV     gate1893  (.A(g2548), .Z(II6001) ) ;
INV     gate1894  (.A(II6001), .Z(g2861) ) ;
INV     gate1895  (.A(g2298), .Z(g2864) ) ;
INV     gate1896  (.A(g2199), .Z(II6007) ) ;
INV     gate1897  (.A(II6007), .Z(g2867) ) ;
INV     gate1898  (.A(g2256), .Z(II6010) ) ;
INV     gate1899  (.A(II6010), .Z(g2868) ) ;
INV     gate1900  (.A(g2200), .Z(II6013) ) ;
INV     gate1901  (.A(II6013), .Z(g2871) ) ;
INV     gate1902  (.A(g2201), .Z(II6016) ) ;
INV     gate1903  (.A(II6016), .Z(g2872) ) ;
INV     gate1904  (.A(g2554), .Z(II6019) ) ;
INV     gate1905  (.A(II6019), .Z(g2873) ) ;
INV     gate1906  (.A(g2258), .Z(II6022) ) ;
INV     gate1907  (.A(II6022), .Z(g2874) ) ;
INV     gate1908  (.A(g2259), .Z(II6025) ) ;
INV     gate1909  (.A(II6025), .Z(g2877) ) ;
INV     gate1910  (.A(g2208), .Z(II6028) ) ;
INV     gate1911  (.A(II6028), .Z(g2880) ) ;
INV     gate1912  (.A(g2209), .Z(II6031) ) ;
INV     gate1913  (.A(II6031), .Z(g2881) ) ;
INV     gate1914  (.A(g2210), .Z(II6034) ) ;
INV     gate1915  (.A(II6034), .Z(g2882) ) ;
INV     gate1916  (.A(g2560), .Z(II6037) ) ;
INV     gate1917  (.A(II6037), .Z(g2883) ) ;
INV     gate1918  (.A(g2216), .Z(II6040) ) ;
INV     gate1919  (.A(II6040), .Z(g2884) ) ;
INV     gate1920  (.A(g2267), .Z(II6043) ) ;
INV     gate1921  (.A(II6043), .Z(g2885) ) ;
INV     gate1922  (.A(g2218), .Z(II6046) ) ;
INV     gate1923  (.A(II6046), .Z(g2888) ) ;
INV     gate1924  (.A(g2219), .Z(II6049) ) ;
INV     gate1925  (.A(II6049), .Z(g2889) ) ;
INV     gate1926  (.A(g2220), .Z(II6052) ) ;
INV     gate1927  (.A(II6052), .Z(g2890) ) ;
INV     gate1928  (.A(g2569), .Z(II6055) ) ;
INV     gate1929  (.A(II6055), .Z(g2891) ) ;
INV     gate1930  (.A(g2356), .Z(g2896) ) ;
INV     gate1931  (.A(g2246), .Z(II6061) ) ;
INV     gate1932  (.A(II6061), .Z(g2902) ) ;
INV     gate1933  (.A(g2166), .Z(g2903) ) ;
INV     gate1934  (.A(g2226), .Z(II6065) ) ;
INV     gate1935  (.A(II6065), .Z(g2904) ) ;
INV     gate1936  (.A(g2227), .Z(II6068) ) ;
INV     gate1937  (.A(II6068), .Z(g2905) ) ;
INV     gate1938  (.A(g2269), .Z(II6071) ) ;
INV     gate1939  (.A(II6071), .Z(g2906) ) ;
INV     gate1940  (.A(g2228), .Z(II6074) ) ;
INV     gate1941  (.A(II6074), .Z(g2907) ) ;
INV     gate1942  (.A(g2349), .Z(II6077) ) ;
INV     gate1943  (.A(II6077), .Z(g2908) ) ;
INV     gate1944  (.A(g2108), .Z(II6080) ) ;
INV     gate1945  (.A(II6080), .Z(g2909) ) ;
INV     gate1946  (.A(g2234), .Z(II6085) ) ;
INV     gate1947  (.A(II6085), .Z(g2912) ) ;
INV     gate1948  (.A(g2235), .Z(II6088) ) ;
INV     gate1949  (.A(II6088), .Z(g2913) ) ;
INV     gate1950  (.A(g2270), .Z(II6091) ) ;
INV     gate1951  (.A(II6091), .Z(g2914) ) ;
INV     gate1952  (.A(g2110), .Z(II6094) ) ;
INV     gate1953  (.A(II6094), .Z(g2915) ) ;
INV     gate1954  (.A(g2391), .Z(II6097) ) ;
INV     gate1955  (.A(II6097), .Z(g2916) ) ;
INV     gate1956  (.A(g2240), .Z(II6102) ) ;
INV     gate1957  (.A(II6102), .Z(g2919) ) ;
INV     gate1958  (.A(g2462), .Z(g2920) ) ;
INV     gate1959  (.A(g2116), .Z(II6106) ) ;
INV     gate1960  (.A(II6106), .Z(g2937) ) ;
INV     gate1961  (.A(g2248), .Z(II6118) ) ;
INV     gate1962  (.A(II6118), .Z(g2941) ) ;
INV     gate1963  (.A(g2121), .Z(II6121) ) ;
INV     gate1964  (.A(II6121), .Z(g2942) ) ;
INV     gate1965  (.A(g2253), .Z(II6133) ) ;
INV     gate1966  (.A(II6133), .Z(g2946) ) ;
INV     gate1967  (.A(g2122), .Z(II6150) ) ;
INV     gate1968  (.A(II6150), .Z(g2949) ) ;
INV     gate1969  (.A(g2455), .Z(g2952) ) ;
INV     gate1970  (.A(g2119), .Z(II6156) ) ;
INV     gate1971  (.A(II6156), .Z(g2955) ) ;
INV     gate1972  (.A(g2123), .Z(II6159) ) ;
INV     gate1973  (.A(II6159), .Z(g2956) ) ;
INV     gate1974  (.A(g2547), .Z(II6163) ) ;
INV     gate1975  (.A(II6163), .Z(g2958) ) ;
INV     gate1976  (.A(g2125), .Z(II6173) ) ;
INV     gate1977  (.A(II6173), .Z(g2960) ) ;
INV     gate1978  (.A(g2131), .Z(II6183) ) ;
INV     gate1979  (.A(II6183), .Z(g2962) ) ;
INV     gate1980  (.A(g2155), .Z(II6193) ) ;
INV     gate1981  (.A(II6193), .Z(g2964) ) ;
INV     gate1982  (.A(g2462), .Z(II6196) ) ;
INV     gate1983  (.A(II6196), .Z(g2965) ) ;
INV     gate1984  (.A(g2046), .Z(g2971) ) ;
INV     gate1985  (.A(g1983), .Z(g2980) ) ;
INV     gate1986  (.A(g2302), .Z(II6217) ) ;
INV     gate1987  (.A(II6217), .Z(g2985) ) ;
INV     gate1988  (.A(g883), .Z(II6220) ) ;
INV     gate1989  (.A(g2135), .Z(g2989) ) ;
INV     gate1990  (.A(g2299), .Z(II6233) ) ;
INV     gate1991  (.A(II6233), .Z(g2991) ) ;
INV     gate1992  (.A(g2057), .Z(g2994) ) ;
INV     gate1993  (.A(g2135), .Z(g2997) ) ;
INV     gate1994  (.A(g2462), .Z(g2998) ) ;
INV     gate1995  (.A(g878), .Z(II6240) ) ;
INV     gate1996  (.A(g2135), .Z(g3009) ) ;
INV     gate1997  (.A(g2462), .Z(II6247) ) ;
INV     gate1998  (.A(II6247), .Z(g3012) ) ;
INV     gate1999  (.A(g2135), .Z(g3037) ) ;
INV     gate2000  (.A(g1982), .Z(g3038) ) ;
NAND2   gate2001  (.A(g591), .B(g605), .Z(g2310) ) ;
INV     gate2002  (.A(g2310), .Z(g3039) ) ;
INV     gate2003  (.A(g2135), .Z(g3040) ) ;
INV     gate2004  (.A(g2462), .Z(II6256) ) ;
INV     gate2005  (.A(II6256), .Z(g3044) ) ;
INV     gate2006  (.A(g2025), .Z(II6260) ) ;
INV     gate2007  (.A(II6260), .Z(g3050) ) ;
INV     gate2008  (.A(g2135), .Z(g3051) ) ;
INV     gate2009  (.A(g2118), .Z(II6264) ) ;
INV     gate2010  (.A(II6264), .Z(g3052) ) ;
INV     gate2011  (.A(g2135), .Z(g3055) ) ;
INV     gate2012  (.A(g2135), .Z(g3060) ) ;
INV     gate2013  (.A(g2135), .Z(g3066) ) ;
INV     gate2014  (.A(g2482), .Z(II6273) ) ;
INV     gate2015  (.A(II6273), .Z(g3067) ) ;
NAND2   gate2016  (.A(II5342), .B(II5343), .Z(g2303) ) ;
INV     gate2017  (.A(g2303), .Z(g3068) ) ;
INV     gate2018  (.A(g1206), .Z(II6277) ) ;
INV     gate2019  (.A(g2231), .Z(II6282) ) ;
INV     gate2020  (.A(II6282), .Z(g3076) ) ;
INV     gate2021  (.A(g2213), .Z(g3077) ) ;
INV     gate2022  (.A(g2276), .Z(g3086) ) ;
INV     gate2023  (.A(g2238), .Z(II6294) ) ;
INV     gate2024  (.A(II6294), .Z(g3088) ) ;
INV     gate2025  (.A(g2181), .Z(g3092) ) ;
INV     gate2026  (.A(g2242), .Z(II6299) ) ;
INV     gate2027  (.A(II6299), .Z(g3093) ) ;
INV     gate2028  (.A(g2243), .Z(II6302) ) ;
INV     gate2029  (.A(II6302), .Z(g3094) ) ;
INV     gate2030  (.A(g2482), .Z(g3095) ) ;
INV     gate2031  (.A(g2482), .Z(g3096) ) ;
INV     gate2032  (.A(g2482), .Z(g3097) ) ;
INV     gate2033  (.A(g2482), .Z(g3102) ) ;
INV     gate2034  (.A(g2391), .Z(g3103) ) ;
INV     gate2035  (.A(g2482), .Z(g3105) ) ;
INV     gate2036  (.A(g2482), .Z(g3109) ) ;
INV     gate2037  (.A(g2482), .Z(g3110) ) ;
INV     gate2038  (.A(g2482), .Z(g3112) ) ;
INV     gate2039  (.A(g1963), .Z(II6343) ) ;
INV     gate2040  (.A(II6343), .Z(g3113) ) ;
INV     gate2041  (.A(g2462), .Z(II6347) ) ;
INV     gate2042  (.A(II6347), .Z(g3119) ) ;
INV     gate2043  (.A(g2462), .Z(g3121) ) ;
NOR4    gate2044  (.A(g1645), .B(g1642), .C(g1651), .D(g1648), .Z(g2459) ) ;
INV     gate2045  (.A(g2459), .Z(II6356) ) ;
INV     gate2046  (.A(II6356), .Z(g3138) ) ;
AND2    gate2047  (.A(II5689), .B(II5690), .Z(g2563) ) ;
INV     gate2048  (.A(g2563), .Z(g3141) ) ;
INV     gate2049  (.A(g2261), .Z(II6360) ) ;
INV     gate2050  (.A(II6360), .Z(g3142) ) ;
INV     gate2051  (.A(g2459), .Z(II6363) ) ;
INV     gate2052  (.A(II6363), .Z(g3143) ) ;
INV     gate2053  (.A(g2462), .Z(g3144) ) ;
INV     gate2054  (.A(g2045), .Z(II6367) ) ;
INV     gate2055  (.A(II6367), .Z(g3161) ) ;
INV     gate2056  (.A(g2356), .Z(II6370) ) ;
INV     gate2057  (.A(II6370), .Z(g3164) ) ;
INV     gate2058  (.A(g2024), .Z(II6373) ) ;
INV     gate2059  (.A(II6373), .Z(g3186) ) ;
INV     gate2060  (.A(g2055), .Z(g3206) ) ;
NAND2   gate2061  (.A(g1814), .B(g1828), .Z(g2439) ) ;
INV     gate2062  (.A(g2439), .Z(g3207) ) ;
NAND2   gate2063  (.A(II5283), .B(II5284), .Z(g2257) ) ;
INV     gate2064  (.A(g2257), .Z(II6381) ) ;
INV     gate2065  (.A(II6381), .Z(g3208) ) ;
NAND2   gate2066  (.A(II5296), .B(II5297), .Z(g2260) ) ;
INV     gate2067  (.A(g2260), .Z(II6385) ) ;
INV     gate2068  (.A(II6385), .Z(g3212) ) ;
INV     gate2069  (.A(g2329), .Z(II6388) ) ;
INV     gate2070  (.A(II6388), .Z(g3213) ) ;
NOR2    gate2071  (.A(g1610), .B(g1737), .Z(g2478) ) ;
INV     gate2072  (.A(g2478), .Z(II6391) ) ;
INV     gate2073  (.A(II6391), .Z(g3214) ) ;
INV     gate2074  (.A(g2334), .Z(II6395) ) ;
INV     gate2075  (.A(II6395), .Z(g3219) ) ;
INV     gate2076  (.A(g2335), .Z(II6398) ) ;
INV     gate2077  (.A(II6398), .Z(g3220) ) ;
INV     gate2078  (.A(g2337), .Z(II6403) ) ;
INV     gate2079  (.A(II6403), .Z(g3226) ) ;
INV     gate2080  (.A(g2339), .Z(II6406) ) ;
INV     gate2081  (.A(II6406), .Z(g3227) ) ;
INV     gate2082  (.A(g2356), .Z(II6409) ) ;
INV     gate2083  (.A(II6409), .Z(g3228) ) ;
INV     gate2084  (.A(g2482), .Z(g3246) ) ;
INV     gate2085  (.A(g2342), .Z(II6414) ) ;
INV     gate2086  (.A(II6414), .Z(g3252) ) ;
INV     gate2087  (.A(g2344), .Z(II6417) ) ;
INV     gate2088  (.A(II6417), .Z(g3253) ) ;
INV     gate2089  (.A(g2322), .Z(g3254) ) ;
INV     gate2090  (.A(g2346), .Z(II6421) ) ;
INV     gate2091  (.A(II6421), .Z(g3255) ) ;
INV     gate2092  (.A(g2462), .Z(II6424) ) ;
INV     gate2093  (.A(II6424), .Z(g3256) ) ;
INV     gate2094  (.A(g2348), .Z(II6428) ) ;
INV     gate2095  (.A(II6428), .Z(g3260) ) ;
INV     gate2096  (.A(g2350), .Z(II6432) ) ;
INV     gate2097  (.A(II6432), .Z(g3262) ) ;
INV     gate2098  (.A(g2351), .Z(II6436) ) ;
INV     gate2099  (.A(II6436), .Z(g3266) ) ;
INV     gate2100  (.A(g2352), .Z(II6439) ) ;
INV     gate2101  (.A(II6439), .Z(g3267) ) ;
INV     gate2102  (.A(g2363), .Z(II6443) ) ;
INV     gate2103  (.A(II6443), .Z(g3271) ) ;
INV     gate2104  (.A(g2450), .Z(g3272) ) ;
INV     gate2105  (.A(g2368), .Z(II6454) ) ;
INV     gate2106  (.A(II6454), .Z(g3274) ) ;
INV     gate2107  (.A(g2261), .Z(II6461) ) ;
INV     gate2108  (.A(II6461), .Z(g3290) ) ;
AND2    gate2109  (.A(II5084), .B(II5085), .Z(g2161) ) ;
INV     gate2110  (.A(g2161), .Z(g3291) ) ;
INV     gate2111  (.A(g2373), .Z(g3292) ) ;
INV     gate2112  (.A(g2297), .Z(II6474) ) ;
INV     gate2113  (.A(II6474), .Z(g3305) ) ;
INV     gate2114  (.A(g2069), .Z(II6477) ) ;
INV     gate2115  (.A(II6477), .Z(g3306) ) ;
INV     gate2116  (.A(g2462), .Z(II6480) ) ;
INV     gate2117  (.A(II6480), .Z(g3307) ) ;
INV     gate2118  (.A(g2245), .Z(g3318) ) ;
INV     gate2119  (.A(g2073), .Z(II6484) ) ;
INV     gate2120  (.A(II6484), .Z(g3321) ) ;
INV     gate2121  (.A(g2157), .Z(g3323) ) ;
INV     gate2122  (.A(g2076), .Z(II6495) ) ;
INV     gate2123  (.A(II6495), .Z(g3326) ) ;
INV     gate2124  (.A(g2958), .Z(II6498) ) ;
INV     gate2125  (.A(g2578), .Z(II6501) ) ;
INV     gate2126  (.A(II6501), .Z(g3328) ) ;
INV     gate2127  (.A(g3214), .Z(II6504) ) ;
INV     gate2128  (.A(g2808), .Z(II6507) ) ;
INV     gate2129  (.A(II6507), .Z(g3330) ) ;
INV     gate2130  (.A(g3267), .Z(II6510) ) ;
INV     gate2131  (.A(II6510), .Z(g3331) ) ;
INV     gate2132  (.A(g2812), .Z(II6513) ) ;
INV     gate2133  (.A(II6513), .Z(g3332) ) ;
INV     gate2134  (.A(g2779), .Z(g3333) ) ;
INV     gate2135  (.A(g3271), .Z(II6517) ) ;
INV     gate2136  (.A(II6517), .Z(g3334) ) ;
INV     gate2137  (.A(g3186), .Z(II6520) ) ;
INV     gate2138  (.A(II6520), .Z(g3335) ) ;
INV     gate2139  (.A(g2819), .Z(II6523) ) ;
INV     gate2140  (.A(II6523), .Z(g3336) ) ;
INV     gate2141  (.A(g2745), .Z(g3337) ) ;
INV     gate2142  (.A(g2779), .Z(g3343) ) ;
INV     gate2143  (.A(g3274), .Z(II6528) ) ;
INV     gate2144  (.A(II6528), .Z(g3344) ) ;
INV     gate2145  (.A(g3186), .Z(II6531) ) ;
INV     gate2146  (.A(II6531), .Z(g3345) ) ;
INV     gate2147  (.A(g2733), .Z(g3348) ) ;
INV     gate2148  (.A(g2826), .Z(II6535) ) ;
INV     gate2149  (.A(II6535), .Z(g3351) ) ;
INV     gate2150  (.A(g2827), .Z(II6538) ) ;
INV     gate2151  (.A(II6538), .Z(g3352) ) ;
INV     gate2152  (.A(g3121), .Z(g3353) ) ;
INV     gate2153  (.A(g3186), .Z(II6543) ) ;
INV     gate2154  (.A(II6543), .Z(g3359) ) ;
NAND2   gate2155  (.A(g2481), .B(g883), .Z(g2987) ) ;
INV     gate2156  (.A(g2987), .Z(II6546) ) ;
INV     gate2157  (.A(II6546), .Z(g3362) ) ;
INV     gate2158  (.A(g2838), .Z(II6549) ) ;
INV     gate2159  (.A(II6549), .Z(g3363) ) ;
INV     gate2160  (.A(g3121), .Z(g3364) ) ;
INV     gate2161  (.A(g3186), .Z(II6553) ) ;
INV     gate2162  (.A(II6553), .Z(g3365) ) ;
INV     gate2163  (.A(g3138), .Z(g3368) ) ;
INV     gate2164  (.A(g3086), .Z(II6557) ) ;
INV     gate2165  (.A(II6557), .Z(g3369) ) ;
INV     gate2166  (.A(g2845), .Z(II6560) ) ;
INV     gate2167  (.A(II6560), .Z(g3370) ) ;
INV     gate2168  (.A(g2837), .Z(g3371) ) ;
INV     gate2169  (.A(g3121), .Z(g3372) ) ;
INV     gate2170  (.A(g2614), .Z(II6565) ) ;
INV     gate2171  (.A(II6565), .Z(g3373) ) ;
INV     gate2172  (.A(g3186), .Z(II6569) ) ;
INV     gate2173  (.A(II6569), .Z(g3375) ) ;
INV     gate2174  (.A(g2853), .Z(II6572) ) ;
INV     gate2175  (.A(II6572), .Z(g3378) ) ;
INV     gate2176  (.A(g3121), .Z(g3379) ) ;
INV     gate2177  (.A(g2617), .Z(II6576) ) ;
INV     gate2178  (.A(II6576), .Z(g3380) ) ;
INV     gate2179  (.A(g3186), .Z(II6580) ) ;
INV     gate2180  (.A(II6580), .Z(g3382) ) ;
INV     gate2181  (.A(g3143), .Z(g3384) ) ;
INV     gate2182  (.A(g3121), .Z(g3385) ) ;
INV     gate2183  (.A(g3144), .Z(g3386) ) ;
INV     gate2184  (.A(g2620), .Z(II6587) ) ;
INV     gate2185  (.A(II6587), .Z(g3387) ) ;
INV     gate2186  (.A(g3186), .Z(II6590) ) ;
INV     gate2187  (.A(II6590), .Z(g3388) ) ;
INV     gate2188  (.A(g3161), .Z(g3390) ) ;
INV     gate2189  (.A(g2896), .Z(g3391) ) ;
INV     gate2190  (.A(g3121), .Z(g3392) ) ;
INV     gate2191  (.A(g3144), .Z(g3393) ) ;
INV     gate2192  (.A(g2623), .Z(II6598) ) ;
INV     gate2193  (.A(II6598), .Z(g3394) ) ;
INV     gate2194  (.A(g3186), .Z(II6601) ) ;
INV     gate2195  (.A(II6601), .Z(g3395) ) ;
INV     gate2196  (.A(g2896), .Z(g3397) ) ;
INV     gate2197  (.A(g2896), .Z(g3398) ) ;
INV     gate2198  (.A(g3121), .Z(g3404) ) ;
INV     gate2199  (.A(g3144), .Z(g3405) ) ;
INV     gate2200  (.A(g2626), .Z(II6611) ) ;
INV     gate2201  (.A(II6611), .Z(g3406) ) ;
AND2    gate2202  (.A(II6330), .B(II6331), .Z(g3108) ) ;
INV     gate2203  (.A(g3108), .Z(g3408) ) ;
INV     gate2204  (.A(g3186), .Z(II6616) ) ;
INV     gate2205  (.A(II6616), .Z(g3411) ) ;
INV     gate2206  (.A(g2896), .Z(g3413) ) ;
INV     gate2207  (.A(g3121), .Z(g3415) ) ;
INV     gate2208  (.A(g3144), .Z(g3416) ) ;
INV     gate2209  (.A(g2629), .Z(II6624) ) ;
INV     gate2210  (.A(II6624), .Z(g3417) ) ;
AND2    gate2211  (.A(II6316), .B(II6317), .Z(g3104) ) ;
INV     gate2212  (.A(g3104), .Z(g3419) ) ;
INV     gate2213  (.A(g2896), .Z(g3424) ) ;
INV     gate2214  (.A(g3121), .Z(g3426) ) ;
INV     gate2215  (.A(g3144), .Z(g3427) ) ;
INV     gate2216  (.A(g2632), .Z(II6639) ) ;
INV     gate2217  (.A(II6639), .Z(g3428) ) ;
NAND2   gate2218  (.A(g2444), .B(g878), .Z(g3008) ) ;
INV     gate2219  (.A(g3008), .Z(II6643) ) ;
INV     gate2220  (.A(II6643), .Z(g3430) ) ;
INV     gate2221  (.A(g3144), .Z(g3432) ) ;
INV     gate2222  (.A(g2635), .Z(II6648) ) ;
INV     gate2223  (.A(II6648), .Z(g3433) ) ;
INV     gate2224  (.A(g3144), .Z(g3436) ) ;
INV     gate2225  (.A(g2952), .Z(II6654) ) ;
INV     gate2226  (.A(II6654), .Z(g3437) ) ;
INV     gate2227  (.A(g3144), .Z(g3439) ) ;
NAND4   gate2228  (.A(g2364), .B(g2399), .C(g2374), .D(g2382), .Z(g3041) ) ;
INV     gate2229  (.A(g3041), .Z(g3440) ) ;
INV     gate2230  (.A(g3144), .Z(g3458) ) ;
INV     gate2231  (.A(g2752), .Z(II6661) ) ;
INV     gate2232  (.A(II6661), .Z(g3459) ) ;
INV     gate2233  (.A(g2757), .Z(II6671) ) ;
INV     gate2234  (.A(II6671), .Z(g3461) ) ;
INV     gate2235  (.A(g3256), .Z(g3463) ) ;
INV     gate2236  (.A(g2759), .Z(II6676) ) ;
INV     gate2237  (.A(II6676), .Z(g3473) ) ;
INV     gate2238  (.A(g2902), .Z(II6679) ) ;
INV     gate2239  (.A(II6679), .Z(g3474) ) ;
NAND2   gate2240  (.A(g2374), .B(g599), .Z(g3056) ) ;
INV     gate2241  (.A(g3056), .Z(g3475) ) ;
INV     gate2242  (.A(g2655), .Z(g3479) ) ;
INV     gate2243  (.A(g2662), .Z(g3485) ) ;
INV     gate2244  (.A(g2669), .Z(g3491) ) ;
AND2    gate2245  (.A(g2028), .B(g2191), .Z(g3015) ) ;
INV     gate2246  (.A(g3015), .Z(II6686) ) ;
INV     gate2247  (.A(II6686), .Z(g3496) ) ;
INV     gate2248  (.A(g2743), .Z(II6690) ) ;
INV     gate2249  (.A(II6690), .Z(g3500) ) ;
INV     gate2250  (.A(g3077), .Z(g3501) ) ;
INV     gate2251  (.A(g2749), .Z(II6694) ) ;
INV     gate2252  (.A(II6694), .Z(g3505) ) ;
INV     gate2253  (.A(g3307), .Z(g3507) ) ;
INV     gate2254  (.A(g2801), .Z(II6702) ) ;
INV     gate2255  (.A(II6702), .Z(g3517) ) ;
INV     gate2256  (.A(g3164), .Z(g3518) ) ;
INV     gate2257  (.A(g3164), .Z(g3519) ) ;
INV     gate2258  (.A(g2779), .Z(g3520) ) ;
INV     gate2259  (.A(g3164), .Z(g3521) ) ;
INV     gate2260  (.A(g3164), .Z(g3522) ) ;
INV     gate2261  (.A(g2971), .Z(g3523) ) ;
INV     gate2262  (.A(g3164), .Z(g3528) ) ;
INV     gate2263  (.A(g2971), .Z(g3531) ) ;
INV     gate2264  (.A(g3164), .Z(g3532) ) ;
INV     gate2265  (.A(g3164), .Z(g3537) ) ;
INV     gate2266  (.A(g3306), .Z(II6726) ) ;
INV     gate2267  (.A(II6726), .Z(g3538) ) ;
INV     gate2268  (.A(g3015), .Z(g3539) ) ;
INV     gate2269  (.A(g3307), .Z(g3540) ) ;
AND2    gate2270  (.A(II6309), .B(II6310), .Z(g3101) ) ;
INV     gate2271  (.A(g3101), .Z(g3543) ) ;
INV     gate2272  (.A(g3164), .Z(g3544) ) ;
INV     gate2273  (.A(g3321), .Z(II6733) ) ;
INV     gate2274  (.A(II6733), .Z(g3545) ) ;
INV     gate2275  (.A(g3307), .Z(g3546) ) ;
INV     gate2276  (.A(g3113), .Z(II6738) ) ;
INV     gate2277  (.A(II6738), .Z(g3566) ) ;
INV     gate2278  (.A(g3164), .Z(g3582) ) ;
INV     gate2279  (.A(g3326), .Z(II6742) ) ;
INV     gate2280  (.A(II6742), .Z(g3583) ) ;
INV     gate2281  (.A(g2906), .Z(II6754) ) ;
INV     gate2282  (.A(II6754), .Z(g3621) ) ;
INV     gate2283  (.A(g2732), .Z(II6757) ) ;
INV     gate2284  (.A(II6757), .Z(g3622) ) ;
INV     gate2285  (.A(g2914), .Z(II6767) ) ;
INV     gate2286  (.A(II6767), .Z(g3624) ) ;
INV     gate2287  (.A(g2742), .Z(II6784) ) ;
INV     gate2288  (.A(II6784), .Z(g3627) ) ;
AND2    gate2289  (.A(II6337), .B(II6338), .Z(g3111) ) ;
INV     gate2290  (.A(g3111), .Z(g3628) ) ;
INV     gate2291  (.A(g3228), .Z(g3629) ) ;
INV     gate2292  (.A(g2748), .Z(II6789) ) ;
INV     gate2293  (.A(II6789), .Z(g3630) ) ;
INV     gate2294  (.A(g2750), .Z(II6799) ) ;
INV     gate2295  (.A(II6799), .Z(g3632) ) ;
INV     gate2296  (.A(g2751), .Z(II6802) ) ;
INV     gate2297  (.A(II6802), .Z(g3633) ) ;
INV     gate2298  (.A(g3290), .Z(II6812) ) ;
INV     gate2299  (.A(II6812), .Z(g3635) ) ;
INV     gate2300  (.A(g2755), .Z(II6815) ) ;
INV     gate2301  (.A(II6815), .Z(g3636) ) ;
INV     gate2302  (.A(g2758), .Z(II6818) ) ;
INV     gate2303  (.A(II6818), .Z(g3637) ) ;
INV     gate2304  (.A(g3015), .Z(II6821) ) ;
INV     gate2305  (.A(II6821), .Z(g3638) ) ;
INV     gate2306  (.A(g2909), .Z(II6832) ) ;
INV     gate2307  (.A(II6832), .Z(g3663) ) ;
NAND4   gate2308  (.A(g2550), .B(g2061), .C(g2564), .D(g2571), .Z(g3209) ) ;
INV     gate2309  (.A(g3209), .Z(g3664) ) ;
INV     gate2310  (.A(g2920), .Z(g3682) ) ;
INV     gate2311  (.A(g2915), .Z(II6844) ) ;
INV     gate2312  (.A(II6844), .Z(g3683) ) ;
INV     gate2313  (.A(g2920), .Z(g3693) ) ;
INV     gate2314  (.A(g2937), .Z(II6851) ) ;
INV     gate2315  (.A(II6851), .Z(g3694) ) ;
INV     gate2316  (.A(g3318), .Z(II6856) ) ;
INV     gate2317  (.A(II6856), .Z(g3697) ) ;
INV     gate2318  (.A(g2920), .Z(g3703) ) ;
INV     gate2319  (.A(g2942), .Z(II6861) ) ;
INV     gate2320  (.A(II6861), .Z(g3704) ) ;
INV     gate2321  (.A(g3113), .Z(g3705) ) ;
INV     gate2322  (.A(g2920), .Z(g3707) ) ;
INV     gate2323  (.A(g2949), .Z(II6867) ) ;
INV     gate2324  (.A(II6867), .Z(g3708) ) ;
INV     gate2325  (.A(g2852), .Z(II6870) ) ;
INV     gate2326  (.A(II6870), .Z(g3709) ) ;
NAND2   gate2327  (.A(g2564), .B(g1822), .Z(g3215) ) ;
INV     gate2328  (.A(g3215), .Z(g3710) ) ;
INV     gate2329  (.A(g2920), .Z(g3715) ) ;
INV     gate2330  (.A(g2956), .Z(II6876) ) ;
INV     gate2331  (.A(II6876), .Z(g3716) ) ;
INV     gate2332  (.A(g2920), .Z(g3719) ) ;
INV     gate2333  (.A(g2960), .Z(II6888) ) ;
INV     gate2334  (.A(II6888), .Z(g3720) ) ;
INV     gate2335  (.A(g2962), .Z(II6891) ) ;
INV     gate2336  (.A(II6891), .Z(g3721) ) ;
INV     gate2337  (.A(g2813), .Z(II6894) ) ;
INV     gate2338  (.A(II6894), .Z(g3722) ) ;
NAND3   gate2339  (.A(g605), .B(g2374), .C(g2382), .Z(g3071) ) ;
INV     gate2340  (.A(g3071), .Z(g3723) ) ;
INV     gate2341  (.A(g2964), .Z(II6898) ) ;
INV     gate2342  (.A(II6898), .Z(g3726) ) ;
INV     gate2343  (.A(g2818), .Z(II6901) ) ;
INV     gate2344  (.A(II6901), .Z(g3727) ) ;
INV     gate2345  (.A(g2820), .Z(II6904) ) ;
INV     gate2346  (.A(II6904), .Z(g3728) ) ;
INV     gate2347  (.A(g2994), .Z(II6907) ) ;
INV     gate2348  (.A(II6907), .Z(g3729) ) ;
INV     gate2349  (.A(g3015), .Z(g3730) ) ;
INV     gate2350  (.A(g2825), .Z(II6911) ) ;
INV     gate2351  (.A(II6911), .Z(g3731) ) ;
INV     gate2352  (.A(g2828), .Z(II6914) ) ;
INV     gate2353  (.A(II6914), .Z(g3732) ) ;
INV     gate2354  (.A(g2832), .Z(II6917) ) ;
INV     gate2355  (.A(II6917), .Z(g3733) ) ;
INV     gate2356  (.A(g2839), .Z(II6921) ) ;
INV     gate2357  (.A(II6921), .Z(g3735) ) ;
INV     gate2358  (.A(g2843), .Z(II6924) ) ;
INV     gate2359  (.A(II6924), .Z(g3736) ) ;
INV     gate2360  (.A(g2834), .Z(g3737) ) ;
NAND3   gate2361  (.A(g2369), .B(g591), .C(g611), .Z(g3062) ) ;
INV     gate2362  (.A(g3062), .Z(g3738) ) ;
INV     gate2363  (.A(g2846), .Z(II6929) ) ;
INV     gate2364  (.A(II6929), .Z(g3742) ) ;
INV     gate2365  (.A(g2850), .Z(II6932) ) ;
INV     gate2366  (.A(II6932), .Z(g3743) ) ;
INV     gate2367  (.A(g3307), .Z(g3744) ) ;
INV     gate2368  (.A(g3015), .Z(g3747) ) ;
INV     gate2369  (.A(g2971), .Z(g3748) ) ;
INV     gate2370  (.A(g2854), .Z(II6938) ) ;
INV     gate2371  (.A(II6938), .Z(g3749) ) ;
INV     gate2372  (.A(g2858), .Z(II6941) ) ;
INV     gate2373  (.A(II6941), .Z(g3750) ) ;
INV     gate2374  (.A(g2859), .Z(II6944) ) ;
INV     gate2375  (.A(II6944), .Z(g3751) ) ;
INV     gate2376  (.A(g2860), .Z(II6947) ) ;
INV     gate2377  (.A(II6947), .Z(g3752) ) ;
INV     gate2378  (.A(g3015), .Z(g3756) ) ;
INV     gate2379  (.A(g2867), .Z(II6952) ) ;
INV     gate2380  (.A(II6952), .Z(g3757) ) ;
INV     gate2381  (.A(g2871), .Z(II6955) ) ;
INV     gate2382  (.A(II6955), .Z(g3758) ) ;
INV     gate2383  (.A(g2872), .Z(II6958) ) ;
INV     gate2384  (.A(II6958), .Z(g3759) ) ;
NAND2   gate2385  (.A(g599), .B(g2399), .Z(g3003) ) ;
INV     gate2386  (.A(g3003), .Z(g3760) ) ;
NOR2    gate2387  (.A(g2187), .B(g750), .Z(g2791) ) ;
INV     gate2388  (.A(g2791), .Z(II6962) ) ;
INV     gate2389  (.A(II6962), .Z(g3761) ) ;
INV     gate2390  (.A(g2880), .Z(II6965) ) ;
INV     gate2391  (.A(II6965), .Z(g3762) ) ;
INV     gate2392  (.A(g2881), .Z(II6968) ) ;
INV     gate2393  (.A(II6968), .Z(g3763) ) ;
INV     gate2394  (.A(g2882), .Z(II6971) ) ;
INV     gate2395  (.A(II6971), .Z(g3764) ) ;
OR2     gate2396  (.A(II6350), .B(II6351), .Z(g3120) ) ;
INV     gate2397  (.A(g3120), .Z(g3765) ) ;
INV     gate2398  (.A(g2884), .Z(II6976) ) ;
INV     gate2399  (.A(II6976), .Z(g3767) ) ;
INV     gate2400  (.A(g2888), .Z(II6979) ) ;
INV     gate2401  (.A(II6979), .Z(g3768) ) ;
INV     gate2402  (.A(g2889), .Z(II6982) ) ;
INV     gate2403  (.A(II6982), .Z(g3769) ) ;
INV     gate2404  (.A(g2890), .Z(II6985) ) ;
INV     gate2405  (.A(II6985), .Z(g3770) ) ;
INV     gate2406  (.A(g2904), .Z(II6996) ) ;
INV     gate2407  (.A(II6996), .Z(g3773) ) ;
INV     gate2408  (.A(g2905), .Z(II6999) ) ;
INV     gate2409  (.A(II6999), .Z(g3774) ) ;
INV     gate2410  (.A(g2907), .Z(II7002) ) ;
INV     gate2411  (.A(II7002), .Z(g3775) ) ;
INV     gate2412  (.A(g2579), .Z(g3776) ) ;
INV     gate2413  (.A(g2912), .Z(II7006) ) ;
INV     gate2414  (.A(II7006), .Z(g3782) ) ;
INV     gate2415  (.A(g2913), .Z(II7009) ) ;
INV     gate2416  (.A(II7009), .Z(g3783) ) ;
INV     gate2417  (.A(g2586), .Z(g3784) ) ;
INV     gate2418  (.A(g3228), .Z(g3790) ) ;
INV     gate2419  (.A(g2919), .Z(II7014) ) ;
INV     gate2420  (.A(II7014), .Z(g3791) ) ;
INV     gate2421  (.A(g3068), .Z(II7017) ) ;
INV     gate2422  (.A(II7017), .Z(g3792) ) ;
INV     gate2423  (.A(g2593), .Z(g3793) ) ;
INV     gate2424  (.A(g3228), .Z(g3798) ) ;
INV     gate2425  (.A(g2941), .Z(II7022) ) ;
INV     gate2426  (.A(II7022), .Z(g3799) ) ;
INV     gate2427  (.A(g3292), .Z(g3800) ) ;
INV     gate2428  (.A(g3228), .Z(g3810) ) ;
INV     gate2429  (.A(g2946), .Z(II7029) ) ;
INV     gate2430  (.A(II7029), .Z(g3811) ) ;
INV     gate2431  (.A(g3228), .Z(g3812) ) ;
INV     gate2432  (.A(g3228), .Z(g3814) ) ;
INV     gate2433  (.A(g3228), .Z(g3815) ) ;
INV     gate2434  (.A(g3228), .Z(g3816) ) ;
INV     gate2435  (.A(g2908), .Z(II7043) ) ;
INV     gate2436  (.A(II7043), .Z(g3817) ) ;
NOR2    gate2437  (.A(g22), .B(g2320), .Z(g2807) ) ;
INV     gate2438  (.A(g2807), .Z(II7048) ) ;
INV     gate2439  (.A(II7048), .Z(g3820) ) ;
INV     gate2440  (.A(g2920), .Z(g3828) ) ;
INV     gate2441  (.A(g3093), .Z(II7054) ) ;
INV     gate2442  (.A(II7054), .Z(g3861) ) ;
INV     gate2443  (.A(g2920), .Z(g3862) ) ;
INV     gate2444  (.A(g2920), .Z(g3874) ) ;
INV     gate2445  (.A(g3050), .Z(II7061) ) ;
INV     gate2446  (.A(II7061), .Z(g3876) ) ;
OR2     gate2447  (.A(g2528), .B(g2522), .Z(g2984) ) ;
INV     gate2448  (.A(g2984), .Z(II7064) ) ;
INV     gate2449  (.A(II7064), .Z(g3877) ) ;
INV     gate2450  (.A(g2920), .Z(g3878) ) ;
INV     gate2451  (.A(g3138), .Z(II7070) ) ;
INV     gate2452  (.A(II7070), .Z(g3903) ) ;
INV     gate2453  (.A(g2920), .Z(g3905) ) ;
INV     gate2454  (.A(g3015), .Z(g3906) ) ;
INV     gate2455  (.A(g2985), .Z(II7076) ) ;
INV     gate2456  (.A(II7076), .Z(g3907) ) ;
INV     gate2457  (.A(g2920), .Z(g3909) ) ;
INV     gate2458  (.A(g3015), .Z(g3910) ) ;
INV     gate2459  (.A(g3015), .Z(g3911) ) ;
INV     gate2460  (.A(g2920), .Z(g3913) ) ;
INV     gate2461  (.A(g3015), .Z(g3914) ) ;
INV     gate2462  (.A(g3142), .Z(II7086) ) ;
INV     gate2463  (.A(II7086), .Z(g3937) ) ;
INV     gate2464  (.A(g2991), .Z(g3938) ) ;
INV     gate2465  (.A(g2920), .Z(g3940) ) ;
INV     gate2466  (.A(g3015), .Z(g3941) ) ;
INV     gate2467  (.A(g2779), .Z(g3943) ) ;
INV     gate2468  (.A(g2920), .Z(g3944) ) ;
INV     gate2469  (.A(g3186), .Z(II7096) ) ;
INV     gate2470  (.A(II7096), .Z(g3945) ) ;
INV     gate2471  (.A(g3228), .Z(II7099) ) ;
INV     gate2472  (.A(II7099), .Z(g3946) ) ;
NAND3   gate2473  (.A(g1828), .B(g2564), .C(g2571), .Z(g3247) ) ;
INV     gate2474  (.A(g3247), .Z(g3967) ) ;
INV     gate2475  (.A(g3186), .Z(II7104) ) ;
INV     gate2476  (.A(II7104), .Z(g3971) ) ;
INV     gate2477  (.A(g3121), .Z(g3975) ) ;
NAND2   gate2478  (.A(II6200), .B(II6201), .Z(g2970) ) ;
INV     gate2479  (.A(g2970), .Z(II7109) ) ;
INV     gate2480  (.A(II7109), .Z(g3976) ) ;
INV     gate2481  (.A(g3186), .Z(II7112) ) ;
INV     gate2482  (.A(II7112), .Z(g3977) ) ;
INV     gate2483  (.A(g3121), .Z(g3980) ) ;
NAND2   gate2484  (.A(II6208), .B(II6209), .Z(g2979) ) ;
INV     gate2485  (.A(g2979), .Z(II7118) ) ;
INV     gate2486  (.A(II7118), .Z(g3981) ) ;
INV     gate2487  (.A(g3052), .Z(g3982) ) ;
NAND3   gate2488  (.A(g2557), .B(g1814), .C(g1834), .Z(g3222) ) ;
INV     gate2489  (.A(g3222), .Z(g3983) ) ;
INV     gate2490  (.A(g3121), .Z(g3988) ) ;
INV     gate2491  (.A(g3121), .Z(g3990) ) ;
INV     gate2492  (.A(g3121), .Z(g3995) ) ;
INV     gate2493  (.A(g3144), .Z(g3996) ) ;
INV     gate2494  (.A(g2640), .Z(II7131) ) ;
INV     gate2495  (.A(II7131), .Z(g3997) ) ;
NAND2   gate2496  (.A(g1822), .B(g2061), .Z(g3200) ) ;
INV     gate2497  (.A(g3200), .Z(g4001) ) ;
INV     gate2498  (.A(g3121), .Z(g4002) ) ;
INV     gate2499  (.A(g3144), .Z(g4003) ) ;
INV     gate2500  (.A(g2641), .Z(II7140) ) ;
INV     gate2501  (.A(II7140), .Z(g4004) ) ;
INV     gate2502  (.A(g2614), .Z(II7143) ) ;
INV     gate2503  (.A(II7143), .Z(g4005) ) ;
INV     gate2504  (.A(g3144), .Z(g4010) ) ;
INV     gate2505  (.A(g2642), .Z(II7151) ) ;
INV     gate2506  (.A(II7151), .Z(g4011) ) ;
INV     gate2507  (.A(g2617), .Z(II7154) ) ;
INV     gate2508  (.A(II7154), .Z(g4012) ) ;
INV     gate2509  (.A(g3015), .Z(II7157) ) ;
INV     gate2510  (.A(II7157), .Z(g4013) ) ;
INV     gate2511  (.A(g3144), .Z(g4049) ) ;
INV     gate2512  (.A(g2643), .Z(II7163) ) ;
INV     gate2513  (.A(II7163), .Z(g4050) ) ;
INV     gate2514  (.A(g2620), .Z(II7166) ) ;
INV     gate2515  (.A(II7166), .Z(g4051) ) ;
INV     gate2516  (.A(g3144), .Z(g4055) ) ;
INV     gate2517  (.A(g2644), .Z(II7173) ) ;
INV     gate2518  (.A(II7173), .Z(g4056) ) ;
INV     gate2519  (.A(g2623), .Z(II7176) ) ;
INV     gate2520  (.A(II7176), .Z(g4057) ) ;
INV     gate2521  (.A(g3144), .Z(g4060) ) ;
INV     gate2522  (.A(g2645), .Z(II7182) ) ;
INV     gate2523  (.A(II7182), .Z(g4061) ) ;
INV     gate2524  (.A(g2626), .Z(II7185) ) ;
INV     gate2525  (.A(II7185), .Z(g4062) ) ;
AND2    gate2526  (.A(II5886), .B(II5887), .Z(g2794) ) ;
INV     gate2527  (.A(g2794), .Z(g4065) ) ;
INV     gate2528  (.A(g2646), .Z(II7191) ) ;
INV     gate2529  (.A(II7191), .Z(g4066) ) ;
INV     gate2530  (.A(g2629), .Z(II7194) ) ;
INV     gate2531  (.A(II7194), .Z(g4067) ) ;
INV     gate2532  (.A(g2647), .Z(II7202) ) ;
INV     gate2533  (.A(II7202), .Z(g4077) ) ;
INV     gate2534  (.A(g2632), .Z(II7205) ) ;
INV     gate2535  (.A(II7205), .Z(g4078) ) ;
INV     gate2536  (.A(g2903), .Z(g4080) ) ;
INV     gate2537  (.A(g2798), .Z(II7210) ) ;
INV     gate2538  (.A(II7210), .Z(g4081) ) ;
INV     gate2539  (.A(g2635), .Z(II7213) ) ;
INV     gate2540  (.A(II7213), .Z(g4082) ) ;
INV     gate2541  (.A(g2952), .Z(II7216) ) ;
INV     gate2542  (.A(II7216), .Z(g4083) ) ;
INV     gate2543  (.A(g3119), .Z(g4084) ) ;
INV     gate2544  (.A(g3213), .Z(II7220) ) ;
INV     gate2545  (.A(II7220), .Z(g4087) ) ;
INV     gate2546  (.A(g2965), .Z(g4093) ) ;
OR2     gate2547  (.A(II5804), .B(II5805), .Z(g2744) ) ;
INV     gate2548  (.A(g2744), .Z(g4094) ) ;
INV     gate2549  (.A(g2817), .Z(II7233) ) ;
INV     gate2550  (.A(II7233), .Z(g4095) ) ;
INV     gate2551  (.A(g3219), .Z(II7236) ) ;
INV     gate2552  (.A(II7236), .Z(g4096) ) ;
INV     gate2553  (.A(g2824), .Z(II7240) ) ;
INV     gate2554  (.A(II7240), .Z(g4098) ) ;
INV     gate2555  (.A(g3226), .Z(II7244) ) ;
INV     gate2556  (.A(II7244), .Z(g4102) ) ;
INV     gate2557  (.A(g2833), .Z(II7249) ) ;
INV     gate2558  (.A(II7249), .Z(g4105) ) ;
INV     gate2559  (.A(g2994), .Z(g4112) ) ;
INV     gate2560  (.A(g3227), .Z(II7255) ) ;
INV     gate2561  (.A(II7255), .Z(g4113) ) ;
INV     gate2562  (.A(g2844), .Z(II7260) ) ;
INV     gate2563  (.A(II7260), .Z(g4116) ) ;
INV     gate2564  (.A(g3252), .Z(II7264) ) ;
INV     gate2565  (.A(II7264), .Z(g4121) ) ;
INV     gate2566  (.A(g2851), .Z(II7269) ) ;
INV     gate2567  (.A(II7269), .Z(g4124) ) ;
INV     gate2568  (.A(g3253), .Z(II7272) ) ;
INV     gate2569  (.A(II7272), .Z(g4125) ) ;
INV     gate2570  (.A(g2861), .Z(II7276) ) ;
INV     gate2571  (.A(II7276), .Z(g4127) ) ;
INV     gate2572  (.A(g3208), .Z(II7280) ) ;
INV     gate2573  (.A(II7280), .Z(g4129) ) ;
INV     gate2574  (.A(g3255), .Z(II7284) ) ;
INV     gate2575  (.A(II7284), .Z(g4140) ) ;
INV     gate2576  (.A(g2873), .Z(II7288) ) ;
INV     gate2577  (.A(II7288), .Z(g4142) ) ;
INV     gate2578  (.A(g3212), .Z(II7291) ) ;
INV     gate2579  (.A(II7291), .Z(g4143) ) ;
INV     gate2580  (.A(g3260), .Z(II7295) ) ;
INV     gate2581  (.A(II7295), .Z(g4156) ) ;
NAND2   gate2582  (.A(II6468), .B(II6469), .Z(g3304) ) ;
INV     gate2583  (.A(g3304), .Z(g4158) ) ;
INV     gate2584  (.A(g2883), .Z(II7300) ) ;
INV     gate2585  (.A(II7300), .Z(g4159) ) ;
INV     gate2586  (.A(g3262), .Z(II7303) ) ;
INV     gate2587  (.A(II7303), .Z(g4160) ) ;
NAND2   gate2588  (.A(g2016), .B(g1206), .Z(g3070) ) ;
INV     gate2589  (.A(g3070), .Z(II7308) ) ;
INV     gate2590  (.A(II7308), .Z(g4163) ) ;
INV     gate2591  (.A(g2803), .Z(II7311) ) ;
INV     gate2592  (.A(II7311), .Z(g4164) ) ;
INV     gate2593  (.A(g3164), .Z(g4165) ) ;
INV     gate2594  (.A(g2891), .Z(II7315) ) ;
INV     gate2595  (.A(II7315), .Z(g4166) ) ;
INV     gate2596  (.A(g3266), .Z(II7318) ) ;
INV     gate2597  (.A(II7318), .Z(g4167) ) ;
INV     gate2598  (.A(g3328), .Z(g4170) ) ;
INV     gate2599  (.A(g3761), .Z(II7330) ) ;
INV     gate2600  (.A(g3729), .Z(II7333) ) ;
INV     gate2601  (.A(g3997), .Z(II7336) ) ;
INV     gate2602  (.A(g4004), .Z(II7339) ) ;
INV     gate2603  (.A(g4011), .Z(II7342) ) ;
INV     gate2604  (.A(g4050), .Z(II7345) ) ;
INV     gate2605  (.A(g4056), .Z(II7348) ) ;
INV     gate2606  (.A(g4061), .Z(II7351) ) ;
INV     gate2607  (.A(g4066), .Z(II7354) ) ;
INV     gate2608  (.A(g4077), .Z(II7357) ) ;
INV     gate2609  (.A(g4081), .Z(II7360) ) ;
INV     gate2610  (.A(g4005), .Z(II7363) ) ;
INV     gate2611  (.A(g4012), .Z(II7366) ) ;
INV     gate2612  (.A(g4051), .Z(II7369) ) ;
INV     gate2613  (.A(g4057), .Z(II7372) ) ;
INV     gate2614  (.A(g4062), .Z(II7375) ) ;
INV     gate2615  (.A(g4067), .Z(II7378) ) ;
INV     gate2616  (.A(g4078), .Z(II7381) ) ;
INV     gate2617  (.A(g4082), .Z(II7384) ) ;
INV     gate2618  (.A(g4083), .Z(II7387) ) ;
INV     gate2619  (.A(g4087), .Z(II7390) ) ;
INV     gate2620  (.A(g4096), .Z(II7393) ) ;
INV     gate2621  (.A(g4102), .Z(II7396) ) ;
INV     gate2622  (.A(g4113), .Z(II7399) ) ;
INV     gate2623  (.A(g4121), .Z(II7402) ) ;
INV     gate2624  (.A(g3861), .Z(II7405) ) ;
INV     gate2625  (.A(g4125), .Z(II7408) ) ;
INV     gate2626  (.A(g4140), .Z(II7411) ) ;
INV     gate2627  (.A(g4156), .Z(II7414) ) ;
INV     gate2628  (.A(g4160), .Z(II7417) ) ;
INV     gate2629  (.A(g4167), .Z(II7420) ) ;
INV     gate2630  (.A(g3331), .Z(II7423) ) ;
INV     gate2631  (.A(g3334), .Z(II7426) ) ;
INV     gate2632  (.A(g3344), .Z(II7429) ) ;
INV     gate2633  (.A(g3663), .Z(II7432) ) ;
INV     gate2634  (.A(g3459), .Z(II7435) ) ;
INV     gate2635  (.A(g3461), .Z(II7438) ) ;
INV     gate2636  (.A(g3473), .Z(II7441) ) ;
INV     gate2637  (.A(g3683), .Z(II7444) ) ;
INV     gate2638  (.A(g3694), .Z(II7447) ) ;
INV     gate2639  (.A(g3704), .Z(II7450) ) ;
INV     gate2640  (.A(g3708), .Z(II7453) ) ;
INV     gate2641  (.A(g3716), .Z(II7456) ) ;
INV     gate2642  (.A(g3720), .Z(II7459) ) ;
INV     gate2643  (.A(g3721), .Z(II7462) ) ;
INV     gate2644  (.A(g3726), .Z(II7465) ) ;
INV     gate2645  (.A(g3697), .Z(II7468) ) ;
INV     gate2646  (.A(g3635), .Z(g4219) ) ;
INV     gate2647  (.A(g3914), .Z(g4221) ) ;
INV     gate2648  (.A(g3638), .Z(g4222) ) ;
INV     gate2649  (.A(g3566), .Z(II7478) ) ;
INV     gate2650  (.A(II7478), .Z(g4225) ) ;
OR2     gate2651  (.A(g3121), .B(g2480), .Z(g3698) ) ;
INV     gate2652  (.A(g3698), .Z(g4226) ) ;
INV     gate2653  (.A(g3914), .Z(g4228) ) ;
INV     gate2654  (.A(g3371), .Z(II7487) ) ;
INV     gate2655  (.A(II7487), .Z(g4232) ) ;
INV     gate2656  (.A(g3698), .Z(g4233) ) ;
INV     gate2657  (.A(g4013), .Z(g4237) ) ;
INV     gate2658  (.A(g3664), .Z(g4240) ) ;
INV     gate2659  (.A(g3664), .Z(g4241) ) ;
INV     gate2660  (.A(g3664), .Z(g4242) ) ;
NAND2   gate2661  (.A(g3209), .B(g3221), .Z(g3524) ) ;
INV     gate2662  (.A(g3524), .Z(g4243) ) ;
INV     gate2663  (.A(g3698), .Z(g4250) ) ;
INV     gate2664  (.A(g4013), .Z(g4254) ) ;
INV     gate2665  (.A(g3664), .Z(g4256) ) ;
INV     gate2666  (.A(g3664), .Z(g4257) ) ;
INV     gate2667  (.A(g3566), .Z(II7509) ) ;
INV     gate2668  (.A(II7509), .Z(g4258) ) ;
NAND2   gate2669  (.A(g2160), .B(g3044), .Z(g4144) ) ;
INV     gate2670  (.A(g4144), .Z(II7513) ) ;
INV     gate2671  (.A(II7513), .Z(g4260) ) ;
INV     gate2672  (.A(g4013), .Z(g4262) ) ;
AND2    gate2673  (.A(g3323), .B(g2191), .Z(g3586) ) ;
INV     gate2674  (.A(g3586), .Z(g4263) ) ;
INV     gate2675  (.A(g3664), .Z(g4265) ) ;
OR2     gate2676  (.A(g3144), .B(g2454), .Z(g3688) ) ;
INV     gate2677  (.A(g3688), .Z(g4266) ) ;
INV     gate2678  (.A(g4095), .Z(II7523) ) ;
INV     gate2679  (.A(II7523), .Z(g4268) ) ;
INV     gate2680  (.A(g4013), .Z(g4270) ) ;
INV     gate2681  (.A(g3971), .Z(g4271) ) ;
INV     gate2682  (.A(g3586), .Z(g4272) ) ;
INV     gate2683  (.A(g4013), .Z(g4273) ) ;
INV     gate2684  (.A(g3664), .Z(g4275) ) ;
INV     gate2685  (.A(g3688), .Z(g4277) ) ;
INV     gate2686  (.A(g4098), .Z(II7536) ) ;
INV     gate2687  (.A(II7536), .Z(g4279) ) ;
INV     gate2688  (.A(g4013), .Z(g4280) ) ;
INV     gate2689  (.A(g3586), .Z(g4281) ) ;
INV     gate2690  (.A(g4013), .Z(g4282) ) ;
INV     gate2691  (.A(g3664), .Z(g4284) ) ;
INV     gate2692  (.A(g3688), .Z(g4285) ) ;
INV     gate2693  (.A(g4105), .Z(II7546) ) ;
INV     gate2694  (.A(II7546), .Z(g4287) ) ;
NAND2   gate2695  (.A(g3044), .B(g2518), .Z(g4130) ) ;
INV     gate2696  (.A(g4130), .Z(g4288) ) ;
INV     gate2697  (.A(g4013), .Z(g4289) ) ;
INV     gate2698  (.A(g3586), .Z(g4290) ) ;
INV     gate2699  (.A(g4013), .Z(g4291) ) ;
AND2    gate2700  (.A(g3323), .B(g2728), .Z(g3863) ) ;
INV     gate2701  (.A(g3863), .Z(g4292) ) ;
INV     gate2702  (.A(g3664), .Z(g4294) ) ;
INV     gate2703  (.A(g4080), .Z(II7556) ) ;
INV     gate2704  (.A(II7556), .Z(g4295) ) ;
INV     gate2705  (.A(g4116), .Z(II7559) ) ;
INV     gate2706  (.A(II7559), .Z(g4296) ) ;
INV     gate2707  (.A(g4130), .Z(g4298) ) ;
INV     gate2708  (.A(g4144), .Z(g4299) ) ;
INV     gate2709  (.A(g4013), .Z(g4305) ) ;
INV     gate2710  (.A(g3586), .Z(g4306) ) ;
INV     gate2711  (.A(g4013), .Z(g4307) ) ;
INV     gate2712  (.A(g3863), .Z(g4308) ) ;
INV     gate2713  (.A(g4124), .Z(II7577) ) ;
INV     gate2714  (.A(II7577), .Z(g4310) ) ;
INV     gate2715  (.A(g4130), .Z(g4311) ) ;
INV     gate2716  (.A(g4144), .Z(g4312) ) ;
INV     gate2717  (.A(g3586), .Z(g4313) ) ;
INV     gate2718  (.A(g4013), .Z(g4314) ) ;
INV     gate2719  (.A(g3863), .Z(g4315) ) ;
INV     gate2720  (.A(g4127), .Z(II7586) ) ;
INV     gate2721  (.A(II7586), .Z(g4317) ) ;
INV     gate2722  (.A(g4130), .Z(g4318) ) ;
INV     gate2723  (.A(g4144), .Z(g4319) ) ;
INV     gate2724  (.A(g4013), .Z(g4320) ) ;
INV     gate2725  (.A(g3863), .Z(g4321) ) ;
INV     gate2726  (.A(g4142), .Z(II7593) ) ;
INV     gate2727  (.A(II7593), .Z(g4322) ) ;
INV     gate2728  (.A(g4130), .Z(g4323) ) ;
INV     gate2729  (.A(g4144), .Z(g4324) ) ;
INV     gate2730  (.A(g3863), .Z(g4326) ) ;
INV     gate2731  (.A(g4159), .Z(II7600) ) ;
INV     gate2732  (.A(II7600), .Z(g4327) ) ;
INV     gate2733  (.A(g4130), .Z(g4328) ) ;
INV     gate2734  (.A(g4144), .Z(g4329) ) ;
INV     gate2735  (.A(g4166), .Z(II7606) ) ;
INV     gate2736  (.A(II7606), .Z(g4331) ) ;
INV     gate2737  (.A(g4130), .Z(g4332) ) ;
INV     gate2738  (.A(g4144), .Z(g4333) ) ;
INV     gate2739  (.A(g3817), .Z(II7612) ) ;
INV     gate2740  (.A(II7612), .Z(g4335) ) ;
INV     gate2741  (.A(g4130), .Z(g4336) ) ;
INV     gate2742  (.A(g4144), .Z(g4337) ) ;
INV     gate2743  (.A(g4144), .Z(g4339) ) ;
INV     gate2744  (.A(g3946), .Z(g4344) ) ;
INV     gate2745  (.A(g4164), .Z(II7625) ) ;
INV     gate2746  (.A(II7625), .Z(g4346) ) ;
AND2    gate2747  (.A(g3186), .B(g2023), .Z(g3880) ) ;
INV     gate2748  (.A(g3880), .Z(g4347) ) ;
INV     gate2749  (.A(g3524), .Z(II7630) ) ;
INV     gate2750  (.A(II7630), .Z(g4351) ) ;
INV     gate2751  (.A(g3474), .Z(II7633) ) ;
INV     gate2752  (.A(II7633), .Z(g4352) ) ;
INV     gate2753  (.A(g3330), .Z(II7636) ) ;
INV     gate2754  (.A(II7636), .Z(g4353) ) ;
INV     gate2755  (.A(g3722), .Z(II7639) ) ;
INV     gate2756  (.A(II7639), .Z(g4354) ) ;
INV     gate2757  (.A(g3440), .Z(II7642) ) ;
INV     gate2758  (.A(II7642), .Z(g4355) ) ;
INV     gate2759  (.A(g3880), .Z(g4359) ) ;
INV     gate2760  (.A(g3727), .Z(II7648) ) ;
INV     gate2761  (.A(II7648), .Z(g4361) ) ;
INV     gate2762  (.A(g3332), .Z(II7651) ) ;
INV     gate2763  (.A(II7651), .Z(g4362) ) ;
INV     gate2764  (.A(g3728), .Z(II7654) ) ;
INV     gate2765  (.A(II7654), .Z(g4363) ) ;
INV     gate2766  (.A(g3880), .Z(g4365) ) ;
INV     gate2767  (.A(g3731), .Z(II7659) ) ;
INV     gate2768  (.A(II7659), .Z(g4366) ) ;
INV     gate2769  (.A(g3336), .Z(II7662) ) ;
INV     gate2770  (.A(II7662), .Z(g4367) ) ;
INV     gate2771  (.A(g3732), .Z(II7665) ) ;
INV     gate2772  (.A(II7665), .Z(g4368) ) ;
INV     gate2773  (.A(g3733), .Z(II7668) ) ;
INV     gate2774  (.A(II7668), .Z(g4369) ) ;
INV     gate2775  (.A(g3351), .Z(II7671) ) ;
INV     gate2776  (.A(II7671), .Z(g4370) ) ;
INV     gate2777  (.A(g3352), .Z(II7674) ) ;
INV     gate2778  (.A(II7674), .Z(g4371) ) ;
INV     gate2779  (.A(g3735), .Z(II7677) ) ;
INV     gate2780  (.A(II7677), .Z(g4372) ) ;
INV     gate2781  (.A(g3736), .Z(II7680) ) ;
INV     gate2782  (.A(II7680), .Z(g4373) ) ;
INV     gate2783  (.A(g3638), .Z(g4375) ) ;
INV     gate2784  (.A(g3363), .Z(II7691) ) ;
INV     gate2785  (.A(II7691), .Z(g4376) ) ;
INV     gate2786  (.A(g3742), .Z(II7694) ) ;
INV     gate2787  (.A(II7694), .Z(g4377) ) ;
INV     gate2788  (.A(g3743), .Z(II7697) ) ;
INV     gate2789  (.A(II7697), .Z(g4378) ) ;
INV     gate2790  (.A(g3698), .Z(g4379) ) ;
OR2     gate2791  (.A(g3118), .B(g2180), .Z(g3513) ) ;
INV     gate2792  (.A(g3513), .Z(II7701) ) ;
INV     gate2793  (.A(II7701), .Z(g4380) ) ;
INV     gate2794  (.A(g3914), .Z(g4381) ) ;
INV     gate2795  (.A(g3638), .Z(g4382) ) ;
INV     gate2796  (.A(g3370), .Z(II7707) ) ;
INV     gate2797  (.A(II7707), .Z(g4384) ) ;
INV     gate2798  (.A(g3749), .Z(II7710) ) ;
INV     gate2799  (.A(II7710), .Z(g4385) ) ;
INV     gate2800  (.A(g3750), .Z(II7713) ) ;
INV     gate2801  (.A(II7713), .Z(g4386) ) ;
INV     gate2802  (.A(g3751), .Z(II7716) ) ;
INV     gate2803  (.A(II7716), .Z(g4387) ) ;
INV     gate2804  (.A(g3752), .Z(II7719) ) ;
INV     gate2805  (.A(II7719), .Z(g4388) ) ;
INV     gate2806  (.A(g3914), .Z(g4390) ) ;
INV     gate2807  (.A(g3638), .Z(g4391) ) ;
INV     gate2808  (.A(g3378), .Z(II7726) ) ;
INV     gate2809  (.A(II7726), .Z(g4393) ) ;
INV     gate2810  (.A(g3757), .Z(II7729) ) ;
INV     gate2811  (.A(II7729), .Z(g4394) ) ;
INV     gate2812  (.A(g3758), .Z(II7732) ) ;
INV     gate2813  (.A(II7732), .Z(g4395) ) ;
INV     gate2814  (.A(g3759), .Z(II7735) ) ;
INV     gate2815  (.A(II7735), .Z(g4396) ) ;
INV     gate2816  (.A(g3914), .Z(g4398) ) ;
INV     gate2817  (.A(g3638), .Z(g4399) ) ;
INV     gate2818  (.A(g3762), .Z(II7743) ) ;
INV     gate2819  (.A(II7743), .Z(g4411) ) ;
INV     gate2820  (.A(g3763), .Z(II7746) ) ;
INV     gate2821  (.A(II7746), .Z(g4412) ) ;
INV     gate2822  (.A(g3764), .Z(II7749) ) ;
INV     gate2823  (.A(II7749), .Z(g4413) ) ;
AND2    gate2824  (.A(g2561), .B(g3012), .Z(g3407) ) ;
INV     gate2825  (.A(g3407), .Z(II7752) ) ;
INV     gate2826  (.A(II7752), .Z(g4414) ) ;
INV     gate2827  (.A(g3914), .Z(g4415) ) ;
INV     gate2828  (.A(g3638), .Z(g4416) ) ;
INV     gate2829  (.A(g3767), .Z(II7757) ) ;
INV     gate2830  (.A(II7757), .Z(g4417) ) ;
INV     gate2831  (.A(g3768), .Z(II7760) ) ;
INV     gate2832  (.A(II7760), .Z(g4418) ) ;
INV     gate2833  (.A(g3769), .Z(II7763) ) ;
INV     gate2834  (.A(II7763), .Z(g4419) ) ;
INV     gate2835  (.A(g3770), .Z(II7766) ) ;
INV     gate2836  (.A(II7766), .Z(g4420) ) ;
INV     gate2837  (.A(g3688), .Z(g4424) ) ;
AND2    gate2838  (.A(g2379), .B(g3012), .Z(g3418) ) ;
INV     gate2839  (.A(g3418), .Z(II7771) ) ;
INV     gate2840  (.A(II7771), .Z(g4425) ) ;
INV     gate2841  (.A(g3914), .Z(g4426) ) ;
INV     gate2842  (.A(g3638), .Z(g4427) ) ;
INV     gate2843  (.A(g3773), .Z(II7776) ) ;
INV     gate2844  (.A(II7776), .Z(g4428) ) ;
INV     gate2845  (.A(g3774), .Z(II7779) ) ;
INV     gate2846  (.A(II7779), .Z(g4429) ) ;
INV     gate2847  (.A(g3775), .Z(II7782) ) ;
INV     gate2848  (.A(II7782), .Z(g4430) ) ;
INV     gate2849  (.A(g3914), .Z(g4435) ) ;
INV     gate2850  (.A(g3638), .Z(g4436) ) ;
INV     gate2851  (.A(g3345), .Z(g4437) ) ;
INV     gate2852  (.A(g3782), .Z(II7790) ) ;
INV     gate2853  (.A(II7790), .Z(g4438) ) ;
INV     gate2854  (.A(g3783), .Z(II7793) ) ;
INV     gate2855  (.A(II7793), .Z(g4439) ) ;
INV     gate2856  (.A(g4130), .Z(g4440) ) ;
INV     gate2857  (.A(g3914), .Z(g4441) ) ;
INV     gate2858  (.A(g3638), .Z(g4442) ) ;
INV     gate2859  (.A(g3359), .Z(g4443) ) ;
INV     gate2860  (.A(g3791), .Z(II7800) ) ;
INV     gate2861  (.A(II7800), .Z(g4444) ) ;
INV     gate2862  (.A(g3820), .Z(II7803) ) ;
INV     gate2863  (.A(II7803), .Z(g4445) ) ;
INV     gate2864  (.A(g4144), .Z(g4449) ) ;
INV     gate2865  (.A(g3914), .Z(g4450) ) ;
INV     gate2866  (.A(g3638), .Z(g4451) ) ;
INV     gate2867  (.A(g3365), .Z(g4452) ) ;
INV     gate2868  (.A(g3799), .Z(II7810) ) ;
INV     gate2869  (.A(II7810), .Z(g4453) ) ;
INV     gate2870  (.A(g3914), .Z(g4454) ) ;
INV     gate2871  (.A(g3375), .Z(g4456) ) ;
AND2    gate2872  (.A(g2028), .B(g2728), .Z(g3829) ) ;
INV     gate2873  (.A(g3829), .Z(g4457) ) ;
OR2     gate2874  (.A(g2918), .B(g2940), .Z(g3399) ) ;
INV     gate2875  (.A(g3399), .Z(II7817) ) ;
INV     gate2876  (.A(II7817), .Z(g4458) ) ;
INV     gate2877  (.A(g3811), .Z(II7820) ) ;
INV     gate2878  (.A(II7820), .Z(g4459) ) ;
INV     gate2879  (.A(g3820), .Z(g4460) ) ;
INV     gate2880  (.A(g3829), .Z(g4461) ) ;
OR2     gate2881  (.A(g2911), .B(g2917), .Z(g3414) ) ;
INV     gate2882  (.A(g3414), .Z(II7825) ) ;
INV     gate2883  (.A(II7825), .Z(g4462) ) ;
INV     gate2884  (.A(g3829), .Z(g4463) ) ;
OR2     gate2885  (.A(g2895), .B(g2910), .Z(g3425) ) ;
INV     gate2886  (.A(g3425), .Z(II7829) ) ;
INV     gate2887  (.A(II7829), .Z(g4464) ) ;
NAND2   gate2888  (.A(II6747), .B(II6748), .Z(g3585) ) ;
INV     gate2889  (.A(g3585), .Z(II7833) ) ;
INV     gate2890  (.A(II7833), .Z(g4466) ) ;
INV     gate2891  (.A(g3829), .Z(g4467) ) ;
INV     gate2892  (.A(g4158), .Z(II7837) ) ;
INV     gate2893  (.A(II7837), .Z(g4468) ) ;
OR2     gate2894  (.A(g2951), .B(g2957), .Z(g3431) ) ;
INV     gate2895  (.A(g3431), .Z(II7840) ) ;
INV     gate2896  (.A(II7840), .Z(g4469) ) ;
INV     gate2897  (.A(g3440), .Z(II7843) ) ;
INV     gate2898  (.A(II7843), .Z(g4470) ) ;
OR2     gate2899  (.A(g2945), .B(g2950), .Z(g3435) ) ;
INV     gate2900  (.A(g3435), .Z(II7847) ) ;
INV     gate2901  (.A(II7847), .Z(g4472) ) ;
INV     gate2902  (.A(g3820), .Z(g4474) ) ;
OR2     gate2903  (.A(g2939), .B(g2944), .Z(g3438) ) ;
INV     gate2904  (.A(g3438), .Z(II7852) ) ;
INV     gate2905  (.A(II7852), .Z(g4475) ) ;
INV     gate2906  (.A(g3820), .Z(g4478) ) ;
NAND2   gate2907  (.A(II6793), .B(II6794), .Z(g3631) ) ;
INV     gate2908  (.A(g3631), .Z(II7858) ) ;
INV     gate2909  (.A(II7858), .Z(g4479) ) ;
INV     gate2910  (.A(g3546), .Z(g4485) ) ;
INV     gate2911  (.A(g3546), .Z(g4491) ) ;
NOR2    gate2912  (.A(g1707), .B(g2864), .Z(g4076) ) ;
INV     gate2913  (.A(g4076), .Z(II7886) ) ;
INV     gate2914  (.A(II7886), .Z(g4495) ) ;
INV     gate2915  (.A(g3373), .Z(II7889) ) ;
INV     gate2916  (.A(II7889), .Z(g4496) ) ;
INV     gate2917  (.A(g3546), .Z(g4499) ) ;
INV     gate2918  (.A(g3946), .Z(g4501) ) ;
INV     gate2919  (.A(g3380), .Z(II7899) ) ;
INV     gate2920  (.A(II7899), .Z(g4504) ) ;
INV     gate2921  (.A(g3546), .Z(g4507) ) ;
INV     gate2922  (.A(g3946), .Z(g4508) ) ;
INV     gate2923  (.A(g3907), .Z(II7906) ) ;
INV     gate2924  (.A(II7906), .Z(g4509) ) ;
INV     gate2925  (.A(g3387), .Z(II7909) ) ;
INV     gate2926  (.A(II7909), .Z(g4510) ) ;
INV     gate2927  (.A(g3586), .Z(g4511) ) ;
INV     gate2928  (.A(g3546), .Z(g4513) ) ;
INV     gate2929  (.A(g3946), .Z(g4514) ) ;
INV     gate2930  (.A(g3664), .Z(II7916) ) ;
INV     gate2931  (.A(II7916), .Z(g4515) ) ;
INV     gate2932  (.A(g3440), .Z(II7920) ) ;
INV     gate2933  (.A(II7920), .Z(g4519) ) ;
INV     gate2934  (.A(g3394), .Z(II7923) ) ;
INV     gate2935  (.A(II7923), .Z(g4520) ) ;
INV     gate2936  (.A(g3586), .Z(g4521) ) ;
INV     gate2937  (.A(g3546), .Z(g4523) ) ;
INV     gate2938  (.A(g3946), .Z(g4524) ) ;
INV     gate2939  (.A(g3880), .Z(g4525) ) ;
INV     gate2940  (.A(g3624), .Z(II7931) ) ;
INV     gate2941  (.A(II7931), .Z(g4526) ) ;
INV     gate2942  (.A(g3440), .Z(II7935) ) ;
INV     gate2943  (.A(II7935), .Z(g4530) ) ;
INV     gate2944  (.A(g3406), .Z(II7938) ) ;
INV     gate2945  (.A(II7938), .Z(g4533) ) ;
INV     gate2946  (.A(g3946), .Z(g4535) ) ;
INV     gate2947  (.A(g3880), .Z(g4536) ) ;
INV     gate2948  (.A(g3417), .Z(II7946) ) ;
INV     gate2949  (.A(II7946), .Z(g4541) ) ;
INV     gate2950  (.A(g3946), .Z(g4543) ) ;
INV     gate2951  (.A(g3880), .Z(g4544) ) ;
INV     gate2952  (.A(g3664), .Z(II7952) ) ;
INV     gate2953  (.A(II7952), .Z(g4545) ) ;
INV     gate2954  (.A(g3428), .Z(II7956) ) ;
INV     gate2955  (.A(II7956), .Z(g4549) ) ;
INV     gate2956  (.A(g3946), .Z(g4551) ) ;
INV     gate2957  (.A(g3880), .Z(g4552) ) ;
INV     gate2958  (.A(g3433), .Z(II7964) ) ;
INV     gate2959  (.A(II7964), .Z(g4555) ) ;
INV     gate2960  (.A(g3946), .Z(g4557) ) ;
INV     gate2961  (.A(g3880), .Z(g4558) ) ;
INV     gate2962  (.A(g3437), .Z(II7973) ) ;
INV     gate2963  (.A(II7973), .Z(g4562) ) ;
INV     gate2964  (.A(g3946), .Z(g4563) ) ;
INV     gate2965  (.A(g3880), .Z(g4564) ) ;
NAND3   gate2966  (.A(g2382), .B(g2364), .C(g2800), .Z(g3753) ) ;
INV     gate2967  (.A(g3753), .Z(g4566) ) ;
AND2    gate2968  (.A(g1231), .B(g3047), .Z(g3374) ) ;
INV     gate2969  (.A(g3374), .Z(g4567) ) ;
INV     gate2970  (.A(g3880), .Z(g4575) ) ;
INV     gate2971  (.A(g3621), .Z(II7984) ) ;
INV     gate2972  (.A(II7984), .Z(g4577) ) ;
INV     gate2973  (.A(g3880), .Z(g4580) ) ;
INV     gate2974  (.A(g3880), .Z(g4583) ) ;
OR2     gate2975  (.A(g1959), .B(g3318), .Z(g4089) ) ;
INV     gate2976  (.A(g4089), .Z(g4586) ) ;
INV     gate2977  (.A(g3829), .Z(g4587) ) ;
NOR2    gate2978  (.A(g2187), .B(g2795), .Z(g3462) ) ;
INV     gate2979  (.A(g3462), .Z(II7996) ) ;
INV     gate2980  (.A(II7996), .Z(g4589) ) ;
AND2    gate2981  (.A(g1351), .B(g3301), .Z(g4114) ) ;
INV     gate2982  (.A(g4114), .Z(II7999) ) ;
INV     gate2983  (.A(II7999), .Z(g4590) ) ;
INV     gate2984  (.A(g3829), .Z(g4591) ) ;
INV     gate2985  (.A(g3829), .Z(g4592) ) ;
INV     gate2986  (.A(g3967), .Z(II8004) ) ;
INV     gate2987  (.A(II8004), .Z(g4593) ) ;
INV     gate2988  (.A(g3829), .Z(II8007) ) ;
INV     gate2989  (.A(II8007), .Z(g4596) ) ;
INV     gate2990  (.A(g3820), .Z(II8011) ) ;
INV     gate2991  (.A(II8011), .Z(g4602) ) ;
INV     gate2992  (.A(g3829), .Z(g4603) ) ;
INV     gate2993  (.A(g3829), .Z(g4606) ) ;
INV     gate2994  (.A(g3829), .Z(g4608) ) ;
INV     gate2995  (.A(g3829), .Z(g4614) ) ;
NAND2   gate2996  (.A(g3041), .B(g3061), .Z(g4117) ) ;
INV     gate2997  (.A(g4117), .Z(II8024) ) ;
INV     gate2998  (.A(II8024), .Z(g4615) ) ;
INV     gate2999  (.A(g3829), .Z(g4618) ) ;
INV     gate3000  (.A(g3540), .Z(II8031) ) ;
INV     gate3001  (.A(II8031), .Z(g4620) ) ;
INV     gate3002  (.A(g3820), .Z(g4631) ) ;
INV     gate3003  (.A(g3820), .Z(II8036) ) ;
INV     gate3004  (.A(II8036), .Z(g4636) ) ;
AND2    gate3005  (.A(g986), .B(g2760), .Z(g3506) ) ;
INV     gate3006  (.A(g3506), .Z(II8039) ) ;
INV     gate3007  (.A(II8039), .Z(g4637) ) ;
OR2     gate3008  (.A(g2920), .B(g2124), .Z(g3354) ) ;
INV     gate3009  (.A(g3354), .Z(g4638) ) ;
INV     gate3010  (.A(g4013), .Z(g4669) ) ;
INV     gate3011  (.A(g3354), .Z(g4671) ) ;
INV     gate3012  (.A(g4013), .Z(g4673) ) ;
INV     gate3013  (.A(g4089), .Z(II8050) ) ;
INV     gate3014  (.A(II8050), .Z(g4674) ) ;
INV     gate3015  (.A(g3354), .Z(g4676) ) ;
INV     gate3016  (.A(g3546), .Z(g4678) ) ;
INV     gate3017  (.A(g4013), .Z(g4679) ) ;
INV     gate3018  (.A(g3829), .Z(g4680) ) ;
INV     gate3019  (.A(g3546), .Z(g4681) ) ;
AND2    gate3020  (.A(g940), .B(g2756), .Z(g3381) ) ;
INV     gate3021  (.A(g3381), .Z(II8061) ) ;
INV     gate3022  (.A(II8061), .Z(g4711) ) ;
INV     gate3023  (.A(g3546), .Z(g4713) ) ;
INV     gate3024  (.A(g3546), .Z(g4716) ) ;
INV     gate3025  (.A(g3829), .Z(g4717) ) ;
INV     gate3026  (.A(g3586), .Z(g4719) ) ;
INV     gate3027  (.A(g3546), .Z(g4721) ) ;
INV     gate3028  (.A(g3586), .Z(g4724) ) ;
INV     gate3029  (.A(g3546), .Z(g4726) ) ;
INV     gate3030  (.A(g3538), .Z(II8080) ) ;
INV     gate3031  (.A(II8080), .Z(g4728) ) ;
INV     gate3032  (.A(g3586), .Z(g4729) ) ;
INV     gate3033  (.A(g3546), .Z(g4730) ) ;
INV     gate3034  (.A(g3664), .Z(II8085) ) ;
INV     gate3035  (.A(II8085), .Z(g4731) ) ;
INV     gate3036  (.A(g3545), .Z(II8089) ) ;
INV     gate3037  (.A(II8089), .Z(g4733) ) ;
INV     gate3038  (.A(g3586), .Z(g4734) ) ;
INV     gate3039  (.A(g3546), .Z(g4735) ) ;
INV     gate3040  (.A(g3440), .Z(g4737) ) ;
INV     gate3041  (.A(g3440), .Z(g4738) ) ;
INV     gate3042  (.A(g4117), .Z(g4739) ) ;
INV     gate3043  (.A(g3583), .Z(II8098) ) ;
INV     gate3044  (.A(II8098), .Z(g4746) ) ;
INV     gate3045  (.A(g3586), .Z(g4747) ) ;
INV     gate3046  (.A(g3546), .Z(g4748) ) ;
INV     gate3047  (.A(g3440), .Z(g4754) ) ;
INV     gate3048  (.A(g3440), .Z(g4755) ) ;
INV     gate3049  (.A(g3440), .Z(g4756) ) ;
INV     gate3050  (.A(g3622), .Z(II8109) ) ;
INV     gate3051  (.A(II8109), .Z(g4757) ) ;
INV     gate3052  (.A(g3586), .Z(g4758) ) ;
INV     gate3053  (.A(g3440), .Z(g4761) ) ;
INV     gate3054  (.A(g3627), .Z(II8116) ) ;
INV     gate3055  (.A(II8116), .Z(g4762) ) ;
INV     gate3056  (.A(g3586), .Z(g4763) ) ;
INV     gate3057  (.A(g3440), .Z(g4766) ) ;
INV     gate3058  (.A(g3630), .Z(II8123) ) ;
INV     gate3059  (.A(II8123), .Z(g4767) ) ;
NAND2   gate3060  (.A(II6826), .B(II6827), .Z(g3662) ) ;
INV     gate3061  (.A(g3662), .Z(II8126) ) ;
INV     gate3062  (.A(II8126), .Z(g4768) ) ;
INV     gate3063  (.A(g3586), .Z(g4769) ) ;
INV     gate3064  (.A(g3440), .Z(g4772) ) ;
INV     gate3065  (.A(g3632), .Z(II8133) ) ;
INV     gate3066  (.A(II8133), .Z(g4773) ) ;
INV     gate3067  (.A(g4144), .Z(II8136) ) ;
INV     gate3068  (.A(II8136), .Z(g4774) ) ;
NAND2   gate3069  (.A(II6837), .B(II6838), .Z(g3681) ) ;
INV     gate3070  (.A(g3681), .Z(II8139) ) ;
INV     gate3071  (.A(II8139), .Z(g4775) ) ;
INV     gate3072  (.A(g3586), .Z(g4776) ) ;
NAND3   gate3073  (.A(g2571), .B(g2550), .C(g2990), .Z(g3992) ) ;
INV     gate3074  (.A(g3992), .Z(g4777) ) ;
INV     gate3075  (.A(g3440), .Z(g4780) ) ;
INV     gate3076  (.A(g3633), .Z(II8147) ) ;
INV     gate3077  (.A(II8147), .Z(g4781) ) ;
INV     gate3078  (.A(g4089), .Z(g4782) ) ;
INV     gate3079  (.A(g3829), .Z(g4783) ) ;
INV     gate3080  (.A(g3337), .Z(g4785) ) ;
INV     gate3081  (.A(g3636), .Z(II8154) ) ;
INV     gate3082  (.A(II8154), .Z(g4786) ) ;
AND2    gate3083  (.A(II6630), .B(II6631), .Z(g3423) ) ;
INV     gate3084  (.A(g3423), .Z(g4787) ) ;
INV     gate3085  (.A(g3337), .Z(g4789) ) ;
INV     gate3086  (.A(g3337), .Z(g4790) ) ;
INV     gate3087  (.A(g3637), .Z(II8161) ) ;
INV     gate3088  (.A(II8161), .Z(g4791) ) ;
INV     gate3089  (.A(g3566), .Z(II8164) ) ;
INV     gate3090  (.A(II8164), .Z(g4794) ) ;
INV     gate3091  (.A(g3337), .Z(g4802) ) ;
INV     gate3092  (.A(g3337), .Z(g4805) ) ;
AND2    gate3093  (.A(g382), .B(g3257), .Z(g3661) ) ;
INV     gate3094  (.A(g3661), .Z(g4811) ) ;
INV     gate3095  (.A(g3354), .Z(g4819) ) ;
AND2    gate3096  (.A(g471), .B(g3268), .Z(g3706) ) ;
INV     gate3097  (.A(g3706), .Z(g4822) ) ;
INV     gate3098  (.A(g3566), .Z(II8192) ) ;
INV     gate3099  (.A(II8192), .Z(g4835) ) ;
INV     gate3100  (.A(g4013), .Z(II8199) ) ;
INV     gate3101  (.A(II8199), .Z(g4840) ) ;
INV     gate3102  (.A(g3976), .Z(II8204) ) ;
INV     gate3103  (.A(II8204), .Z(g4867) ) ;
INV     gate3104  (.A(g3566), .Z(II8211) ) ;
INV     gate3105  (.A(II8211), .Z(g4872) ) ;
INV     gate3106  (.A(g3981), .Z(II8215) ) ;
INV     gate3107  (.A(II8215), .Z(g4874) ) ;
INV     gate3108  (.A(g3638), .Z(g4880) ) ;
INV     gate3109  (.A(g4468), .Z(II8228) ) ;
INV     gate3110  (.A(g4170), .Z(II8231) ) ;
INV     gate3111  (.A(II8231), .Z(g4886) ) ;
INV     gate3112  (.A(g4232), .Z(II8234) ) ;
INV     gate3113  (.A(g4295), .Z(II8237) ) ;
INV     gate3114  (.A(g4380), .Z(II8240) ) ;
INV     gate3115  (.A(II8240), .Z(g4889) ) ;
INV     gate3116  (.A(g4615), .Z(II8247) ) ;
INV     gate3117  (.A(g4589), .Z(II8250) ) ;
INV     gate3118  (.A(g4637), .Z(II8253) ) ;
INV     gate3119  (.A(g4711), .Z(II8256) ) ;
INV     gate3120  (.A(g4590), .Z(II8259) ) ;
INV     gate3121  (.A(g4636), .Z(II8262) ) ;
INV     gate3122  (.A(g4602), .Z(II8265) ) ;
INV     gate3123  (.A(g4674), .Z(II8268) ) ;
INV     gate3124  (.A(g4351), .Z(II8275) ) ;
INV     gate3125  (.A(g4495), .Z(II8278) ) ;
INV     gate3126  (.A(g4396), .Z(g4908) ) ;
AND2    gate3127  (.A(g416), .B(g3415), .Z(g4770) ) ;
INV     gate3128  (.A(g4770), .Z(II8282) ) ;
INV     gate3129  (.A(II8282), .Z(g4912) ) ;
AND2    gate3130  (.A(g496), .B(g3416), .Z(g4771) ) ;
INV     gate3131  (.A(g4771), .Z(II8285) ) ;
INV     gate3132  (.A(II8285), .Z(g4913) ) ;
INV     gate3133  (.A(g4413), .Z(g4915) ) ;
AND2    gate3134  (.A(g421), .B(g3426), .Z(g4778) ) ;
INV     gate3135  (.A(g4778), .Z(II8290) ) ;
INV     gate3136  (.A(II8290), .Z(g4919) ) ;
AND2    gate3137  (.A(g501), .B(g3427), .Z(g4779) ) ;
INV     gate3138  (.A(g4779), .Z(II8293) ) ;
INV     gate3139  (.A(II8293), .Z(g4920) ) ;
INV     gate3140  (.A(g4437), .Z(II8298) ) ;
INV     gate3141  (.A(II8298), .Z(g4933) ) ;
INV     gate3142  (.A(g4243), .Z(g4934) ) ;
INV     gate3143  (.A(g4420), .Z(g4935) ) ;
AND2    gate3144  (.A(g506), .B(g3432), .Z(g4784) ) ;
INV     gate3145  (.A(g4784), .Z(II8303) ) ;
INV     gate3146  (.A(II8303), .Z(g4939) ) ;
INV     gate3147  (.A(g4443), .Z(II8308) ) ;
INV     gate3148  (.A(II8308), .Z(g4942) ) ;
INV     gate3149  (.A(g4794), .Z(II8311) ) ;
INV     gate3150  (.A(II8311), .Z(g4943) ) ;
INV     gate3151  (.A(g4430), .Z(g4944) ) ;
AND2    gate3152  (.A(g511), .B(g3436), .Z(g4788) ) ;
INV     gate3153  (.A(g4788), .Z(II8315) ) ;
INV     gate3154  (.A(II8315), .Z(g4948) ) ;
INV     gate3155  (.A(g4452), .Z(II8320) ) ;
INV     gate3156  (.A(II8320), .Z(g4951) ) ;
INV     gate3157  (.A(g4794), .Z(II8324) ) ;
INV     gate3158  (.A(II8324), .Z(g4953) ) ;
INV     gate3159  (.A(g4509), .Z(g4954) ) ;
AND2    gate3160  (.A(g516), .B(g3439), .Z(g4801) ) ;
INV     gate3161  (.A(g4801), .Z(II8328) ) ;
INV     gate3162  (.A(II8328), .Z(g4958) ) ;
INV     gate3163  (.A(g4456), .Z(II8333) ) ;
INV     gate3164  (.A(II8333), .Z(g4961) ) ;
INV     gate3165  (.A(g4352), .Z(II8337) ) ;
INV     gate3166  (.A(II8337), .Z(g4963) ) ;
AND2    gate3167  (.A(g476), .B(g3458), .Z(g4804) ) ;
INV     gate3168  (.A(g4804), .Z(II8340) ) ;
INV     gate3169  (.A(II8340), .Z(g4966) ) ;
INV     gate3170  (.A(g4411), .Z(g4970) ) ;
INV     gate3171  (.A(g4794), .Z(II8351) ) ;
INV     gate3172  (.A(II8351), .Z(g4975) ) ;
INV     gate3173  (.A(g4794), .Z(II8358) ) ;
INV     gate3174  (.A(II8358), .Z(g4988) ) ;
OR2     gate3175  (.A(g3991), .B(g3998), .Z(g4231) ) ;
INV     gate3176  (.A(g4231), .Z(II8379) ) ;
INV     gate3177  (.A(II8379), .Z(g5007) ) ;
OR2     gate3178  (.A(g3999), .B(g4007), .Z(g4238) ) ;
INV     gate3179  (.A(g4238), .Z(II8385) ) ;
INV     gate3180  (.A(II8385), .Z(g5011) ) ;
OR2     gate3181  (.A(g4000), .B(g4008), .Z(g4239) ) ;
INV     gate3182  (.A(g4239), .Z(II8388) ) ;
INV     gate3183  (.A(II8388), .Z(g5012) ) ;
OR2     gate3184  (.A(g4009), .B(g4047), .Z(g4255) ) ;
INV     gate3185  (.A(g4255), .Z(II8396) ) ;
INV     gate3186  (.A(II8396), .Z(g5027) ) ;
OR2     gate3187  (.A(g4048), .B(g4053), .Z(g4264) ) ;
INV     gate3188  (.A(g4264), .Z(II8403) ) ;
INV     gate3189  (.A(II8403), .Z(g5032) ) ;
OR2     gate3190  (.A(g4054), .B(g4058), .Z(g4274) ) ;
INV     gate3191  (.A(g4274), .Z(II8406) ) ;
INV     gate3192  (.A(II8406), .Z(g5033) ) ;
OR2     gate3193  (.A(g4059), .B(g4063), .Z(g4283) ) ;
INV     gate3194  (.A(g4283), .Z(II8410) ) ;
INV     gate3195  (.A(II8410), .Z(g5035) ) ;
OR2     gate3196  (.A(g4064), .B(g4068), .Z(g4293) ) ;
INV     gate3197  (.A(g4293), .Z(II8414) ) ;
INV     gate3198  (.A(II8414), .Z(g5037) ) ;
INV     gate3199  (.A(g4794), .Z(II8418) ) ;
INV     gate3200  (.A(II8418), .Z(g5039) ) ;
OR2     gate3201  (.A(g4069), .B(g4079), .Z(g4309) ) ;
INV     gate3202  (.A(g4309), .Z(II8421) ) ;
INV     gate3203  (.A(II8421), .Z(g5040) ) ;
INV     gate3204  (.A(g4840), .Z(g5042) ) ;
INV     gate3205  (.A(g4840), .Z(g5043) ) ;
INV     gate3206  (.A(g4354), .Z(g5047) ) ;
INV     gate3207  (.A(g4458), .Z(II8429) ) ;
INV     gate3208  (.A(II8429), .Z(g5050) ) ;
INV     gate3209  (.A(g4394), .Z(g5052) ) ;
INV     gate3210  (.A(g4840), .Z(g5062) ) ;
INV     gate3211  (.A(g4363), .Z(g5063) ) ;
INV     gate3212  (.A(g4462), .Z(II8436) ) ;
INV     gate3213  (.A(II8436), .Z(g5066) ) ;
INV     gate3214  (.A(g4840), .Z(g5068) ) ;
INV     gate3215  (.A(g4368), .Z(g5069) ) ;
INV     gate3216  (.A(g4464), .Z(II8442) ) ;
INV     gate3217  (.A(II8442), .Z(g5072) ) ;
INV     gate3218  (.A(g4840), .Z(g5073) ) ;
INV     gate3219  (.A(g4439), .Z(g5075) ) ;
INV     gate3220  (.A(g4372), .Z(g5078) ) ;
INV     gate3221  (.A(g4469), .Z(II8449) ) ;
INV     gate3222  (.A(II8449), .Z(g5081) ) ;
INV     gate3223  (.A(g4840), .Z(g5082) ) ;
INV     gate3224  (.A(g4377), .Z(g5085) ) ;
INV     gate3225  (.A(g4472), .Z(II8456) ) ;
INV     gate3226  (.A(II8456), .Z(g5088) ) ;
INV     gate3227  (.A(g4840), .Z(g5089) ) ;
INV     gate3228  (.A(g4385), .Z(g5091) ) ;
INV     gate3229  (.A(g4475), .Z(II8462) ) ;
INV     gate3230  (.A(II8462), .Z(g5094) ) ;
AND3    gate3231  (.A(g3015), .B(g1289), .C(g3937), .Z(g4807) ) ;
INV     gate3232  (.A(g4807), .Z(II8465) ) ;
INV     gate3233  (.A(II8465), .Z(g5095) ) ;
INV     gate3234  (.A(g4840), .Z(g5096) ) ;
INV     gate3235  (.A(g4840), .Z(g5098) ) ;
INV     gate3236  (.A(g4577), .Z(II8473) ) ;
INV     gate3237  (.A(g4577), .Z(II8476) ) ;
INV     gate3238  (.A(II8476), .Z(g5102) ) ;
INV     gate3239  (.A(g4526), .Z(II8487) ) ;
INV     gate3240  (.A(g4526), .Z(II8490) ) ;
INV     gate3241  (.A(II8490), .Z(g5106) ) ;
INV     gate3242  (.A(g4459), .Z(g5107) ) ;
AND2    gate3243  (.A(g1166), .B(g3682), .Z(g4325) ) ;
INV     gate3244  (.A(g4325), .Z(II8495) ) ;
INV     gate3245  (.A(II8495), .Z(g5109) ) ;
AND2    gate3246  (.A(g1163), .B(g3693), .Z(g4330) ) ;
INV     gate3247  (.A(g4330), .Z(II8499) ) ;
INV     gate3248  (.A(II8499), .Z(g5111) ) ;
OR3     gate3249  (.A(g3563), .B(g3348), .C(g1570), .Z(g4682) ) ;
INV     gate3250  (.A(g4682), .Z(g5112) ) ;
INV     gate3251  (.A(g4445), .Z(II8503) ) ;
INV     gate3252  (.A(II8503), .Z(g5113) ) ;
AND2    gate3253  (.A(g1160), .B(g3703), .Z(g4334) ) ;
INV     gate3254  (.A(g4334), .Z(II8506) ) ;
INV     gate3255  (.A(II8506), .Z(g5114) ) ;
INV     gate3256  (.A(g4682), .Z(g5116) ) ;
INV     gate3257  (.A(g4682), .Z(g5117) ) ;
AND2    gate3258  (.A(g1157), .B(g3707), .Z(g4338) ) ;
INV     gate3259  (.A(g4338), .Z(II8520) ) ;
INV     gate3260  (.A(II8520), .Z(g5120) ) ;
INV     gate3261  (.A(g4682), .Z(g5121) ) ;
INV     gate3262  (.A(g4682), .Z(g5122) ) ;
INV     gate3263  (.A(g4596), .Z(g5124) ) ;
AND2    gate3264  (.A(g1153), .B(g3715), .Z(g4340) ) ;
INV     gate3265  (.A(g4340), .Z(II8535) ) ;
INV     gate3266  (.A(II8535), .Z(g5127) ) ;
INV     gate3267  (.A(g4682), .Z(g5143) ) ;
INV     gate3268  (.A(g4682), .Z(g5144) ) ;
INV     gate3269  (.A(g4596), .Z(g5146) ) ;
AND2    gate3270  (.A(g1149), .B(g3719), .Z(g4342) ) ;
INV     gate3271  (.A(g4342), .Z(II8551) ) ;
INV     gate3272  (.A(II8551), .Z(g5149) ) ;
INV     gate3273  (.A(g4682), .Z(g5166) ) ;
INV     gate3274  (.A(g4682), .Z(g5167) ) ;
INV     gate3275  (.A(g4596), .Z(g5169) ) ;
INV     gate3276  (.A(g4682), .Z(g5175) ) ;
INV     gate3277  (.A(g4682), .Z(g5176) ) ;
INV     gate3278  (.A(g4596), .Z(g5177) ) ;
OR3     gate3279  (.A(g3348), .B(g3563), .C(g1527), .Z(g4640) ) ;
INV     gate3280  (.A(g4640), .Z(g5183) ) ;
INV     gate3281  (.A(g4682), .Z(g5184) ) ;
INV     gate3282  (.A(g4682), .Z(g5185) ) ;
INV     gate3283  (.A(g4640), .Z(g5191) ) ;
INV     gate3284  (.A(g4640), .Z(g5192) ) ;
INV     gate3285  (.A(g4682), .Z(g5193) ) ;
INV     gate3286  (.A(g4453), .Z(g5195) ) ;
INV     gate3287  (.A(g4562), .Z(II8611) ) ;
INV     gate3288  (.A(II8611), .Z(g5197) ) ;
INV     gate3289  (.A(g4414), .Z(II8614) ) ;
INV     gate3290  (.A(II8614), .Z(g5198) ) ;
INV     gate3291  (.A(g4567), .Z(g5200) ) ;
INV     gate3292  (.A(g4640), .Z(g5202) ) ;
INV     gate3293  (.A(g4640), .Z(g5203) ) ;
INV     gate3294  (.A(g4366), .Z(g5205) ) ;
INV     gate3295  (.A(g4425), .Z(II8631) ) ;
INV     gate3296  (.A(II8631), .Z(g5210) ) ;
INV     gate3297  (.A(g4640), .Z(g5213) ) ;
INV     gate3298  (.A(g4640), .Z(g5214) ) ;
INV     gate3299  (.A(g4445), .Z(g5216) ) ;
INV     gate3300  (.A(g4219), .Z(II8647) ) ;
INV     gate3301  (.A(II8647), .Z(g5218) ) ;
INV     gate3302  (.A(g4640), .Z(g5222) ) ;
INV     gate3303  (.A(g4640), .Z(g5223) ) ;
INV     gate3304  (.A(g4640), .Z(g5231) ) ;
INV     gate3305  (.A(g4640), .Z(g5232) ) ;
INV     gate3306  (.A(g4361), .Z(g5236) ) ;
INV     gate3307  (.A(g4386), .Z(g5241) ) ;
INV     gate3308  (.A(g4369), .Z(g5245) ) ;
INV     gate3309  (.A(g4640), .Z(g5251) ) ;
INV     gate3310  (.A(g4640), .Z(g5252) ) ;
INV     gate3311  (.A(g4346), .Z(g5253) ) ;
INV     gate3312  (.A(g4640), .Z(g5261) ) ;
INV     gate3313  (.A(g4353), .Z(g5262) ) ;
INV     gate3314  (.A(g4362), .Z(g5265) ) ;
INV     gate3315  (.A(g4530), .Z(II8711) ) ;
INV     gate3316  (.A(II8711), .Z(g5267) ) ;
INV     gate3317  (.A(g4367), .Z(g5270) ) ;
INV     gate3318  (.A(g4791), .Z(II8724) ) ;
INV     gate3319  (.A(II8724), .Z(g5272) ) ;
INV     gate3320  (.A(g4371), .Z(g5275) ) ;
INV     gate3321  (.A(g4428), .Z(g5281) ) ;
INV     gate3322  (.A(g4376), .Z(g5284) ) ;
INV     gate3323  (.A(g4355), .Z(g5285) ) ;
INV     gate3324  (.A(g4438), .Z(g5288) ) ;
INV     gate3325  (.A(g4384), .Z(g5291) ) ;
INV     gate3326  (.A(g4445), .Z(g5292) ) ;
INV     gate3327  (.A(g4444), .Z(g5296) ) ;
INV     gate3328  (.A(g4393), .Z(g5299) ) ;
INV     gate3329  (.A(g4373), .Z(g5301) ) ;
INV     gate3330  (.A(g4378), .Z(g5305) ) ;
INV     gate3331  (.A(g4387), .Z(g5314) ) ;
INV     gate3332  (.A(g4418), .Z(g5320) ) ;
AND2    gate3333  (.A(g1117), .B(g3828), .Z(g4465) ) ;
INV     gate3334  (.A(g4465), .Z(II8811) ) ;
INV     gate3335  (.A(II8811), .Z(g5344) ) ;
AND2    gate3336  (.A(g1121), .B(g3862), .Z(g4471) ) ;
INV     gate3337  (.A(g4471), .Z(II8815) ) ;
INV     gate3338  (.A(II8815), .Z(g5348) ) ;
AND2    gate3339  (.A(g1125), .B(g3874), .Z(g4473) ) ;
INV     gate3340  (.A(g4473), .Z(II8820) ) ;
INV     gate3341  (.A(II8820), .Z(g5353) ) ;
AND2    gate3342  (.A(g1129), .B(g3878), .Z(g4477) ) ;
INV     gate3343  (.A(g4477), .Z(II8827) ) ;
INV     gate3344  (.A(II8827), .Z(g5391) ) ;
AND2    gate3345  (.A(g1133), .B(g3905), .Z(g4480) ) ;
INV     gate3346  (.A(g4480), .Z(II8831) ) ;
INV     gate3347  (.A(II8831), .Z(g5395) ) ;
INV     gate3348  (.A(g4791), .Z(II8835) ) ;
INV     gate3349  (.A(II8835), .Z(g5397) ) ;
AND2    gate3350  (.A(g1137), .B(g3909), .Z(g4484) ) ;
INV     gate3351  (.A(g4484), .Z(II8839) ) ;
INV     gate3352  (.A(II8839), .Z(g5401) ) ;
OR2     gate3353  (.A(g3536), .B(g2916), .Z(g4556) ) ;
INV     gate3354  (.A(g4556), .Z(II8842) ) ;
INV     gate3355  (.A(II8842), .Z(g5402) ) ;
AND2    gate3356  (.A(g1141), .B(g3913), .Z(g4490) ) ;
INV     gate3357  (.A(g4490), .Z(II8848) ) ;
INV     gate3358  (.A(II8848), .Z(g5415) ) ;
AND2    gate3359  (.A(g1145), .B(g3940), .Z(g4498) ) ;
INV     gate3360  (.A(g4498), .Z(II8851) ) ;
INV     gate3361  (.A(II8851), .Z(g5416) ) ;
AND2    gate3362  (.A(g1357), .B(g3941), .Z(g4500) ) ;
INV     gate3363  (.A(g4500), .Z(II8854) ) ;
INV     gate3364  (.A(II8854), .Z(g5417) ) ;
AND2    gate3365  (.A(g1113), .B(g3944), .Z(g4506) ) ;
INV     gate3366  (.A(g4506), .Z(II8858) ) ;
INV     gate3367  (.A(II8858), .Z(g5419) ) ;
OR2     gate3368  (.A(g3546), .B(g2391), .Z(g4300) ) ;
INV     gate3369  (.A(g4300), .Z(g5420) ) ;
INV     gate3370  (.A(g4470), .Z(g5422) ) ;
INV     gate3371  (.A(g4300), .Z(g5423) ) ;
AND2    gate3372  (.A(g452), .B(g3975), .Z(g4518) ) ;
INV     gate3373  (.A(g4518), .Z(II8865) ) ;
INV     gate3374  (.A(II8865), .Z(g5424) ) ;
INV     gate3375  (.A(g4300), .Z(g5425) ) ;
AND2    gate3376  (.A(g4112), .B(g2980), .Z(g4421) ) ;
INV     gate3377  (.A(g4421), .Z(II8869) ) ;
INV     gate3378  (.A(II8869), .Z(g5426) ) ;
AND2    gate3379  (.A(g448), .B(g3980), .Z(g4529) ) ;
INV     gate3380  (.A(g4529), .Z(II8872) ) ;
INV     gate3381  (.A(II8872), .Z(g5443) ) ;
INV     gate3382  (.A(g4421), .Z(II8877) ) ;
INV     gate3383  (.A(II8877), .Z(g5446) ) ;
AND2    gate3384  (.A(g444), .B(g3988), .Z(g4537) ) ;
INV     gate3385  (.A(g4537), .Z(II8880) ) ;
INV     gate3386  (.A(II8880), .Z(g5469) ) ;
INV     gate3387  (.A(g4370), .Z(g5471) ) ;
AND2    gate3388  (.A(g440), .B(g3990), .Z(g4548) ) ;
INV     gate3389  (.A(g4548), .Z(II8885) ) ;
INV     gate3390  (.A(II8885), .Z(g5472) ) ;
AND2    gate3391  (.A(g435), .B(g3995), .Z(g4553) ) ;
INV     gate3392  (.A(g4553), .Z(II8889) ) ;
INV     gate3393  (.A(II8889), .Z(g5474) ) ;
AND2    gate3394  (.A(g542), .B(g3996), .Z(g4554) ) ;
INV     gate3395  (.A(g4554), .Z(II8892) ) ;
INV     gate3396  (.A(II8892), .Z(g5475) ) ;
AND2    gate3397  (.A(g431), .B(g4002), .Z(g4560) ) ;
INV     gate3398  (.A(g4560), .Z(II8900) ) ;
INV     gate3399  (.A(II8900), .Z(g5481) ) ;
AND2    gate3400  (.A(g538), .B(g4003), .Z(g4561) ) ;
INV     gate3401  (.A(g4561), .Z(II8903) ) ;
INV     gate3402  (.A(II8903), .Z(g5482) ) ;
INV     gate3403  (.A(g4395), .Z(g5486) ) ;
AND2    gate3404  (.A(g534), .B(g4010), .Z(g4565) ) ;
INV     gate3405  (.A(g4565), .Z(II8911) ) ;
INV     gate3406  (.A(II8911), .Z(g5490) ) ;
INV     gate3407  (.A(g4412), .Z(g5494) ) ;
AND2    gate3408  (.A(g530), .B(g4049), .Z(g4576) ) ;
INV     gate3409  (.A(g4576), .Z(II8919) ) ;
INV     gate3410  (.A(II8919), .Z(g5498) ) ;
INV     gate3411  (.A(g4515), .Z(g5503) ) ;
INV     gate3412  (.A(g4419), .Z(g5504) ) ;
AND2    gate3413  (.A(g525), .B(g4055), .Z(g4582) ) ;
INV     gate3414  (.A(g4582), .Z(II8929) ) ;
INV     gate3415  (.A(II8929), .Z(g5508) ) ;
INV     gate3416  (.A(g4739), .Z(g5509) ) ;
INV     gate3417  (.A(g4271), .Z(II8934) ) ;
INV     gate3418  (.A(II8934), .Z(g5511) ) ;
INV     gate3419  (.A(g4429), .Z(g5515) ) ;
INV     gate3420  (.A(g4811), .Z(g5519) ) ;
AND2    gate3421  (.A(g521), .B(g4060), .Z(g4585) ) ;
INV     gate3422  (.A(g4585), .Z(II8943) ) ;
INV     gate3423  (.A(II8943), .Z(g5520) ) ;
INV     gate3424  (.A(g4530), .Z(g5521) ) ;
INV     gate3425  (.A(g4545), .Z(g5534) ) ;
NAND2   gate3426  (.A(II7864), .B(II7865), .Z(g4482) ) ;
INV     gate3427  (.A(g4482), .Z(II8967) ) ;
INV     gate3428  (.A(II8967), .Z(g5542) ) ;
NAND2   gate3429  (.A(II7876), .B(II7877), .Z(g4488) ) ;
INV     gate3430  (.A(g4488), .Z(II8973) ) ;
INV     gate3431  (.A(II8973), .Z(g5546) ) ;
INV     gate3432  (.A(g4728), .Z(II8982) ) ;
INV     gate3433  (.A(II8982), .Z(g5567) ) ;
INV     gate3434  (.A(g4733), .Z(II8985) ) ;
INV     gate3435  (.A(II8985), .Z(g5568) ) ;
INV     gate3436  (.A(g4746), .Z(II8989) ) ;
INV     gate3437  (.A(II8989), .Z(g5572) ) ;
INV     gate3438  (.A(g4300), .Z(g5574) ) ;
INV     gate3439  (.A(g4757), .Z(II8996) ) ;
INV     gate3440  (.A(II8996), .Z(g5586) ) ;
INV     gate3441  (.A(g4762), .Z(II9001) ) ;
INV     gate3442  (.A(II9001), .Z(g5589) ) ;
INV     gate3443  (.A(g4767), .Z(II9013) ) ;
INV     gate3444  (.A(II9013), .Z(g5593) ) ;
AND2    gate3445  (.A(g426), .B(g3353), .Z(g4722) ) ;
INV     gate3446  (.A(g4722), .Z(II9016) ) ;
INV     gate3447  (.A(II9016), .Z(g5594) ) ;
INV     gate3448  (.A(g4773), .Z(II9020) ) ;
INV     gate3449  (.A(II9020), .Z(g5596) ) ;
AND2    gate3450  (.A(g386), .B(g3364), .Z(g4727) ) ;
INV     gate3451  (.A(g4727), .Z(II9023) ) ;
INV     gate3452  (.A(II9023), .Z(g5597) ) ;
INV     gate3453  (.A(g4781), .Z(II9029) ) ;
INV     gate3454  (.A(II9029), .Z(g5603) ) ;
AND2    gate3455  (.A(g391), .B(g3372), .Z(g4732) ) ;
INV     gate3456  (.A(g4732), .Z(II9032) ) ;
INV     gate3457  (.A(II9032), .Z(g5604) ) ;
INV     gate3458  (.A(g4840), .Z(g5613) ) ;
INV     gate3459  (.A(g4794), .Z(II9040) ) ;
INV     gate3460  (.A(II9040), .Z(g5614) ) ;
INV     gate3461  (.A(g4786), .Z(II9043) ) ;
INV     gate3462  (.A(II9043), .Z(g5615) ) ;
AND2    gate3463  (.A(g396), .B(g3379), .Z(g4736) ) ;
INV     gate3464  (.A(g4736), .Z(II9046) ) ;
INV     gate3465  (.A(II9046), .Z(g5616) ) ;
INV     gate3466  (.A(g4840), .Z(g5619) ) ;
INV     gate3467  (.A(g4417), .Z(g5620) ) ;
AND2    gate3468  (.A(g401), .B(g3385), .Z(g4752) ) ;
INV     gate3469  (.A(g4752), .Z(II9053) ) ;
INV     gate3470  (.A(II9053), .Z(g5623) ) ;
AND2    gate3471  (.A(g481), .B(g3386), .Z(g4753) ) ;
INV     gate3472  (.A(g4753), .Z(II9056) ) ;
INV     gate3473  (.A(II9056), .Z(g5624) ) ;
INV     gate3474  (.A(g4840), .Z(g5627) ) ;
AND2    gate3475  (.A(g406), .B(g3392), .Z(g4759) ) ;
INV     gate3476  (.A(g4759), .Z(II9062) ) ;
INV     gate3477  (.A(II9062), .Z(g5628) ) ;
AND2    gate3478  (.A(g486), .B(g3393), .Z(g4760) ) ;
INV     gate3479  (.A(g4760), .Z(II9065) ) ;
INV     gate3480  (.A(II9065), .Z(g5629) ) ;
INV     gate3481  (.A(g4768), .Z(II9068) ) ;
INV     gate3482  (.A(II9068), .Z(g5630) ) ;
INV     gate3483  (.A(g4388), .Z(g5633) ) ;
AND2    gate3484  (.A(g411), .B(g3404), .Z(g4764) ) ;
INV     gate3485  (.A(g4764), .Z(II9074) ) ;
INV     gate3486  (.A(II9074), .Z(g5637) ) ;
AND2    gate3487  (.A(g491), .B(g3405), .Z(g4765) ) ;
INV     gate3488  (.A(g4765), .Z(II9077) ) ;
INV     gate3489  (.A(II9077), .Z(g5638) ) ;
INV     gate3490  (.A(g4775), .Z(II9080) ) ;
INV     gate3491  (.A(II9080), .Z(g5639) ) ;
INV     gate3492  (.A(g4886), .Z(II9084) ) ;
INV     gate3493  (.A(II9084), .Z(g5641) ) ;
INV     gate3494  (.A(g5113), .Z(II9087) ) ;
INV     gate3495  (.A(g5567), .Z(II9090) ) ;
INV     gate3496  (.A(g5397), .Z(II9093) ) ;
INV     gate3497  (.A(g5568), .Z(II9096) ) ;
INV     gate3498  (.A(g5572), .Z(II9099) ) ;
INV     gate3499  (.A(g5586), .Z(II9102) ) ;
INV     gate3500  (.A(g5589), .Z(II9105) ) ;
INV     gate3501  (.A(g5593), .Z(II9108) ) ;
INV     gate3502  (.A(g5596), .Z(II9111) ) ;
INV     gate3503  (.A(g5603), .Z(II9114) ) ;
INV     gate3504  (.A(g5615), .Z(II9117) ) ;
INV     gate3505  (.A(g5218), .Z(II9120) ) ;
AND2    gate3506  (.A(g630), .B(g4739), .Z(g4890) ) ;
INV     gate3507  (.A(g4890), .Z(II9123) ) ;
AND2    gate3508  (.A(g631), .B(g4739), .Z(g4891) ) ;
INV     gate3509  (.A(g4891), .Z(II9126) ) ;
AND2    gate3510  (.A(g632), .B(g4739), .Z(g4892) ) ;
INV     gate3511  (.A(g4892), .Z(II9129) ) ;
AND2    gate3512  (.A(g635), .B(g4739), .Z(g4893) ) ;
INV     gate3513  (.A(g4893), .Z(II9132) ) ;
INV     gate3514  (.A(g5198), .Z(II9135) ) ;
INV     gate3515  (.A(g5210), .Z(II9138) ) ;
INV     gate3516  (.A(g5402), .Z(II9141) ) ;
INV     gate3517  (.A(g5007), .Z(II9144) ) ;
INV     gate3518  (.A(g5011), .Z(II9147) ) ;
INV     gate3519  (.A(g5012), .Z(II9150) ) ;
INV     gate3520  (.A(g5027), .Z(II9153) ) ;
INV     gate3521  (.A(g5032), .Z(II9156) ) ;
INV     gate3522  (.A(g5033), .Z(II9159) ) ;
INV     gate3523  (.A(g5035), .Z(II9162) ) ;
INV     gate3524  (.A(g5037), .Z(II9165) ) ;
INV     gate3525  (.A(g5040), .Z(II9168) ) ;
AND2    gate3526  (.A(g1848), .B(g4243), .Z(g4902) ) ;
INV     gate3527  (.A(g4902), .Z(II9171) ) ;
AND2    gate3528  (.A(g1849), .B(g4243), .Z(g4903) ) ;
INV     gate3529  (.A(g4903), .Z(II9174) ) ;
AND2    gate3530  (.A(g1850), .B(g4243), .Z(g4904) ) ;
INV     gate3531  (.A(g4904), .Z(II9177) ) ;
AND2    gate3532  (.A(g1853), .B(g4243), .Z(g4905) ) ;
INV     gate3533  (.A(g4905), .Z(II9180) ) ;
INV     gate3534  (.A(g4915), .Z(II9185) ) ;
INV     gate3535  (.A(II9185), .Z(g5676) ) ;
INV     gate3536  (.A(g4908), .Z(II9188) ) ;
INV     gate3537  (.A(II9188), .Z(g5677) ) ;
INV     gate3538  (.A(g5546), .Z(II9191) ) ;
INV     gate3539  (.A(II9191), .Z(g5678) ) ;
INV     gate3540  (.A(g5236), .Z(II9194) ) ;
INV     gate3541  (.A(II9194), .Z(g5679) ) ;
INV     gate3542  (.A(g4935), .Z(II9199) ) ;
INV     gate3543  (.A(II9199), .Z(g5682) ) ;
INV     gate3544  (.A(g4915), .Z(II9202) ) ;
INV     gate3545  (.A(II9202), .Z(g5683) ) ;
OR2     gate3546  (.A(g3664), .B(g4401), .Z(g5309) ) ;
INV     gate3547  (.A(g5309), .Z(II9205) ) ;
INV     gate3548  (.A(II9205), .Z(g5684) ) ;
INV     gate3549  (.A(g5047), .Z(II9208) ) ;
INV     gate3550  (.A(II9208), .Z(g5685) ) ;
INV     gate3551  (.A(g4944), .Z(II9213) ) ;
INV     gate3552  (.A(II9213), .Z(g5688) ) ;
INV     gate3553  (.A(g4935), .Z(II9216) ) ;
INV     gate3554  (.A(II9216), .Z(g5689) ) ;
INV     gate3555  (.A(g5236), .Z(g5691) ) ;
INV     gate3556  (.A(g5236), .Z(II9221) ) ;
INV     gate3557  (.A(II9221), .Z(g5692) ) ;
INV     gate3558  (.A(g5063), .Z(II9224) ) ;
INV     gate3559  (.A(II9224), .Z(g5693) ) ;
INV     gate3560  (.A(g4954), .Z(II9229) ) ;
INV     gate3561  (.A(II9229), .Z(g5696) ) ;
INV     gate3562  (.A(g4944), .Z(II9232) ) ;
INV     gate3563  (.A(II9232), .Z(g5697) ) ;
INV     gate3564  (.A(g5205), .Z(II9237) ) ;
INV     gate3565  (.A(II9237), .Z(g5700) ) ;
INV     gate3566  (.A(g5069), .Z(II9240) ) ;
INV     gate3567  (.A(II9240), .Z(g5701) ) ;
INV     gate3568  (.A(g5245), .Z(II9243) ) ;
INV     gate3569  (.A(II9243), .Z(g5702) ) ;
INV     gate3570  (.A(g4954), .Z(II9248) ) ;
INV     gate3571  (.A(II9248), .Z(g5705) ) ;
INV     gate3572  (.A(g5052), .Z(II9253) ) ;
INV     gate3573  (.A(II9253), .Z(g5708) ) ;
INV     gate3574  (.A(g5078), .Z(II9256) ) ;
INV     gate3575  (.A(II9256), .Z(g5718) ) ;
INV     gate3576  (.A(g5301), .Z(II9259) ) ;
INV     gate3577  (.A(II9259), .Z(g5719) ) ;
INV     gate3578  (.A(g5085), .Z(II9265) ) ;
INV     gate3579  (.A(II9265), .Z(g5723) ) ;
INV     gate3580  (.A(g5305), .Z(II9268) ) ;
INV     gate3581  (.A(II9268), .Z(g5724) ) ;
INV     gate3582  (.A(g5091), .Z(II9273) ) ;
INV     gate3583  (.A(II9273), .Z(g5727) ) ;
INV     gate3584  (.A(g5241), .Z(II9276) ) ;
INV     gate3585  (.A(II9276), .Z(g5728) ) ;
INV     gate3586  (.A(g5314), .Z(II9279) ) ;
INV     gate3587  (.A(II9279), .Z(g5729) ) ;
INV     gate3588  (.A(g5633), .Z(II9282) ) ;
INV     gate3589  (.A(II9282), .Z(g5730) ) ;
OR2     gate3590  (.A(g4675), .B(g3664), .Z(g5576) ) ;
INV     gate3591  (.A(g5576), .Z(II9287) ) ;
INV     gate3592  (.A(II9287), .Z(g5733) ) ;
INV     gate3593  (.A(g5052), .Z(II9290) ) ;
INV     gate3594  (.A(II9290), .Z(g5734) ) ;
INV     gate3595  (.A(g5486), .Z(II9293) ) ;
INV     gate3596  (.A(II9293), .Z(g5735) ) ;
INV     gate3597  (.A(g4908), .Z(II9296) ) ;
INV     gate3598  (.A(II9296), .Z(g5736) ) ;
INV     gate3599  (.A(g5576), .Z(II9302) ) ;
INV     gate3600  (.A(II9302), .Z(g5740) ) ;
INV     gate3601  (.A(g4970), .Z(II9305) ) ;
INV     gate3602  (.A(II9305), .Z(g5741) ) ;
INV     gate3603  (.A(g5494), .Z(II9308) ) ;
INV     gate3604  (.A(II9308), .Z(g5742) ) ;
INV     gate3605  (.A(g4915), .Z(II9311) ) ;
INV     gate3606  (.A(II9311), .Z(g5743) ) ;
INV     gate3607  (.A(g5576), .Z(II9317) ) ;
INV     gate3608  (.A(II9317), .Z(g5747) ) ;
NAND3   gate3609  (.A(g4749), .B(g3247), .C(g3205), .Z(g5013) ) ;
INV     gate3610  (.A(g5013), .Z(II9320) ) ;
INV     gate3611  (.A(II9320), .Z(g5748) ) ;
INV     gate3612  (.A(g5620), .Z(II9323) ) ;
INV     gate3613  (.A(II9323), .Z(g5751) ) ;
INV     gate3614  (.A(g5320), .Z(II9326) ) ;
INV     gate3615  (.A(II9326), .Z(g5752) ) ;
INV     gate3616  (.A(g5504), .Z(II9329) ) ;
INV     gate3617  (.A(II9329), .Z(g5753) ) ;
INV     gate3618  (.A(g4935), .Z(II9332) ) ;
INV     gate3619  (.A(II9332), .Z(g5754) ) ;
INV     gate3620  (.A(g5576), .Z(II9338) ) ;
INV     gate3621  (.A(II9338), .Z(g5758) ) ;
INV     gate3622  (.A(g5013), .Z(II9341) ) ;
INV     gate3623  (.A(II9341), .Z(g5759) ) ;
INV     gate3624  (.A(g5281), .Z(II9346) ) ;
INV     gate3625  (.A(II9346), .Z(g5766) ) ;
INV     gate3626  (.A(g5515), .Z(II9349) ) ;
INV     gate3627  (.A(II9349), .Z(g5767) ) ;
INV     gate3628  (.A(g4944), .Z(II9352) ) ;
INV     gate3629  (.A(II9352), .Z(g5768) ) ;
INV     gate3630  (.A(g5576), .Z(II9359) ) ;
INV     gate3631  (.A(II9359), .Z(g5773) ) ;
INV     gate3632  (.A(g5013), .Z(II9362) ) ;
INV     gate3633  (.A(II9362), .Z(g5774) ) ;
NOR2    gate3634  (.A(g3369), .B(g4258), .Z(g5392) ) ;
INV     gate3635  (.A(g5392), .Z(II9365) ) ;
INV     gate3636  (.A(II9365), .Z(g5777) ) ;
INV     gate3637  (.A(g5288), .Z(II9368) ) ;
INV     gate3638  (.A(II9368), .Z(g5778) ) ;
INV     gate3639  (.A(g5075), .Z(II9371) ) ;
INV     gate3640  (.A(II9371), .Z(g5779) ) ;
INV     gate3641  (.A(g5576), .Z(II9377) ) ;
INV     gate3642  (.A(II9377), .Z(g5783) ) ;
INV     gate3643  (.A(g5013), .Z(II9380) ) ;
INV     gate3644  (.A(II9380), .Z(g5784) ) ;
INV     gate3645  (.A(g5296), .Z(II9383) ) ;
INV     gate3646  (.A(II9383), .Z(g5787) ) ;
INV     gate3647  (.A(g5576), .Z(II9388) ) ;
INV     gate3648  (.A(II9388), .Z(g5790) ) ;
INV     gate3649  (.A(g5013), .Z(II9391) ) ;
INV     gate3650  (.A(II9391), .Z(g5791) ) ;
INV     gate3651  (.A(g5195), .Z(II9394) ) ;
INV     gate3652  (.A(II9394), .Z(g5794) ) ;
INV     gate3653  (.A(g5013), .Z(II9399) ) ;
INV     gate3654  (.A(II9399), .Z(g5797) ) ;
INV     gate3655  (.A(g5107), .Z(II9402) ) ;
INV     gate3656  (.A(II9402), .Z(g5800) ) ;
INV     gate3657  (.A(g5320), .Z(g5801) ) ;
INV     gate3658  (.A(g5013), .Z(II9409) ) ;
INV     gate3659  (.A(II9409), .Z(g5805) ) ;
INV     gate3660  (.A(g5320), .Z(g5808) ) ;
INV     gate3661  (.A(g5047), .Z(II9415) ) ;
INV     gate3662  (.A(II9415), .Z(g5811) ) ;
INV     gate3663  (.A(g5320), .Z(g5812) ) ;
INV     gate3664  (.A(g5063), .Z(II9421) ) ;
INV     gate3665  (.A(II9421), .Z(g5815) ) ;
INV     gate3666  (.A(g4963), .Z(II9424) ) ;
INV     gate3667  (.A(g4963), .Z(II9427) ) ;
INV     gate3668  (.A(II9427), .Z(g5817) ) ;
INV     gate3669  (.A(g5320), .Z(g5818) ) ;
INV     gate3670  (.A(g5069), .Z(II9433) ) ;
INV     gate3671  (.A(II9433), .Z(g5821) ) ;
INV     gate3672  (.A(g5320), .Z(g5822) ) ;
INV     gate3673  (.A(g5078), .Z(II9440) ) ;
INV     gate3674  (.A(II9440), .Z(g5826) ) ;
NAND3   gate3675  (.A(g4538), .B(g3071), .C(g3011), .Z(g5557) ) ;
INV     gate3676  (.A(g5557), .Z(II9443) ) ;
INV     gate3677  (.A(II9443), .Z(g5827) ) ;
INV     gate3678  (.A(g5052), .Z(II9446) ) ;
INV     gate3679  (.A(II9446), .Z(g5830) ) ;
INV     gate3680  (.A(g5320), .Z(g5836) ) ;
INV     gate3681  (.A(g5085), .Z(II9452) ) ;
INV     gate3682  (.A(II9452), .Z(g5839) ) ;
INV     gate3683  (.A(g5320), .Z(g5840) ) ;
INV     gate3684  (.A(g5091), .Z(II9458) ) ;
INV     gate3685  (.A(II9458), .Z(g5843) ) ;
AND2    gate3686  (.A(g3500), .B(g4440), .Z(g4940) ) ;
INV     gate3687  (.A(g4940), .Z(II9461) ) ;
INV     gate3688  (.A(II9461), .Z(g5844) ) ;
INV     gate3689  (.A(g5320), .Z(g5845) ) ;
INV     gate3690  (.A(g5320), .Z(g5850) ) ;
INV     gate3691  (.A(g5245), .Z(g5856) ) ;
AND3    gate3692  (.A(g4631), .B(g3875), .C(g2733), .Z(g5445) ) ;
INV     gate3693  (.A(g5445), .Z(II9475) ) ;
INV     gate3694  (.A(II9475), .Z(g5858) ) ;
INV     gate3695  (.A(g4954), .Z(II9479) ) ;
INV     gate3696  (.A(II9479), .Z(g5862) ) ;
INV     gate3697  (.A(g5050), .Z(II9483) ) ;
INV     gate3698  (.A(II9483), .Z(g5864) ) ;
INV     gate3699  (.A(g5066), .Z(II9486) ) ;
INV     gate3700  (.A(II9486), .Z(g5865) ) ;
OR3     gate3701  (.A(g4316), .B(g4093), .C(g126), .Z(g5361) ) ;
INV     gate3702  (.A(g5361), .Z(g5866) ) ;
INV     gate3703  (.A(g5072), .Z(II9491) ) ;
INV     gate3704  (.A(II9491), .Z(g5874) ) ;
INV     gate3705  (.A(g5361), .Z(g5875) ) ;
INV     gate3706  (.A(g5361), .Z(g5876) ) ;
INV     gate3707  (.A(g5309), .Z(g5878) ) ;
INV     gate3708  (.A(g5081), .Z(II9498) ) ;
INV     gate3709  (.A(II9498), .Z(g5879) ) ;
INV     gate3710  (.A(g5361), .Z(g5880) ) ;
INV     gate3711  (.A(g5361), .Z(g5881) ) ;
INV     gate3712  (.A(g5309), .Z(g5883) ) ;
INV     gate3713  (.A(g5088), .Z(II9505) ) ;
INV     gate3714  (.A(II9505), .Z(g5884) ) ;
INV     gate3715  (.A(g5361), .Z(g5885) ) ;
INV     gate3716  (.A(g5361), .Z(g5886) ) ;
AND3    gate3717  (.A(g4631), .B(g2733), .C(g3819), .Z(g5421) ) ;
INV     gate3718  (.A(g5421), .Z(II9510) ) ;
INV     gate3719  (.A(II9510), .Z(g5887) ) ;
INV     gate3720  (.A(g5102), .Z(g5888) ) ;
INV     gate3721  (.A(g5094), .Z(II9514) ) ;
INV     gate3722  (.A(II9514), .Z(g5889) ) ;
INV     gate3723  (.A(g5361), .Z(g5890) ) ;
INV     gate3724  (.A(g5361), .Z(g5891) ) ;
AND2    gate3725  (.A(g1304), .B(g4485), .Z(g4998) ) ;
INV     gate3726  (.A(g4998), .Z(II9519) ) ;
INV     gate3727  (.A(II9519), .Z(g5892) ) ;
INV     gate3728  (.A(g5106), .Z(g5893) ) ;
INV     gate3729  (.A(g5361), .Z(g5894) ) ;
INV     gate3730  (.A(g5361), .Z(g5895) ) ;
AND2    gate3731  (.A(g1300), .B(g4491), .Z(g5001) ) ;
INV     gate3732  (.A(g5001), .Z(II9525) ) ;
INV     gate3733  (.A(II9525), .Z(g5896) ) ;
INV     gate3734  (.A(g5361), .Z(g5898) ) ;
INV     gate3735  (.A(g5361), .Z(g5899) ) ;
AND2    gate3736  (.A(g1296), .B(g4499), .Z(g5004) ) ;
INV     gate3737  (.A(g5004), .Z(II9531) ) ;
INV     gate3738  (.A(II9531), .Z(g5900) ) ;
INV     gate3739  (.A(g5361), .Z(g5901) ) ;
AND2    gate3740  (.A(g1292), .B(g4507), .Z(g5008) ) ;
INV     gate3741  (.A(g5008), .Z(II9536) ) ;
INV     gate3742  (.A(II9536), .Z(g5903) ) ;
AND2    gate3743  (.A(g2733), .B(g4460), .Z(g5354) ) ;
INV     gate3744  (.A(g5354), .Z(II9539) ) ;
INV     gate3745  (.A(II9539), .Z(g5904) ) ;
AND2    gate3746  (.A(g1284), .B(g4513), .Z(g5024) ) ;
INV     gate3747  (.A(g5024), .Z(II9544) ) ;
INV     gate3748  (.A(II9544), .Z(g5912) ) ;
AND2    gate3749  (.A(g1280), .B(g4523), .Z(g5030) ) ;
INV     gate3750  (.A(g5030), .Z(II9550) ) ;
INV     gate3751  (.A(II9550), .Z(g5916) ) ;
INV     gate3752  (.A(g5109), .Z(II9564) ) ;
INV     gate3753  (.A(II9564), .Z(g5936) ) ;
NOR4    gate3754  (.A(g4787), .B(g2695), .C(g2299), .D(g2031), .Z(g5556) ) ;
INV     gate3755  (.A(g5556), .Z(II9567) ) ;
INV     gate3756  (.A(II9567), .Z(g5937) ) ;
INV     gate3757  (.A(g5509), .Z(II9571) ) ;
INV     gate3758  (.A(II9571), .Z(g5941) ) ;
INV     gate3759  (.A(g5111), .Z(II9581) ) ;
INV     gate3760  (.A(II9581), .Z(g5943) ) ;
INV     gate3761  (.A(g5241), .Z(II9585) ) ;
INV     gate3762  (.A(II9585), .Z(g5947) ) ;
INV     gate3763  (.A(g5114), .Z(II9588) ) ;
INV     gate3764  (.A(II9588), .Z(g5948) ) ;
INV     gate3765  (.A(g5095), .Z(II9591) ) ;
INV     gate3766  (.A(II9591), .Z(g5949) ) ;
AND2    gate3767  (.A(g3709), .B(g4586), .Z(g5083) ) ;
INV     gate3768  (.A(g5083), .Z(II9594) ) ;
INV     gate3769  (.A(II9594), .Z(g5980) ) ;
INV     gate3770  (.A(g5120), .Z(II9598) ) ;
INV     gate3771  (.A(II9598), .Z(g5982) ) ;
INV     gate3772  (.A(g5013), .Z(II9602) ) ;
INV     gate3773  (.A(II9602), .Z(g5984) ) ;
INV     gate3774  (.A(g5620), .Z(II9605) ) ;
INV     gate3775  (.A(II9605), .Z(g5987) ) ;
INV     gate3776  (.A(g5127), .Z(II9608) ) ;
INV     gate3777  (.A(II9608), .Z(g5992) ) ;
INV     gate3778  (.A(g5149), .Z(II9612) ) ;
INV     gate3779  (.A(II9612), .Z(g5994) ) ;
OR2     gate3780  (.A(g4476), .B(g3440), .Z(g5405) ) ;
INV     gate3781  (.A(g5405), .Z(II9617) ) ;
INV     gate3782  (.A(II9617), .Z(g5997) ) ;
OR2     gate3783  (.A(g4345), .B(g3496), .Z(g5189) ) ;
INV     gate3784  (.A(g5189), .Z(II9620) ) ;
INV     gate3785  (.A(II9620), .Z(g5998) ) ;
INV     gate3786  (.A(g5405), .Z(II9625) ) ;
INV     gate3787  (.A(II9625), .Z(g6001) ) ;
INV     gate3788  (.A(g5309), .Z(g6014) ) ;
INV     gate3789  (.A(g5557), .Z(II9632) ) ;
INV     gate3790  (.A(II9632), .Z(g6016) ) ;
AND2    gate3791  (.A(g3076), .B(g4638), .Z(g5126) ) ;
INV     gate3792  (.A(g5126), .Z(II9639) ) ;
INV     gate3793  (.A(II9639), .Z(g6030) ) ;
OR2     gate3794  (.A(g4364), .B(g3516), .Z(g5229) ) ;
INV     gate3795  (.A(g5229), .Z(II9642) ) ;
INV     gate3796  (.A(II9642), .Z(g6031) ) ;
AND2    gate3797  (.A(g3088), .B(g4671), .Z(g5148) ) ;
INV     gate3798  (.A(g5148), .Z(II9647) ) ;
INV     gate3799  (.A(II9647), .Z(g6036) ) ;
INV     gate3800  (.A(g5426), .Z(II9652) ) ;
INV     gate3801  (.A(II9652), .Z(g6039) ) ;
AND2    gate3802  (.A(g3094), .B(g4676), .Z(g5173) ) ;
INV     gate3803  (.A(g5173), .Z(II9655) ) ;
INV     gate3804  (.A(II9655), .Z(g6040) ) ;
AND2    gate3805  (.A(g1275), .B(g4678), .Z(g5150) ) ;
INV     gate3806  (.A(g5150), .Z(II9658) ) ;
INV     gate3807  (.A(II9658), .Z(g6041) ) ;
NAND2   gate3808  (.A(II8804), .B(II8805), .Z(g5319) ) ;
INV     gate3809  (.A(g5319), .Z(II9662) ) ;
INV     gate3810  (.A(II9662), .Z(g6043) ) ;
AND2    gate3811  (.A(g1235), .B(g4681), .Z(g5174) ) ;
INV     gate3812  (.A(g5174), .Z(II9665) ) ;
INV     gate3813  (.A(II9665), .Z(g6044) ) ;
INV     gate3814  (.A(g5426), .Z(II9669) ) ;
INV     gate3815  (.A(II9669), .Z(g6046) ) ;
AND2    gate3816  (.A(g1240), .B(g4713), .Z(g5182) ) ;
INV     gate3817  (.A(g5182), .Z(II9673) ) ;
INV     gate3818  (.A(II9673), .Z(g6048) ) ;
AND2    gate3819  (.A(g1245), .B(g4716), .Z(g5190) ) ;
INV     gate3820  (.A(g5190), .Z(II9677) ) ;
INV     gate3821  (.A(II9677), .Z(g6050) ) ;
AND2    gate3822  (.A(g1610), .B(g4717), .Z(g5194) ) ;
INV     gate3823  (.A(g5194), .Z(II9680) ) ;
INV     gate3824  (.A(II9680), .Z(g6051) ) ;
INV     gate3825  (.A(g5426), .Z(g6052) ) ;
INV     gate3826  (.A(g5426), .Z(II9684) ) ;
INV     gate3827  (.A(II9684), .Z(g6053) ) ;
AND2    gate3828  (.A(g1250), .B(g4721), .Z(g5201) ) ;
INV     gate3829  (.A(g5201), .Z(II9688) ) ;
INV     gate3830  (.A(II9688), .Z(g6055) ) ;
INV     gate3831  (.A(g5426), .Z(g6056) ) ;
INV     gate3832  (.A(g5446), .Z(g6057) ) ;
AND2    gate3833  (.A(g1255), .B(g4726), .Z(g5212) ) ;
INV     gate3834  (.A(g5212), .Z(II9695) ) ;
INV     gate3835  (.A(II9695), .Z(g6060) ) ;
INV     gate3836  (.A(g5426), .Z(II9699) ) ;
INV     gate3837  (.A(II9699), .Z(g6062) ) ;
INV     gate3838  (.A(g5446), .Z(g6063) ) ;
AND2    gate3839  (.A(g1260), .B(g4730), .Z(g5221) ) ;
INV     gate3840  (.A(g5221), .Z(II9706) ) ;
INV     gate3841  (.A(II9706), .Z(g6069) ) ;
AND2    gate3842  (.A(g4567), .B(g4807), .Z(g4977) ) ;
INV     gate3843  (.A(g4977), .Z(g6072) ) ;
AND2    gate3844  (.A(g1265), .B(g4735), .Z(g5230) ) ;
INV     gate3845  (.A(g5230), .Z(II9712) ) ;
INV     gate3846  (.A(II9712), .Z(g6073) ) ;
INV     gate3847  (.A(g5426), .Z(II9717) ) ;
INV     gate3848  (.A(II9717), .Z(g6076) ) ;
AND2    gate3849  (.A(g673), .B(g4738), .Z(g5248) ) ;
INV     gate3850  (.A(g5248), .Z(II9720) ) ;
INV     gate3851  (.A(II9720), .Z(g6077) ) ;
INV     gate3852  (.A(g4977), .Z(g6081) ) ;
AND2    gate3853  (.A(g1270), .B(g4748), .Z(g5250) ) ;
INV     gate3854  (.A(g5250), .Z(II9727) ) ;
INV     gate3855  (.A(II9727), .Z(g6082) ) ;
AND2    gate3856  (.A(g682), .B(g4754), .Z(g5255) ) ;
INV     gate3857  (.A(g5255), .Z(II9731) ) ;
INV     gate3858  (.A(II9731), .Z(g6084) ) ;
AND2    gate3859  (.A(g691), .B(g4755), .Z(g5257) ) ;
INV     gate3860  (.A(g5257), .Z(II9734) ) ;
INV     gate3861  (.A(II9734), .Z(g6085) ) ;
AND2    gate3862  (.A(g700), .B(g4756), .Z(g5258) ) ;
INV     gate3863  (.A(g5258), .Z(II9737) ) ;
INV     gate3864  (.A(II9737), .Z(g6086) ) ;
INV     gate3865  (.A(g4977), .Z(g6089) ) ;
AND2    gate3866  (.A(g709), .B(g4761), .Z(g5263) ) ;
INV     gate3867  (.A(g5263), .Z(II9744) ) ;
INV     gate3868  (.A(II9744), .Z(g6091) ) ;
AND2    gate3869  (.A(g718), .B(g4766), .Z(g5266) ) ;
INV     gate3870  (.A(g5266), .Z(II9749) ) ;
INV     gate3871  (.A(II9749), .Z(g6094) ) ;
AND2    gate3872  (.A(g727), .B(g4772), .Z(g5271) ) ;
INV     gate3873  (.A(g5271), .Z(II9754) ) ;
INV     gate3874  (.A(II9754), .Z(g6097) ) ;
INV     gate3875  (.A(g5344), .Z(II9759) ) ;
INV     gate3876  (.A(II9759), .Z(g6100) ) ;
AND2    gate3877  (.A(g736), .B(g4780), .Z(g5276) ) ;
INV     gate3878  (.A(g5276), .Z(II9762) ) ;
INV     gate3879  (.A(II9762), .Z(g6101) ) ;
INV     gate3880  (.A(g5348), .Z(II9766) ) ;
INV     gate3881  (.A(II9766), .Z(g6103) ) ;
AND2    gate3882  (.A(g3876), .B(g4782), .Z(g5287) ) ;
INV     gate3883  (.A(g5287), .Z(II9769) ) ;
INV     gate3884  (.A(II9769), .Z(g6104) ) ;
INV     gate3885  (.A(g4934), .Z(II9773) ) ;
INV     gate3886  (.A(II9773), .Z(g6106) ) ;
INV     gate3887  (.A(g5353), .Z(II9776) ) ;
INV     gate3888  (.A(II9776), .Z(g6107) ) ;
INV     gate3889  (.A(g5391), .Z(II9779) ) ;
INV     gate3890  (.A(II9779), .Z(g6108) ) ;
INV     gate3891  (.A(g5052), .Z(g6109) ) ;
INV     gate3892  (.A(g5395), .Z(II9783) ) ;
INV     gate3893  (.A(II9783), .Z(g6110) ) ;
OR2     gate3894  (.A(g4481), .B(g3684), .Z(g5396) ) ;
INV     gate3895  (.A(g5396), .Z(II9786) ) ;
INV     gate3896  (.A(II9786), .Z(g6111) ) ;
INV     gate3897  (.A(g5401), .Z(II9789) ) ;
INV     gate3898  (.A(II9789), .Z(g6112) ) ;
OR2     gate3899  (.A(g4486), .B(g3695), .Z(g5403) ) ;
INV     gate3900  (.A(g5403), .Z(II9792) ) ;
INV     gate3901  (.A(II9792), .Z(g6113) ) ;
OR2     gate3902  (.A(g4487), .B(g3696), .Z(g5404) ) ;
INV     gate3903  (.A(g5404), .Z(II9795) ) ;
INV     gate3904  (.A(II9795), .Z(g6114) ) ;
INV     gate3905  (.A(g5415), .Z(II9798) ) ;
INV     gate3906  (.A(II9798), .Z(g6115) ) ;
INV     gate3907  (.A(g5416), .Z(II9801) ) ;
INV     gate3908  (.A(II9801), .Z(g6116) ) ;
INV     gate3909  (.A(g5417), .Z(II9804) ) ;
INV     gate3910  (.A(II9804), .Z(g6117) ) ;
INV     gate3911  (.A(g5419), .Z(II9807) ) ;
INV     gate3912  (.A(II9807), .Z(g6118) ) ;
INV     gate3913  (.A(g5576), .Z(II9810) ) ;
INV     gate3914  (.A(II9810), .Z(g6119) ) ;
INV     gate3915  (.A(g5241), .Z(II9813) ) ;
INV     gate3916  (.A(II9813), .Z(g6120) ) ;
INV     gate3917  (.A(g5576), .Z(II9816) ) ;
INV     gate3918  (.A(II9816), .Z(g6121) ) ;
NAND2   gate3919  (.A(II8651), .B(II8652), .Z(g5219) ) ;
INV     gate3920  (.A(g5219), .Z(II9822) ) ;
INV     gate3921  (.A(II9822), .Z(g6125) ) ;
AND2    gate3922  (.A(g3220), .B(g4819), .Z(g5390) ) ;
INV     gate3923  (.A(g5390), .Z(II9826) ) ;
INV     gate3924  (.A(II9826), .Z(g6127) ) ;
INV     gate3925  (.A(g5013), .Z(II9829) ) ;
INV     gate3926  (.A(II9829), .Z(g6128) ) ;
NAND2   gate3927  (.A(g1840), .B(g4401), .Z(g5548) ) ;
INV     gate3928  (.A(g5548), .Z(g6131) ) ;
INV     gate3929  (.A(g5197), .Z(II9833) ) ;
INV     gate3930  (.A(II9833), .Z(g6132) ) ;
INV     gate3931  (.A(g5405), .Z(II9836) ) ;
INV     gate3932  (.A(II9836), .Z(g6133) ) ;
NAND2   gate3933  (.A(II8670), .B(II8671), .Z(g5226) ) ;
INV     gate3934  (.A(g5226), .Z(II9839) ) ;
INV     gate3935  (.A(II9839), .Z(g6134) ) ;
INV     gate3936  (.A(g5405), .Z(II9842) ) ;
INV     gate3937  (.A(II9842), .Z(g6135) ) ;
INV     gate3938  (.A(g5405), .Z(II9845) ) ;
INV     gate3939  (.A(II9845), .Z(g6136) ) ;
INV     gate3940  (.A(g5557), .Z(II9848) ) ;
INV     gate3941  (.A(II9848), .Z(g6137) ) ;
INV     gate3942  (.A(g5405), .Z(II9851) ) ;
INV     gate3943  (.A(II9851), .Z(g6140) ) ;
INV     gate3944  (.A(g5557), .Z(II9854) ) ;
INV     gate3945  (.A(II9854), .Z(g6141) ) ;
NAND2   gate3946  (.A(II8716), .B(II8717), .Z(g5269) ) ;
INV     gate3947  (.A(g5269), .Z(II9857) ) ;
INV     gate3948  (.A(II9857), .Z(g6144) ) ;
INV     gate3949  (.A(g5405), .Z(II9860) ) ;
INV     gate3950  (.A(II9860), .Z(g6145) ) ;
INV     gate3951  (.A(g5557), .Z(II9863) ) ;
INV     gate3952  (.A(II9863), .Z(g6146) ) ;
NAND2   gate3953  (.A(II8729), .B(II8730), .Z(g5274) ) ;
INV     gate3954  (.A(g5274), .Z(II9866) ) ;
INV     gate3955  (.A(II9866), .Z(g6149) ) ;
INV     gate3956  (.A(g5405), .Z(II9869) ) ;
INV     gate3957  (.A(II9869), .Z(g6150) ) ;
INV     gate3958  (.A(g5557), .Z(II9872) ) ;
INV     gate3959  (.A(II9872), .Z(g6151) ) ;
NAND2   gate3960  (.A(II8739), .B(II8740), .Z(g5278) ) ;
INV     gate3961  (.A(g5278), .Z(II9875) ) ;
INV     gate3962  (.A(II9875), .Z(g6154) ) ;
INV     gate3963  (.A(g5426), .Z(g6156) ) ;
INV     gate3964  (.A(g5405), .Z(II9880) ) ;
INV     gate3965  (.A(II9880), .Z(g6157) ) ;
INV     gate3966  (.A(g5557), .Z(II9883) ) ;
INV     gate3967  (.A(II9883), .Z(g6158) ) ;
NAND2   gate3968  (.A(II8751), .B(II8752), .Z(g5286) ) ;
INV     gate3969  (.A(g5286), .Z(II9886) ) ;
INV     gate3970  (.A(II9886), .Z(g6161) ) ;
INV     gate3971  (.A(g5426), .Z(g6164) ) ;
INV     gate3972  (.A(g5446), .Z(g6165) ) ;
INV     gate3973  (.A(g5557), .Z(II9893) ) ;
INV     gate3974  (.A(II9893), .Z(g6166) ) ;
NAND2   gate3975  (.A(II8762), .B(II8763), .Z(g5295) ) ;
INV     gate3976  (.A(g5295), .Z(II9896) ) ;
INV     gate3977  (.A(II9896), .Z(g6169) ) ;
INV     gate3978  (.A(g5426), .Z(g6170) ) ;
INV     gate3979  (.A(g5446), .Z(g6171) ) ;
INV     gate3980  (.A(g5557), .Z(II9901) ) ;
INV     gate3981  (.A(II9901), .Z(g6172) ) ;
INV     gate3982  (.A(g5320), .Z(g6175) ) ;
NAND2   gate3983  (.A(II8771), .B(II8772), .Z(g5300) ) ;
INV     gate3984  (.A(g5300), .Z(II9905) ) ;
INV     gate3985  (.A(II9905), .Z(g6176) ) ;
INV     gate3986  (.A(g4977), .Z(g6178) ) ;
INV     gate3987  (.A(g5426), .Z(g6181) ) ;
INV     gate3988  (.A(g5446), .Z(g6182) ) ;
INV     gate3989  (.A(g5320), .Z(g6183) ) ;
NAND2   gate3990  (.A(II8779), .B(II8780), .Z(g5304) ) ;
INV     gate3991  (.A(g5304), .Z(II9915) ) ;
INV     gate3992  (.A(II9915), .Z(g6184) ) ;
INV     gate3993  (.A(g5426), .Z(g6190) ) ;
INV     gate3994  (.A(g5446), .Z(g6191) ) ;
NAND2   gate3995  (.A(II8787), .B(II8788), .Z(g5308) ) ;
INV     gate3996  (.A(g5308), .Z(II9923) ) ;
INV     gate3997  (.A(II9923), .Z(g6192) ) ;
INV     gate3998  (.A(g5426), .Z(g6195) ) ;
INV     gate3999  (.A(g5446), .Z(g6196) ) ;
NAND2   gate4000  (.A(II8796), .B(II8797), .Z(g5317) ) ;
INV     gate4001  (.A(g5317), .Z(II9930) ) ;
INV     gate4002  (.A(II9930), .Z(g6197) ) ;
AND2    gate4003  (.A(g1887), .B(g4241), .Z(g5477) ) ;
INV     gate4004  (.A(g5477), .Z(II9935) ) ;
INV     gate4005  (.A(II9935), .Z(g6200) ) ;
AND2    gate4006  (.A(g1905), .B(g4242), .Z(g5478) ) ;
INV     gate4007  (.A(g5478), .Z(II9938) ) ;
INV     gate4008  (.A(II9938), .Z(g6201) ) ;
INV     gate4009  (.A(g5426), .Z(g6202) ) ;
INV     gate4010  (.A(g5446), .Z(g6203) ) ;
AND2    gate4011  (.A(g1896), .B(g4256), .Z(g5484) ) ;
INV     gate4012  (.A(g5484), .Z(II9953) ) ;
INV     gate4013  (.A(II9953), .Z(g6208) ) ;
AND2    gate4014  (.A(g1914), .B(g4257), .Z(g5485) ) ;
INV     gate4015  (.A(g5485), .Z(II9956) ) ;
INV     gate4016  (.A(II9956), .Z(g6209) ) ;
INV     gate4017  (.A(g5205), .Z(g6210) ) ;
INV     gate4018  (.A(g5426), .Z(g6213) ) ;
INV     gate4019  (.A(g5446), .Z(g6214) ) ;
AND2    gate4020  (.A(g1923), .B(g4265), .Z(g5493) ) ;
INV     gate4021  (.A(g5493), .Z(II9965) ) ;
INV     gate4022  (.A(II9965), .Z(g6218) ) ;
INV     gate4023  (.A(g5426), .Z(g6219) ) ;
INV     gate4024  (.A(g5446), .Z(g6220) ) ;
AND2    gate4025  (.A(g1932), .B(g4275), .Z(g5502) ) ;
INV     gate4026  (.A(g5502), .Z(II9973) ) ;
INV     gate4027  (.A(II9973), .Z(g6226) ) ;
INV     gate4028  (.A(g5446), .Z(g6227) ) ;
AND2    gate4029  (.A(g1941), .B(g4284), .Z(g5514) ) ;
INV     gate4030  (.A(g5514), .Z(II9981) ) ;
INV     gate4031  (.A(II9981), .Z(g6236) ) ;
AND2    gate4032  (.A(g4129), .B(g4288), .Z(g5529) ) ;
INV     gate4033  (.A(g5529), .Z(II9984) ) ;
INV     gate4034  (.A(II9984), .Z(g6237) ) ;
AND2    gate4035  (.A(g1950), .B(g4294), .Z(g5526) ) ;
INV     gate4036  (.A(g5526), .Z(II9988) ) ;
INV     gate4037  (.A(II9988), .Z(g6239) ) ;
INV     gate4038  (.A(g5633), .Z(II9992) ) ;
INV     gate4039  (.A(II9992), .Z(g6241) ) ;
AND2    gate4040  (.A(g4867), .B(g4298), .Z(g5536) ) ;
INV     gate4041  (.A(g5536), .Z(II9995) ) ;
INV     gate4042  (.A(II9995), .Z(g6242) ) ;
INV     gate4043  (.A(g4908), .Z(II10003) ) ;
INV     gate4044  (.A(II10003), .Z(g6248) ) ;
INV     gate4045  (.A(g5633), .Z(II10006) ) ;
INV     gate4046  (.A(II10006), .Z(g6249) ) ;
INV     gate4047  (.A(g5542), .Z(II10009) ) ;
INV     gate4048  (.A(II10009), .Z(g6250) ) ;
AND2    gate4049  (.A(g4874), .B(g4312), .Z(g5543) ) ;
INV     gate4050  (.A(g5543), .Z(II10012) ) ;
INV     gate4051  (.A(II10012), .Z(g6251) ) ;
INV     gate4052  (.A(g5641), .Z(II10015) ) ;
INV     gate4053  (.A(II10015), .Z(g6252) ) ;
INV     gate4054  (.A(g5862), .Z(II10018) ) ;
INV     gate4055  (.A(g5692), .Z(II10021) ) ;
INV     gate4056  (.A(g5700), .Z(II10024) ) ;
INV     gate4057  (.A(g5751), .Z(II10027) ) ;
INV     gate4058  (.A(g5685), .Z(II10030) ) ;
INV     gate4059  (.A(g5693), .Z(II10033) ) ;
INV     gate4060  (.A(g5701), .Z(II10036) ) ;
INV     gate4061  (.A(g5718), .Z(II10039) ) ;
INV     gate4062  (.A(g5723), .Z(II10042) ) ;
INV     gate4063  (.A(g5727), .Z(II10045) ) ;
INV     gate4064  (.A(g5734), .Z(II10048) ) ;
INV     gate4065  (.A(g5702), .Z(II10051) ) ;
INV     gate4066  (.A(g5728), .Z(II10054) ) ;
INV     gate4067  (.A(g5741), .Z(II10057) ) ;
INV     gate4068  (.A(g5752), .Z(II10060) ) ;
INV     gate4069  (.A(g5766), .Z(II10063) ) ;
INV     gate4070  (.A(g5778), .Z(II10066) ) ;
INV     gate4071  (.A(g5787), .Z(II10069) ) ;
INV     gate4072  (.A(g5719), .Z(II10072) ) ;
INV     gate4073  (.A(g5724), .Z(II10075) ) ;
INV     gate4074  (.A(g5729), .Z(II10078) ) ;
INV     gate4075  (.A(g5735), .Z(II10081) ) ;
INV     gate4076  (.A(g5742), .Z(II10084) ) ;
INV     gate4077  (.A(g5753), .Z(II10087) ) ;
INV     gate4078  (.A(g5767), .Z(II10090) ) ;
INV     gate4079  (.A(g5779), .Z(II10093) ) ;
INV     gate4080  (.A(g5794), .Z(II10096) ) ;
INV     gate4081  (.A(g5800), .Z(II10099) ) ;
INV     gate4082  (.A(g5730), .Z(II10102) ) ;
INV     gate4083  (.A(g5736), .Z(II10105) ) ;
INV     gate4084  (.A(g5743), .Z(II10108) ) ;
INV     gate4085  (.A(g5754), .Z(II10111) ) ;
INV     gate4086  (.A(g5768), .Z(II10114) ) ;
INV     gate4087  (.A(g6241), .Z(II10117) ) ;
INV     gate4088  (.A(g6248), .Z(II10120) ) ;
INV     gate4089  (.A(g5676), .Z(II10123) ) ;
INV     gate4090  (.A(g5682), .Z(II10126) ) ;
INV     gate4091  (.A(g5688), .Z(II10129) ) ;
INV     gate4092  (.A(g5696), .Z(II10132) ) ;
INV     gate4093  (.A(g6249), .Z(II10135) ) ;
INV     gate4094  (.A(g5677), .Z(II10138) ) ;
INV     gate4095  (.A(g5683), .Z(II10141) ) ;
INV     gate4096  (.A(g5689), .Z(II10144) ) ;
INV     gate4097  (.A(g5697), .Z(II10147) ) ;
INV     gate4098  (.A(g5705), .Z(II10150) ) ;
INV     gate4099  (.A(g5947), .Z(II10153) ) ;
INV     gate4100  (.A(g6100), .Z(II10156) ) ;
INV     gate4101  (.A(g5936), .Z(II10159) ) ;
INV     gate4102  (.A(g5943), .Z(II10162) ) ;
INV     gate4103  (.A(g5948), .Z(II10165) ) ;
INV     gate4104  (.A(g5982), .Z(II10168) ) ;
INV     gate4105  (.A(g5992), .Z(II10171) ) ;
INV     gate4106  (.A(g5994), .Z(II10174) ) ;
INV     gate4107  (.A(g6103), .Z(II10177) ) ;
INV     gate4108  (.A(g6107), .Z(II10180) ) ;
INV     gate4109  (.A(g6108), .Z(II10183) ) ;
INV     gate4110  (.A(g6110), .Z(II10186) ) ;
INV     gate4111  (.A(g6112), .Z(II10189) ) ;
INV     gate4112  (.A(g6115), .Z(II10192) ) ;
INV     gate4113  (.A(g6116), .Z(II10195) ) ;
INV     gate4114  (.A(g6118), .Z(II10198) ) ;
INV     gate4115  (.A(g5998), .Z(II10201) ) ;
INV     gate4116  (.A(g6031), .Z(II10204) ) ;
INV     gate4117  (.A(g6117), .Z(II10221) ) ;
INV     gate4118  (.A(g6113), .Z(II10228) ) ;
INV     gate4119  (.A(g6111), .Z(II10231) ) ;
INV     gate4120  (.A(g6114), .Z(II10234) ) ;
INV     gate4121  (.A(g6120), .Z(II10237) ) ;
INV     gate4122  (.A(g5937), .Z(II10240) ) ;
AND3    gate4123  (.A(g2965), .B(g5292), .C(g4609), .Z(g5918) ) ;
INV     gate4124  (.A(g5918), .Z(II10243) ) ;
INV     gate4125  (.A(II10243), .Z(g6340) ) ;
INV     gate4126  (.A(g6125), .Z(II10248) ) ;
INV     gate4127  (.A(II10248), .Z(g6343) ) ;
AND2    gate4128  (.A(g5639), .B(g4319), .Z(g6126) ) ;
INV     gate4129  (.A(g6126), .Z(II10251) ) ;
INV     gate4130  (.A(II10251), .Z(g6344) ) ;
INV     gate4131  (.A(g6134), .Z(II10258) ) ;
INV     gate4132  (.A(II10258), .Z(g6349) ) ;
OR2     gate4133  (.A(g3440), .B(g4921), .Z(g5867) ) ;
INV     gate4134  (.A(g5867), .Z(g6354) ) ;
INV     gate4135  (.A(g5867), .Z(g6361) ) ;
INV     gate4136  (.A(g5811), .Z(II10274) ) ;
INV     gate4137  (.A(II10274), .Z(g6365) ) ;
INV     gate4138  (.A(g5987), .Z(g6368) ) ;
INV     gate4139  (.A(g5815), .Z(II10278) ) ;
INV     gate4140  (.A(II10278), .Z(g6382) ) ;
INV     gate4141  (.A(g6119), .Z(g6385) ) ;
AND2    gate4142  (.A(g4572), .B(g5354), .Z(g6163) ) ;
INV     gate4143  (.A(g6163), .Z(II10282) ) ;
INV     gate4144  (.A(II10282), .Z(g6386) ) ;
INV     gate4145  (.A(g6121), .Z(g6387) ) ;
INV     gate4146  (.A(g6237), .Z(II10286) ) ;
INV     gate4147  (.A(II10286), .Z(g6388) ) ;
NAND2   gate4148  (.A(g5552), .B(g5548), .Z(g6003) ) ;
INV     gate4149  (.A(g6003), .Z(II10289) ) ;
INV     gate4150  (.A(II10289), .Z(g6389) ) ;
AND2    gate4151  (.A(g5272), .B(g2173), .Z(g5863) ) ;
INV     gate4152  (.A(g5863), .Z(II10293) ) ;
INV     gate4153  (.A(II10293), .Z(g6395) ) ;
INV     gate4154  (.A(g6242), .Z(II10296) ) ;
INV     gate4155  (.A(II10296), .Z(g6396) ) ;
OR2     gate4156  (.A(g5537), .B(g4774), .Z(g6243) ) ;
INV     gate4157  (.A(g6243), .Z(II10299) ) ;
INV     gate4158  (.A(II10299), .Z(g6397) ) ;
AND2    gate4159  (.A(g5115), .B(g5354), .Z(g6179) ) ;
INV     gate4160  (.A(g6179), .Z(II10302) ) ;
INV     gate4161  (.A(II10302), .Z(g6398) ) ;
AND2    gate4162  (.A(g2190), .B(g5128), .Z(g6180) ) ;
INV     gate4163  (.A(g6180), .Z(II10305) ) ;
INV     gate4164  (.A(II10305), .Z(g6399) ) ;
INV     gate4165  (.A(g6003), .Z(II10308) ) ;
INV     gate4166  (.A(II10308), .Z(g6400) ) ;
INV     gate4167  (.A(g6128), .Z(g6403) ) ;
INV     gate4168  (.A(g6133), .Z(g6405) ) ;
INV     gate4169  (.A(g6251), .Z(II10314) ) ;
INV     gate4170  (.A(II10314), .Z(g6406) ) ;
INV     gate4171  (.A(g6003), .Z(II10317) ) ;
INV     gate4172  (.A(II10317), .Z(g6407) ) ;
INV     gate4173  (.A(g6135), .Z(g6411) ) ;
AND2    gate4174  (.A(g2206), .B(g5151), .Z(g6193) ) ;
INV     gate4175  (.A(g6193), .Z(II10322) ) ;
INV     gate4176  (.A(II10322), .Z(g6412) ) ;
INV     gate4177  (.A(g6003), .Z(II10325) ) ;
INV     gate4178  (.A(II10325), .Z(g6413) ) ;
INV     gate4179  (.A(g6136), .Z(g6417) ) ;
INV     gate4180  (.A(g6137), .Z(g6418) ) ;
AND2    gate4181  (.A(g1499), .B(g5128), .Z(g6198) ) ;
INV     gate4182  (.A(g6198), .Z(II10331) ) ;
INV     gate4183  (.A(II10331), .Z(g6419) ) ;
INV     gate4184  (.A(g6003), .Z(II10334) ) ;
INV     gate4185  (.A(II10334), .Z(g6420) ) ;
INV     gate4186  (.A(g6140), .Z(g6424) ) ;
INV     gate4187  (.A(g6141), .Z(g6425) ) ;
AND2    gate4188  (.A(g1515), .B(g5151), .Z(g6205) ) ;
INV     gate4189  (.A(g6205), .Z(II10340) ) ;
INV     gate4190  (.A(II10340), .Z(g6426) ) ;
INV     gate4191  (.A(g6003), .Z(II10343) ) ;
INV     gate4192  (.A(II10343), .Z(g6427) ) ;
INV     gate4193  (.A(g6145), .Z(g6431) ) ;
INV     gate4194  (.A(g6146), .Z(g6432) ) ;
AND2    gate4195  (.A(g1504), .B(g5128), .Z(g6215) ) ;
INV     gate4196  (.A(g6215), .Z(II10349) ) ;
INV     gate4197  (.A(II10349), .Z(g6433) ) ;
AND2    gate4198  (.A(g2232), .B(g5151), .Z(g6216) ) ;
INV     gate4199  (.A(g6216), .Z(II10352) ) ;
INV     gate4200  (.A(II10352), .Z(g6434) ) ;
INV     gate4201  (.A(g6003), .Z(II10355) ) ;
INV     gate4202  (.A(II10355), .Z(g6435) ) ;
INV     gate4203  (.A(g6150), .Z(g6440) ) ;
INV     gate4204  (.A(g6151), .Z(g6441) ) ;
AND2    gate4205  (.A(g1520), .B(g5151), .Z(g6224) ) ;
INV     gate4206  (.A(g6224), .Z(II10362) ) ;
INV     gate4207  (.A(II10362), .Z(g6442) ) ;
INV     gate4208  (.A(g6157), .Z(g6443) ) ;
INV     gate4209  (.A(g6158), .Z(g6444) ) ;
AND2    gate4210  (.A(g2244), .B(g5151), .Z(g6234) ) ;
INV     gate4211  (.A(g6234), .Z(II10367) ) ;
INV     gate4212  (.A(II10367), .Z(g6445) ) ;
OR2     gate4213  (.A(g5418), .B(g4670), .Z(g5857) ) ;
INV     gate4214  (.A(g5857), .Z(II10370) ) ;
INV     gate4215  (.A(II10370), .Z(g6446) ) ;
INV     gate4216  (.A(g6166), .Z(g6447) ) ;
OR2     gate4217  (.A(g5632), .B(g4883), .Z(g5852) ) ;
INV     gate4218  (.A(g5852), .Z(II10374) ) ;
INV     gate4219  (.A(II10374), .Z(g6448) ) ;
INV     gate4220  (.A(g6172), .Z(g6449) ) ;
AND2    gate4221  (.A(g2255), .B(g5151), .Z(g6244) ) ;
INV     gate4222  (.A(g6244), .Z(II10378) ) ;
INV     gate4223  (.A(II10378), .Z(g6450) ) ;
OR2     gate4224  (.A(g5626), .B(g4877), .Z(g5847) ) ;
INV     gate4225  (.A(g5847), .Z(II10381) ) ;
INV     gate4226  (.A(II10381), .Z(g6451) ) ;
OR2     gate4227  (.A(g5618), .B(g4870), .Z(g5842) ) ;
INV     gate4228  (.A(g5842), .Z(II10384) ) ;
INV     gate4229  (.A(II10384), .Z(g6452) ) ;
INV     gate4230  (.A(g5817), .Z(g6453) ) ;
INV     gate4231  (.A(g5830), .Z(II10388) ) ;
INV     gate4232  (.A(II10388), .Z(g6454) ) ;
OR2     gate4233  (.A(g5612), .B(g4866), .Z(g5838) ) ;
INV     gate4234  (.A(g5838), .Z(II10391) ) ;
INV     gate4235  (.A(II10391), .Z(g6461) ) ;
OR2     gate4236  (.A(g5602), .B(g4839), .Z(g5824) ) ;
INV     gate4237  (.A(g5824), .Z(II10394) ) ;
INV     gate4238  (.A(II10394), .Z(g6462) ) ;
OR2     gate4239  (.A(g5595), .B(g4834), .Z(g5820) ) ;
INV     gate4240  (.A(g5820), .Z(II10398) ) ;
INV     gate4241  (.A(II10398), .Z(g6464) ) ;
INV     gate4242  (.A(g5987), .Z(g6475) ) ;
INV     gate4243  (.A(g5821), .Z(II10412) ) ;
INV     gate4244  (.A(II10412), .Z(g6482) ) ;
INV     gate4245  (.A(g5867), .Z(g6499) ) ;
INV     gate4246  (.A(g5826), .Z(II10421) ) ;
INV     gate4247  (.A(II10421), .Z(g6503) ) ;
INV     gate4248  (.A(g5839), .Z(II10427) ) ;
INV     gate4249  (.A(II10427), .Z(g6509) ) ;
INV     gate4250  (.A(g5843), .Z(II10434) ) ;
INV     gate4251  (.A(II10434), .Z(g6517) ) ;
AND2    gate4252  (.A(g5103), .B(g5354), .Z(g5755) ) ;
INV     gate4253  (.A(g5755), .Z(II10437) ) ;
INV     gate4254  (.A(II10437), .Z(g6521) ) ;
AND2    gate4255  (.A(g4466), .B(g5128), .Z(g5770) ) ;
INV     gate4256  (.A(g5770), .Z(II10445) ) ;
INV     gate4257  (.A(II10445), .Z(g6527) ) ;
INV     gate4258  (.A(g5844), .Z(II10456) ) ;
INV     gate4259  (.A(II10456), .Z(g6536) ) ;
OR2     gate4260  (.A(g4949), .B(g4260), .Z(g5849) ) ;
INV     gate4261  (.A(g5849), .Z(II10461) ) ;
INV     gate4262  (.A(II10461), .Z(g6539) ) ;
INV     gate4263  (.A(g5888), .Z(g6543) ) ;
INV     gate4264  (.A(g5893), .Z(g6547) ) ;
INV     gate4265  (.A(g5733), .Z(g6552) ) ;
OR2     gate4266  (.A(g5254), .B(g3718), .Z(g6049) ) ;
INV     gate4267  (.A(g6049), .Z(II10477) ) ;
INV     gate4268  (.A(II10477), .Z(g6553) ) ;
INV     gate4269  (.A(g5740), .Z(g6555) ) ;
INV     gate4270  (.A(g5747), .Z(g6556) ) ;
INV     gate4271  (.A(g5748), .Z(g6557) ) ;
NOR2    gate4272  (.A(g4974), .B(g2864), .Z(g6155) ) ;
INV     gate4273  (.A(g6155), .Z(II10484) ) ;
INV     gate4274  (.A(II10484), .Z(g6558) ) ;
INV     gate4275  (.A(g5758), .Z(g6559) ) ;
INV     gate4276  (.A(g5759), .Z(g6560) ) ;
INV     gate4277  (.A(g5773), .Z(g6561) ) ;
INV     gate4278  (.A(g5774), .Z(g6562) ) ;
INV     gate4279  (.A(g5783), .Z(g6563) ) ;
INV     gate4280  (.A(g5784), .Z(g6564) ) ;
INV     gate4281  (.A(g5790), .Z(g6565) ) ;
INV     gate4282  (.A(g5791), .Z(g6566) ) ;
INV     gate4283  (.A(g6144), .Z(II10495) ) ;
INV     gate4284  (.A(II10495), .Z(g6567) ) ;
INV     gate4285  (.A(g5797), .Z(g6568) ) ;
INV     gate4286  (.A(g6149), .Z(II10499) ) ;
INV     gate4287  (.A(II10499), .Z(g6569) ) ;
INV     gate4288  (.A(g5949), .Z(g6570) ) ;
INV     gate4289  (.A(g5858), .Z(II10503) ) ;
INV     gate4290  (.A(II10503), .Z(g6571) ) ;
INV     gate4291  (.A(g5805), .Z(g6572) ) ;
INV     gate4292  (.A(g6154), .Z(II10514) ) ;
INV     gate4293  (.A(II10514), .Z(g6574) ) ;
INV     gate4294  (.A(g5949), .Z(g6575) ) ;
INV     gate4295  (.A(g6161), .Z(II10526) ) ;
INV     gate4296  (.A(II10526), .Z(g6578) ) ;
INV     gate4297  (.A(g5949), .Z(g6579) ) ;
INV     gate4298  (.A(g6169), .Z(II10531) ) ;
INV     gate4299  (.A(II10531), .Z(g6581) ) ;
INV     gate4300  (.A(g5949), .Z(g6582) ) ;
INV     gate4301  (.A(g5867), .Z(II10535) ) ;
INV     gate4302  (.A(II10535), .Z(g6583) ) ;
OR2     gate4303  (.A(g5023), .B(g4341), .Z(g5910) ) ;
INV     gate4304  (.A(g5910), .Z(II10538) ) ;
INV     gate4305  (.A(II10538), .Z(g6584) ) ;
INV     gate4306  (.A(g6176), .Z(II10541) ) ;
INV     gate4307  (.A(II10541), .Z(g6585) ) ;
INV     gate4308  (.A(g5949), .Z(g6586) ) ;
INV     gate4309  (.A(g5827), .Z(g6587) ) ;
OR2     gate4310  (.A(g5029), .B(g4343), .Z(g5914) ) ;
INV     gate4311  (.A(g5914), .Z(II10546) ) ;
INV     gate4312  (.A(II10546), .Z(g6588) ) ;
INV     gate4313  (.A(g6184), .Z(II10549) ) ;
INV     gate4314  (.A(II10549), .Z(g6589) ) ;
INV     gate4315  (.A(g5949), .Z(g6590) ) ;
INV     gate4316  (.A(g6192), .Z(II10553) ) ;
INV     gate4317  (.A(II10553), .Z(g6591) ) ;
INV     gate4318  (.A(g6197), .Z(II10557) ) ;
INV     gate4319  (.A(II10557), .Z(g6593) ) ;
INV     gate4320  (.A(g5887), .Z(II10560) ) ;
INV     gate4321  (.A(II10560), .Z(g6594) ) ;
INV     gate4322  (.A(g6043), .Z(II10563) ) ;
INV     gate4323  (.A(II10563), .Z(g6595) ) ;
INV     gate4324  (.A(g5904), .Z(II10566) ) ;
INV     gate4325  (.A(II10566), .Z(g6596) ) ;
NAND2   gate4326  (.A(g617), .B(g4921), .Z(g6019) ) ;
INV     gate4327  (.A(g6019), .Z(g6617) ) ;
INV     gate4328  (.A(g5980), .Z(II10573) ) ;
INV     gate4329  (.A(II10573), .Z(g6620) ) ;
INV     gate4330  (.A(g5864), .Z(II10584) ) ;
INV     gate4331  (.A(II10584), .Z(g6629) ) ;
NOR2    gate4332  (.A(g5350), .B(g5345), .Z(g5763) ) ;
INV     gate4333  (.A(g5763), .Z(II10589) ) ;
INV     gate4334  (.A(II10589), .Z(g6634) ) ;
INV     gate4335  (.A(g5865), .Z(II10592) ) ;
INV     gate4336  (.A(II10592), .Z(g6635) ) ;
INV     gate4337  (.A(g5874), .Z(II10598) ) ;
INV     gate4338  (.A(II10598), .Z(g6641) ) ;
OR2     gate4339  (.A(g5473), .B(g3908), .Z(g5996) ) ;
INV     gate4340  (.A(g5996), .Z(II10601) ) ;
INV     gate4341  (.A(II10601), .Z(g6644) ) ;
INV     gate4342  (.A(g5763), .Z(II10607) ) ;
INV     gate4343  (.A(II10607), .Z(g6648) ) ;
INV     gate4344  (.A(g5879), .Z(II10610) ) ;
INV     gate4345  (.A(II10610), .Z(g6649) ) ;
OR2     gate4346  (.A(g5480), .B(g3912), .Z(g6000) ) ;
INV     gate4347  (.A(g6000), .Z(II10613) ) ;
INV     gate4348  (.A(II10613), .Z(g6652) ) ;
INV     gate4349  (.A(g5884), .Z(II10620) ) ;
INV     gate4350  (.A(II10620), .Z(g6657) ) ;
OR2     gate4351  (.A(g5489), .B(g3939), .Z(g6002) ) ;
INV     gate4352  (.A(g6002), .Z(II10623) ) ;
INV     gate4353  (.A(II10623), .Z(g6660) ) ;
INV     gate4354  (.A(g5889), .Z(II10630) ) ;
INV     gate4355  (.A(II10630), .Z(g6667) ) ;
OR2     gate4356  (.A(g5497), .B(g3942), .Z(g6015) ) ;
INV     gate4357  (.A(g6015), .Z(II10633) ) ;
INV     gate4358  (.A(II10633), .Z(g6670) ) ;
INV     gate4359  (.A(g5830), .Z(II10639) ) ;
INV     gate4360  (.A(II10639), .Z(g6674) ) ;
OR2     gate4361  (.A(g5507), .B(g3970), .Z(g6026) ) ;
INV     gate4362  (.A(g6026), .Z(II10643) ) ;
INV     gate4363  (.A(II10643), .Z(g6680) ) ;
INV     gate4364  (.A(g5830), .Z(g6681) ) ;
INV     gate4365  (.A(g6030), .Z(II10648) ) ;
INV     gate4366  (.A(II10648), .Z(g6685) ) ;
OR2     gate4367  (.A(g5518), .B(g3974), .Z(g6035) ) ;
INV     gate4368  (.A(g6035), .Z(II10651) ) ;
INV     gate4369  (.A(II10651), .Z(g6686) ) ;
INV     gate4370  (.A(g6036), .Z(II10655) ) ;
INV     gate4371  (.A(II10655), .Z(g6688) ) ;
INV     gate4372  (.A(g5830), .Z(g6689) ) ;
OR2     gate4373  (.A(g5528), .B(g3979), .Z(g6038) ) ;
INV     gate4374  (.A(g6038), .Z(II10659) ) ;
INV     gate4375  (.A(II10659), .Z(g6692) ) ;
INV     gate4376  (.A(g6040), .Z(II10663) ) ;
INV     gate4377  (.A(II10663), .Z(g6694) ) ;
OR2     gate4378  (.A(g5535), .B(g3987), .Z(g6042) ) ;
INV     gate4379  (.A(g6042), .Z(II10666) ) ;
INV     gate4380  (.A(II10666), .Z(g6695) ) ;
INV     gate4381  (.A(g5949), .Z(g6697) ) ;
OR2     gate4382  (.A(g5541), .B(g3989), .Z(g6045) ) ;
INV     gate4383  (.A(g6045), .Z(II10671) ) ;
INV     gate4384  (.A(II10671), .Z(g6698) ) ;
INV     gate4385  (.A(g5949), .Z(g6700) ) ;
INV     gate4386  (.A(g5949), .Z(g6702) ) ;
INV     gate4387  (.A(g5777), .Z(II10678) ) ;
INV     gate4388  (.A(II10678), .Z(g6703) ) ;
INV     gate4389  (.A(g5949), .Z(g6704) ) ;
INV     gate4390  (.A(g6051), .Z(II10682) ) ;
INV     gate4391  (.A(II10682), .Z(g6705) ) ;
OR2     gate4392  (.A(g5199), .B(g4483), .Z(g6054) ) ;
INV     gate4393  (.A(g6054), .Z(II10685) ) ;
INV     gate4394  (.A(II10685), .Z(g6706) ) ;
INV     gate4395  (.A(g5949), .Z(g6707) ) ;
OR2     gate4396  (.A(g5211), .B(g4489), .Z(g6059) ) ;
INV     gate4397  (.A(g6059), .Z(II10689) ) ;
INV     gate4398  (.A(II10689), .Z(g6708) ) ;
INV     gate4399  (.A(g5949), .Z(g6709) ) ;
OR2     gate4400  (.A(g5220), .B(g4497), .Z(g6068) ) ;
INV     gate4401  (.A(g6068), .Z(II10693) ) ;
INV     gate4402  (.A(II10693), .Z(g6710) ) ;
INV     gate4403  (.A(g5949), .Z(g6711) ) ;
INV     gate4404  (.A(g5984), .Z(g6712) ) ;
INV     gate4405  (.A(g5856), .Z(II10698) ) ;
INV     gate4406  (.A(II10698), .Z(g6713) ) ;
INV     gate4407  (.A(g5867), .Z(g6714) ) ;
OR2     gate4408  (.A(g5228), .B(g4505), .Z(g6071) ) ;
INV     gate4409  (.A(g6071), .Z(II10702) ) ;
INV     gate4410  (.A(II10702), .Z(g6715) ) ;
INV     gate4411  (.A(g5949), .Z(g6716) ) ;
OR2     gate4412  (.A(g5249), .B(g4512), .Z(g6080) ) ;
INV     gate4413  (.A(g6080), .Z(II10706) ) ;
INV     gate4414  (.A(II10706), .Z(g6717) ) ;
INV     gate4415  (.A(g5949), .Z(g6718) ) ;
OR2     gate4416  (.A(g5260), .B(g4522), .Z(g6088) ) ;
INV     gate4417  (.A(g6088), .Z(II10710) ) ;
INV     gate4418  (.A(II10710), .Z(g6719) ) ;
INV     gate4419  (.A(g6003), .Z(II10713) ) ;
INV     gate4420  (.A(II10713), .Z(g6720) ) ;
OR2     gate4421  (.A(g5264), .B(g4534), .Z(g6093) ) ;
INV     gate4422  (.A(g6093), .Z(II10716) ) ;
INV     gate4423  (.A(II10716), .Z(g6723) ) ;
INV     gate4424  (.A(g6003), .Z(II10719) ) ;
INV     gate4425  (.A(II10719), .Z(g6724) ) ;
INV     gate4426  (.A(g5997), .Z(g6727) ) ;
OR2     gate4427  (.A(g5268), .B(g4542), .Z(g6096) ) ;
INV     gate4428  (.A(g6096), .Z(II10724) ) ;
INV     gate4429  (.A(II10724), .Z(g6729) ) ;
INV     gate4430  (.A(g6001), .Z(g6731) ) ;
NAND2   gate4431  (.A(II9558), .B(II9559), .Z(g5935) ) ;
INV     gate4432  (.A(g5935), .Z(II10729) ) ;
INV     gate4433  (.A(II10729), .Z(g6732) ) ;
OR2     gate4434  (.A(g5273), .B(g4550), .Z(g6099) ) ;
INV     gate4435  (.A(g6099), .Z(II10733) ) ;
INV     gate4436  (.A(II10733), .Z(g6734) ) ;
INV     gate4437  (.A(g6104), .Z(II10736) ) ;
INV     gate4438  (.A(II10736), .Z(g6735) ) ;
NAND2   gate4439  (.A(II9575), .B(II9576), .Z(g5942) ) ;
INV     gate4440  (.A(g5942), .Z(II10739) ) ;
INV     gate4441  (.A(II10739), .Z(g6736) ) ;
INV     gate4442  (.A(g6016), .Z(g6737) ) ;
INV     gate4443  (.A(g5830), .Z(g6742) ) ;
OR2     gate4444  (.A(g5591), .B(g4827), .Z(g5814) ) ;
INV     gate4445  (.A(g5814), .Z(II10753) ) ;
INV     gate4446  (.A(II10753), .Z(g6748) ) ;
OR2     gate4447  (.A(g5588), .B(g4823), .Z(g5810) ) ;
INV     gate4448  (.A(g5810), .Z(II10756) ) ;
INV     gate4449  (.A(II10756), .Z(g6749) ) ;
OR2     gate4450  (.A(g5575), .B(g4820), .Z(g5803) ) ;
INV     gate4451  (.A(g5803), .Z(II10759) ) ;
INV     gate4452  (.A(II10759), .Z(g6750) ) ;
INV     gate4453  (.A(g6127), .Z(II10762) ) ;
INV     gate4454  (.A(II10762), .Z(g6751) ) ;
INV     gate4455  (.A(g5987), .Z(g6764) ) ;
INV     gate4456  (.A(g5987), .Z(g6778) ) ;
INV     gate4457  (.A(g5867), .Z(II10789) ) ;
INV     gate4458  (.A(II10789), .Z(g6789) ) ;
AND2    gate4459  (.A(g5630), .B(g4311), .Z(g6123) ) ;
INV     gate4460  (.A(g6123), .Z(II10795) ) ;
INV     gate4461  (.A(II10795), .Z(g6793) ) ;
INV     gate4462  (.A(g6252), .Z(g6796) ) ;
INV     gate4463  (.A(g6536), .Z(II10801) ) ;
INV     gate4464  (.A(g6388), .Z(II10804) ) ;
INV     gate4465  (.A(g6396), .Z(II10807) ) ;
INV     gate4466  (.A(g6539), .Z(II10810) ) ;
INV     gate4467  (.A(g6397), .Z(II10813) ) ;
INV     gate4468  (.A(g6406), .Z(II10816) ) ;
INV     gate4469  (.A(g6706), .Z(II10819) ) ;
INV     gate4470  (.A(g6584), .Z(II10822) ) ;
INV     gate4471  (.A(g6588), .Z(II10825) ) ;
INV     gate4472  (.A(g6708), .Z(II10828) ) ;
INV     gate4473  (.A(g6710), .Z(II10831) ) ;
INV     gate4474  (.A(g6715), .Z(II10834) ) ;
INV     gate4475  (.A(g6717), .Z(II10837) ) ;
INV     gate4476  (.A(g6719), .Z(II10840) ) ;
INV     gate4477  (.A(g6723), .Z(II10843) ) ;
INV     gate4478  (.A(g6729), .Z(II10846) ) ;
INV     gate4479  (.A(g6734), .Z(II10849) ) ;
INV     gate4480  (.A(g6751), .Z(II10852) ) ;
INV     gate4481  (.A(g6685), .Z(II10855) ) ;
INV     gate4482  (.A(g6688), .Z(II10858) ) ;
INV     gate4483  (.A(g6694), .Z(II10861) ) ;
INV     gate4484  (.A(g6634), .Z(II10864) ) ;
AND2    gate4485  (.A(g201), .B(g5904), .Z(g6331) ) ;
INV     gate4486  (.A(g6331), .Z(II10873) ) ;
AND2    gate4487  (.A(g1374), .B(g5904), .Z(g6332) ) ;
INV     gate4488  (.A(g6332), .Z(II10885) ) ;
AND2    gate4489  (.A(g197), .B(g5904), .Z(g6333) ) ;
INV     gate4490  (.A(g6333), .Z(II10888) ) ;
AND2    gate4491  (.A(g1389), .B(g5904), .Z(g6334) ) ;
INV     gate4492  (.A(g6334), .Z(II10891) ) ;
INV     gate4493  (.A(g6735), .Z(II10898) ) ;
INV     gate4494  (.A(g6620), .Z(II10901) ) ;
INV     gate4495  (.A(g6558), .Z(II10904) ) ;
INV     gate4496  (.A(g6705), .Z(II10907) ) ;
INV     gate4497  (.A(g6703), .Z(II10910) ) ;
INV     gate4498  (.A(g6482), .Z(g6847) ) ;
AND2    gate4499  (.A(g6250), .B(g4318), .Z(g6728) ) ;
INV     gate4500  (.A(g6728), .Z(II10914) ) ;
INV     gate4501  (.A(II10914), .Z(g6852) ) ;
INV     gate4502  (.A(g6732), .Z(II10917) ) ;
INV     gate4503  (.A(II10917), .Z(g6853) ) ;
AND2    gate4504  (.A(g5678), .B(g4324), .Z(g6733) ) ;
INV     gate4505  (.A(g6733), .Z(II10920) ) ;
INV     gate4506  (.A(II10920), .Z(g6854) ) ;
INV     gate4507  (.A(g6736), .Z(II10924) ) ;
INV     gate4508  (.A(II10924), .Z(g6856) ) ;
OR2     gate4509  (.A(g6106), .B(g5479), .Z(g6755) ) ;
INV     gate4510  (.A(g6755), .Z(II10927) ) ;
INV     gate4511  (.A(II10927), .Z(g6857) ) ;
INV     gate4512  (.A(g6552), .Z(II10937) ) ;
INV     gate4513  (.A(II10937), .Z(g6859) ) ;
INV     gate4514  (.A(g6475), .Z(g6860) ) ;
INV     gate4515  (.A(g6555), .Z(II10941) ) ;
INV     gate4516  (.A(II10941), .Z(g6861) ) ;
INV     gate4517  (.A(g6720), .Z(g6862) ) ;
NAND2   gate4518  (.A(g6131), .B(g2550), .Z(g6740) ) ;
INV     gate4519  (.A(g6740), .Z(g6863) ) ;
NAND3   gate4520  (.A(g6132), .B(g6124), .C(g6122), .Z(g6548) ) ;
INV     gate4521  (.A(g6548), .Z(II10946) ) ;
INV     gate4522  (.A(II10946), .Z(g6868) ) ;
AND2    gate4523  (.A(g2214), .B(g5897), .Z(g6747) ) ;
INV     gate4524  (.A(g6747), .Z(II10949) ) ;
INV     gate4525  (.A(II10949), .Z(g6869) ) ;
INV     gate4526  (.A(g6556), .Z(II10952) ) ;
INV     gate4527  (.A(II10952), .Z(g6870) ) ;
INV     gate4528  (.A(g6724), .Z(g6871) ) ;
INV     gate4529  (.A(g6559), .Z(II10958) ) ;
INV     gate4530  (.A(II10958), .Z(g6874) ) ;
INV     gate4531  (.A(g6793), .Z(II10963) ) ;
INV     gate4532  (.A(II10963), .Z(g6877) ) ;
INV     gate4533  (.A(g6561), .Z(II10966) ) ;
INV     gate4534  (.A(II10966), .Z(g6878) ) ;
INV     gate4535  (.A(g6344), .Z(II10971) ) ;
INV     gate4536  (.A(II10971), .Z(g6881) ) ;
INV     gate4537  (.A(g6563), .Z(II10974) ) ;
INV     gate4538  (.A(II10974), .Z(g6882) ) ;
INV     gate4539  (.A(g6565), .Z(II10979) ) ;
INV     gate4540  (.A(II10979), .Z(g6885) ) ;
AND2    gate4541  (.A(g2221), .B(g5919), .Z(g6757) ) ;
INV     gate4542  (.A(g6757), .Z(II10984) ) ;
INV     gate4543  (.A(II10984), .Z(g6888) ) ;
AND2    gate4544  (.A(g148), .B(g5919), .Z(g6759) ) ;
INV     gate4545  (.A(g6759), .Z(II10991) ) ;
INV     gate4546  (.A(II10991), .Z(g6893) ) ;
AND2    gate4547  (.A(g178), .B(g5919), .Z(g6786) ) ;
INV     gate4548  (.A(g6786), .Z(II10996) ) ;
INV     gate4549  (.A(II10996), .Z(g6896) ) ;
INV     gate4550  (.A(g6386), .Z(II11005) ) ;
INV     gate4551  (.A(II11005), .Z(g6903) ) ;
AND2    gate4552  (.A(g5036), .B(g5878), .Z(g6795) ) ;
INV     gate4553  (.A(g6795), .Z(II11008) ) ;
INV     gate4554  (.A(II11008), .Z(g6904) ) ;
INV     gate4555  (.A(g6340), .Z(II11011) ) ;
INV     gate4556  (.A(II11011), .Z(g6905) ) ;
INV     gate4557  (.A(g6398), .Z(II11021) ) ;
INV     gate4558  (.A(II11021), .Z(g6913) ) ;
INV     gate4559  (.A(g6399), .Z(II11024) ) ;
INV     gate4560  (.A(II11024), .Z(g6914) ) ;
OR2     gate4561  (.A(g5848), .B(g5067), .Z(g6485) ) ;
INV     gate4562  (.A(g6485), .Z(II11029) ) ;
INV     gate4563  (.A(II11029), .Z(g6917) ) ;
INV     gate4564  (.A(g6453), .Z(g6919) ) ;
INV     gate4565  (.A(g6629), .Z(II11034) ) ;
INV     gate4566  (.A(g6629), .Z(II11037) ) ;
INV     gate4567  (.A(II11037), .Z(g6921) ) ;
INV     gate4568  (.A(g6412), .Z(II11043) ) ;
INV     gate4569  (.A(II11043), .Z(g6925) ) ;
INV     gate4570  (.A(g6635), .Z(II11046) ) ;
INV     gate4571  (.A(g6635), .Z(II11049) ) ;
INV     gate4572  (.A(II11049), .Z(g6927) ) ;
INV     gate4573  (.A(g6419), .Z(II11055) ) ;
INV     gate4574  (.A(II11055), .Z(g6931) ) ;
INV     gate4575  (.A(g6641), .Z(II11058) ) ;
INV     gate4576  (.A(g6641), .Z(II11061) ) ;
INV     gate4577  (.A(II11061), .Z(g6933) ) ;
INV     gate4578  (.A(g6750), .Z(II11065) ) ;
INV     gate4579  (.A(II11065), .Z(g6935) ) ;
INV     gate4580  (.A(g6426), .Z(II11068) ) ;
INV     gate4581  (.A(II11068), .Z(g6938) ) ;
AND3    gate4582  (.A(g2733), .B(g6061), .C(g4631), .Z(g6656) ) ;
INV     gate4583  (.A(g6656), .Z(II11071) ) ;
INV     gate4584  (.A(II11071), .Z(g6939) ) ;
INV     gate4585  (.A(g6503), .Z(g6941) ) ;
INV     gate4586  (.A(g6649), .Z(II11076) ) ;
INV     gate4587  (.A(g6649), .Z(II11079) ) ;
INV     gate4588  (.A(II11079), .Z(g6943) ) ;
INV     gate4589  (.A(g6749), .Z(II11082) ) ;
INV     gate4590  (.A(II11082), .Z(g6944) ) ;
INV     gate4591  (.A(g6433), .Z(II11085) ) ;
INV     gate4592  (.A(II11085), .Z(g6947) ) ;
INV     gate4593  (.A(g6434), .Z(II11088) ) ;
INV     gate4594  (.A(II11088), .Z(g6948) ) ;
INV     gate4595  (.A(g6657), .Z(II11091) ) ;
INV     gate4596  (.A(g6657), .Z(II11094) ) ;
INV     gate4597  (.A(II11094), .Z(g6950) ) ;
INV     gate4598  (.A(g6748), .Z(II11097) ) ;
INV     gate4599  (.A(II11097), .Z(g6951) ) ;
INV     gate4600  (.A(g6442), .Z(II11100) ) ;
INV     gate4601  (.A(II11100), .Z(g6954) ) ;
INV     gate4602  (.A(g6667), .Z(II11103) ) ;
INV     gate4603  (.A(g6667), .Z(II11106) ) ;
INV     gate4604  (.A(II11106), .Z(g6956) ) ;
INV     gate4605  (.A(g6464), .Z(II11109) ) ;
INV     gate4606  (.A(II11109), .Z(g6957) ) ;
INV     gate4607  (.A(g6445), .Z(II11112) ) ;
INV     gate4608  (.A(II11112), .Z(g6960) ) ;
INV     gate4609  (.A(g6462), .Z(II11115) ) ;
INV     gate4610  (.A(II11115), .Z(g6961) ) ;
INV     gate4611  (.A(g6509), .Z(g6964) ) ;
INV     gate4612  (.A(g6461), .Z(II11119) ) ;
INV     gate4613  (.A(II11119), .Z(g6967) ) ;
INV     gate4614  (.A(g6450), .Z(II11122) ) ;
INV     gate4615  (.A(II11122), .Z(g6970) ) ;
INV     gate4616  (.A(g6517), .Z(g6971) ) ;
INV     gate4617  (.A(g6365), .Z(g6974) ) ;
INV     gate4618  (.A(g6452), .Z(II11127) ) ;
INV     gate4619  (.A(II11127), .Z(g6980) ) ;
INV     gate4620  (.A(g6382), .Z(g6984) ) ;
INV     gate4621  (.A(g6451), .Z(II11132) ) ;
INV     gate4622  (.A(II11132), .Z(g6990) ) ;
AND3    gate4623  (.A(g4631), .B(g6074), .C(g2733), .Z(g6679) ) ;
INV     gate4624  (.A(g6679), .Z(II11135) ) ;
INV     gate4625  (.A(II11135), .Z(g6993) ) ;
INV     gate4626  (.A(g6482), .Z(g6995) ) ;
INV     gate4627  (.A(g6448), .Z(II11140) ) ;
INV     gate4628  (.A(II11140), .Z(g7001) ) ;
INV     gate4629  (.A(g6446), .Z(II11143) ) ;
INV     gate4630  (.A(II11143), .Z(g7004) ) ;
AND2    gate4631  (.A(g4479), .B(g5919), .Z(g6439) ) ;
INV     gate4632  (.A(g6439), .Z(II11146) ) ;
INV     gate4633  (.A(II11146), .Z(g7007) ) ;
OR2     gate4634  (.A(g5690), .B(g4950), .Z(g6468) ) ;
INV     gate4635  (.A(g6468), .Z(II11149) ) ;
INV     gate4636  (.A(II11149), .Z(g7008) ) ;
OR2     gate4637  (.A(g5698), .B(g4959), .Z(g6469) ) ;
INV     gate4638  (.A(g6469), .Z(II11152) ) ;
INV     gate4639  (.A(II11152), .Z(g7009) ) ;
OR2     gate4640  (.A(g5699), .B(g4960), .Z(g6470) ) ;
INV     gate4641  (.A(g6470), .Z(II11155) ) ;
INV     gate4642  (.A(II11155), .Z(g7010) ) ;
INV     gate4643  (.A(g6503), .Z(g7011) ) ;
OR2     gate4644  (.A(g5706), .B(g4967), .Z(g6478) ) ;
INV     gate4645  (.A(g6478), .Z(II11159) ) ;
INV     gate4646  (.A(II11159), .Z(g7020) ) ;
OR2     gate4647  (.A(g5707), .B(g4968), .Z(g6479) ) ;
INV     gate4648  (.A(g6479), .Z(II11162) ) ;
INV     gate4649  (.A(II11162), .Z(g7021) ) ;
INV     gate4650  (.A(g6389), .Z(g7022) ) ;
OR2     gate4651  (.A(g5721), .B(g4971), .Z(g6480) ) ;
INV     gate4652  (.A(g6480), .Z(II11166) ) ;
INV     gate4653  (.A(II11166), .Z(g7023) ) ;
OR2     gate4654  (.A(g5722), .B(g4972), .Z(g6481) ) ;
INV     gate4655  (.A(g6481), .Z(II11169) ) ;
INV     gate4656  (.A(II11169), .Z(g7024) ) ;
INV     gate4657  (.A(g6400), .Z(g7025) ) ;
OR2     gate4658  (.A(g5725), .B(g4986), .Z(g6500) ) ;
INV     gate4659  (.A(g6500), .Z(II11173) ) ;
INV     gate4660  (.A(II11173), .Z(g7026) ) ;
OR2     gate4661  (.A(g5726), .B(g4987), .Z(g6501) ) ;
INV     gate4662  (.A(g6501), .Z(II11176) ) ;
INV     gate4663  (.A(II11176), .Z(g7027) ) ;
INV     gate4664  (.A(g6407), .Z(g7028) ) ;
OR2     gate4665  (.A(g5731), .B(g4989), .Z(g6506) ) ;
INV     gate4666  (.A(g6506), .Z(II11180) ) ;
INV     gate4667  (.A(II11180), .Z(g7029) ) ;
OR2     gate4668  (.A(g5732), .B(g4990), .Z(g6507) ) ;
INV     gate4669  (.A(g6507), .Z(II11183) ) ;
INV     gate4670  (.A(II11183), .Z(g7030) ) ;
INV     gate4671  (.A(g6413), .Z(g7031) ) ;
OR2     gate4672  (.A(g5737), .B(g4991), .Z(g6513) ) ;
INV     gate4673  (.A(g6513), .Z(II11188) ) ;
INV     gate4674  (.A(II11188), .Z(g7033) ) ;
OR2     gate4675  (.A(g5738), .B(g4992), .Z(g6514) ) ;
INV     gate4676  (.A(g6514), .Z(II11191) ) ;
INV     gate4677  (.A(II11191), .Z(g7034) ) ;
OR2     gate4678  (.A(g5739), .B(g4993), .Z(g6515) ) ;
INV     gate4679  (.A(g6515), .Z(II11194) ) ;
INV     gate4680  (.A(II11194), .Z(g7035) ) ;
INV     gate4681  (.A(g6420), .Z(g7036) ) ;
INV     gate4682  (.A(g6521), .Z(II11198) ) ;
INV     gate4683  (.A(II11198), .Z(g7037) ) ;
OR2     gate4684  (.A(g5744), .B(g4994), .Z(g6522) ) ;
INV     gate4685  (.A(g6522), .Z(II11201) ) ;
INV     gate4686  (.A(II11201), .Z(g7038) ) ;
OR2     gate4687  (.A(g5745), .B(g4995), .Z(g6523) ) ;
INV     gate4688  (.A(g6523), .Z(II11204) ) ;
INV     gate4689  (.A(II11204), .Z(g7039) ) ;
OR2     gate4690  (.A(g5746), .B(g4996), .Z(g6524) ) ;
INV     gate4691  (.A(g6524), .Z(II11207) ) ;
INV     gate4692  (.A(II11207), .Z(g7040) ) ;
INV     gate4693  (.A(g6427), .Z(g7041) ) ;
INV     gate4694  (.A(g6527), .Z(II11211) ) ;
INV     gate4695  (.A(II11211), .Z(g7042) ) ;
OR2     gate4696  (.A(g5756), .B(g4999), .Z(g6528) ) ;
INV     gate4697  (.A(g6528), .Z(II11214) ) ;
INV     gate4698  (.A(II11214), .Z(g7043) ) ;
OR2     gate4699  (.A(g5757), .B(g5000), .Z(g6529) ) ;
INV     gate4700  (.A(g6529), .Z(II11217) ) ;
INV     gate4701  (.A(II11217), .Z(g7044) ) ;
INV     gate4702  (.A(g6435), .Z(g7045) ) ;
OR2     gate4703  (.A(g5771), .B(g5002), .Z(g6533) ) ;
INV     gate4704  (.A(g6533), .Z(II11222) ) ;
INV     gate4705  (.A(II11222), .Z(g7047) ) ;
OR2     gate4706  (.A(g5772), .B(g5003), .Z(g6534) ) ;
INV     gate4707  (.A(g6534), .Z(II11225) ) ;
INV     gate4708  (.A(II11225), .Z(g7048) ) ;
AND2    gate4709  (.A(g5224), .B(g6014), .Z(g6471) ) ;
INV     gate4710  (.A(g6471), .Z(II11228) ) ;
INV     gate4711  (.A(II11228), .Z(g7049) ) ;
OR2     gate4712  (.A(g5781), .B(g5005), .Z(g6537) ) ;
INV     gate4713  (.A(g6537), .Z(II11232) ) ;
INV     gate4714  (.A(II11232), .Z(g7051) ) ;
OR2     gate4715  (.A(g5782), .B(g5006), .Z(g6538) ) ;
INV     gate4716  (.A(g6538), .Z(II11235) ) ;
INV     gate4717  (.A(II11235), .Z(g7052) ) ;
INV     gate4718  (.A(g6543), .Z(II11238) ) ;
INV     gate4719  (.A(II11238), .Z(g7053) ) ;
OR2     gate4720  (.A(g5788), .B(g5009), .Z(g6541) ) ;
INV     gate4721  (.A(g6541), .Z(II11249) ) ;
INV     gate4722  (.A(II11249), .Z(g7056) ) ;
OR2     gate4723  (.A(g5789), .B(g5010), .Z(g6542) ) ;
INV     gate4724  (.A(g6542), .Z(II11252) ) ;
INV     gate4725  (.A(II11252), .Z(g7057) ) ;
INV     gate4726  (.A(g6547), .Z(II11255) ) ;
INV     gate4727  (.A(II11255), .Z(g7058) ) ;
OR2     gate4728  (.A(g5795), .B(g5025), .Z(g6545) ) ;
INV     gate4729  (.A(g6545), .Z(II11269) ) ;
INV     gate4730  (.A(II11269), .Z(g7064) ) ;
OR2     gate4731  (.A(g5796), .B(g5026), .Z(g6546) ) ;
INV     gate4732  (.A(g6546), .Z(II11272) ) ;
INV     gate4733  (.A(II11272), .Z(g7065) ) ;
AND2    gate4734  (.A(g5981), .B(g3095), .Z(g6502) ) ;
INV     gate4735  (.A(g6502), .Z(II11275) ) ;
INV     gate4736  (.A(II11275), .Z(g7066) ) ;
OR2     gate4737  (.A(g5804), .B(g5031), .Z(g6551) ) ;
INV     gate4738  (.A(g6551), .Z(II11286) ) ;
INV     gate4739  (.A(II11286), .Z(g7069) ) ;
AND2    gate4740  (.A(g5983), .B(g3096), .Z(g6508) ) ;
INV     gate4741  (.A(g6508), .Z(II11289) ) ;
INV     gate4742  (.A(II11289), .Z(g7070) ) ;
AND2    gate4743  (.A(g5993), .B(g3097), .Z(g6516) ) ;
INV     gate4744  (.A(g6516), .Z(II11293) ) ;
INV     gate4745  (.A(II11293), .Z(g7072) ) ;
AND2    gate4746  (.A(g5995), .B(g3102), .Z(g6525) ) ;
INV     gate4747  (.A(g6525), .Z(II11296) ) ;
INV     gate4748  (.A(II11296), .Z(g7073) ) ;
INV     gate4749  (.A(g6727), .Z(II11299) ) ;
INV     gate4750  (.A(II11299), .Z(g7074) ) ;
AND2    gate4751  (.A(g76), .B(g6052), .Z(g6526) ) ;
INV     gate4752  (.A(g6526), .Z(II11303) ) ;
INV     gate4753  (.A(II11303), .Z(g7076) ) ;
INV     gate4754  (.A(g6731), .Z(II11306) ) ;
INV     gate4755  (.A(II11306), .Z(g7077) ) ;
AND2    gate4756  (.A(g79), .B(g6056), .Z(g6531) ) ;
INV     gate4757  (.A(g6531), .Z(II11309) ) ;
INV     gate4758  (.A(II11309), .Z(g7078) ) ;
NAND2   gate4759  (.A(g6027), .B(g6019), .Z(g6488) ) ;
INV     gate4760  (.A(g6488), .Z(II11312) ) ;
INV     gate4761  (.A(II11312), .Z(g7079) ) ;
INV     gate4762  (.A(g6644), .Z(II11315) ) ;
INV     gate4763  (.A(II11315), .Z(g7082) ) ;
INV     gate4764  (.A(g6488), .Z(II11318) ) ;
INV     gate4765  (.A(II11318), .Z(g7085) ) ;
INV     gate4766  (.A(g6652), .Z(II11322) ) ;
INV     gate4767  (.A(II11322), .Z(g7089) ) ;
INV     gate4768  (.A(g6660), .Z(II11326) ) ;
INV     gate4769  (.A(II11326), .Z(g7093) ) ;
INV     gate4770  (.A(g6571), .Z(II11330) ) ;
INV     gate4771  (.A(II11330), .Z(g7097) ) ;
INV     gate4772  (.A(g6670), .Z(II11333) ) ;
INV     gate4773  (.A(II11333), .Z(g7098) ) ;
INV     gate4774  (.A(g6680), .Z(II11338) ) ;
INV     gate4775  (.A(II11338), .Z(g7103) ) ;
INV     gate4776  (.A(g6686), .Z(II11342) ) ;
INV     gate4777  (.A(II11342), .Z(g7107) ) ;
INV     gate4778  (.A(g6692), .Z(II11345) ) ;
INV     gate4779  (.A(II11345), .Z(g7110) ) ;
INV     gate4780  (.A(g6695), .Z(II11348) ) ;
INV     gate4781  (.A(II11348), .Z(g7113) ) ;
INV     gate4782  (.A(g6698), .Z(II11351) ) ;
INV     gate4783  (.A(II11351), .Z(g7116) ) ;
INV     gate4784  (.A(g6553), .Z(II11354) ) ;
INV     gate4785  (.A(II11354), .Z(g7119) ) ;
INV     gate4786  (.A(g6594), .Z(II11357) ) ;
INV     gate4787  (.A(II11357), .Z(g7122) ) ;
AND2    gate4788  (.A(g6210), .B(g5052), .Z(g6351) ) ;
INV     gate4789  (.A(g6351), .Z(II11360) ) ;
INV     gate4790  (.A(II11360), .Z(g7123) ) ;
INV     gate4791  (.A(g6595), .Z(II11363) ) ;
INV     gate4792  (.A(II11363), .Z(g7124) ) ;
NOR2    gate4793  (.A(g5859), .B(g5938), .Z(g6392) ) ;
INV     gate4794  (.A(g6392), .Z(II11367) ) ;
INV     gate4795  (.A(II11367), .Z(g7126) ) ;
INV     gate4796  (.A(g6385), .Z(II11383) ) ;
INV     gate4797  (.A(II11383), .Z(g7142) ) ;
OR2     gate4798  (.A(g5941), .B(g5259), .Z(g6672) ) ;
INV     gate4799  (.A(g6672), .Z(II11387) ) ;
INV     gate4800  (.A(II11387), .Z(g7144) ) ;
INV     gate4801  (.A(g6387), .Z(II11391) ) ;
INV     gate4802  (.A(II11391), .Z(g7146) ) ;
AND2    gate4803  (.A(g52), .B(g6164), .Z(g6621) ) ;
INV     gate4804  (.A(g6621), .Z(II11394) ) ;
INV     gate4805  (.A(II11394), .Z(g7147) ) ;
INV     gate4806  (.A(g6713), .Z(II11397) ) ;
INV     gate4807  (.A(II11397), .Z(g7148) ) ;
AND2    gate4808  (.A(g58), .B(g6181), .Z(g6627) ) ;
INV     gate4809  (.A(g6627), .Z(II11405) ) ;
INV     gate4810  (.A(II11405), .Z(g7187) ) ;
INV     gate4811  (.A(g6405), .Z(II11408) ) ;
INV     gate4812  (.A(II11408), .Z(g7188) ) ;
INV     gate4813  (.A(g6411), .Z(II11412) ) ;
INV     gate4814  (.A(II11412), .Z(g7190) ) ;
INV     gate4815  (.A(g6742), .Z(g7192) ) ;
AND2    gate4816  (.A(g64), .B(g6195), .Z(g6638) ) ;
INV     gate4817  (.A(g6638), .Z(II11417) ) ;
INV     gate4818  (.A(II11417), .Z(g7195) ) ;
INV     gate4819  (.A(g6417), .Z(II11420) ) ;
INV     gate4820  (.A(II11420), .Z(g7196) ) ;
INV     gate4821  (.A(g6488), .Z(II11423) ) ;
INV     gate4822  (.A(II11423), .Z(g7197) ) ;
NAND2   gate4823  (.A(II10508), .B(II10509), .Z(g6573) ) ;
INV     gate4824  (.A(g6573), .Z(II11427) ) ;
INV     gate4825  (.A(II11427), .Z(g7201) ) ;
INV     gate4826  (.A(g6424), .Z(II11433) ) ;
INV     gate4827  (.A(II11433), .Z(g7205) ) ;
INV     gate4828  (.A(g6488), .Z(II11436) ) ;
INV     gate4829  (.A(II11436), .Z(g7206) ) ;
NAND2   gate4830  (.A(II10520), .B(II10521), .Z(g6577) ) ;
INV     gate4831  (.A(g6577), .Z(II11440) ) ;
INV     gate4832  (.A(II11440), .Z(g7210) ) ;
AND2    gate4833  (.A(g70), .B(g6213), .Z(g6653) ) ;
INV     gate4834  (.A(g6653), .Z(II11444) ) ;
INV     gate4835  (.A(II11444), .Z(g7212) ) ;
INV     gate4836  (.A(g6431), .Z(II11447) ) ;
INV     gate4837  (.A(II11447), .Z(g7213) ) ;
INV     gate4838  (.A(g6488), .Z(II11450) ) ;
INV     gate4839  (.A(II11450), .Z(g7214) ) ;
INV     gate4840  (.A(g6440), .Z(II11456) ) ;
INV     gate4841  (.A(II11456), .Z(g7220) ) ;
INV     gate4842  (.A(g6488), .Z(II11459) ) ;
INV     gate4843  (.A(II11459), .Z(g7221) ) ;
INV     gate4844  (.A(g6443), .Z(II11464) ) ;
INV     gate4845  (.A(II11464), .Z(g7226) ) ;
INV     gate4846  (.A(g6488), .Z(II11467) ) ;
INV     gate4847  (.A(II11467), .Z(g7227) ) ;
INV     gate4848  (.A(g6488), .Z(II11472) ) ;
INV     gate4849  (.A(II11472), .Z(g7232) ) ;
INV     gate4850  (.A(g6488), .Z(II11477) ) ;
INV     gate4851  (.A(II11477), .Z(g7237) ) ;
INV     gate4852  (.A(g6567), .Z(II11483) ) ;
INV     gate4853  (.A(II11483), .Z(g7243) ) ;
INV     gate4854  (.A(g6569), .Z(II11489) ) ;
INV     gate4855  (.A(II11489), .Z(g7256) ) ;
INV     gate4856  (.A(g6574), .Z(II11494) ) ;
INV     gate4857  (.A(II11494), .Z(g7259) ) ;
INV     gate4858  (.A(g6578), .Z(II11498) ) ;
INV     gate4859  (.A(II11498), .Z(g7263) ) ;
INV     gate4860  (.A(g6581), .Z(II11501) ) ;
INV     gate4861  (.A(II11501), .Z(g7264) ) ;
INV     gate4862  (.A(g6585), .Z(II11505) ) ;
INV     gate4863  (.A(II11505), .Z(g7268) ) ;
INV     gate4864  (.A(g6589), .Z(II11515) ) ;
INV     gate4865  (.A(II11515), .Z(g7270) ) ;
INV     gate4866  (.A(g6591), .Z(II11519) ) ;
INV     gate4867  (.A(II11519), .Z(g7272) ) ;
INV     gate4868  (.A(g6365), .Z(g7273) ) ;
INV     gate4869  (.A(g6593), .Z(II11524) ) ;
INV     gate4870  (.A(II11524), .Z(g7278) ) ;
INV     gate4871  (.A(g6382), .Z(g7279) ) ;
INV     gate4872  (.A(g6796), .Z(II11528) ) ;
INV     gate4873  (.A(II11528), .Z(g7284) ) ;
INV     gate4874  (.A(g7126), .Z(II11531) ) ;
INV     gate4875  (.A(g6917), .Z(II11534) ) ;
INV     gate4876  (.A(II11534), .Z(g7286) ) ;
INV     gate4877  (.A(g7144), .Z(II11537) ) ;
INV     gate4878  (.A(g6877), .Z(II11540) ) ;
INV     gate4879  (.A(g6881), .Z(II11543) ) ;
INV     gate4880  (.A(g7037), .Z(II11560) ) ;
AND2    gate4881  (.A(g243), .B(g6596), .Z(g6819) ) ;
INV     gate4882  (.A(g6819), .Z(II11563) ) ;
AND2    gate4883  (.A(g1362), .B(g6596), .Z(g6820) ) ;
INV     gate4884  (.A(g6820), .Z(II11566) ) ;
AND2    gate4885  (.A(g237), .B(g6596), .Z(g6821) ) ;
INV     gate4886  (.A(g6821), .Z(II11569) ) ;
AND2    gate4887  (.A(g231), .B(g6596), .Z(g6822) ) ;
INV     gate4888  (.A(g6822), .Z(II11572) ) ;
AND2    gate4889  (.A(g1368), .B(g6596), .Z(g6823) ) ;
INV     gate4890  (.A(g6823), .Z(II11575) ) ;
AND2    gate4891  (.A(g1371), .B(g6596), .Z(g6824) ) ;
INV     gate4892  (.A(g6824), .Z(II11578) ) ;
AND2    gate4893  (.A(g225), .B(g6596), .Z(g6826) ) ;
INV     gate4894  (.A(g6826), .Z(II11581) ) ;
AND2    gate4895  (.A(g219), .B(g6596), .Z(g6827) ) ;
INV     gate4896  (.A(g6827), .Z(II11584) ) ;
AND2    gate4897  (.A(g1377), .B(g6596), .Z(g6828) ) ;
INV     gate4898  (.A(g6828), .Z(II11587) ) ;
AND2    gate4899  (.A(g213), .B(g6596), .Z(g6829) ) ;
INV     gate4900  (.A(g6829), .Z(II11590) ) ;
AND2    gate4901  (.A(g1380), .B(g6596), .Z(g6830) ) ;
INV     gate4902  (.A(g6830), .Z(II11593) ) ;
AND2    gate4903  (.A(g207), .B(g6596), .Z(g6831) ) ;
INV     gate4904  (.A(g6831), .Z(II11596) ) ;
AND2    gate4905  (.A(g1383), .B(g6596), .Z(g6832) ) ;
INV     gate4906  (.A(g6832), .Z(II11599) ) ;
AND2    gate4907  (.A(g186), .B(g6596), .Z(g6833) ) ;
INV     gate4908  (.A(g6833), .Z(II11602) ) ;
AND2    gate4909  (.A(g1365), .B(g6596), .Z(g6834) ) ;
INV     gate4910  (.A(g6834), .Z(II11605) ) ;
INV     gate4911  (.A(g6903), .Z(II11608) ) ;
INV     gate4912  (.A(g6913), .Z(II11611) ) ;
AND2    gate4913  (.A(g192), .B(g6596), .Z(g6838) ) ;
INV     gate4914  (.A(g6838), .Z(II11614) ) ;
AND2    gate4915  (.A(g1397), .B(g6596), .Z(g6839) ) ;
INV     gate4916  (.A(g6839), .Z(II11617) ) ;
AND2    gate4917  (.A(g248), .B(g6596), .Z(g6840) ) ;
INV     gate4918  (.A(g6840), .Z(II11620) ) ;
AND2    gate4919  (.A(g1400), .B(g6596), .Z(g6841) ) ;
INV     gate4920  (.A(g6841), .Z(II11623) ) ;
INV     gate4921  (.A(g7042), .Z(II11626) ) ;
INV     gate4922  (.A(g6914), .Z(II11629) ) ;
INV     gate4923  (.A(g6931), .Z(II11632) ) ;
INV     gate4924  (.A(g6947), .Z(II11635) ) ;
INV     gate4925  (.A(g6948), .Z(II11638) ) ;
INV     gate4926  (.A(g6960), .Z(II11641) ) ;
INV     gate4927  (.A(g6970), .Z(II11644) ) ;
INV     gate4928  (.A(g6925), .Z(II11647) ) ;
INV     gate4929  (.A(g6938), .Z(II11650) ) ;
INV     gate4930  (.A(g6954), .Z(II11653) ) ;
INV     gate4931  (.A(g7122), .Z(II11656) ) ;
INV     gate4932  (.A(g7097), .Z(II11659) ) ;
INV     gate4933  (.A(g7033), .Z(II11662) ) ;
INV     gate4934  (.A(g7038), .Z(II11665) ) ;
INV     gate4935  (.A(g7043), .Z(II11668) ) ;
INV     gate4936  (.A(g7047), .Z(II11671) ) ;
INV     gate4937  (.A(g7051), .Z(II11674) ) ;
INV     gate4938  (.A(g7056), .Z(II11677) ) ;
INV     gate4939  (.A(g7064), .Z(II11680) ) ;
INV     gate4940  (.A(g7069), .Z(II11683) ) ;
INV     gate4941  (.A(g7039), .Z(II11686) ) ;
INV     gate4942  (.A(g7044), .Z(II11689) ) ;
INV     gate4943  (.A(g7048), .Z(II11692) ) ;
INV     gate4944  (.A(g7052), .Z(II11695) ) ;
INV     gate4945  (.A(g7057), .Z(II11698) ) ;
INV     gate4946  (.A(g7065), .Z(II11701) ) ;
INV     gate4947  (.A(g7008), .Z(II11704) ) ;
INV     gate4948  (.A(g7009), .Z(II11707) ) ;
INV     gate4949  (.A(g7020), .Z(II11710) ) ;
INV     gate4950  (.A(g7023), .Z(II11713) ) ;
INV     gate4951  (.A(g7026), .Z(II11716) ) ;
INV     gate4952  (.A(g7029), .Z(II11719) ) ;
INV     gate4953  (.A(g7034), .Z(II11722) ) ;
INV     gate4954  (.A(g7040), .Z(II11725) ) ;
INV     gate4955  (.A(g7010), .Z(II11728) ) ;
INV     gate4956  (.A(g7021), .Z(II11731) ) ;
INV     gate4957  (.A(g7024), .Z(II11734) ) ;
INV     gate4958  (.A(g7027), .Z(II11737) ) ;
INV     gate4959  (.A(g7030), .Z(II11740) ) ;
INV     gate4960  (.A(g7035), .Z(II11743) ) ;
INV     gate4961  (.A(g6857), .Z(II11746) ) ;
INV     gate4962  (.A(g7273), .Z(g7369) ) ;
AND3    gate4963  (.A(g2965), .B(g6626), .C(g5292), .Z(g7032) ) ;
INV     gate4964  (.A(g7032), .Z(II11752) ) ;
INV     gate4965  (.A(II11752), .Z(g7374) ) ;
AND2    gate4966  (.A(g6343), .B(g4323), .Z(g7191) ) ;
INV     gate4967  (.A(g7191), .Z(II11756) ) ;
INV     gate4968  (.A(II11756), .Z(g7376) ) ;
OR2     gate4969  (.A(g6699), .B(g4720), .Z(g7244) ) ;
INV     gate4970  (.A(g7244), .Z(II11759) ) ;
INV     gate4971  (.A(II11759), .Z(g7377) ) ;
INV     gate4972  (.A(g6863), .Z(g7379) ) ;
INV     gate4973  (.A(g7279), .Z(g7380) ) ;
INV     gate4974  (.A(g7201), .Z(II11767) ) ;
INV     gate4975  (.A(II11767), .Z(g7386) ) ;
AND2    gate4976  (.A(g6349), .B(g4329), .Z(g7202) ) ;
INV     gate4977  (.A(g7202), .Z(II11770) ) ;
INV     gate4978  (.A(II11770), .Z(g7387) ) ;
OR2     gate4979  (.A(g6701), .B(g4725), .Z(g7257) ) ;
INV     gate4980  (.A(g7257), .Z(II11773) ) ;
INV     gate4981  (.A(II11773), .Z(g7388) ) ;
INV     gate4982  (.A(g6847), .Z(g7390) ) ;
INV     gate4983  (.A(g7210), .Z(II11778) ) ;
INV     gate4984  (.A(II11778), .Z(g7394) ) ;
INV     gate4985  (.A(g6941), .Z(g7395) ) ;
INV     gate4986  (.A(g6860), .Z(g7402) ) ;
OR2     gate4987  (.A(g6465), .B(g6003), .Z(g7246) ) ;
INV     gate4988  (.A(g7246), .Z(II11783) ) ;
INV     gate4989  (.A(II11783), .Z(g7403) ) ;
INV     gate4990  (.A(g7246), .Z(II11786) ) ;
INV     gate4991  (.A(II11786), .Z(g7406) ) ;
INV     gate4992  (.A(g7246), .Z(II11790) ) ;
INV     gate4993  (.A(II11790), .Z(g7410) ) ;
INV     gate4994  (.A(g7197), .Z(g7413) ) ;
INV     gate4995  (.A(g7188), .Z(II11794) ) ;
INV     gate4996  (.A(II11794), .Z(g7414) ) ;
INV     gate4997  (.A(g6852), .Z(II11797) ) ;
INV     gate4998  (.A(II11797), .Z(g7415) ) ;
INV     gate4999  (.A(g7246), .Z(II11800) ) ;
INV     gate5000  (.A(II11800), .Z(g7416) ) ;
INV     gate5001  (.A(g7206), .Z(g7419) ) ;
INV     gate5002  (.A(g7190), .Z(II11804) ) ;
INV     gate5003  (.A(II11804), .Z(g7420) ) ;
INV     gate5004  (.A(g6854), .Z(II11807) ) ;
INV     gate5005  (.A(II11807), .Z(g7421) ) ;
INV     gate5006  (.A(g7246), .Z(II11810) ) ;
INV     gate5007  (.A(II11810), .Z(g7422) ) ;
INV     gate5008  (.A(g7214), .Z(g7425) ) ;
INV     gate5009  (.A(g7196), .Z(II11814) ) ;
INV     gate5010  (.A(II11814), .Z(g7426) ) ;
INV     gate5011  (.A(g7246), .Z(II11817) ) ;
INV     gate5012  (.A(II11817), .Z(g7427) ) ;
INV     gate5013  (.A(g7221), .Z(g7430) ) ;
INV     gate5014  (.A(g7205), .Z(II11821) ) ;
INV     gate5015  (.A(II11821), .Z(g7431) ) ;
INV     gate5016  (.A(g7246), .Z(II11824) ) ;
INV     gate5017  (.A(II11824), .Z(g7432) ) ;
INV     gate5018  (.A(g7227), .Z(g7436) ) ;
INV     gate5019  (.A(g7213), .Z(II11829) ) ;
INV     gate5020  (.A(II11829), .Z(g7437) ) ;
INV     gate5021  (.A(g7232), .Z(g7438) ) ;
INV     gate5022  (.A(g7077), .Z(II11833) ) ;
INV     gate5023  (.A(II11833), .Z(g7439) ) ;
INV     gate5024  (.A(g7220), .Z(II11836) ) ;
INV     gate5025  (.A(II11836), .Z(g7440) ) ;
INV     gate5026  (.A(g7237), .Z(g7442) ) ;
INV     gate5027  (.A(g7226), .Z(II11841) ) ;
INV     gate5028  (.A(II11841), .Z(g7443) ) ;
INV     gate5029  (.A(g6869), .Z(II11845) ) ;
INV     gate5030  (.A(II11845), .Z(g7445) ) ;
INV     gate5031  (.A(g7148), .Z(g7446) ) ;
INV     gate5032  (.A(g7148), .Z(g7450) ) ;
INV     gate5033  (.A(g7148), .Z(g7454) ) ;
INV     gate5034  (.A(g7123), .Z(g7458) ) ;
INV     gate5035  (.A(g7148), .Z(g7460) ) ;
INV     gate5036  (.A(g6921), .Z(g7463) ) ;
INV     gate5037  (.A(g6888), .Z(II11858) ) ;
INV     gate5038  (.A(II11858), .Z(g7464) ) ;
INV     gate5039  (.A(g7148), .Z(g7467) ) ;
INV     gate5040  (.A(g6927), .Z(g7470) ) ;
INV     gate5041  (.A(g7148), .Z(g7473) ) ;
INV     gate5042  (.A(g6933), .Z(g7476) ) ;
OR2     gate5043  (.A(g6763), .B(g4868), .Z(g6894) ) ;
INV     gate5044  (.A(g6894), .Z(II11869) ) ;
INV     gate5045  (.A(II11869), .Z(g7477) ) ;
INV     gate5046  (.A(g6863), .Z(II11873) ) ;
INV     gate5047  (.A(II11873), .Z(g7479) ) ;
INV     gate5048  (.A(g7148), .Z(g7497) ) ;
INV     gate5049  (.A(g6943), .Z(g7500) ) ;
INV     gate5050  (.A(g6893), .Z(II11879) ) ;
INV     gate5051  (.A(II11879), .Z(g7501) ) ;
OR2     gate5052  (.A(g6776), .B(g4875), .Z(g6895) ) ;
INV     gate5053  (.A(g6895), .Z(II11882) ) ;
INV     gate5054  (.A(II11882), .Z(g7502) ) ;
INV     gate5055  (.A(g7148), .Z(g7505) ) ;
INV     gate5056  (.A(g6950), .Z(g7508) ) ;
OR2     gate5057  (.A(g6790), .B(g4881), .Z(g6898) ) ;
INV     gate5058  (.A(g6898), .Z(II11889) ) ;
INV     gate5059  (.A(II11889), .Z(g7509) ) ;
INV     gate5060  (.A(g7148), .Z(g7512) ) ;
INV     gate5061  (.A(g7148), .Z(g7516) ) ;
INV     gate5062  (.A(g6956), .Z(g7519) ) ;
INV     gate5063  (.A(g6896), .Z(II11898) ) ;
INV     gate5064  (.A(II11898), .Z(g7520) ) ;
OR2     gate5065  (.A(g6771), .B(g6240), .Z(g6897) ) ;
INV     gate5066  (.A(g6897), .Z(II11901) ) ;
INV     gate5067  (.A(II11901), .Z(g7521) ) ;
OR2     gate5068  (.A(g6794), .B(g4223), .Z(g6902) ) ;
INV     gate5069  (.A(g6902), .Z(II11904) ) ;
INV     gate5070  (.A(II11904), .Z(g7522) ) ;
INV     gate5071  (.A(g6904), .Z(II11921) ) ;
INV     gate5072  (.A(II11921), .Z(g7525) ) ;
INV     gate5073  (.A(g7148), .Z(g7527) ) ;
OR2     gate5074  (.A(g6787), .B(g6246), .Z(g6900) ) ;
INV     gate5075  (.A(g6900), .Z(II11926) ) ;
INV     gate5076  (.A(II11926), .Z(g7530) ) ;
OR2     gate5077  (.A(g6788), .B(g6247), .Z(g6901) ) ;
INV     gate5078  (.A(g6901), .Z(II11929) ) ;
INV     gate5079  (.A(II11929), .Z(g7531) ) ;
OR2     gate5080  (.A(g6345), .B(g4229), .Z(g6908) ) ;
INV     gate5081  (.A(g6908), .Z(II11932) ) ;
INV     gate5082  (.A(II11932), .Z(g7532) ) ;
OR2     gate5083  (.A(g6346), .B(g5684), .Z(g6909) ) ;
INV     gate5084  (.A(g6909), .Z(II11942) ) ;
INV     gate5085  (.A(II11942), .Z(g7534) ) ;
INV     gate5086  (.A(g6905), .Z(II11947) ) ;
INV     gate5087  (.A(II11947), .Z(g7537) ) ;
OR2     gate5088  (.A(g6791), .B(g5674), .Z(g6906) ) ;
INV     gate5089  (.A(g6906), .Z(II11950) ) ;
INV     gate5090  (.A(II11950), .Z(g7538) ) ;
OR2     gate5091  (.A(g6792), .B(g5675), .Z(g6907) ) ;
INV     gate5092  (.A(g6907), .Z(II11953) ) ;
INV     gate5093  (.A(II11953), .Z(g7539) ) ;
OR2     gate5094  (.A(g6350), .B(g4235), .Z(g6912) ) ;
INV     gate5095  (.A(g6912), .Z(II11956) ) ;
INV     gate5096  (.A(II11956), .Z(g7540) ) ;
INV     gate5097  (.A(g7053), .Z(II11961) ) ;
INV     gate5098  (.A(II11961), .Z(g7543) ) ;
OR2     gate5099  (.A(g6341), .B(g5680), .Z(g6910) ) ;
INV     gate5100  (.A(g6910), .Z(II11964) ) ;
INV     gate5101  (.A(II11964), .Z(g7544) ) ;
OR2     gate5102  (.A(g6342), .B(g5681), .Z(g6911) ) ;
INV     gate5103  (.A(g6911), .Z(II11967) ) ;
INV     gate5104  (.A(II11967), .Z(g7545) ) ;
OR2     gate5105  (.A(g6358), .B(g4252), .Z(g6918) ) ;
INV     gate5106  (.A(g6918), .Z(II11970) ) ;
INV     gate5107  (.A(II11970), .Z(g7546) ) ;
INV     gate5108  (.A(g6974), .Z(g7550) ) ;
INV     gate5109  (.A(g6919), .Z(II11989) ) ;
INV     gate5110  (.A(II11989), .Z(g7555) ) ;
INV     gate5111  (.A(g7058), .Z(II11992) ) ;
INV     gate5112  (.A(II11992), .Z(g7556) ) ;
OR2     gate5113  (.A(g6347), .B(g5686), .Z(g6915) ) ;
INV     gate5114  (.A(g6915), .Z(II12009) ) ;
INV     gate5115  (.A(II12009), .Z(g7559) ) ;
OR2     gate5116  (.A(g6348), .B(g5687), .Z(g6916) ) ;
INV     gate5117  (.A(g6916), .Z(II12012) ) ;
INV     gate5118  (.A(II12012), .Z(g7560) ) ;
OR2     gate5119  (.A(g6362), .B(g4261), .Z(g6924) ) ;
INV     gate5120  (.A(g6924), .Z(II12015) ) ;
INV     gate5121  (.A(II12015), .Z(g7561) ) ;
INV     gate5122  (.A(g6984), .Z(g7562) ) ;
INV     gate5123  (.A(g7119), .Z(II12026) ) ;
INV     gate5124  (.A(II12026), .Z(g7568) ) ;
OR2     gate5125  (.A(g6352), .B(g5694), .Z(g6922) ) ;
INV     gate5126  (.A(g6922), .Z(II12029) ) ;
INV     gate5127  (.A(II12029), .Z(g7569) ) ;
OR2     gate5128  (.A(g6353), .B(g5695), .Z(g6923) ) ;
INV     gate5129  (.A(g6923), .Z(II12032) ) ;
INV     gate5130  (.A(II12032), .Z(g7570) ) ;
OR2     gate5131  (.A(g6364), .B(g4269), .Z(g6930) ) ;
INV     gate5132  (.A(g6930), .Z(II12035) ) ;
INV     gate5133  (.A(II12035), .Z(g7571) ) ;
INV     gate5134  (.A(g6995), .Z(g7574) ) ;
OR2     gate5135  (.A(g6359), .B(g5703), .Z(g6928) ) ;
INV     gate5136  (.A(g6928), .Z(II12053) ) ;
INV     gate5137  (.A(II12053), .Z(g7579) ) ;
OR2     gate5138  (.A(g6360), .B(g5704), .Z(g6929) ) ;
INV     gate5139  (.A(g6929), .Z(II12056) ) ;
INV     gate5140  (.A(II12056), .Z(g7580) ) ;
OR2     gate5141  (.A(g6363), .B(g5720), .Z(g6934) ) ;
INV     gate5142  (.A(g6934), .Z(II12081) ) ;
INV     gate5143  (.A(II12081), .Z(g7585) ) ;
OR2     gate5144  (.A(g6549), .B(g5913), .Z(g7258) ) ;
INV     gate5145  (.A(g7258), .Z(II12099) ) ;
INV     gate5146  (.A(II12099), .Z(g7589) ) ;
INV     gate5147  (.A(g6859), .Z(II12103) ) ;
INV     gate5148  (.A(II12103), .Z(g7591) ) ;
OR2     gate5149  (.A(g6554), .B(g5917), .Z(g7106) ) ;
INV     gate5150  (.A(g7106), .Z(II12120) ) ;
INV     gate5151  (.A(II12120), .Z(g7594) ) ;
INV     gate5152  (.A(g6861), .Z(II12123) ) ;
INV     gate5153  (.A(II12123), .Z(g7595) ) ;
INV     gate5154  (.A(g6870), .Z(II12133) ) ;
INV     gate5155  (.A(II12133), .Z(g7597) ) ;
INV     gate5156  (.A(g7074), .Z(II12150) ) ;
INV     gate5157  (.A(II12150), .Z(g7600) ) ;
INV     gate5158  (.A(g6874), .Z(II12153) ) ;
INV     gate5159  (.A(II12153), .Z(g7601) ) ;
INV     gate5160  (.A(g6878), .Z(II12156) ) ;
INV     gate5161  (.A(II12156), .Z(g7602) ) ;
INV     gate5162  (.A(g7243), .Z(II12159) ) ;
INV     gate5163  (.A(II12159), .Z(g7603) ) ;
INV     gate5164  (.A(g7146), .Z(II12162) ) ;
INV     gate5165  (.A(II12162), .Z(g7604) ) ;
INV     gate5166  (.A(g6882), .Z(II12165) ) ;
INV     gate5167  (.A(II12165), .Z(g7605) ) ;
INV     gate5168  (.A(g7256), .Z(II12168) ) ;
INV     gate5169  (.A(II12168), .Z(g7606) ) ;
INV     gate5170  (.A(g6885), .Z(II12171) ) ;
INV     gate5171  (.A(II12171), .Z(g7607) ) ;
INV     gate5172  (.A(g6939), .Z(II12174) ) ;
INV     gate5173  (.A(II12174), .Z(g7608) ) ;
INV     gate5174  (.A(g7259), .Z(II12177) ) ;
INV     gate5175  (.A(II12177), .Z(g7609) ) ;
INV     gate5176  (.A(g7263), .Z(II12180) ) ;
INV     gate5177  (.A(II12180), .Z(g7610) ) ;
INV     gate5178  (.A(g7007), .Z(II12183) ) ;
INV     gate5179  (.A(II12183), .Z(g7611) ) ;
INV     gate5180  (.A(g7264), .Z(II12186) ) ;
INV     gate5181  (.A(II12186), .Z(g7612) ) ;
INV     gate5182  (.A(g7268), .Z(II12190) ) ;
INV     gate5183  (.A(II12190), .Z(g7614) ) ;
INV     gate5184  (.A(g7270), .Z(II12193) ) ;
INV     gate5185  (.A(II12193), .Z(g7615) ) ;
INV     gate5186  (.A(g7272), .Z(II12196) ) ;
INV     gate5187  (.A(II12196), .Z(g7616) ) ;
INV     gate5188  (.A(g7278), .Z(II12199) ) ;
INV     gate5189  (.A(II12199), .Z(g7617) ) ;
AND2    gate5190  (.A(g6592), .B(g3105), .Z(g6983) ) ;
INV     gate5191  (.A(g6983), .Z(II12202) ) ;
INV     gate5192  (.A(II12202), .Z(g7618) ) ;
INV     gate5193  (.A(g6993), .Z(II12205) ) ;
INV     gate5194  (.A(II12205), .Z(g7619) ) ;
INV     gate5195  (.A(g7124), .Z(II12208) ) ;
INV     gate5196  (.A(II12208), .Z(g7620) ) ;
NAND2   gate5197  (.A(II11279), .B(II11280), .Z(g7067) ) ;
INV     gate5198  (.A(g7067), .Z(g7622) ) ;
INV     gate5199  (.A(g7049), .Z(II12223) ) ;
INV     gate5200  (.A(II12223), .Z(g7627) ) ;
INV     gate5201  (.A(g7066), .Z(II12226) ) ;
INV     gate5202  (.A(II12226), .Z(g7628) ) ;
INV     gate5203  (.A(g7070), .Z(II12229) ) ;
INV     gate5204  (.A(II12229), .Z(g7629) ) ;
INV     gate5205  (.A(g7072), .Z(II12232) ) ;
INV     gate5206  (.A(II12232), .Z(g7630) ) ;
INV     gate5207  (.A(g7082), .Z(II12235) ) ;
INV     gate5208  (.A(II12235), .Z(g7631) ) ;
INV     gate5209  (.A(g7073), .Z(II12239) ) ;
INV     gate5210  (.A(II12239), .Z(g7633) ) ;
INV     gate5211  (.A(g7089), .Z(II12242) ) ;
INV     gate5212  (.A(II12242), .Z(g7634) ) ;
INV     gate5213  (.A(g7093), .Z(II12245) ) ;
INV     gate5214  (.A(II12245), .Z(g7635) ) ;
INV     gate5215  (.A(g7098), .Z(II12248) ) ;
INV     gate5216  (.A(II12248), .Z(g7636) ) ;
INV     gate5217  (.A(g7076), .Z(II12251) ) ;
INV     gate5218  (.A(II12251), .Z(g7637) ) ;
OR2     gate5219  (.A(g6640), .B(g6058), .Z(g7203) ) ;
INV     gate5220  (.A(g7203), .Z(II12255) ) ;
INV     gate5221  (.A(II12255), .Z(g7648) ) ;
INV     gate5222  (.A(g7103), .Z(II12258) ) ;
INV     gate5223  (.A(II12258), .Z(g7649) ) ;
INV     gate5224  (.A(g7078), .Z(II12261) ) ;
INV     gate5225  (.A(II12261), .Z(g7650) ) ;
OR2     gate5226  (.A(g6647), .B(g6067), .Z(g7211) ) ;
INV     gate5227  (.A(g7211), .Z(II12265) ) ;
INV     gate5228  (.A(II12265), .Z(g7656) ) ;
INV     gate5229  (.A(g7107), .Z(II12268) ) ;
INV     gate5230  (.A(II12268), .Z(g7657) ) ;
OR2     gate5231  (.A(g6655), .B(g6070), .Z(g7218) ) ;
INV     gate5232  (.A(g7218), .Z(II12271) ) ;
INV     gate5233  (.A(II12271), .Z(g7658) ) ;
INV     gate5234  (.A(g7110), .Z(II12274) ) ;
INV     gate5235  (.A(II12274), .Z(g7659) ) ;
OR2     gate5236  (.A(g6666), .B(g6079), .Z(g7225) ) ;
INV     gate5237  (.A(g7225), .Z(II12279) ) ;
INV     gate5238  (.A(II12279), .Z(g7662) ) ;
INV     gate5239  (.A(g7113), .Z(II12282) ) ;
INV     gate5240  (.A(II12282), .Z(g7663) ) ;
OR2     gate5241  (.A(g6673), .B(g6087), .Z(g7231) ) ;
INV     gate5242  (.A(g7231), .Z(II12286) ) ;
INV     gate5243  (.A(II12286), .Z(g7669) ) ;
INV     gate5244  (.A(g7142), .Z(II12289) ) ;
INV     gate5245  (.A(II12289), .Z(g7670) ) ;
INV     gate5246  (.A(g7116), .Z(II12293) ) ;
INV     gate5247  (.A(II12293), .Z(g7672) ) ;
OR2     gate5248  (.A(g6684), .B(g6092), .Z(g7236) ) ;
INV     gate5249  (.A(g7236), .Z(II12296) ) ;
INV     gate5250  (.A(II12296), .Z(g7673) ) ;
OR2     gate5251  (.A(g6687), .B(g6095), .Z(g7240) ) ;
INV     gate5252  (.A(g7240), .Z(II12300) ) ;
INV     gate5253  (.A(II12300), .Z(g7675) ) ;
OR2     gate5254  (.A(g6693), .B(g6098), .Z(g7242) ) ;
INV     gate5255  (.A(g7242), .Z(II12303) ) ;
INV     gate5256  (.A(II12303), .Z(g7676) ) ;
INV     gate5257  (.A(g7148), .Z(g7677) ) ;
OR2     gate5258  (.A(g6696), .B(g6102), .Z(g7245) ) ;
INV     gate5259  (.A(g7245), .Z(II12307) ) ;
INV     gate5260  (.A(II12307), .Z(g7678) ) ;
INV     gate5261  (.A(g7148), .Z(g7680) ) ;
INV     gate5262  (.A(g7148), .Z(g7681) ) ;
INV     gate5263  (.A(g7148), .Z(g7682) ) ;
INV     gate5264  (.A(g7148), .Z(g7683) ) ;
INV     gate5265  (.A(g7148), .Z(g7684) ) ;
INV     gate5266  (.A(g7148), .Z(g7685) ) ;
INV     gate5267  (.A(g7148), .Z(g7686) ) ;
INV     gate5268  (.A(g6862), .Z(II12318) ) ;
INV     gate5269  (.A(II12318), .Z(g7687) ) ;
INV     gate5270  (.A(g7148), .Z(g7688) ) ;
INV     gate5271  (.A(g7246), .Z(II12322) ) ;
INV     gate5272  (.A(II12322), .Z(g7689) ) ;
INV     gate5273  (.A(g7148), .Z(g7692) ) ;
INV     gate5274  (.A(g7246), .Z(II12326) ) ;
INV     gate5275  (.A(II12326), .Z(g7693) ) ;
INV     gate5276  (.A(g7148), .Z(g7696) ) ;
NAND2   gate5277  (.A(g6617), .B(g2364), .Z(g7101) ) ;
INV     gate5278  (.A(g7101), .Z(g7697) ) ;
INV     gate5279  (.A(g7079), .Z(g7702) ) ;
INV     gate5280  (.A(g7085), .Z(g7703) ) ;
OR2     gate5281  (.A(g6616), .B(g3067), .Z(g7133) ) ;
INV     gate5282  (.A(g7133), .Z(II12335) ) ;
INV     gate5283  (.A(II12335), .Z(g7706) ) ;
NAND2   gate5284  (.A(II11242), .B(II11243), .Z(g7054) ) ;
INV     gate5285  (.A(g7054), .Z(II12339) ) ;
INV     gate5286  (.A(II12339), .Z(g7708) ) ;
NAND2   gate5287  (.A(II11262), .B(II11263), .Z(g7062) ) ;
INV     gate5288  (.A(g7062), .Z(II12344) ) ;
INV     gate5289  (.A(II12344), .Z(g7711) ) ;
OR2     gate5290  (.A(g6619), .B(g6039), .Z(g7143) ) ;
INV     gate5291  (.A(g7143), .Z(II12354) ) ;
INV     gate5292  (.A(II12354), .Z(g7723) ) ;
INV     gate5293  (.A(g7147), .Z(II12357) ) ;
INV     gate5294  (.A(II12357), .Z(g7724) ) ;
OR2     gate5295  (.A(g6623), .B(g6046), .Z(g7183) ) ;
INV     gate5296  (.A(g7183), .Z(II12360) ) ;
INV     gate5297  (.A(II12360), .Z(g7725) ) ;
INV     gate5298  (.A(g7187), .Z(II12363) ) ;
INV     gate5299  (.A(II12363), .Z(g7726) ) ;
AND2    gate5300  (.A(g5587), .B(g6354), .Z(g7134) ) ;
INV     gate5301  (.A(g7134), .Z(II12366) ) ;
INV     gate5302  (.A(II12366), .Z(g7727) ) ;
OR2     gate5303  (.A(g6632), .B(g6053), .Z(g7189) ) ;
INV     gate5304  (.A(g7189), .Z(II12369) ) ;
INV     gate5305  (.A(II12369), .Z(g7728) ) ;
AND2    gate5306  (.A(g5590), .B(g6361), .Z(g7137) ) ;
INV     gate5307  (.A(g7137), .Z(II12372) ) ;
INV     gate5308  (.A(II12372), .Z(g7729) ) ;
INV     gate5309  (.A(g7195), .Z(II12376) ) ;
INV     gate5310  (.A(II12376), .Z(g7731) ) ;
OR2     gate5311  (.A(g6645), .B(g6062), .Z(g7204) ) ;
INV     gate5312  (.A(g7204), .Z(II12380) ) ;
INV     gate5313  (.A(II12380), .Z(g7733) ) ;
INV     gate5314  (.A(g7212), .Z(II12384) ) ;
INV     gate5315  (.A(II12384), .Z(g7735) ) ;
OR2     gate5316  (.A(g6661), .B(g6076), .Z(g7219) ) ;
INV     gate5317  (.A(g7219), .Z(II12388) ) ;
INV     gate5318  (.A(II12388), .Z(g7737) ) ;
INV     gate5319  (.A(g7284), .Z(II12397) ) ;
INV     gate5320  (.A(g7537), .Z(II12400) ) ;
INV     gate5321  (.A(g7611), .Z(II12403) ) ;
INV     gate5322  (.A(g7464), .Z(II12406) ) ;
INV     gate5323  (.A(g7501), .Z(II12409) ) ;
INV     gate5324  (.A(g7520), .Z(II12412) ) ;
INV     gate5325  (.A(g7631), .Z(II12415) ) ;
INV     gate5326  (.A(g7568), .Z(II12418) ) ;
INV     gate5327  (.A(g7634), .Z(II12421) ) ;
INV     gate5328  (.A(g7635), .Z(II12424) ) ;
INV     gate5329  (.A(g7636), .Z(II12427) ) ;
INV     gate5330  (.A(g7649), .Z(II12430) ) ;
INV     gate5331  (.A(g7657), .Z(II12433) ) ;
INV     gate5332  (.A(g7659), .Z(II12436) ) ;
INV     gate5333  (.A(g7663), .Z(II12439) ) ;
INV     gate5334  (.A(g7672), .Z(II12442) ) ;
INV     gate5335  (.A(g7521), .Z(II12445) ) ;
INV     gate5336  (.A(g7530), .Z(II12448) ) ;
INV     gate5337  (.A(g7538), .Z(II12451) ) ;
INV     gate5338  (.A(g7544), .Z(II12454) ) ;
INV     gate5339  (.A(g7559), .Z(II12457) ) ;
INV     gate5340  (.A(g7569), .Z(II12460) ) ;
INV     gate5341  (.A(g7579), .Z(II12463) ) ;
INV     gate5342  (.A(g7585), .Z(II12466) ) ;
INV     gate5343  (.A(g7531), .Z(II12469) ) ;
INV     gate5344  (.A(g7539), .Z(II12472) ) ;
INV     gate5345  (.A(g7545), .Z(II12475) ) ;
INV     gate5346  (.A(g7560), .Z(II12478) ) ;
INV     gate5347  (.A(g7570), .Z(II12481) ) ;
INV     gate5348  (.A(g7580), .Z(II12484) ) ;
INV     gate5349  (.A(g7723), .Z(II12487) ) ;
INV     gate5350  (.A(g7637), .Z(II12490) ) ;
INV     gate5351  (.A(g7650), .Z(II12493) ) ;
INV     gate5352  (.A(g7724), .Z(II12496) ) ;
INV     gate5353  (.A(g7725), .Z(II12499) ) ;
INV     gate5354  (.A(g7726), .Z(II12502) ) ;
INV     gate5355  (.A(g7728), .Z(II12505) ) ;
INV     gate5356  (.A(g7731), .Z(II12508) ) ;
INV     gate5357  (.A(g7733), .Z(II12511) ) ;
INV     gate5358  (.A(g7735), .Z(II12514) ) ;
INV     gate5359  (.A(g7737), .Z(II12517) ) ;
INV     gate5360  (.A(g7415), .Z(II12520) ) ;
INV     gate5361  (.A(g7421), .Z(II12523) ) ;
INV     gate5362  (.A(g7648), .Z(II12526) ) ;
INV     gate5363  (.A(g7589), .Z(II12529) ) ;
INV     gate5364  (.A(g7594), .Z(II12532) ) ;
INV     gate5365  (.A(g7656), .Z(II12535) ) ;
INV     gate5366  (.A(g7658), .Z(II12538) ) ;
INV     gate5367  (.A(g7662), .Z(II12541) ) ;
INV     gate5368  (.A(g7669), .Z(II12544) ) ;
INV     gate5369  (.A(g7673), .Z(II12547) ) ;
INV     gate5370  (.A(g7675), .Z(II12550) ) ;
INV     gate5371  (.A(g7676), .Z(II12553) ) ;
INV     gate5372  (.A(g7678), .Z(II12556) ) ;
INV     gate5373  (.A(g7477), .Z(II12559) ) ;
INV     gate5374  (.A(g7377), .Z(II12562) ) ;
INV     gate5375  (.A(g7388), .Z(II12565) ) ;
INV     gate5376  (.A(g7502), .Z(II12568) ) ;
INV     gate5377  (.A(g7509), .Z(II12571) ) ;
INV     gate5378  (.A(g7522), .Z(II12574) ) ;
INV     gate5379  (.A(g7532), .Z(II12577) ) ;
INV     gate5380  (.A(g7540), .Z(II12580) ) ;
INV     gate5381  (.A(g7546), .Z(II12583) ) ;
INV     gate5382  (.A(g7561), .Z(II12586) ) ;
INV     gate5383  (.A(g7571), .Z(II12589) ) ;
INV     gate5384  (.A(g7445), .Z(II12592) ) ;
INV     gate5385  (.A(g7706), .Z(II12595) ) ;
INV     gate5386  (.A(g7628), .Z(II12598) ) ;
INV     gate5387  (.A(g7629), .Z(II12601) ) ;
INV     gate5388  (.A(g7630), .Z(II12604) ) ;
INV     gate5389  (.A(g7633), .Z(II12607) ) ;
INV     gate5390  (.A(g7627), .Z(II12610) ) ;
INV     gate5391  (.A(g7525), .Z(II12613) ) ;
INV     gate5392  (.A(g7534), .Z(II12616) ) ;
INV     gate5393  (.A(g7697), .Z(II12627) ) ;
INV     gate5394  (.A(II12627), .Z(g7826) ) ;
AND2    gate5395  (.A(g6853), .B(g4328), .Z(g7705) ) ;
INV     gate5396  (.A(g7705), .Z(II12631) ) ;
INV     gate5397  (.A(II12631), .Z(g7844) ) ;
INV     gate5398  (.A(g7727), .Z(II12634) ) ;
INV     gate5399  (.A(II12634), .Z(g7845) ) ;
INV     gate5400  (.A(g7708), .Z(II12638) ) ;
INV     gate5401  (.A(II12638), .Z(g7847) ) ;
AND2    gate5402  (.A(g6856), .B(g4333), .Z(g7709) ) ;
INV     gate5403  (.A(g7709), .Z(II12641) ) ;
INV     gate5404  (.A(II12641), .Z(g7848) ) ;
INV     gate5405  (.A(g7729), .Z(II12644) ) ;
INV     gate5406  (.A(II12644), .Z(g7849) ) ;
INV     gate5407  (.A(g7711), .Z(II12647) ) ;
INV     gate5408  (.A(II12647), .Z(g7850) ) ;
INV     gate5409  (.A(g7479), .Z(g7851) ) ;
INV     gate5410  (.A(g7479), .Z(g7852) ) ;
INV     gate5411  (.A(g7458), .Z(II12652) ) ;
INV     gate5412  (.A(II12652), .Z(g7853) ) ;
INV     gate5413  (.A(g7402), .Z(II12655) ) ;
INV     gate5414  (.A(II12655), .Z(g7872) ) ;
INV     gate5415  (.A(g7479), .Z(g7877) ) ;
INV     gate5416  (.A(g7479), .Z(g7878) ) ;
INV     gate5417  (.A(g7479), .Z(g7880) ) ;
INV     gate5418  (.A(g7479), .Z(g7882) ) ;
INV     gate5419  (.A(g7689), .Z(g7883) ) ;
INV     gate5420  (.A(g7479), .Z(g7886) ) ;
INV     gate5421  (.A(g7693), .Z(g7887) ) ;
INV     gate5422  (.A(g7479), .Z(g7890) ) ;
INV     gate5423  (.A(g7376), .Z(II12678) ) ;
INV     gate5424  (.A(II12678), .Z(g7896) ) ;
OR2     gate5425  (.A(g7125), .B(g3540), .Z(g7712) ) ;
INV     gate5426  (.A(g7712), .Z(g7897) ) ;
INV     gate5427  (.A(g7387), .Z(II12683) ) ;
INV     gate5428  (.A(II12683), .Z(g7899) ) ;
INV     gate5429  (.A(g7712), .Z(g7900) ) ;
INV     gate5430  (.A(g7712), .Z(g7901) ) ;
INV     gate5431  (.A(g7446), .Z(g7903) ) ;
INV     gate5432  (.A(g7555), .Z(II12690) ) ;
INV     gate5433  (.A(II12690), .Z(g7904) ) ;
INV     gate5434  (.A(g7450), .Z(g7905) ) ;
INV     gate5435  (.A(g7374), .Z(II12694) ) ;
INV     gate5436  (.A(II12694), .Z(g7906) ) ;
OR2     gate5437  (.A(g6855), .B(g4084), .Z(g7664) ) ;
INV     gate5438  (.A(g7664), .Z(g7907) ) ;
INV     gate5439  (.A(g7454), .Z(g7908) ) ;
INV     gate5440  (.A(g7664), .Z(g7909) ) ;
INV     gate5441  (.A(g7460), .Z(g7910) ) ;
INV     gate5442  (.A(g7664), .Z(g7911) ) ;
OR2     gate5443  (.A(g7135), .B(g4084), .Z(g7651) ) ;
INV     gate5444  (.A(g7651), .Z(g7912) ) ;
INV     gate5445  (.A(g7467), .Z(g7913) ) ;
INV     gate5446  (.A(g7651), .Z(g7914) ) ;
INV     gate5447  (.A(g7473), .Z(g7915) ) ;
INV     gate5448  (.A(g7651), .Z(g7916) ) ;
INV     gate5449  (.A(g7497), .Z(g7917) ) ;
INV     gate5450  (.A(g7505), .Z(g7918) ) ;
INV     gate5451  (.A(g7512), .Z(g7919) ) ;
INV     gate5452  (.A(g7516), .Z(g7920) ) ;
INV     gate5453  (.A(g7463), .Z(g7921) ) ;
OR2     gate5454  (.A(g7271), .B(g6789), .Z(g7441) ) ;
INV     gate5455  (.A(g7441), .Z(II12712) ) ;
INV     gate5456  (.A(II12712), .Z(g7922) ) ;
INV     gate5457  (.A(g7527), .Z(g7923) ) ;
INV     gate5458  (.A(g7470), .Z(g7924) ) ;
INV     gate5459  (.A(g7476), .Z(g7925) ) ;
INV     gate5460  (.A(g7500), .Z(g7927) ) ;
INV     gate5461  (.A(g7508), .Z(g7928) ) ;
INV     gate5462  (.A(g7519), .Z(g7929) ) ;
INV     gate5463  (.A(g7712), .Z(g7936) ) ;
INV     gate5464  (.A(g7403), .Z(g7938) ) ;
INV     gate5465  (.A(g7406), .Z(g7941) ) ;
INV     gate5466  (.A(g7410), .Z(g7944) ) ;
INV     gate5467  (.A(g7416), .Z(g7946) ) ;
INV     gate5468  (.A(g7422), .Z(g7949) ) ;
INV     gate5469  (.A(g7427), .Z(g7952) ) ;
INV     gate5470  (.A(g7432), .Z(g7956) ) ;
OR2     gate5471  (.A(g7060), .B(g5267), .Z(g7626) ) ;
INV     gate5472  (.A(g7626), .Z(II12751) ) ;
INV     gate5473  (.A(II12751), .Z(g7959) ) ;
INV     gate5474  (.A(g7664), .Z(g7961) ) ;
INV     gate5475  (.A(g7651), .Z(g7964) ) ;
INV     gate5476  (.A(g7702), .Z(II12759) ) ;
INV     gate5477  (.A(II12759), .Z(g7965) ) ;
AND2    gate5478  (.A(g7075), .B(g3109), .Z(g7541) ) ;
INV     gate5479  (.A(g7541), .Z(II12762) ) ;
INV     gate5480  (.A(II12762), .Z(g7966) ) ;
OR2     gate5481  (.A(g7265), .B(g6488), .Z(g7638) ) ;
INV     gate5482  (.A(g7638), .Z(II12765) ) ;
INV     gate5483  (.A(II12765), .Z(g7967) ) ;
INV     gate5484  (.A(g7638), .Z(II12770) ) ;
INV     gate5485  (.A(II12770), .Z(g7972) ) ;
AND2    gate5486  (.A(g7092), .B(g5420), .Z(g7581) ) ;
INV     gate5487  (.A(g7581), .Z(II12773) ) ;
INV     gate5488  (.A(II12773), .Z(g7975) ) ;
AND2    gate5489  (.A(g7096), .B(g5423), .Z(g7586) ) ;
INV     gate5490  (.A(g7586), .Z(II12776) ) ;
INV     gate5491  (.A(II12776), .Z(g7976) ) ;
INV     gate5492  (.A(g7608), .Z(II12779) ) ;
INV     gate5493  (.A(II12779), .Z(g7977) ) ;
AND2    gate5494  (.A(g7102), .B(g5425), .Z(g7590) ) ;
INV     gate5495  (.A(g7590), .Z(II12783) ) ;
INV     gate5496  (.A(II12783), .Z(g7979) ) ;
INV     gate5497  (.A(g7622), .Z(II12786) ) ;
INV     gate5498  (.A(II12786), .Z(g7980) ) ;
NAND2   gate5499  (.A(II12215), .B(II12216), .Z(g7624) ) ;
INV     gate5500  (.A(g7624), .Z(g7981) ) ;
INV     gate5501  (.A(g7618), .Z(II12790) ) ;
INV     gate5502  (.A(II12790), .Z(g7982) ) ;
INV     gate5503  (.A(g7619), .Z(II12793) ) ;
INV     gate5504  (.A(II12793), .Z(g7983) ) ;
INV     gate5505  (.A(g7543), .Z(II12796) ) ;
INV     gate5506  (.A(II12796), .Z(g7984) ) ;
INV     gate5507  (.A(g7556), .Z(II12799) ) ;
INV     gate5508  (.A(II12799), .Z(g7985) ) ;
INV     gate5509  (.A(g7684), .Z(II12805) ) ;
INV     gate5510  (.A(II12805), .Z(g7989) ) ;
INV     gate5511  (.A(g7686), .Z(II12809) ) ;
INV     gate5512  (.A(II12809), .Z(g7991) ) ;
INV     gate5513  (.A(g7688), .Z(II12813) ) ;
INV     gate5514  (.A(II12813), .Z(g7993) ) ;
INV     gate5515  (.A(g7692), .Z(II12817) ) ;
INV     gate5516  (.A(II12817), .Z(g7995) ) ;
INV     gate5517  (.A(g7697), .Z(g7997) ) ;
INV     gate5518  (.A(g7677), .Z(II12822) ) ;
INV     gate5519  (.A(II12822), .Z(g7998) ) ;
INV     gate5520  (.A(g7696), .Z(II12825) ) ;
INV     gate5521  (.A(II12825), .Z(g7999) ) ;
INV     gate5522  (.A(g7680), .Z(II12829) ) ;
INV     gate5523  (.A(II12829), .Z(g8001) ) ;
INV     gate5524  (.A(g7681), .Z(II12832) ) ;
INV     gate5525  (.A(II12832), .Z(g8002) ) ;
OR2     gate5526  (.A(g7059), .B(g6583), .Z(g7660) ) ;
INV     gate5527  (.A(g7660), .Z(II12835) ) ;
INV     gate5528  (.A(II12835), .Z(g8003) ) ;
INV     gate5529  (.A(g7682), .Z(II12838) ) ;
INV     gate5530  (.A(II12838), .Z(g8004) ) ;
INV     gate5531  (.A(g7683), .Z(II12843) ) ;
INV     gate5532  (.A(II12843), .Z(g8007) ) ;
INV     gate5533  (.A(g7685), .Z(II12846) ) ;
INV     gate5534  (.A(II12846), .Z(g8008) ) ;
AND2    gate5535  (.A(g7184), .B(g5574), .Z(g7632) ) ;
INV     gate5536  (.A(g7632), .Z(II12849) ) ;
INV     gate5537  (.A(II12849), .Z(g8009) ) ;
INV     gate5538  (.A(g7638), .Z(II12853) ) ;
INV     gate5539  (.A(II12853), .Z(g8011) ) ;
INV     gate5540  (.A(g7638), .Z(II12857) ) ;
INV     gate5541  (.A(II12857), .Z(g8015) ) ;
INV     gate5542  (.A(g7638), .Z(II12862) ) ;
INV     gate5543  (.A(II12862), .Z(g8020) ) ;
INV     gate5544  (.A(g7638), .Z(II12867) ) ;
INV     gate5545  (.A(II12867), .Z(g8025) ) ;
INV     gate5546  (.A(g7638), .Z(II12871) ) ;
INV     gate5547  (.A(II12871), .Z(g8029) ) ;
INV     gate5548  (.A(g7638), .Z(II12875) ) ;
INV     gate5549  (.A(II12875), .Z(g8033) ) ;
INV     gate5550  (.A(g7638), .Z(II12878) ) ;
INV     gate5551  (.A(II12878), .Z(g8036) ) ;
NAND4   gate5552  (.A(g7011), .B(g6995), .C(g6984), .D(g6974), .Z(g7671) ) ;
INV     gate5553  (.A(g7671), .Z(g8056) ) ;
INV     gate5554  (.A(g7984), .Z(II12901) ) ;
INV     gate5555  (.A(g7985), .Z(II12904) ) ;
INV     gate5556  (.A(g7959), .Z(II12907) ) ;
INV     gate5557  (.A(g7922), .Z(II12910) ) ;
INV     gate5558  (.A(g7845), .Z(II12913) ) ;
INV     gate5559  (.A(g7849), .Z(II12916) ) ;
INV     gate5560  (.A(g8003), .Z(II12919) ) ;
INV     gate5561  (.A(g7896), .Z(II12930) ) ;
INV     gate5562  (.A(g7899), .Z(II12933) ) ;
INV     gate5563  (.A(g7983), .Z(II12936) ) ;
INV     gate5564  (.A(g7977), .Z(II12939) ) ;
INV     gate5565  (.A(g7982), .Z(II12942) ) ;
NAND4   gate5566  (.A(g7011), .B(g7574), .C(g7562), .D(g7550), .Z(g8000) ) ;
INV     gate5567  (.A(g8000), .Z(g8081) ) ;
NAND4   gate5568  (.A(g7395), .B(g6847), .C(g7279), .D(g7273), .Z(g7932) ) ;
INV     gate5569  (.A(g7932), .Z(g8085) ) ;
NAND4   gate5570  (.A(g7395), .B(g6847), .C(g7279), .D(g7369), .Z(g7934) ) ;
INV     gate5571  (.A(g7934), .Z(g8089) ) ;
AND2    gate5572  (.A(g7386), .B(g4332), .Z(g8019) ) ;
INV     gate5573  (.A(g8019), .Z(II12948) ) ;
INV     gate5574  (.A(II12948), .Z(g8093) ) ;
NAND4   gate5575  (.A(g7011), .B(g6995), .C(g7562), .D(g6974), .Z(g7987) ) ;
INV     gate5576  (.A(g7987), .Z(g8094) ) ;
NAND4   gate5577  (.A(g7395), .B(g6847), .C(g7380), .D(g7369), .Z(g7942) ) ;
INV     gate5578  (.A(g7942), .Z(g8095) ) ;
AND2    gate5579  (.A(g7394), .B(g4337), .Z(g8024) ) ;
INV     gate5580  (.A(g8024), .Z(II12953) ) ;
INV     gate5581  (.A(II12953), .Z(g8096) ) ;
NAND4   gate5582  (.A(g7011), .B(g6995), .C(g7562), .D(g7550), .Z(g7990) ) ;
INV     gate5583  (.A(g7990), .Z(g8099) ) ;
NAND4   gate5584  (.A(g7395), .B(g7390), .C(g7279), .D(g7369), .Z(g7947) ) ;
INV     gate5585  (.A(g7947), .Z(g8100) ) ;
NAND4   gate5586  (.A(g7011), .B(g7574), .C(g6984), .D(g7550), .Z(g7994) ) ;
INV     gate5587  (.A(g7994), .Z(g8103) ) ;
NAND4   gate5588  (.A(g7011), .B(g7574), .C(g6984), .D(g6974), .Z(g7992) ) ;
INV     gate5589  (.A(g7992), .Z(g8105) ) ;
NAND4   gate5590  (.A(g7395), .B(g7390), .C(g7380), .D(g7273), .Z(g7950) ) ;
INV     gate5591  (.A(g7950), .Z(g8106) ) ;
NAND4   gate5592  (.A(g7011), .B(g7574), .C(g7562), .D(g6974), .Z(g7996) ) ;
INV     gate5593  (.A(g7996), .Z(g8110) ) ;
NAND4   gate5594  (.A(g7395), .B(g7390), .C(g7380), .D(g7369), .Z(g7953) ) ;
INV     gate5595  (.A(g7953), .Z(g8115) ) ;
AND2    gate5596  (.A(g7587), .B(g5128), .Z(g8039) ) ;
INV     gate5597  (.A(g8039), .Z(II12971) ) ;
INV     gate5598  (.A(II12971), .Z(g8116) ) ;
AND2    gate5599  (.A(g7523), .B(g5128), .Z(g8040) ) ;
INV     gate5600  (.A(g8040), .Z(II12978) ) ;
INV     gate5601  (.A(II12978), .Z(g8121) ) ;
AND2    gate5602  (.A(g7524), .B(g5128), .Z(g8041) ) ;
INV     gate5603  (.A(g8041), .Z(II12981) ) ;
INV     gate5604  (.A(II12981), .Z(g8122) ) ;
INV     gate5605  (.A(g8011), .Z(g8124) ) ;
AND2    gate5606  (.A(g7533), .B(g5128), .Z(g8042) ) ;
INV     gate5607  (.A(g8042), .Z(II12986) ) ;
INV     gate5608  (.A(II12986), .Z(g8125) ) ;
AND2    gate5609  (.A(g7582), .B(g5128), .Z(g8043) ) ;
INV     gate5610  (.A(g8043), .Z(II12989) ) ;
INV     gate5611  (.A(II12989), .Z(g8126) ) ;
AND2    gate5612  (.A(g7598), .B(g5919), .Z(g8044) ) ;
INV     gate5613  (.A(g8044), .Z(II12993) ) ;
INV     gate5614  (.A(II12993), .Z(g8128) ) ;
INV     gate5615  (.A(g8015), .Z(g8129) ) ;
INV     gate5616  (.A(g8020), .Z(g8131) ) ;
INV     gate5617  (.A(g7844), .Z(II12999) ) ;
INV     gate5618  (.A(II12999), .Z(g8132) ) ;
AND2    gate5619  (.A(g7547), .B(g5128), .Z(g8045) ) ;
INV     gate5620  (.A(g8045), .Z(II13002) ) ;
INV     gate5621  (.A(II13002), .Z(g8133) ) ;
AND2    gate5622  (.A(g7548), .B(g5128), .Z(g8046) ) ;
INV     gate5623  (.A(g8046), .Z(II13005) ) ;
INV     gate5624  (.A(II13005), .Z(g8134) ) ;
AND2    gate5625  (.A(g7557), .B(g5919), .Z(g8047) ) ;
INV     gate5626  (.A(g8047), .Z(II13010) ) ;
INV     gate5627  (.A(II13010), .Z(g8137) ) ;
AND2    gate5628  (.A(g7558), .B(g5919), .Z(g8048) ) ;
INV     gate5629  (.A(g8048), .Z(II13013) ) ;
INV     gate5630  (.A(II13013), .Z(g8138) ) ;
INV     gate5631  (.A(g8025), .Z(g8139) ) ;
INV     gate5632  (.A(g7848), .Z(II13017) ) ;
INV     gate5633  (.A(II13017), .Z(g8140) ) ;
AND2    gate5634  (.A(g7567), .B(g5919), .Z(g8049) ) ;
INV     gate5635  (.A(g8049), .Z(II13020) ) ;
INV     gate5636  (.A(II13020), .Z(g8141) ) ;
AND2    gate5637  (.A(g7596), .B(g5919), .Z(g8050) ) ;
INV     gate5638  (.A(g8050), .Z(II13023) ) ;
INV     gate5639  (.A(II13023), .Z(g8142) ) ;
INV     gate5640  (.A(g8029), .Z(g8143) ) ;
AND2    gate5641  (.A(g7572), .B(g5128), .Z(g8051) ) ;
INV     gate5642  (.A(g8051), .Z(II13027) ) ;
INV     gate5643  (.A(II13027), .Z(g8144) ) ;
AND2    gate5644  (.A(g7573), .B(g5128), .Z(g8052) ) ;
INV     gate5645  (.A(g8052), .Z(II13030) ) ;
INV     gate5646  (.A(II13030), .Z(g8145) ) ;
INV     gate5647  (.A(g8033), .Z(g8146) ) ;
AND2    gate5648  (.A(g7583), .B(g5919), .Z(g8053) ) ;
INV     gate5649  (.A(g8053), .Z(II13036) ) ;
INV     gate5650  (.A(II13036), .Z(g8149) ) ;
AND2    gate5651  (.A(g7584), .B(g5919), .Z(g8054) ) ;
INV     gate5652  (.A(g8054), .Z(II13039) ) ;
INV     gate5653  (.A(II13039), .Z(g8150) ) ;
INV     gate5654  (.A(g8036), .Z(g8151) ) ;
AND2    gate5655  (.A(g7588), .B(g5128), .Z(g8055) ) ;
INV     gate5656  (.A(g8055), .Z(II13043) ) ;
INV     gate5657  (.A(II13043), .Z(g8152) ) ;
AND2    gate5658  (.A(g7592), .B(g5919), .Z(g8059) ) ;
INV     gate5659  (.A(g8059), .Z(II13048) ) ;
INV     gate5660  (.A(II13048), .Z(g8155) ) ;
AND2    gate5661  (.A(g7593), .B(g5919), .Z(g8060) ) ;
INV     gate5662  (.A(g8060), .Z(II13051) ) ;
INV     gate5663  (.A(II13051), .Z(g8156) ) ;
AND2    gate5664  (.A(g7599), .B(g5919), .Z(g7843) ) ;
INV     gate5665  (.A(g7843), .Z(II13057) ) ;
INV     gate5666  (.A(II13057), .Z(g8160) ) ;
INV     gate5667  (.A(g7872), .Z(g8164) ) ;
INV     gate5668  (.A(g7906), .Z(II13068) ) ;
INV     gate5669  (.A(II13068), .Z(g8171) ) ;
INV     gate5670  (.A(g7921), .Z(II13083) ) ;
INV     gate5671  (.A(II13083), .Z(g8178) ) ;
INV     gate5672  (.A(g7924), .Z(II13086) ) ;
INV     gate5673  (.A(II13086), .Z(g8179) ) ;
INV     gate5674  (.A(g7925), .Z(II13096) ) ;
INV     gate5675  (.A(II13096), .Z(g8181) ) ;
INV     gate5676  (.A(g7927), .Z(II13099) ) ;
INV     gate5677  (.A(II13099), .Z(g8182) ) ;
INV     gate5678  (.A(g7928), .Z(II13102) ) ;
INV     gate5679  (.A(II13102), .Z(g8183) ) ;
INV     gate5680  (.A(g7929), .Z(II13105) ) ;
INV     gate5681  (.A(II13105), .Z(g8184) ) ;
INV     gate5682  (.A(g7981), .Z(II13109) ) ;
INV     gate5683  (.A(II13109), .Z(g8186) ) ;
AND2    gate5684  (.A(g7621), .B(g3110), .Z(g7930) ) ;
INV     gate5685  (.A(g7930), .Z(II13114) ) ;
INV     gate5686  (.A(II13114), .Z(g8191) ) ;
INV     gate5687  (.A(g7904), .Z(II13117) ) ;
INV     gate5688  (.A(II13117), .Z(g8192) ) ;
INV     gate5689  (.A(g7966), .Z(II13122) ) ;
INV     gate5690  (.A(II13122), .Z(g8195) ) ;
INV     gate5691  (.A(g7975), .Z(II13125) ) ;
INV     gate5692  (.A(II13125), .Z(g8196) ) ;
INV     gate5693  (.A(g7976), .Z(II13128) ) ;
INV     gate5694  (.A(II13128), .Z(g8197) ) ;
INV     gate5695  (.A(g7979), .Z(II13131) ) ;
INV     gate5696  (.A(II13131), .Z(g8198) ) ;
INV     gate5697  (.A(g7826), .Z(g8213) ) ;
INV     gate5698  (.A(g7826), .Z(g8218) ) ;
INV     gate5699  (.A(g7826), .Z(g8219) ) ;
INV     gate5700  (.A(g7826), .Z(g8220) ) ;
INV     gate5701  (.A(g7826), .Z(g8225) ) ;
INV     gate5702  (.A(g7826), .Z(g8229) ) ;
INV     gate5703  (.A(g7872), .Z(g8233) ) ;
INV     gate5704  (.A(g7826), .Z(g8234) ) ;
INV     gate5705  (.A(g7967), .Z(g8235) ) ;
INV     gate5706  (.A(g7826), .Z(g8239) ) ;
INV     gate5707  (.A(g7972), .Z(g8240) ) ;
INV     gate5708  (.A(g8009), .Z(II13166) ) ;
INV     gate5709  (.A(II13166), .Z(g8251) ) ;
NAND4   gate5710  (.A(g7011), .B(g6995), .C(g6984), .D(g7550), .Z(g7986) ) ;
INV     gate5711  (.A(g7986), .Z(g8255) ) ;
INV     gate5712  (.A(g8192), .Z(II13185) ) ;
INV     gate5713  (.A(g8171), .Z(II13188) ) ;
INV     gate5714  (.A(g8132), .Z(II13191) ) ;
INV     gate5715  (.A(g8140), .Z(II13194) ) ;
INV     gate5716  (.A(g8186), .Z(II13197) ) ;
INV     gate5717  (.A(g8251), .Z(II13200) ) ;
INV     gate5718  (.A(g8196), .Z(II13203) ) ;
INV     gate5719  (.A(g8197), .Z(II13206) ) ;
INV     gate5720  (.A(g8198), .Z(II13209) ) ;
INV     gate5721  (.A(g8195), .Z(II13212) ) ;
OR2     gate5722  (.A(g7876), .B(g3383), .Z(g8261) ) ;
INV     gate5723  (.A(g8261), .Z(II13224) ) ;
INV     gate5724  (.A(II13224), .Z(g8290) ) ;
OR2     gate5725  (.A(g7879), .B(g3389), .Z(g8264) ) ;
INV     gate5726  (.A(g8264), .Z(II13227) ) ;
INV     gate5727  (.A(II13227), .Z(g8291) ) ;
AND2    gate5728  (.A(g7847), .B(g4336), .Z(g8244) ) ;
INV     gate5729  (.A(g8244), .Z(II13230) ) ;
INV     gate5730  (.A(II13230), .Z(g8292) ) ;
OR2     gate5731  (.A(g7881), .B(g3396), .Z(g8265) ) ;
INV     gate5732  (.A(g8265), .Z(II13233) ) ;
INV     gate5733  (.A(II13233), .Z(g8293) ) ;
AND2    gate5734  (.A(g7850), .B(g4339), .Z(g8245) ) ;
INV     gate5735  (.A(g8245), .Z(II13236) ) ;
INV     gate5736  (.A(II13236), .Z(g8294) ) ;
OR2     gate5737  (.A(g7885), .B(g3412), .Z(g8266) ) ;
INV     gate5738  (.A(g8266), .Z(II13239) ) ;
INV     gate5739  (.A(II13239), .Z(g8295) ) ;
OR2     gate5740  (.A(g7889), .B(g3422), .Z(g8267) ) ;
INV     gate5741  (.A(g8267), .Z(II13242) ) ;
INV     gate5742  (.A(II13242), .Z(g8296) ) ;
OR2     gate5743  (.A(g7892), .B(g3429), .Z(g8269) ) ;
INV     gate5744  (.A(g8269), .Z(II13245) ) ;
INV     gate5745  (.A(II13245), .Z(g8297) ) ;
OR2     gate5746  (.A(g7894), .B(g3434), .Z(g8270) ) ;
INV     gate5747  (.A(g8270), .Z(II13255) ) ;
INV     gate5748  (.A(II13255), .Z(g8299) ) ;
AND2    gate5749  (.A(g2771), .B(g7907), .Z(g8250) ) ;
INV     gate5750  (.A(g8250), .Z(II13280) ) ;
INV     gate5751  (.A(II13280), .Z(g8304) ) ;
AND2    gate5752  (.A(g2773), .B(g7909), .Z(g8254) ) ;
INV     gate5753  (.A(g8254), .Z(II13290) ) ;
INV     gate5754  (.A(II13290), .Z(g8306) ) ;
AND2    gate5755  (.A(g2775), .B(g7911), .Z(g8260) ) ;
INV     gate5756  (.A(g8260), .Z(II13314) ) ;
INV     gate5757  (.A(II13314), .Z(g8310) ) ;
INV     gate5758  (.A(g8093), .Z(II13317) ) ;
INV     gate5759  (.A(II13317), .Z(g8311) ) ;
INV     gate5760  (.A(g8096), .Z(II13320) ) ;
INV     gate5761  (.A(II13320), .Z(g8312) ) ;
OR2     gate5762  (.A(g7453), .B(g7999), .Z(g8203) ) ;
INV     gate5763  (.A(g8203), .Z(II13323) ) ;
INV     gate5764  (.A(g8203), .Z(II13326) ) ;
INV     gate5765  (.A(II13326), .Z(g8314) ) ;
INV     gate5766  (.A(g8116), .Z(II13329) ) ;
INV     gate5767  (.A(II13329), .Z(g8315) ) ;
OR2     gate5768  (.A(g7459), .B(g8007), .Z(g8206) ) ;
INV     gate5769  (.A(g8206), .Z(II13332) ) ;
INV     gate5770  (.A(g8206), .Z(II13335) ) ;
INV     gate5771  (.A(II13335), .Z(g8317) ) ;
OR2     gate5772  (.A(g7466), .B(g7995), .Z(g8210) ) ;
INV     gate5773  (.A(g8210), .Z(II13338) ) ;
INV     gate5774  (.A(g8210), .Z(II13341) ) ;
INV     gate5775  (.A(II13341), .Z(g8319) ) ;
INV     gate5776  (.A(g8121), .Z(II13344) ) ;
INV     gate5777  (.A(II13344), .Z(g8320) ) ;
INV     gate5778  (.A(g8122), .Z(II13347) ) ;
INV     gate5779  (.A(II13347), .Z(g8321) ) ;
OR2     gate5780  (.A(g7472), .B(g8004), .Z(g8214) ) ;
INV     gate5781  (.A(g8214), .Z(II13351) ) ;
INV     gate5782  (.A(g8214), .Z(II13354) ) ;
INV     gate5783  (.A(II13354), .Z(g8324) ) ;
INV     gate5784  (.A(g8125), .Z(II13357) ) ;
INV     gate5785  (.A(II13357), .Z(g8325) ) ;
INV     gate5786  (.A(g8126), .Z(II13360) ) ;
INV     gate5787  (.A(II13360), .Z(g8326) ) ;
INV     gate5788  (.A(g8164), .Z(g8327) ) ;
OR2     gate5789  (.A(g7496), .B(g7993), .Z(g8221) ) ;
INV     gate5790  (.A(g8221), .Z(II13364) ) ;
INV     gate5791  (.A(g8221), .Z(II13367) ) ;
INV     gate5792  (.A(II13367), .Z(g8329) ) ;
INV     gate5793  (.A(g8128), .Z(II13370) ) ;
INV     gate5794  (.A(II13370), .Z(g8330) ) ;
OR2     gate5795  (.A(g7504), .B(g8002), .Z(g8226) ) ;
INV     gate5796  (.A(g8226), .Z(II13373) ) ;
INV     gate5797  (.A(g8226), .Z(II13376) ) ;
INV     gate5798  (.A(II13376), .Z(g8332) ) ;
INV     gate5799  (.A(g8133), .Z(II13379) ) ;
INV     gate5800  (.A(II13379), .Z(g8333) ) ;
INV     gate5801  (.A(g8134), .Z(II13382) ) ;
INV     gate5802  (.A(II13382), .Z(g8334) ) ;
OR2     gate5803  (.A(g7515), .B(g7991), .Z(g8230) ) ;
INV     gate5804  (.A(g8230), .Z(II13385) ) ;
INV     gate5805  (.A(g8230), .Z(II13388) ) ;
INV     gate5806  (.A(II13388), .Z(g8336) ) ;
INV     gate5807  (.A(g8178), .Z(II13391) ) ;
INV     gate5808  (.A(II13391), .Z(g8337) ) ;
INV     gate5809  (.A(g8137), .Z(II13394) ) ;
INV     gate5810  (.A(II13394), .Z(g8338) ) ;
INV     gate5811  (.A(g8138), .Z(II13397) ) ;
INV     gate5812  (.A(II13397), .Z(g8339) ) ;
OR2     gate5813  (.A(g7526), .B(g8001), .Z(g8236) ) ;
INV     gate5814  (.A(g8236), .Z(II13400) ) ;
INV     gate5815  (.A(g8236), .Z(II13403) ) ;
INV     gate5816  (.A(II13403), .Z(g8341) ) ;
INV     gate5817  (.A(g8179), .Z(II13406) ) ;
INV     gate5818  (.A(II13406), .Z(g8342) ) ;
INV     gate5819  (.A(g8141), .Z(II13409) ) ;
INV     gate5820  (.A(II13409), .Z(g8343) ) ;
INV     gate5821  (.A(g8142), .Z(II13412) ) ;
INV     gate5822  (.A(II13412), .Z(g8344) ) ;
INV     gate5823  (.A(g8144), .Z(II13415) ) ;
INV     gate5824  (.A(II13415), .Z(g8345) ) ;
INV     gate5825  (.A(g8145), .Z(II13418) ) ;
INV     gate5826  (.A(II13418), .Z(g8346) ) ;
OR2     gate5827  (.A(g7535), .B(g8008), .Z(g8200) ) ;
INV     gate5828  (.A(g8200), .Z(II13421) ) ;
INV     gate5829  (.A(g8200), .Z(II13424) ) ;
INV     gate5830  (.A(II13424), .Z(g8348) ) ;
OR2     gate5831  (.A(g7536), .B(g7989), .Z(g8241) ) ;
INV     gate5832  (.A(g8241), .Z(II13427) ) ;
INV     gate5833  (.A(g8241), .Z(II13430) ) ;
INV     gate5834  (.A(II13430), .Z(g8350) ) ;
INV     gate5835  (.A(g8181), .Z(II13433) ) ;
INV     gate5836  (.A(II13433), .Z(g8351) ) ;
OR2     gate5837  (.A(g7542), .B(g7998), .Z(g8187) ) ;
INV     gate5838  (.A(g8187), .Z(II13436) ) ;
INV     gate5839  (.A(g8187), .Z(II13439) ) ;
INV     gate5840  (.A(II13439), .Z(g8353) ) ;
INV     gate5841  (.A(g8182), .Z(II13442) ) ;
INV     gate5842  (.A(II13442), .Z(g8354) ) ;
INV     gate5843  (.A(g8149), .Z(II13445) ) ;
INV     gate5844  (.A(II13445), .Z(g8355) ) ;
INV     gate5845  (.A(g8150), .Z(II13448) ) ;
INV     gate5846  (.A(II13448), .Z(g8356) ) ;
INV     gate5847  (.A(g8152), .Z(II13451) ) ;
INV     gate5848  (.A(II13451), .Z(g8357) ) ;
INV     gate5849  (.A(g8183), .Z(II13454) ) ;
INV     gate5850  (.A(II13454), .Z(g8358) ) ;
INV     gate5851  (.A(g8184), .Z(II13457) ) ;
INV     gate5852  (.A(II13457), .Z(g8359) ) ;
INV     gate5853  (.A(g8155), .Z(II13460) ) ;
INV     gate5854  (.A(II13460), .Z(g8360) ) ;
INV     gate5855  (.A(g8156), .Z(II13463) ) ;
INV     gate5856  (.A(II13463), .Z(g8361) ) ;
INV     gate5857  (.A(g8160), .Z(II13466) ) ;
INV     gate5858  (.A(II13466), .Z(g8362) ) ;
AND2    gate5859  (.A(g2955), .B(g7961), .Z(g8147) ) ;
INV     gate5860  (.A(g8147), .Z(II13469) ) ;
INV     gate5861  (.A(II13469), .Z(g8363) ) ;
AND2    gate5862  (.A(g7971), .B(g3112), .Z(g8173) ) ;
INV     gate5863  (.A(g8173), .Z(II13475) ) ;
INV     gate5864  (.A(II13475), .Z(g8375) ) ;
INV     gate5865  (.A(g8191), .Z(II13478) ) ;
INV     gate5866  (.A(II13478), .Z(g8376) ) ;
OR2     gate5867  (.A(g5145), .B(g7937), .Z(g8193) ) ;
INV     gate5868  (.A(g8193), .Z(II13482) ) ;
INV     gate5869  (.A(II13482), .Z(g8378) ) ;
OR2     gate5870  (.A(g5168), .B(g7940), .Z(g8194) ) ;
INV     gate5871  (.A(g8194), .Z(II13485) ) ;
INV     gate5872  (.A(II13485), .Z(g8379) ) ;
INV     gate5873  (.A(g8233), .Z(II13489) ) ;
INV     gate5874  (.A(II13489), .Z(g8381) ) ;
INV     gate5875  (.A(g8343), .Z(II13568) ) ;
INV     gate5876  (.A(g8355), .Z(II13571) ) ;
INV     gate5877  (.A(g8360), .Z(II13574) ) ;
INV     gate5878  (.A(g8330), .Z(II13577) ) ;
INV     gate5879  (.A(g8338), .Z(II13580) ) ;
INV     gate5880  (.A(g8344), .Z(II13583) ) ;
INV     gate5881  (.A(g8356), .Z(II13586) ) ;
INV     gate5882  (.A(g8361), .Z(II13589) ) ;
INV     gate5883  (.A(g8362), .Z(II13592) ) ;
INV     gate5884  (.A(g8339), .Z(II13595) ) ;
INV     gate5885  (.A(g8311), .Z(II13606) ) ;
INV     gate5886  (.A(g8312), .Z(II13609) ) ;
INV     gate5887  (.A(g8325), .Z(II13612) ) ;
INV     gate5888  (.A(g8333), .Z(II13615) ) ;
INV     gate5889  (.A(g8345), .Z(II13618) ) ;
INV     gate5890  (.A(g8315), .Z(II13621) ) ;
INV     gate5891  (.A(g8320), .Z(II13624) ) ;
INV     gate5892  (.A(g8326), .Z(II13627) ) ;
INV     gate5893  (.A(g8334), .Z(II13630) ) ;
INV     gate5894  (.A(g8346), .Z(II13633) ) ;
INV     gate5895  (.A(g8357), .Z(II13636) ) ;
INV     gate5896  (.A(g8321), .Z(II13639) ) ;
INV     gate5897  (.A(g8378), .Z(II13642) ) ;
INV     gate5898  (.A(g8379), .Z(II13645) ) ;
INV     gate5899  (.A(g8376), .Z(II13648) ) ;
AND3    gate5900  (.A(g6777), .B(g8109), .C(g6475), .Z(g8289) ) ;
INV     gate5901  (.A(g8289), .Z(g8465) ) ;
INV     gate5902  (.A(g8292), .Z(II13666) ) ;
INV     gate5903  (.A(II13666), .Z(g8472) ) ;
INV     gate5904  (.A(g8294), .Z(II13669) ) ;
INV     gate5905  (.A(II13669), .Z(g8473) ) ;
INV     gate5906  (.A(g8314), .Z(g8475) ) ;
INV     gate5907  (.A(g8304), .Z(II13674) ) ;
INV     gate5908  (.A(II13674), .Z(g8476) ) ;
INV     gate5909  (.A(g8317), .Z(g8477) ) ;
INV     gate5910  (.A(g8306), .Z(II13678) ) ;
INV     gate5911  (.A(II13678), .Z(g8478) ) ;
INV     gate5912  (.A(g8319), .Z(g8479) ) ;
INV     gate5913  (.A(g8310), .Z(II13682) ) ;
INV     gate5914  (.A(II13682), .Z(g8480) ) ;
INV     gate5915  (.A(g8324), .Z(g8481) ) ;
INV     gate5916  (.A(g8329), .Z(g8482) ) ;
INV     gate5917  (.A(g8332), .Z(g8483) ) ;
INV     gate5918  (.A(g8336), .Z(g8484) ) ;
INV     gate5919  (.A(g8341), .Z(g8485) ) ;
INV     gate5920  (.A(g8348), .Z(g8486) ) ;
INV     gate5921  (.A(g8350), .Z(g8487) ) ;
INV     gate5922  (.A(g8353), .Z(g8498) ) ;
INV     gate5923  (.A(g8363), .Z(II13695) ) ;
INV     gate5924  (.A(II13695), .Z(g8500) ) ;
AND2    gate5925  (.A(g8199), .B(g7265), .Z(g8366) ) ;
INV     gate5926  (.A(g8366), .Z(g8509) ) ;
INV     gate5927  (.A(g8337), .Z(II13708) ) ;
INV     gate5928  (.A(II13708), .Z(g8513) ) ;
INV     gate5929  (.A(g8342), .Z(II13711) ) ;
INV     gate5930  (.A(II13711), .Z(g8514) ) ;
INV     gate5931  (.A(g8351), .Z(II13714) ) ;
INV     gate5932  (.A(II13714), .Z(g8515) ) ;
INV     gate5933  (.A(g8354), .Z(II13717) ) ;
INV     gate5934  (.A(II13717), .Z(g8516) ) ;
INV     gate5935  (.A(g8358), .Z(II13720) ) ;
INV     gate5936  (.A(II13720), .Z(g8517) ) ;
INV     gate5937  (.A(g8359), .Z(II13723) ) ;
INV     gate5938  (.A(II13723), .Z(g8518) ) ;
INV     gate5939  (.A(g8375), .Z(II13726) ) ;
INV     gate5940  (.A(II13726), .Z(g8519) ) ;
INV     gate5941  (.A(g8290), .Z(II13729) ) ;
INV     gate5942  (.A(II13729), .Z(g8520) ) ;
INV     gate5943  (.A(g8291), .Z(II13732) ) ;
INV     gate5944  (.A(II13732), .Z(g8523) ) ;
INV     gate5945  (.A(g8293), .Z(II13735) ) ;
INV     gate5946  (.A(II13735), .Z(g8526) ) ;
INV     gate5947  (.A(g8295), .Z(II13738) ) ;
INV     gate5948  (.A(II13738), .Z(g8529) ) ;
INV     gate5949  (.A(g8296), .Z(II13741) ) ;
INV     gate5950  (.A(II13741), .Z(g8532) ) ;
INV     gate5951  (.A(g8297), .Z(II13744) ) ;
INV     gate5952  (.A(II13744), .Z(g8535) ) ;
INV     gate5953  (.A(g8299), .Z(II13747) ) ;
INV     gate5954  (.A(II13747), .Z(g8538) ) ;
AND2    gate5955  (.A(g8268), .B(g6465), .Z(g8390) ) ;
INV     gate5956  (.A(g8390), .Z(g8548) ) ;
AND2    gate5957  (.A(g8180), .B(g3397), .Z(g8384) ) ;
INV     gate5958  (.A(g8384), .Z(II13773) ) ;
INV     gate5959  (.A(II13773), .Z(g8560) ) ;
INV     gate5960  (.A(g8513), .Z(II13776) ) ;
INV     gate5961  (.A(g8514), .Z(II13779) ) ;
INV     gate5962  (.A(g8515), .Z(II13782) ) ;
INV     gate5963  (.A(g8516), .Z(II13785) ) ;
INV     gate5964  (.A(g8517), .Z(II13788) ) ;
INV     gate5965  (.A(g8518), .Z(II13791) ) ;
INV     gate5966  (.A(g8472), .Z(II13794) ) ;
INV     gate5967  (.A(g8473), .Z(II13797) ) ;
INV     gate5968  (.A(g8500), .Z(II13800) ) ;
INV     gate5969  (.A(g8476), .Z(II13803) ) ;
INV     gate5970  (.A(g8478), .Z(II13806) ) ;
INV     gate5971  (.A(g8480), .Z(II13809) ) ;
INV     gate5972  (.A(g8519), .Z(II13812) ) ;
OR2     gate5973  (.A(g8380), .B(g4731), .Z(g8559) ) ;
INV     gate5974  (.A(g8559), .Z(II13816) ) ;
INV     gate5975  (.A(II13816), .Z(g8575) ) ;
OR2     gate5976  (.A(g3664), .B(g8390), .Z(g8488) ) ;
INV     gate5977  (.A(g8488), .Z(II13819) ) ;
INV     gate5978  (.A(II13819), .Z(g8576) ) ;
INV     gate5979  (.A(g8488), .Z(II13822) ) ;
INV     gate5980  (.A(II13822), .Z(g8579) ) ;
INV     gate5981  (.A(g8488), .Z(II13825) ) ;
INV     gate5982  (.A(II13825), .Z(g8582) ) ;
INV     gate5983  (.A(g8488), .Z(II13828) ) ;
INV     gate5984  (.A(II13828), .Z(g8585) ) ;
INV     gate5985  (.A(g8560), .Z(II13831) ) ;
INV     gate5986  (.A(II13831), .Z(g8588) ) ;
INV     gate5987  (.A(g8488), .Z(II13834) ) ;
INV     gate5988  (.A(II13834), .Z(g8589) ) ;
INV     gate5989  (.A(g8488), .Z(II13837) ) ;
INV     gate5990  (.A(II13837), .Z(g8592) ) ;
INV     gate5991  (.A(g8488), .Z(II13840) ) ;
INV     gate5992  (.A(II13840), .Z(g8595) ) ;
NAND2   gate5993  (.A(g3983), .B(g8390), .Z(g8546) ) ;
INV     gate5994  (.A(g8546), .Z(g8599) ) ;
INV     gate5995  (.A(g8475), .Z(g8600) ) ;
INV     gate5996  (.A(g8477), .Z(g8601) ) ;
INV     gate5997  (.A(g8479), .Z(g8604) ) ;
INV     gate5998  (.A(g8481), .Z(g8606) ) ;
INV     gate5999  (.A(g8482), .Z(g8608) ) ;
INV     gate6000  (.A(g8483), .Z(g8610) ) ;
INV     gate6001  (.A(g8484), .Z(g8613) ) ;
INV     gate6002  (.A(g8465), .Z(g8617) ) ;
INV     gate6003  (.A(g8485), .Z(g8622) ) ;
INV     gate6004  (.A(g8486), .Z(g8624) ) ;
INV     gate6005  (.A(g8487), .Z(g8625) ) ;
INV     gate6006  (.A(g8498), .Z(g8626) ) ;
OR2     gate6007  (.A(g3440), .B(g8366), .Z(g8451) ) ;
INV     gate6008  (.A(g8451), .Z(II13915) ) ;
INV     gate6009  (.A(II13915), .Z(g8632) ) ;
INV     gate6010  (.A(g8451), .Z(II13918) ) ;
INV     gate6011  (.A(II13918), .Z(g8635) ) ;
NAND2   gate6012  (.A(g3723), .B(g8366), .Z(g8512) ) ;
INV     gate6013  (.A(g8512), .Z(g8640) ) ;
AND2    gate6014  (.A(g8309), .B(g4789), .Z(g8505) ) ;
INV     gate6015  (.A(g8505), .Z(II13933) ) ;
INV     gate6016  (.A(II13933), .Z(g8650) ) ;
INV     gate6017  (.A(g8488), .Z(II13941) ) ;
INV     gate6018  (.A(II13941), .Z(g8656) ) ;
INV     gate6019  (.A(g8488), .Z(II13945) ) ;
INV     gate6020  (.A(II13945), .Z(g8660) ) ;
INV     gate6021  (.A(g8451), .Z(II13949) ) ;
INV     gate6022  (.A(II13949), .Z(g8664) ) ;
INV     gate6023  (.A(g8451), .Z(II13952) ) ;
INV     gate6024  (.A(II13952), .Z(g8667) ) ;
NAND2   gate6025  (.A(g3967), .B(g8390), .Z(g8551) ) ;
INV     gate6026  (.A(g8551), .Z(g8670) ) ;
INV     gate6027  (.A(g8451), .Z(II13956) ) ;
INV     gate6028  (.A(II13956), .Z(g8671) ) ;
INV     gate6029  (.A(g8451), .Z(II13959) ) ;
INV     gate6030  (.A(II13959), .Z(g8674) ) ;
INV     gate6031  (.A(g8451), .Z(II13962) ) ;
INV     gate6032  (.A(II13962), .Z(g8677) ) ;
INV     gate6033  (.A(g8451), .Z(II13965) ) ;
INV     gate6034  (.A(II13965), .Z(g8680) ) ;
INV     gate6035  (.A(g8451), .Z(II13969) ) ;
INV     gate6036  (.A(II13969), .Z(g8684) ) ;
NAND2   gate6037  (.A(g3738), .B(g8366), .Z(g8507) ) ;
INV     gate6038  (.A(g8507), .Z(g8688) ) ;
INV     gate6039  (.A(g8588), .Z(II13975) ) ;
INV     gate6040  (.A(g8575), .Z(II13978) ) ;
INV     gate6041  (.A(g8656), .Z(g8696) ) ;
INV     gate6042  (.A(g8660), .Z(g8697) ) ;
OR3     gate6043  (.A(g5679), .B(g7853), .C(g8465), .Z(g8574) ) ;
INV     gate6044  (.A(g8574), .Z(g8700) ) ;
INV     gate6045  (.A(g8664), .Z(g8702) ) ;
INV     gate6046  (.A(g8667), .Z(g8704) ) ;
INV     gate6047  (.A(g8671), .Z(g8707) ) ;
INV     gate6048  (.A(g8674), .Z(g8709) ) ;
INV     gate6049  (.A(g8677), .Z(g8711) ) ;
INV     gate6050  (.A(g8680), .Z(g8712) ) ;
INV     gate6051  (.A(g8684), .Z(g8713) ) ;
OR2     gate6052  (.A(g8474), .B(g7449), .Z(g8631) ) ;
INV     gate6053  (.A(g8631), .Z(II14005) ) ;
INV     gate6054  (.A(II14005), .Z(g8714) ) ;
INV     gate6055  (.A(g8576), .Z(g8716) ) ;
OR3     gate6056  (.A(g5236), .B(g5205), .C(g8465), .Z(g8642) ) ;
INV     gate6057  (.A(g8642), .Z(II14010) ) ;
INV     gate6058  (.A(II14010), .Z(g8717) ) ;
INV     gate6059  (.A(g8579), .Z(g8719) ) ;
INV     gate6060  (.A(g8582), .Z(g8721) ) ;
INV     gate6061  (.A(g8585), .Z(g8723) ) ;
INV     gate6062  (.A(g8589), .Z(g8725) ) ;
INV     gate6063  (.A(g8592), .Z(g8727) ) ;
INV     gate6064  (.A(g8595), .Z(g8729) ) ;
INV     gate6065  (.A(g8640), .Z(g8739) ) ;
OR2     gate6066  (.A(g8499), .B(g4519), .Z(g8649) ) ;
INV     gate6067  (.A(g8649), .Z(II14040) ) ;
INV     gate6068  (.A(II14040), .Z(g8747) ) ;
AND2    gate6069  (.A(g3983), .B(g8548), .Z(g8603) ) ;
INV     gate6070  (.A(g8603), .Z(II14045) ) ;
INV     gate6071  (.A(II14045), .Z(g8750) ) ;
INV     gate6072  (.A(g8632), .Z(g8751) ) ;
INV     gate6073  (.A(g8635), .Z(g8752) ) ;
INV     gate6074  (.A(g8650), .Z(II14055) ) ;
INV     gate6075  (.A(II14055), .Z(g8758) ) ;
INV     gate6076  (.A(g8670), .Z(g8760) ) ;
INV     gate6077  (.A(g8758), .Z(II14077) ) ;
INV     gate6078  (.A(g8714), .Z(II14080) ) ;
INV     gate6079  (.A(g8747), .Z(II14083) ) ;
NAND3   gate6080  (.A(g8617), .B(g6517), .C(g6509), .Z(g8746) ) ;
INV     gate6081  (.A(g8746), .Z(g8783) ) ;
OR2     gate6082  (.A(g5476), .B(g8651), .Z(g8770) ) ;
INV     gate6083  (.A(g8770), .Z(II14087) ) ;
INV     gate6084  (.A(II14087), .Z(g8784) ) ;
OR2     gate6085  (.A(g5483), .B(g8652), .Z(g8771) ) ;
INV     gate6086  (.A(g8771), .Z(II14090) ) ;
INV     gate6087  (.A(II14090), .Z(g8785) ) ;
INV     gate6088  (.A(g8700), .Z(II14094) ) ;
INV     gate6089  (.A(II14094), .Z(g8787) ) ;
OR2     gate6090  (.A(g5491), .B(g8653), .Z(g8773) ) ;
INV     gate6091  (.A(g8773), .Z(II14097) ) ;
INV     gate6092  (.A(II14097), .Z(g8788) ) ;
OR2     gate6093  (.A(g5499), .B(g8654), .Z(g8774) ) ;
INV     gate6094  (.A(g8774), .Z(II14101) ) ;
INV     gate6095  (.A(II14101), .Z(g8790) ) ;
OR2     gate6096  (.A(g5510), .B(g8655), .Z(g8776) ) ;
INV     gate6097  (.A(g8776), .Z(II14105) ) ;
INV     gate6098  (.A(II14105), .Z(g8792) ) ;
AND2    gate6099  (.A(g8630), .B(g5151), .Z(g8765) ) ;
INV     gate6100  (.A(g8765), .Z(II14109) ) ;
INV     gate6101  (.A(II14109), .Z(g8794) ) ;
OR2     gate6102  (.A(g5522), .B(g8659), .Z(g8777) ) ;
INV     gate6103  (.A(g8777), .Z(II14112) ) ;
INV     gate6104  (.A(II14112), .Z(g8795) ) ;
AND2    gate6105  (.A(g8612), .B(g5151), .Z(g8766) ) ;
INV     gate6106  (.A(g8766), .Z(II14116) ) ;
INV     gate6107  (.A(II14116), .Z(g8797) ) ;
OR2     gate6108  (.A(g5530), .B(g8663), .Z(g8779) ) ;
INV     gate6109  (.A(g8779), .Z(II14119) ) ;
INV     gate6110  (.A(II14119), .Z(g8798) ) ;
AND2    gate6111  (.A(g8616), .B(g5151), .Z(g8767) ) ;
INV     gate6112  (.A(g8767), .Z(II14123) ) ;
INV     gate6113  (.A(II14123), .Z(g8800) ) ;
AND2    gate6114  (.A(g8623), .B(g5151), .Z(g8768) ) ;
INV     gate6115  (.A(g8768), .Z(II14127) ) ;
INV     gate6116  (.A(II14127), .Z(g8802) ) ;
AND2    gate6117  (.A(g8629), .B(g5151), .Z(g8769) ) ;
INV     gate6118  (.A(g8769), .Z(II14130) ) ;
INV     gate6119  (.A(II14130), .Z(g8803) ) ;
AND2    gate6120  (.A(g8627), .B(g5151), .Z(g8772) ) ;
INV     gate6121  (.A(g8772), .Z(II14133) ) ;
INV     gate6122  (.A(II14133), .Z(g8804) ) ;
AND2    gate6123  (.A(g8628), .B(g5151), .Z(g8775) ) ;
INV     gate6124  (.A(g8775), .Z(II14136) ) ;
INV     gate6125  (.A(II14136), .Z(g8805) ) ;
INV     gate6126  (.A(g8717), .Z(II14140) ) ;
INV     gate6127  (.A(II14140), .Z(g8807) ) ;
NAND3   gate6128  (.A(g8617), .B(g6509), .C(g6971), .Z(g8744) ) ;
INV     gate6129  (.A(g8744), .Z(g8828) ) ;
NAND3   gate6130  (.A(g8617), .B(g6517), .C(g6964), .Z(g8745) ) ;
INV     gate6131  (.A(g8745), .Z(g8849) ) ;
NAND3   gate6132  (.A(g8617), .B(g6971), .C(g6964), .Z(g8743) ) ;
INV     gate6133  (.A(g8743), .Z(g8858) ) ;
INV     gate6134  (.A(g8784), .Z(II14176) ) ;
INV     gate6135  (.A(g8785), .Z(II14179) ) ;
INV     gate6136  (.A(g8788), .Z(II14182) ) ;
INV     gate6137  (.A(g8790), .Z(II14185) ) ;
INV     gate6138  (.A(g8792), .Z(II14188) ) ;
INV     gate6139  (.A(g8795), .Z(II14191) ) ;
INV     gate6140  (.A(g8798), .Z(II14194) ) ;
INV     gate6141  (.A(g8794), .Z(II14224) ) ;
INV     gate6142  (.A(II14224), .Z(g8884) ) ;
INV     gate6143  (.A(g8797), .Z(II14228) ) ;
INV     gate6144  (.A(II14228), .Z(g8886) ) ;
INV     gate6145  (.A(g8800), .Z(II14232) ) ;
INV     gate6146  (.A(II14232), .Z(g8888) ) ;
INV     gate6147  (.A(g8802), .Z(II14236) ) ;
INV     gate6148  (.A(II14236), .Z(g8890) ) ;
INV     gate6149  (.A(g8803), .Z(II14239) ) ;
INV     gate6150  (.A(II14239), .Z(g8891) ) ;
INV     gate6151  (.A(g8787), .Z(II14242) ) ;
INV     gate6152  (.A(II14242), .Z(g8892) ) ;
INV     gate6153  (.A(g8804), .Z(II14249) ) ;
INV     gate6154  (.A(II14249), .Z(g8924) ) ;
INV     gate6155  (.A(g8783), .Z(II14252) ) ;
INV     gate6156  (.A(II14252), .Z(g8925) ) ;
INV     gate6157  (.A(g8805), .Z(II14257) ) ;
INV     gate6158  (.A(II14257), .Z(g8928) ) ;
OR2     gate6159  (.A(g7931), .B(g8718), .Z(g8806) ) ;
INV     gate6160  (.A(g8806), .Z(II14295) ) ;
INV     gate6161  (.A(II14295), .Z(g8946) ) ;
OR2     gate6162  (.A(g7933), .B(g8720), .Z(g8810) ) ;
INV     gate6163  (.A(g8810), .Z(II14299) ) ;
INV     gate6164  (.A(II14299), .Z(g8948) ) ;
OR2     gate6165  (.A(g7935), .B(g8722), .Z(g8811) ) ;
INV     gate6166  (.A(g8811), .Z(II14303) ) ;
INV     gate6167  (.A(II14303), .Z(g8950) ) ;
OR2     gate6168  (.A(g7939), .B(g8724), .Z(g8812) ) ;
INV     gate6169  (.A(g8812), .Z(II14306) ) ;
INV     gate6170  (.A(II14306), .Z(g8951) ) ;
OR2     gate6171  (.A(g7943), .B(g8726), .Z(g8813) ) ;
INV     gate6172  (.A(g8813), .Z(II14309) ) ;
INV     gate6173  (.A(II14309), .Z(g8952) ) ;
OR2     gate6174  (.A(g7945), .B(g8728), .Z(g8814) ) ;
INV     gate6175  (.A(g8814), .Z(II14312) ) ;
INV     gate6176  (.A(II14312), .Z(g8953) ) ;
OR2     gate6177  (.A(g7948), .B(g8730), .Z(g8815) ) ;
INV     gate6178  (.A(g8815), .Z(II14315) ) ;
INV     gate6179  (.A(II14315), .Z(g8954) ) ;
OR2     gate6180  (.A(g7951), .B(g8731), .Z(g8816) ) ;
INV     gate6181  (.A(g8816), .Z(II14319) ) ;
INV     gate6182  (.A(II14319), .Z(g8956) ) ;
OR2     gate6183  (.A(g7954), .B(g8732), .Z(g8817) ) ;
INV     gate6184  (.A(g8817), .Z(II14323) ) ;
INV     gate6185  (.A(II14323), .Z(g8958) ) ;
OR2     gate6186  (.A(g7955), .B(g8733), .Z(g8818) ) ;
INV     gate6187  (.A(g8818), .Z(II14326) ) ;
INV     gate6188  (.A(II14326), .Z(g8959) ) ;
OR2     gate6189  (.A(g7957), .B(g8734), .Z(g8819) ) ;
INV     gate6190  (.A(g8819), .Z(II14330) ) ;
INV     gate6191  (.A(II14330), .Z(g8961) ) ;
AND2    gate6192  (.A(g8705), .B(g5422), .Z(g8820) ) ;
INV     gate6193  (.A(g8820), .Z(II14340) ) ;
INV     gate6194  (.A(II14340), .Z(g8969) ) ;
INV     gate6195  (.A(g8958), .Z(II14349) ) ;
INV     gate6196  (.A(g8946), .Z(II14352) ) ;
INV     gate6197  (.A(g8948), .Z(II14355) ) ;
INV     gate6198  (.A(g8950), .Z(II14358) ) ;
INV     gate6199  (.A(g8951), .Z(II14361) ) ;
INV     gate6200  (.A(g8952), .Z(II14364) ) ;
INV     gate6201  (.A(g8953), .Z(II14367) ) ;
INV     gate6202  (.A(g8954), .Z(II14370) ) ;
INV     gate6203  (.A(g8956), .Z(II14373) ) ;
INV     gate6204  (.A(g8959), .Z(II14376) ) ;
INV     gate6205  (.A(g8961), .Z(II14379) ) ;
INV     gate6206  (.A(g8886), .Z(II14382) ) ;
INV     gate6207  (.A(g8890), .Z(II14385) ) ;
INV     gate6208  (.A(g8924), .Z(II14388) ) ;
INV     gate6209  (.A(g8928), .Z(II14391) ) ;
INV     gate6210  (.A(g8884), .Z(II14394) ) ;
INV     gate6211  (.A(g8888), .Z(II14397) ) ;
INV     gate6212  (.A(g8891), .Z(II14400) ) ;
OR2     gate6213  (.A(g8786), .B(g8698), .Z(g8937) ) ;
INV     gate6214  (.A(g8937), .Z(II14405) ) ;
INV     gate6215  (.A(II14405), .Z(g9009) ) ;
OR2     gate6216  (.A(g8789), .B(g8699), .Z(g8938) ) ;
INV     gate6217  (.A(g8938), .Z(II14409) ) ;
INV     gate6218  (.A(II14409), .Z(g9024) ) ;
OR2     gate6219  (.A(g8791), .B(g8701), .Z(g8939) ) ;
INV     gate6220  (.A(g8939), .Z(II14412) ) ;
INV     gate6221  (.A(II14412), .Z(g9025) ) ;
OR2     gate6222  (.A(g8793), .B(g8703), .Z(g8940) ) ;
INV     gate6223  (.A(g8940), .Z(II14415) ) ;
INV     gate6224  (.A(II14415), .Z(g9026) ) ;
OR2     gate6225  (.A(g8796), .B(g8706), .Z(g8941) ) ;
INV     gate6226  (.A(g8941), .Z(II14418) ) ;
INV     gate6227  (.A(II14418), .Z(g9027) ) ;
OR2     gate6228  (.A(g8799), .B(g8708), .Z(g8944) ) ;
INV     gate6229  (.A(g8944), .Z(II14421) ) ;
INV     gate6230  (.A(II14421), .Z(g9028) ) ;
OR2     gate6231  (.A(g8801), .B(g8710), .Z(g8945) ) ;
INV     gate6232  (.A(g8945), .Z(II14424) ) ;
INV     gate6233  (.A(II14424), .Z(g9029) ) ;
INV     gate6234  (.A(g8892), .Z(g9076) ) ;
INV     gate6235  (.A(g8892), .Z(g9079) ) ;
INV     gate6236  (.A(g8892), .Z(g9082) ) ;
INV     gate6237  (.A(g8892), .Z(g9085) ) ;
INV     gate6238  (.A(g8892), .Z(g9091) ) ;
INV     gate6239  (.A(g8892), .Z(g9094) ) ;
INV     gate6240  (.A(g8892), .Z(g9097) ) ;
INV     gate6241  (.A(g8892), .Z(g9100) ) ;
INV     gate6242  (.A(g8892), .Z(g9103) ) ;
INV     gate6243  (.A(g8969), .Z(II14439) ) ;
INV     gate6244  (.A(II14439), .Z(g9106) ) ;
OR2     gate6245  (.A(g8821), .B(g8735), .Z(g8973) ) ;
INV     gate6246  (.A(g8973), .Z(II14449) ) ;
INV     gate6247  (.A(II14449), .Z(g9108) ) ;
OR2     gate6248  (.A(g8822), .B(g8736), .Z(g8922) ) ;
INV     gate6249  (.A(g8922), .Z(II14452) ) ;
INV     gate6250  (.A(II14452), .Z(g9109) ) ;
INV     gate6251  (.A(g8892), .Z(g9258) ) ;
INV     gate6252  (.A(g8892), .Z(g9259) ) ;
INV     gate6253  (.A(g8892), .Z(g9260) ) ;
INV     gate6254  (.A(g8892), .Z(g9261) ) ;
OR2     gate6255  (.A(g8827), .B(g8748), .Z(g8921) ) ;
INV     gate6256  (.A(g8921), .Z(II14473) ) ;
INV     gate6257  (.A(II14473), .Z(g9262) ) ;
INV     gate6258  (.A(g8892), .Z(g9263) ) ;
OR2     gate6259  (.A(g8837), .B(g8749), .Z(g8943) ) ;
INV     gate6260  (.A(g8943), .Z(II14477) ) ;
INV     gate6261  (.A(II14477), .Z(g9264) ) ;
INV     gate6262  (.A(g8892), .Z(g9265) ) ;
INV     gate6263  (.A(g8892), .Z(g9267) ) ;
OR2     gate6264  (.A(g8838), .B(g8753), .Z(g8883) ) ;
INV     gate6265  (.A(g8883), .Z(II14485) ) ;
INV     gate6266  (.A(II14485), .Z(g9270) ) ;
OR2     gate6267  (.A(g8841), .B(g8754), .Z(g8885) ) ;
INV     gate6268  (.A(g8885), .Z(II14490) ) ;
INV     gate6269  (.A(II14490), .Z(g9273) ) ;
OR2     gate6270  (.A(g8842), .B(g8755), .Z(g8887) ) ;
INV     gate6271  (.A(g8887), .Z(II14494) ) ;
INV     gate6272  (.A(II14494), .Z(g9290) ) ;
INV     gate6273  (.A(g8892), .Z(g9291) ) ;
OR2     gate6274  (.A(g8844), .B(g8756), .Z(g8889) ) ;
INV     gate6275  (.A(g8889), .Z(II14499) ) ;
INV     gate6276  (.A(II14499), .Z(g9308) ) ;
INV     gate6277  (.A(g8892), .Z(g9309) ) ;
OR2     gate6278  (.A(g8845), .B(g8759), .Z(g8920) ) ;
INV     gate6279  (.A(g8920), .Z(II14503) ) ;
INV     gate6280  (.A(II14503), .Z(g9310) ) ;
OR2     gate6281  (.A(g8846), .B(g8763), .Z(g8923) ) ;
INV     gate6282  (.A(g8923), .Z(II14506) ) ;
INV     gate6283  (.A(II14506), .Z(g9311) ) ;
OR2     gate6284  (.A(g8848), .B(g8764), .Z(g8926) ) ;
INV     gate6285  (.A(g8926), .Z(II14509) ) ;
INV     gate6286  (.A(II14509), .Z(g9312) ) ;
INV     gate6287  (.A(g9106), .Z(II14519) ) ;
INV     gate6288  (.A(g9108), .Z(II14522) ) ;
INV     gate6289  (.A(g9109), .Z(II14525) ) ;
INV     gate6290  (.A(g9270), .Z(II14528) ) ;
INV     gate6291  (.A(g9273), .Z(II14531) ) ;
INV     gate6292  (.A(g9290), .Z(II14534) ) ;
INV     gate6293  (.A(g9308), .Z(II14537) ) ;
INV     gate6294  (.A(g9310), .Z(II14540) ) ;
INV     gate6295  (.A(g9311), .Z(II14543) ) ;
INV     gate6296  (.A(g9312), .Z(II14546) ) ;
INV     gate6297  (.A(g9262), .Z(II14549) ) ;
INV     gate6298  (.A(g9264), .Z(II14552) ) ;
INV     gate6299  (.A(g9009), .Z(II14555) ) ;
INV     gate6300  (.A(g9024), .Z(II14558) ) ;
INV     gate6301  (.A(g9025), .Z(II14561) ) ;
INV     gate6302  (.A(g9026), .Z(II14564) ) ;
INV     gate6303  (.A(g9027), .Z(II14567) ) ;
INV     gate6304  (.A(g9028), .Z(II14570) ) ;
INV     gate6305  (.A(g9029), .Z(II14573) ) ;
AND2    gate6306  (.A(g8934), .B(g3424), .Z(g9272) ) ;
INV     gate6307  (.A(g9272), .Z(II14579) ) ;
INV     gate6308  (.A(II14579), .Z(g9360) ) ;
INV     gate6309  (.A(g9076), .Z(g9424) ) ;
INV     gate6310  (.A(g9079), .Z(g9427) ) ;
INV     gate6311  (.A(g9082), .Z(g9429) ) ;
INV     gate6312  (.A(g9085), .Z(g9431) ) ;
AND2    gate6313  (.A(g8876), .B(g5708), .Z(g9313) ) ;
INV     gate6314  (.A(g9313), .Z(g9432) ) ;
INV     gate6315  (.A(g9091), .Z(g9448) ) ;
INV     gate6316  (.A(g9094), .Z(g9449) ) ;
INV     gate6317  (.A(g9097), .Z(g9450) ) ;
OR2     gate6318  (.A(g8927), .B(g8381), .Z(g9088) ) ;
INV     gate6319  (.A(g9088), .Z(II14642) ) ;
INV     gate6320  (.A(g9088), .Z(II14645) ) ;
INV     gate6321  (.A(II14645), .Z(g9452) ) ;
INV     gate6322  (.A(g9100), .Z(g9453) ) ;
INV     gate6323  (.A(g9103), .Z(g9473) ) ;
AND2    gate6324  (.A(g8972), .B(g5708), .Z(g9331) ) ;
INV     gate6325  (.A(g9331), .Z(g9474) ) ;
AND2    gate6326  (.A(g8879), .B(g5708), .Z(g9324) ) ;
INV     gate6327  (.A(g9324), .Z(g9490) ) ;
AND2    gate6328  (.A(g8936), .B(g7192), .Z(g9052) ) ;
INV     gate6329  (.A(g9052), .Z(g9505) ) ;
AND2    gate6330  (.A(g6681), .B(g8947), .Z(g9268) ) ;
INV     gate6331  (.A(g9268), .Z(g9507) ) ;
AND2    gate6332  (.A(g6681), .B(g8949), .Z(g9271) ) ;
INV     gate6333  (.A(g9271), .Z(g9508) ) ;
AND2    gate6334  (.A(g6689), .B(g8964), .Z(g9257) ) ;
INV     gate6335  (.A(g9257), .Z(g9525) ) ;
AND2    gate6336  (.A(g6689), .B(g8963), .Z(g9256) ) ;
INV     gate6337  (.A(g9256), .Z(g9526) ) ;
INV     gate6338  (.A(g9309), .Z(II14668) ) ;
INV     gate6339  (.A(II14668), .Z(g9527) ) ;
INV     gate6340  (.A(g9261), .Z(II14672) ) ;
INV     gate6341  (.A(II14672), .Z(g9529) ) ;
INV     gate6342  (.A(g9263), .Z(II14675) ) ;
INV     gate6343  (.A(II14675), .Z(g9530) ) ;
INV     gate6344  (.A(g9265), .Z(II14678) ) ;
INV     gate6345  (.A(II14678), .Z(g9531) ) ;
AND2    gate6346  (.A(g8880), .B(g4790), .Z(g9110) ) ;
INV     gate6347  (.A(g9110), .Z(II14681) ) ;
INV     gate6348  (.A(II14681), .Z(g9532) ) ;
AND2    gate6349  (.A(g8881), .B(g4802), .Z(g9124) ) ;
INV     gate6350  (.A(g9124), .Z(II14684) ) ;
INV     gate6351  (.A(II14684), .Z(g9533) ) ;
INV     gate6352  (.A(g9258), .Z(II14687) ) ;
INV     gate6353  (.A(II14687), .Z(g9534) ) ;
AND2    gate6354  (.A(g8882), .B(g4805), .Z(g9150) ) ;
INV     gate6355  (.A(g9150), .Z(II14690) ) ;
INV     gate6356  (.A(II14690), .Z(g9535) ) ;
INV     gate6357  (.A(g9259), .Z(II14694) ) ;
INV     gate6358  (.A(II14694), .Z(g9553) ) ;
INV     gate6359  (.A(g9260), .Z(II14697) ) ;
INV     gate6360  (.A(II14697), .Z(g9554) ) ;
INV     gate6361  (.A(g9291), .Z(II14701) ) ;
INV     gate6362  (.A(II14701), .Z(g9556) ) ;
INV     gate6363  (.A(g9267), .Z(II14709) ) ;
INV     gate6364  (.A(II14709), .Z(g9572) ) ;
INV     gate6365  (.A(g9052), .Z(II14713) ) ;
INV     gate6366  (.A(II14713), .Z(g9576) ) ;
AND2    gate6367  (.A(g8932), .B(g3398), .Z(g9266) ) ;
INV     gate6368  (.A(g9266), .Z(II14786) ) ;
INV     gate6369  (.A(II14786), .Z(g9661) ) ;
AND2    gate6370  (.A(g8933), .B(g3413), .Z(g9269) ) ;
INV     gate6371  (.A(g9269), .Z(II14793) ) ;
INV     gate6372  (.A(II14793), .Z(g9666) ) ;
INV     gate6373  (.A(g9490), .Z(g9668) ) ;
INV     gate6374  (.A(g9661), .Z(II14799) ) ;
INV     gate6375  (.A(II14799), .Z(g9670) ) ;
INV     gate6376  (.A(g9666), .Z(II14802) ) ;
INV     gate6377  (.A(II14802), .Z(g9671) ) ;
INV     gate6378  (.A(g9360), .Z(II14805) ) ;
INV     gate6379  (.A(II14805), .Z(g9672) ) ;
INV     gate6380  (.A(g9452), .Z(g9679) ) ;
INV     gate6381  (.A(g9525), .Z(II14873) ) ;
INV     gate6382  (.A(II14873), .Z(g9732) ) ;
INV     gate6383  (.A(g9526), .Z(II14876) ) ;
INV     gate6384  (.A(II14876), .Z(g9733) ) ;
AND2    gate6385  (.A(g8994), .B(g5708), .Z(g9454) ) ;
INV     gate6386  (.A(g9454), .Z(II14884) ) ;
INV     gate6387  (.A(II14884), .Z(g9739) ) ;
INV     gate6388  (.A(g9454), .Z(II14888) ) ;
INV     gate6389  (.A(II14888), .Z(g9741) ) ;
INV     gate6390  (.A(g9454), .Z(g9745) ) ;
INV     gate6391  (.A(g9454), .Z(g9760) ) ;
INV     gate6392  (.A(g9454), .Z(g9761) ) ;
INV     gate6393  (.A(g9507), .Z(II14903) ) ;
INV     gate6394  (.A(II14903), .Z(g9762) ) ;
INV     gate6395  (.A(g9508), .Z(II14906) ) ;
INV     gate6396  (.A(II14906), .Z(g9763) ) ;
INV     gate6397  (.A(g9432), .Z(g9764) ) ;
INV     gate6398  (.A(g9532), .Z(II14910) ) ;
INV     gate6399  (.A(II14910), .Z(g9765) ) ;
INV     gate6400  (.A(g9432), .Z(g9766) ) ;
INV     gate6401  (.A(g9533), .Z(II14914) ) ;
INV     gate6402  (.A(II14914), .Z(g9767) ) ;
INV     gate6403  (.A(g9432), .Z(g9768) ) ;
INV     gate6404  (.A(g9535), .Z(II14918) ) ;
INV     gate6405  (.A(II14918), .Z(g9769) ) ;
INV     gate6406  (.A(g9432), .Z(g9770) ) ;
INV     gate6407  (.A(g9432), .Z(g9771) ) ;
INV     gate6408  (.A(g9432), .Z(g9772) ) ;
INV     gate6409  (.A(g9474), .Z(g9773) ) ;
INV     gate6410  (.A(g9474), .Z(g9774) ) ;
INV     gate6411  (.A(g9474), .Z(g9775) ) ;
INV     gate6412  (.A(g9474), .Z(g9777) ) ;
INV     gate6413  (.A(g9474), .Z(g9778) ) ;
INV     gate6414  (.A(g9474), .Z(g9780) ) ;
INV     gate6415  (.A(g9454), .Z(II14933) ) ;
INV     gate6416  (.A(II14933), .Z(g9782) ) ;
INV     gate6417  (.A(g9490), .Z(g9802) ) ;
INV     gate6418  (.A(g9454), .Z(II14939) ) ;
INV     gate6419  (.A(II14939), .Z(g9804) ) ;
INV     gate6420  (.A(g9490), .Z(g9807) ) ;
INV     gate6421  (.A(g9454), .Z(II14944) ) ;
INV     gate6422  (.A(II14944), .Z(g9809) ) ;
INV     gate6423  (.A(g9490), .Z(g9812) ) ;
AND2    gate6424  (.A(g9107), .B(g3391), .Z(g9555) ) ;
INV     gate6425  (.A(g9555), .Z(II14948) ) ;
INV     gate6426  (.A(II14948), .Z(g9813) ) ;
INV     gate6427  (.A(g9490), .Z(g9814) ) ;
INV     gate6428  (.A(g9490), .Z(g9816) ) ;
INV     gate6429  (.A(g9765), .Z(II14955) ) ;
INV     gate6430  (.A(g9767), .Z(II14958) ) ;
INV     gate6431  (.A(g9769), .Z(II14961) ) ;
INV     gate6432  (.A(g9762), .Z(II14964) ) ;
INV     gate6433  (.A(g9763), .Z(II14967) ) ;
INV     gate6434  (.A(g9732), .Z(II14970) ) ;
INV     gate6435  (.A(g9733), .Z(II14973) ) ;
INV     gate6436  (.A(g9670), .Z(II14976) ) ;
INV     gate6437  (.A(g9671), .Z(II14979) ) ;
INV     gate6438  (.A(g9672), .Z(II14982) ) ;
INV     gate6439  (.A(g9813), .Z(II14989) ) ;
INV     gate6440  (.A(II14989), .Z(g9832) ) ;
INV     gate6441  (.A(g9679), .Z(g9845) ) ;
AND2    gate6442  (.A(g9413), .B(g4785), .Z(g9721) ) ;
INV     gate6443  (.A(g9721), .Z(II15036) ) ;
INV     gate6444  (.A(II15036), .Z(g9875) ) ;
AND2    gate6445  (.A(g281), .B(g9432), .Z(g9696) ) ;
INV     gate6446  (.A(g9696), .Z(II15060) ) ;
INV     gate6447  (.A(II15060), .Z(g9883) ) ;
AND2    gate6448  (.A(g284), .B(g9432), .Z(g9699) ) ;
INV     gate6449  (.A(g9699), .Z(II15063) ) ;
INV     gate6450  (.A(II15063), .Z(g9884) ) ;
AND2    gate6451  (.A(g1586), .B(g9474), .Z(g9710) ) ;
INV     gate6452  (.A(g9710), .Z(II15068) ) ;
INV     gate6453  (.A(II15068), .Z(g9887) ) ;
AND2    gate6454  (.A(g1589), .B(g9474), .Z(g9713) ) ;
INV     gate6455  (.A(g9713), .Z(II15072) ) ;
INV     gate6456  (.A(II15072), .Z(g9889) ) ;
INV     gate6457  (.A(g9761), .Z(II15075) ) ;
INV     gate6458  (.A(II15075), .Z(g9890) ) ;
INV     gate6459  (.A(g9745), .Z(II15079) ) ;
INV     gate6460  (.A(II15079), .Z(g9892) ) ;
AND2    gate6461  (.A(g1543), .B(g9490), .Z(g9719) ) ;
INV     gate6462  (.A(g9719), .Z(II15082) ) ;
INV     gate6463  (.A(II15082), .Z(g9893) ) ;
AND2    gate6464  (.A(g1546), .B(g9490), .Z(g9720) ) ;
INV     gate6465  (.A(g9720), .Z(II15085) ) ;
INV     gate6466  (.A(II15085), .Z(g9894) ) ;
INV     gate6467  (.A(g9832), .Z(II15088) ) ;
INV     gate6468  (.A(g9875), .Z(II15114) ) ;
INV     gate6469  (.A(II15114), .Z(g9919) ) ;
INV     gate6470  (.A(g9919), .Z(II15127) ) ;
OR2     gate6471  (.A(g8931), .B(g9900), .Z(g9931) ) ;
INV     gate6472  (.A(g9931), .Z(II15157) ) ;
INV     gate6473  (.A(II15157), .Z(g9958) ) ;
INV     gate6474  (.A(g9958), .Z(II15162) ) ;
OR2     gate6475  (.A(II15171), .B(II15172), .Z(g9968) ) ;
INV     gate6476  (.A(g9968), .Z(II15181) ) ;
INV     gate6477  (.A(II15181), .Z(g9980) ) ;
OR2     gate6478  (.A(II15176), .B(II15177), .Z(g9974) ) ;
INV     gate6479  (.A(g9974), .Z(II15184) ) ;
INV     gate6480  (.A(II15184), .Z(g9984) ) ;
INV     gate6481  (.A(g9968), .Z(II15187) ) ;
INV     gate6482  (.A(II15187), .Z(g9987) ) ;
INV     gate6483  (.A(g9974), .Z(II15190) ) ;
INV     gate6484  (.A(II15190), .Z(g9990) ) ;
INV     gate6485  (.A(g9968), .Z(II15193) ) ;
INV     gate6486  (.A(II15193), .Z(g9993) ) ;
INV     gate6487  (.A(g9974), .Z(II15196) ) ;
INV     gate6488  (.A(II15196), .Z(g9994) ) ;
INV     gate6489  (.A(g9968), .Z(II15229) ) ;
INV     gate6490  (.A(II15229), .Z(g10031) ) ;
INV     gate6491  (.A(g9974), .Z(II15232) ) ;
INV     gate6492  (.A(II15232), .Z(g10032) ) ;
INV     gate6493  (.A(g9968), .Z(II15235) ) ;
INV     gate6494  (.A(II15235), .Z(g10033) ) ;
INV     gate6495  (.A(g9974), .Z(II15238) ) ;
INV     gate6496  (.A(II15238), .Z(g10034) ) ;
OR2     gate6497  (.A(II15214), .B(II15215), .Z(g10013) ) ;
INV     gate6498  (.A(g10013), .Z(II15241) ) ;
INV     gate6499  (.A(II15241), .Z(g10035) ) ;
INV     gate6500  (.A(g10031), .Z(II15244) ) ;
INV     gate6501  (.A(II15244), .Z(g10039) ) ;
INV     gate6502  (.A(g10032), .Z(II15247) ) ;
INV     gate6503  (.A(II15247), .Z(g10040) ) ;
INV     gate6504  (.A(g9980), .Z(II15250) ) ;
INV     gate6505  (.A(II15250), .Z(g10041) ) ;
INV     gate6506  (.A(g9987), .Z(II15253) ) ;
INV     gate6507  (.A(II15253), .Z(g10042) ) ;
OR2     gate6508  (.A(II15199), .B(II15200), .Z(g9995) ) ;
INV     gate6509  (.A(g9995), .Z(II15263) ) ;
INV     gate6510  (.A(II15263), .Z(g10044) ) ;
OR2     gate6511  (.A(II15204), .B(II15205), .Z(g10001) ) ;
INV     gate6512  (.A(g10001), .Z(II15266) ) ;
INV     gate6513  (.A(II15266), .Z(g10047) ) ;
INV     gate6514  (.A(g9993), .Z(II15269) ) ;
INV     gate6515  (.A(II15269), .Z(g10050) ) ;
OR2     gate6516  (.A(II15219), .B(II15220), .Z(g10019) ) ;
INV     gate6517  (.A(g10019), .Z(II15272) ) ;
INV     gate6518  (.A(II15272), .Z(g10051) ) ;
INV     gate6519  (.A(g9994), .Z(II15275) ) ;
INV     gate6520  (.A(II15275), .Z(g10056) ) ;
INV     gate6521  (.A(g10033), .Z(II15278) ) ;
INV     gate6522  (.A(II15278), .Z(g10057) ) ;
OR2     gate6523  (.A(II15224), .B(II15225), .Z(g10025) ) ;
INV     gate6524  (.A(g10025), .Z(II15281) ) ;
INV     gate6525  (.A(II15281), .Z(g10058) ) ;
INV     gate6526  (.A(g10034), .Z(II15284) ) ;
INV     gate6527  (.A(II15284), .Z(g10062) ) ;
INV     gate6528  (.A(g9980), .Z(II15287) ) ;
INV     gate6529  (.A(II15287), .Z(g10063) ) ;
INV     gate6530  (.A(g9984), .Z(II15290) ) ;
INV     gate6531  (.A(II15290), .Z(g10064) ) ;
INV     gate6532  (.A(g10001), .Z(II15293) ) ;
INV     gate6533  (.A(II15293), .Z(g10065) ) ;
INV     gate6534  (.A(g9995), .Z(II15296) ) ;
INV     gate6535  (.A(II15296), .Z(g10069) ) ;
INV     gate6536  (.A(g9995), .Z(II15299) ) ;
INV     gate6537  (.A(II15299), .Z(g10074) ) ;
OR2     gate6538  (.A(II15209), .B(II15210), .Z(g10007) ) ;
INV     gate6539  (.A(g10007), .Z(II15302) ) ;
INV     gate6540  (.A(II15302), .Z(g10075) ) ;
INV     gate6541  (.A(g10001), .Z(II15305) ) ;
INV     gate6542  (.A(II15305), .Z(g10079) ) ;
INV     gate6543  (.A(g10019), .Z(II15308) ) ;
INV     gate6544  (.A(II15308), .Z(g10080) ) ;
INV     gate6545  (.A(g10013), .Z(II15311) ) ;
INV     gate6546  (.A(II15311), .Z(g10083) ) ;
INV     gate6547  (.A(g10007), .Z(II15314) ) ;
INV     gate6548  (.A(II15314), .Z(g10087) ) ;
INV     gate6549  (.A(g10025), .Z(II15317) ) ;
INV     gate6550  (.A(II15317), .Z(g10088) ) ;
INV     gate6551  (.A(g10013), .Z(II15320) ) ;
INV     gate6552  (.A(II15320), .Z(g10091) ) ;
INV     gate6553  (.A(g10019), .Z(II15323) ) ;
INV     gate6554  (.A(II15323), .Z(g10092) ) ;
INV     gate6555  (.A(g10025), .Z(II15326) ) ;
INV     gate6556  (.A(II15326), .Z(g10093) ) ;
INV     gate6557  (.A(g9995), .Z(II15329) ) ;
INV     gate6558  (.A(II15329), .Z(g10094) ) ;
INV     gate6559  (.A(g10001), .Z(II15332) ) ;
INV     gate6560  (.A(II15332), .Z(g10098) ) ;
INV     gate6561  (.A(g10007), .Z(II15335) ) ;
INV     gate6562  (.A(II15335), .Z(g10101) ) ;
INV     gate6563  (.A(g10013), .Z(II15338) ) ;
INV     gate6564  (.A(II15338), .Z(g10104) ) ;
INV     gate6565  (.A(g10019), .Z(II15341) ) ;
INV     gate6566  (.A(II15341), .Z(g10107) ) ;
INV     gate6567  (.A(g10025), .Z(II15344) ) ;
INV     gate6568  (.A(II15344), .Z(g10110) ) ;
INV     gate6569  (.A(g9995), .Z(II15347) ) ;
INV     gate6570  (.A(II15347), .Z(g10111) ) ;
INV     gate6571  (.A(g10001), .Z(II15350) ) ;
INV     gate6572  (.A(II15350), .Z(g10114) ) ;
INV     gate6573  (.A(g10007), .Z(II15353) ) ;
INV     gate6574  (.A(II15353), .Z(g10115) ) ;
INV     gate6575  (.A(g10013), .Z(II15356) ) ;
INV     gate6576  (.A(II15356), .Z(g10116) ) ;
INV     gate6577  (.A(g10019), .Z(II15359) ) ;
INV     gate6578  (.A(II15359), .Z(g10117) ) ;
INV     gate6579  (.A(g9987), .Z(II15362) ) ;
INV     gate6580  (.A(II15362), .Z(g10118) ) ;
INV     gate6581  (.A(g10025), .Z(II15365) ) ;
INV     gate6582  (.A(II15365), .Z(g10119) ) ;
INV     gate6583  (.A(g9990), .Z(II15368) ) ;
INV     gate6584  (.A(II15368), .Z(g10120) ) ;
INV     gate6585  (.A(g9990), .Z(II15371) ) ;
INV     gate6586  (.A(II15371), .Z(g10121) ) ;
INV     gate6587  (.A(g10007), .Z(II15374) ) ;
INV     gate6588  (.A(II15374), .Z(g10122) ) ;
INV     gate6589  (.A(g10104), .Z(II15377) ) ;
INV     gate6590  (.A(II15377), .Z(g10125) ) ;
INV     gate6591  (.A(g10098), .Z(II15380) ) ;
INV     gate6592  (.A(II15380), .Z(g10126) ) ;
INV     gate6593  (.A(g10107), .Z(II15383) ) ;
INV     gate6594  (.A(II15383), .Z(g10127) ) ;
INV     gate6595  (.A(g10101), .Z(II15386) ) ;
INV     gate6596  (.A(II15386), .Z(g10128) ) ;
INV     gate6597  (.A(g10110), .Z(II15389) ) ;
INV     gate6598  (.A(II15389), .Z(g10129) ) ;
INV     gate6599  (.A(g10104), .Z(II15392) ) ;
INV     gate6600  (.A(II15392), .Z(g10130) ) ;
INV     gate6601  (.A(g10058), .Z(II15395) ) ;
INV     gate6602  (.A(II15395), .Z(g10131) ) ;
INV     gate6603  (.A(g10063), .Z(g10132) ) ;
INV     gate6604  (.A(g10064), .Z(g10133) ) ;
INV     gate6605  (.A(g10069), .Z(II15400) ) ;
INV     gate6606  (.A(II15400), .Z(g10134) ) ;
INV     gate6607  (.A(g10069), .Z(II15403) ) ;
INV     gate6608  (.A(II15403), .Z(g10135) ) ;
INV     gate6609  (.A(g10065), .Z(II15406) ) ;
INV     gate6610  (.A(II15406), .Z(g10136) ) ;
INV     gate6611  (.A(g10065), .Z(II15409) ) ;
INV     gate6612  (.A(II15409), .Z(g10137) ) ;
INV     gate6613  (.A(g10075), .Z(II15412) ) ;
INV     gate6614  (.A(II15412), .Z(g10138) ) ;
INV     gate6615  (.A(g10075), .Z(II15415) ) ;
INV     gate6616  (.A(II15415), .Z(g10139) ) ;
INV     gate6617  (.A(g10083), .Z(II15418) ) ;
INV     gate6618  (.A(II15418), .Z(g10140) ) ;
INV     gate6619  (.A(g10083), .Z(II15421) ) ;
INV     gate6620  (.A(II15421), .Z(g10141) ) ;
INV     gate6621  (.A(g10080), .Z(II15424) ) ;
INV     gate6622  (.A(II15424), .Z(g10142) ) ;
INV     gate6623  (.A(g10088), .Z(II15427) ) ;
INV     gate6624  (.A(II15427), .Z(g10143) ) ;
INV     gate6625  (.A(g10050), .Z(II15437) ) ;
INV     gate6626  (.A(II15437), .Z(g10145) ) ;
INV     gate6627  (.A(g10121), .Z(g10148) ) ;
INV     gate6628  (.A(g10056), .Z(II15448) ) ;
INV     gate6629  (.A(II15448), .Z(g10150) ) ;
INV     gate6630  (.A(g10069), .Z(II15458) ) ;
INV     gate6631  (.A(II15458), .Z(g10154) ) ;
INV     gate6632  (.A(g10074), .Z(II15461) ) ;
INV     gate6633  (.A(II15461), .Z(g10155) ) ;
INV     gate6634  (.A(g10094), .Z(II15464) ) ;
INV     gate6635  (.A(II15464), .Z(g10156) ) ;
INV     gate6636  (.A(g10079), .Z(II15467) ) ;
INV     gate6637  (.A(II15467), .Z(g10157) ) ;
INV     gate6638  (.A(g10111), .Z(II15470) ) ;
INV     gate6639  (.A(II15470), .Z(g10158) ) ;
INV     gate6640  (.A(g10087), .Z(II15473) ) ;
INV     gate6641  (.A(II15473), .Z(g10159) ) ;
INV     gate6642  (.A(g10114), .Z(II15476) ) ;
INV     gate6643  (.A(II15476), .Z(g10160) ) ;
INV     gate6644  (.A(g10091), .Z(II15479) ) ;
INV     gate6645  (.A(II15479), .Z(g10161) ) ;
INV     gate6646  (.A(g10115), .Z(II15482) ) ;
INV     gate6647  (.A(II15482), .Z(g10162) ) ;
INV     gate6648  (.A(g10092), .Z(II15485) ) ;
INV     gate6649  (.A(II15485), .Z(g10163) ) ;
INV     gate6650  (.A(g10116), .Z(II15488) ) ;
INV     gate6651  (.A(II15488), .Z(g10164) ) ;
INV     gate6652  (.A(g10093), .Z(II15491) ) ;
INV     gate6653  (.A(II15491), .Z(g10165) ) ;
INV     gate6654  (.A(g10117), .Z(II15494) ) ;
INV     gate6655  (.A(II15494), .Z(g10166) ) ;
INV     gate6656  (.A(g10119), .Z(II15497) ) ;
INV     gate6657  (.A(II15497), .Z(g10167) ) ;
INV     gate6658  (.A(g10051), .Z(II15500) ) ;
INV     gate6659  (.A(II15500), .Z(g10168) ) ;
INV     gate6660  (.A(g10044), .Z(II15503) ) ;
INV     gate6661  (.A(II15503), .Z(g10169) ) ;
INV     gate6662  (.A(g10118), .Z(g10170) ) ;
INV     gate6663  (.A(g10047), .Z(II15507) ) ;
INV     gate6664  (.A(II15507), .Z(g10171) ) ;
INV     gate6665  (.A(g10035), .Z(II15510) ) ;
INV     gate6666  (.A(II15510), .Z(g10172) ) ;
INV     gate6667  (.A(g10120), .Z(g10173) ) ;
INV     gate6668  (.A(g10122), .Z(II15514) ) ;
INV     gate6669  (.A(II15514), .Z(g10174) ) ;
INV     gate6670  (.A(g10051), .Z(II15517) ) ;
INV     gate6671  (.A(II15517), .Z(g10175) ) ;
INV     gate6672  (.A(g10035), .Z(II15520) ) ;
INV     gate6673  (.A(II15520), .Z(g10176) ) ;
INV     gate6674  (.A(g10058), .Z(II15523) ) ;
INV     gate6675  (.A(II15523), .Z(g10177) ) ;
INV     gate6676  (.A(g10051), .Z(II15526) ) ;
INV     gate6677  (.A(II15526), .Z(g10178) ) ;
INV     gate6678  (.A(g10041), .Z(g10179) ) ;
INV     gate6679  (.A(g10107), .Z(II15530) ) ;
INV     gate6680  (.A(II15530), .Z(g10182) ) ;
INV     gate6681  (.A(g10042), .Z(g10183) ) ;
INV     gate6682  (.A(g10039), .Z(g10184) ) ;
INV     gate6683  (.A(g10040), .Z(g10185) ) ;
INV     gate6684  (.A(g10111), .Z(II15536) ) ;
INV     gate6685  (.A(II15536), .Z(g10186) ) ;
INV     gate6686  (.A(g10069), .Z(II15539) ) ;
INV     gate6687  (.A(II15539), .Z(g10187) ) ;
INV     gate6688  (.A(g10065), .Z(II15542) ) ;
INV     gate6689  (.A(II15542), .Z(g10188) ) ;
INV     gate6690  (.A(g10075), .Z(II15545) ) ;
INV     gate6691  (.A(II15545), .Z(g10189) ) ;
INV     gate6692  (.A(g10083), .Z(II15548) ) ;
INV     gate6693  (.A(II15548), .Z(g10190) ) ;
INV     gate6694  (.A(g10080), .Z(II15551) ) ;
INV     gate6695  (.A(II15551), .Z(g10191) ) ;
INV     gate6696  (.A(g10088), .Z(II15554) ) ;
INV     gate6697  (.A(II15554), .Z(g10192) ) ;
INV     gate6698  (.A(g10057), .Z(g10193) ) ;
INV     gate6699  (.A(g10062), .Z(g10194) ) ;
INV     gate6700  (.A(g10094), .Z(II15559) ) ;
INV     gate6701  (.A(II15559), .Z(g10195) ) ;
INV     gate6702  (.A(g10098), .Z(II15562) ) ;
INV     gate6703  (.A(II15562), .Z(g10196) ) ;
INV     gate6704  (.A(g10101), .Z(II15565) ) ;
INV     gate6705  (.A(II15565), .Z(g10197) ) ;
INV     gate6706  (.A(g10094), .Z(II15568) ) ;
INV     gate6707  (.A(II15568), .Z(g10198) ) ;
INV     gate6708  (.A(g10172), .Z(g10199) ) ;
INV     gate6709  (.A(g10169), .Z(g10200) ) ;
INV     gate6710  (.A(g10175), .Z(g10201) ) ;
INV     gate6711  (.A(g10171), .Z(g10202) ) ;
INV     gate6712  (.A(g10177), .Z(g10203) ) ;
INV     gate6713  (.A(g10174), .Z(g10204) ) ;
INV     gate6714  (.A(g10176), .Z(g10205) ) ;
INV     gate6715  (.A(g10178), .Z(g10206) ) ;
INV     gate6716  (.A(g10186), .Z(g10207) ) ;
INV     gate6717  (.A(g10155), .Z(II15580) ) ;
INV     gate6718  (.A(II15580), .Z(g10208) ) ;
INV     gate6719  (.A(g10157), .Z(II15583) ) ;
INV     gate6720  (.A(II15583), .Z(g10211) ) ;
INV     gate6721  (.A(g10159), .Z(II15586) ) ;
INV     gate6722  (.A(II15586), .Z(g10214) ) ;
INV     gate6723  (.A(g10161), .Z(II15589) ) ;
INV     gate6724  (.A(II15589), .Z(g10217) ) ;
INV     gate6725  (.A(g10163), .Z(II15592) ) ;
INV     gate6726  (.A(II15592), .Z(g10220) ) ;
INV     gate6727  (.A(g10165), .Z(II15595) ) ;
INV     gate6728  (.A(II15595), .Z(g10223) ) ;
INV     gate6729  (.A(g10170), .Z(II15598) ) ;
INV     gate6730  (.A(II15598), .Z(g10226) ) ;
INV     gate6731  (.A(g10173), .Z(II15601) ) ;
INV     gate6732  (.A(II15601), .Z(g10227) ) ;
INV     gate6733  (.A(g10148), .Z(II15604) ) ;
INV     gate6734  (.A(II15604), .Z(g10228) ) ;
INV     gate6735  (.A(g10187), .Z(g10233) ) ;
INV     gate6736  (.A(g10188), .Z(g10234) ) ;
INV     gate6737  (.A(g10189), .Z(g10235) ) ;
INV     gate6738  (.A(g10190), .Z(g10236) ) ;
INV     gate6739  (.A(g10191), .Z(g10238) ) ;
INV     gate6740  (.A(g10192), .Z(g10241) ) ;
INV     gate6741  (.A(g10184), .Z(II15632) ) ;
INV     gate6742  (.A(II15632), .Z(g10242) ) ;
INV     gate6743  (.A(g10185), .Z(II15635) ) ;
INV     gate6744  (.A(II15635), .Z(g10243) ) ;
INV     gate6745  (.A(g10131), .Z(g10244) ) ;
INV     gate6746  (.A(g10179), .Z(II15639) ) ;
INV     gate6747  (.A(II15639), .Z(g10247) ) ;
INV     gate6748  (.A(g10134), .Z(g10248) ) ;
INV     gate6749  (.A(g10135), .Z(g10249) ) ;
INV     gate6750  (.A(g10136), .Z(g10250) ) ;
INV     gate6751  (.A(g10195), .Z(g10251) ) ;
INV     gate6752  (.A(g10137), .Z(g10252) ) ;
INV     gate6753  (.A(g10138), .Z(g10253) ) ;
INV     gate6754  (.A(g10196), .Z(g10254) ) ;
INV     gate6755  (.A(g10139), .Z(g10255) ) ;
INV     gate6756  (.A(g10140), .Z(g10256) ) ;
INV     gate6757  (.A(g10197), .Z(g10257) ) ;
INV     gate6758  (.A(g10198), .Z(g10258) ) ;
INV     gate6759  (.A(g10141), .Z(g10259) ) ;
INV     gate6760  (.A(g10125), .Z(g10260) ) ;
INV     gate6761  (.A(g10126), .Z(g10261) ) ;
INV     gate6762  (.A(g10142), .Z(g10262) ) ;
INV     gate6763  (.A(g10127), .Z(g10263) ) ;
INV     gate6764  (.A(g10128), .Z(g10264) ) ;
INV     gate6765  (.A(g10143), .Z(g10265) ) ;
INV     gate6766  (.A(g10129), .Z(g10266) ) ;
INV     gate6767  (.A(g10130), .Z(g10267) ) ;
INV     gate6768  (.A(g10154), .Z(g10269) ) ;
INV     gate6769  (.A(g10156), .Z(g10270) ) ;
INV     gate6770  (.A(g10193), .Z(II15665) ) ;
INV     gate6771  (.A(II15665), .Z(g10271) ) ;
INV     gate6772  (.A(g10168), .Z(g10272) ) ;
INV     gate6773  (.A(g10194), .Z(II15669) ) ;
INV     gate6774  (.A(II15669), .Z(g10275) ) ;
INV     gate6775  (.A(g10132), .Z(II15672) ) ;
INV     gate6776  (.A(II15672), .Z(g10276) ) ;
INV     gate6777  (.A(g10133), .Z(II15675) ) ;
INV     gate6778  (.A(II15675), .Z(g10277) ) ;
INV     gate6779  (.A(g10182), .Z(g10278) ) ;
INV     gate6780  (.A(g10158), .Z(g10279) ) ;
INV     gate6781  (.A(g10160), .Z(g10280) ) ;
INV     gate6782  (.A(g10162), .Z(g10281) ) ;
INV     gate6783  (.A(g10164), .Z(g10282) ) ;
INV     gate6784  (.A(g10166), .Z(g10283) ) ;
INV     gate6785  (.A(g10167), .Z(g10284) ) ;
INV     gate6786  (.A(g10207), .Z(II15688) ) ;
INV     gate6787  (.A(II15688), .Z(g10288) ) ;
INV     gate6788  (.A(g10233), .Z(II15691) ) ;
INV     gate6789  (.A(II15691), .Z(g10289) ) ;
INV     gate6790  (.A(g10234), .Z(II15694) ) ;
INV     gate6791  (.A(II15694), .Z(g10290) ) ;
INV     gate6792  (.A(g10235), .Z(II15698) ) ;
INV     gate6793  (.A(II15698), .Z(g10292) ) ;
INV     gate6794  (.A(g10236), .Z(II15701) ) ;
INV     gate6795  (.A(II15701), .Z(g10293) ) ;
INV     gate6796  (.A(g10238), .Z(II15704) ) ;
INV     gate6797  (.A(II15704), .Z(g10294) ) ;
INV     gate6798  (.A(g10241), .Z(II15708) ) ;
INV     gate6799  (.A(II15708), .Z(g10296) ) ;
INV     gate6800  (.A(g10251), .Z(II15725) ) ;
INV     gate6801  (.A(II15725), .Z(g10305) ) ;
INV     gate6802  (.A(g10254), .Z(II15729) ) ;
INV     gate6803  (.A(II15729), .Z(g10307) ) ;
INV     gate6804  (.A(g10257), .Z(II15733) ) ;
INV     gate6805  (.A(II15733), .Z(g10309) ) ;
INV     gate6806  (.A(g10258), .Z(II15736) ) ;
INV     gate6807  (.A(II15736), .Z(g10310) ) ;
INV     gate6808  (.A(g10242), .Z(g10311) ) ;
INV     gate6809  (.A(g10260), .Z(II15741) ) ;
INV     gate6810  (.A(II15741), .Z(g10313) ) ;
INV     gate6811  (.A(g10261), .Z(II15744) ) ;
INV     gate6812  (.A(II15744), .Z(g10314) ) ;
INV     gate6813  (.A(g10243), .Z(g10315) ) ;
INV     gate6814  (.A(g10263), .Z(II15749) ) ;
INV     gate6815  (.A(II15749), .Z(g10317) ) ;
INV     gate6816  (.A(g10264), .Z(II15752) ) ;
INV     gate6817  (.A(II15752), .Z(g10318) ) ;
INV     gate6818  (.A(g10270), .Z(g10319) ) ;
INV     gate6819  (.A(g10266), .Z(II15756) ) ;
INV     gate6820  (.A(II15756), .Z(g10320) ) ;
INV     gate6821  (.A(g10267), .Z(II15759) ) ;
INV     gate6822  (.A(II15759), .Z(g10321) ) ;
INV     gate6823  (.A(g10244), .Z(II15763) ) ;
INV     gate6824  (.A(II15763), .Z(g10323) ) ;
INV     gate6825  (.A(g10249), .Z(II15768) ) ;
INV     gate6826  (.A(II15768), .Z(g10326) ) ;
INV     gate6827  (.A(g10250), .Z(II15771) ) ;
INV     gate6828  (.A(II15771), .Z(g10327) ) ;
INV     gate6829  (.A(g10253), .Z(II15775) ) ;
INV     gate6830  (.A(II15775), .Z(g10329) ) ;
INV     gate6831  (.A(g10255), .Z(II15778) ) ;
INV     gate6832  (.A(II15778), .Z(g10330) ) ;
INV     gate6833  (.A(g10259), .Z(II15782) ) ;
INV     gate6834  (.A(II15782), .Z(g10332) ) ;
INV     gate6835  (.A(g10269), .Z(II15787) ) ;
INV     gate6836  (.A(II15787), .Z(g10335) ) ;
INV     gate6837  (.A(g10279), .Z(II15792) ) ;
INV     gate6838  (.A(II15792), .Z(g10342) ) ;
INV     gate6839  (.A(g10280), .Z(II15795) ) ;
INV     gate6840  (.A(II15795), .Z(g10343) ) ;
INV     gate6841  (.A(g10281), .Z(II15798) ) ;
INV     gate6842  (.A(II15798), .Z(g10344) ) ;
INV     gate6843  (.A(g10282), .Z(II15801) ) ;
INV     gate6844  (.A(II15801), .Z(g10345) ) ;
INV     gate6845  (.A(g10283), .Z(II15804) ) ;
INV     gate6846  (.A(II15804), .Z(g10346) ) ;
INV     gate6847  (.A(g10284), .Z(II15807) ) ;
INV     gate6848  (.A(II15807), .Z(g10347) ) ;
INV     gate6849  (.A(g10200), .Z(II15811) ) ;
INV     gate6850  (.A(II15811), .Z(g10349) ) ;
INV     gate6851  (.A(g10202), .Z(II15814) ) ;
INV     gate6852  (.A(II15814), .Z(g10350) ) ;
INV     gate6853  (.A(g10199), .Z(II15817) ) ;
INV     gate6854  (.A(II15817), .Z(g10351) ) ;
INV     gate6855  (.A(g10204), .Z(II15820) ) ;
INV     gate6856  (.A(II15820), .Z(g10352) ) ;
INV     gate6857  (.A(g10201), .Z(II15823) ) ;
INV     gate6858  (.A(II15823), .Z(g10353) ) ;
INV     gate6859  (.A(g10205), .Z(II15826) ) ;
INV     gate6860  (.A(II15826), .Z(g10354) ) ;
INV     gate6861  (.A(g10203), .Z(II15829) ) ;
INV     gate6862  (.A(II15829), .Z(g10355) ) ;
INV     gate6863  (.A(g10206), .Z(II15832) ) ;
INV     gate6864  (.A(II15832), .Z(g10356) ) ;
AND2    gate6865  (.A(g10183), .B(g3307), .Z(g10268) ) ;
INV     gate6866  (.A(g10268), .Z(g10361) ) ;
OR2     gate6867  (.A(g10230), .B(g9572), .Z(g10336) ) ;
INV     gate6868  (.A(g10336), .Z(II15855) ) ;
INV     gate6869  (.A(g10336), .Z(II15858) ) ;
INV     gate6870  (.A(II15858), .Z(g10378) ) ;
OR2     gate6871  (.A(g10232), .B(g9556), .Z(g10339) ) ;
INV     gate6872  (.A(g10339), .Z(II15861) ) ;
INV     gate6873  (.A(g10339), .Z(II15864) ) ;
INV     gate6874  (.A(II15864), .Z(g10380) ) ;
AND2    gate6875  (.A(g10278), .B(g2462), .Z(g10357) ) ;
INV     gate6876  (.A(g10357), .Z(g10387) ) ;
INV     gate6877  (.A(g10305), .Z(g10388) ) ;
INV     gate6878  (.A(g10307), .Z(g10389) ) ;
INV     gate6879  (.A(g10309), .Z(g10390) ) ;
INV     gate6880  (.A(g10313), .Z(g10391) ) ;
INV     gate6881  (.A(g10317), .Z(g10393) ) ;
INV     gate6882  (.A(g10320), .Z(g10395) ) ;
AND2    gate6883  (.A(g10272), .B(g3705), .Z(g10348) ) ;
INV     gate6884  (.A(g10348), .Z(g10400) ) ;
AND2    gate6885  (.A(g10256), .B(g3307), .Z(g10331) ) ;
INV     gate6886  (.A(g10331), .Z(g10421) ) ;
AND2    gate6887  (.A(g10252), .B(g3307), .Z(g10328) ) ;
INV     gate6888  (.A(g10328), .Z(g10431) ) ;
AND2    gate6889  (.A(g10262), .B(g3307), .Z(g10333) ) ;
INV     gate6890  (.A(g10333), .Z(g10437) ) ;
AND2    gate6891  (.A(g10265), .B(g3307), .Z(g10334) ) ;
INV     gate6892  (.A(g10334), .Z(g10439) ) ;
AND2    gate6893  (.A(g10248), .B(g3307), .Z(g10325) ) ;
INV     gate6894  (.A(g10325), .Z(g10444) ) ;
OR2     gate6895  (.A(g10295), .B(g9554), .Z(g10402) ) ;
INV     gate6896  (.A(g10402), .Z(II15956) ) ;
INV     gate6897  (.A(g10402), .Z(II15959) ) ;
INV     gate6898  (.A(II15959), .Z(g10456) ) ;
OR2     gate6899  (.A(g10297), .B(g9530), .Z(g10405) ) ;
INV     gate6900  (.A(g10405), .Z(II15962) ) ;
INV     gate6901  (.A(g10405), .Z(II15965) ) ;
INV     gate6902  (.A(II15965), .Z(g10458) ) ;
OR2     gate6903  (.A(g10298), .B(g9553), .Z(g10408) ) ;
INV     gate6904  (.A(g10408), .Z(II15968) ) ;
INV     gate6905  (.A(g10408), .Z(II15971) ) ;
INV     gate6906  (.A(II15971), .Z(g10460) ) ;
OR2     gate6907  (.A(g10299), .B(g9529), .Z(g10411) ) ;
INV     gate6908  (.A(g10411), .Z(II15974) ) ;
INV     gate6909  (.A(g10411), .Z(II15977) ) ;
INV     gate6910  (.A(II15977), .Z(g10462) ) ;
OR2     gate6911  (.A(g10300), .B(g9534), .Z(g10414) ) ;
INV     gate6912  (.A(g10414), .Z(II15980) ) ;
INV     gate6913  (.A(g10414), .Z(II15983) ) ;
INV     gate6914  (.A(II15983), .Z(g10464) ) ;
OR2     gate6915  (.A(g10301), .B(g9527), .Z(g10417) ) ;
INV     gate6916  (.A(g10417), .Z(II15986) ) ;
INV     gate6917  (.A(g10417), .Z(II15989) ) ;
INV     gate6918  (.A(II15989), .Z(g10466) ) ;
INV     gate6919  (.A(g10378), .Z(g10471) ) ;
INV     gate6920  (.A(g10380), .Z(g10473) ) ;
OR2     gate6921  (.A(g9317), .B(g10291), .Z(g10401) ) ;
INV     gate6922  (.A(g10401), .Z(II16095) ) ;
INV     gate6923  (.A(II16095), .Z(g10486) ) ;
AND2    gate6924  (.A(g10361), .B(g3382), .Z(g10369) ) ;
INV     gate6925  (.A(g10369), .Z(II16098) ) ;
INV     gate6926  (.A(II16098), .Z(g10487) ) ;
NOR2    gate6927  (.A(g10310), .B(g2998), .Z(g10381) ) ;
INV     gate6928  (.A(g10381), .Z(II16101) ) ;
INV     gate6929  (.A(II16101), .Z(g10488) ) ;
NOR2    gate6930  (.A(g10314), .B(g2998), .Z(g10382) ) ;
INV     gate6931  (.A(g10382), .Z(II16105) ) ;
INV     gate6932  (.A(II16105), .Z(g10490) ) ;
NOR2    gate6933  (.A(g10318), .B(g2998), .Z(g10383) ) ;
INV     gate6934  (.A(g10383), .Z(II16108) ) ;
INV     gate6935  (.A(II16108), .Z(g10491) ) ;
NOR2    gate6936  (.A(g10321), .B(g2998), .Z(g10385) ) ;
INV     gate6937  (.A(g10385), .Z(II16111) ) ;
INV     gate6938  (.A(II16111), .Z(g10492) ) ;
INV     gate6939  (.A(g10387), .Z(II16114) ) ;
INV     gate6940  (.A(II16114), .Z(g10493) ) ;
NAND2   gate6941  (.A(II15907), .B(II15908), .Z(g10396) ) ;
INV     gate6942  (.A(g10396), .Z(II16121) ) ;
INV     gate6943  (.A(II16121), .Z(g10498) ) ;
INV     gate6944  (.A(g10396), .Z(II16124) ) ;
INV     gate6945  (.A(II16124), .Z(g10499) ) ;
INV     gate6946  (.A(g10456), .Z(g10523) ) ;
INV     gate6947  (.A(g10458), .Z(g10524) ) ;
INV     gate6948  (.A(g10499), .Z(g10525) ) ;
INV     gate6949  (.A(g10460), .Z(g10526) ) ;
INV     gate6950  (.A(g10462), .Z(g10527) ) ;
INV     gate6951  (.A(g10464), .Z(g10528) ) ;
INV     gate6952  (.A(g10466), .Z(g10530) ) ;
INV     gate6953  (.A(g10471), .Z(g10531) ) ;
INV     gate6954  (.A(g10473), .Z(g10532) ) ;
AND2    gate6955  (.A(g10421), .B(g3335), .Z(g10448) ) ;
INV     gate6956  (.A(g10448), .Z(II16169) ) ;
INV     gate6957  (.A(II16169), .Z(g10534) ) ;
INV     gate6958  (.A(g10498), .Z(II16172) ) ;
INV     gate6959  (.A(II16172), .Z(g10535) ) ;
INV     gate6960  (.A(g10488), .Z(II16175) ) ;
INV     gate6961  (.A(II16175), .Z(g10536) ) ;
INV     gate6962  (.A(g10490), .Z(II16178) ) ;
INV     gate6963  (.A(II16178), .Z(g10537) ) ;
INV     gate6964  (.A(g10491), .Z(II16181) ) ;
INV     gate6965  (.A(II16181), .Z(g10538) ) ;
OR2     gate6966  (.A(g9317), .B(g10400), .Z(g10484) ) ;
INV     gate6967  (.A(g10484), .Z(II16184) ) ;
INV     gate6968  (.A(II16184), .Z(g10539) ) ;
INV     gate6969  (.A(g10492), .Z(II16187) ) ;
INV     gate6970  (.A(II16187), .Z(g10540) ) ;
INV     gate6971  (.A(g10493), .Z(II16190) ) ;
INV     gate6972  (.A(II16190), .Z(g10541) ) ;
OR2     gate6973  (.A(g9317), .B(g10376), .Z(g10485) ) ;
INV     gate6974  (.A(g10485), .Z(II16193) ) ;
INV     gate6975  (.A(II16193), .Z(g10542) ) ;
AND2    gate6976  (.A(g10429), .B(g3977), .Z(g10496) ) ;
INV     gate6977  (.A(g10496), .Z(II16196) ) ;
INV     gate6978  (.A(II16196), .Z(g10543) ) ;
AND2    gate6979  (.A(g10433), .B(g3945), .Z(g10494) ) ;
INV     gate6980  (.A(g10494), .Z(II16200) ) ;
INV     gate6981  (.A(II16200), .Z(g10545) ) ;
AND2    gate6982  (.A(g10435), .B(g3411), .Z(g10454) ) ;
INV     gate6983  (.A(g10454), .Z(II16203) ) ;
INV     gate6984  (.A(II16203), .Z(g10546) ) ;
AND2    gate6985  (.A(g10437), .B(g3395), .Z(g10453) ) ;
INV     gate6986  (.A(g10453), .Z(II16206) ) ;
INV     gate6987  (.A(II16206), .Z(g10547) ) ;
AND2    gate6988  (.A(g10439), .B(g3388), .Z(g10452) ) ;
INV     gate6989  (.A(g10452), .Z(II16209) ) ;
INV     gate6990  (.A(II16209), .Z(g10548) ) ;
OR2     gate6991  (.A(g4157), .B(g10442), .Z(g10500) ) ;
INV     gate6992  (.A(g10500), .Z(II16214) ) ;
INV     gate6993  (.A(II16214), .Z(g10551) ) ;
OR2     gate6994  (.A(g4161), .B(g10445), .Z(g10501) ) ;
INV     gate6995  (.A(g10501), .Z(II16217) ) ;
INV     gate6996  (.A(II16217), .Z(g10552) ) ;
OR2     gate6997  (.A(g4169), .B(g10365), .Z(g10502) ) ;
INV     gate6998  (.A(g10502), .Z(II16220) ) ;
INV     gate6999  (.A(II16220), .Z(g10553) ) ;
INV     gate7000  (.A(g10535), .Z(II16236) ) ;
INV     gate7001  (.A(II16236), .Z(g10571) ) ;
INV     gate7002  (.A(g10525), .Z(II16239) ) ;
INV     gate7003  (.A(II16239), .Z(g10574) ) ;
INV     gate7004  (.A(g10523), .Z(g10575) ) ;
INV     gate7005  (.A(g10524), .Z(g10576) ) ;
INV     gate7006  (.A(g10526), .Z(g10577) ) ;
INV     gate7007  (.A(g10527), .Z(g10578) ) ;
INV     gate7008  (.A(g10528), .Z(g10579) ) ;
INV     gate7009  (.A(g10530), .Z(g10580) ) ;
NOR2    gate7010  (.A(g10486), .B(g10239), .Z(g10522) ) ;
INV     gate7011  (.A(g10522), .Z(g10584) ) ;
AND3    gate7012  (.A(g10505), .B(g10469), .C(II16142), .Z(g10515) ) ;
INV     gate7013  (.A(g10515), .Z(II16252) ) ;
INV     gate7014  (.A(II16252), .Z(g10589) ) ;
OR2     gate7015  (.A(g4097), .B(g10503), .Z(g10554) ) ;
INV     gate7016  (.A(g10554), .Z(II16255) ) ;
INV     gate7017  (.A(II16255), .Z(g10590) ) ;
OR2     gate7018  (.A(g4103), .B(g10504), .Z(g10555) ) ;
INV     gate7019  (.A(g10555), .Z(II16258) ) ;
INV     gate7020  (.A(II16258), .Z(g10591) ) ;
OR2     gate7021  (.A(g4115), .B(g10506), .Z(g10556) ) ;
INV     gate7022  (.A(g10556), .Z(II16261) ) ;
INV     gate7023  (.A(II16261), .Z(g10592) ) ;
OR2     gate7024  (.A(g4123), .B(g10508), .Z(g10557) ) ;
INV     gate7025  (.A(g10557), .Z(II16264) ) ;
INV     gate7026  (.A(II16264), .Z(g10593) ) ;
OR2     gate7027  (.A(g4126), .B(g10510), .Z(g10558) ) ;
INV     gate7028  (.A(g10558), .Z(II16269) ) ;
INV     gate7029  (.A(II16269), .Z(g10596) ) ;
OR2     gate7030  (.A(g4141), .B(g10512), .Z(g10559) ) ;
INV     gate7031  (.A(g10559), .Z(II16273) ) ;
INV     gate7032  (.A(II16273), .Z(g10598) ) ;
INV     gate7033  (.A(g10536), .Z(II16277) ) ;
INV     gate7034  (.A(II16277), .Z(g10600) ) ;
INV     gate7035  (.A(g10537), .Z(II16280) ) ;
INV     gate7036  (.A(II16280), .Z(g10604) ) ;
INV     gate7037  (.A(g10538), .Z(II16283) ) ;
INV     gate7038  (.A(II16283), .Z(g10608) ) ;
INV     gate7039  (.A(g10540), .Z(II16286) ) ;
INV     gate7040  (.A(II16286), .Z(g10612) ) ;
INV     gate7041  (.A(g10541), .Z(II16289) ) ;
INV     gate7042  (.A(II16289), .Z(g10616) ) ;
INV     gate7043  (.A(g10551), .Z(II16292) ) ;
INV     gate7044  (.A(II16292), .Z(g10619) ) ;
INV     gate7045  (.A(g10552), .Z(II16295) ) ;
INV     gate7046  (.A(II16295), .Z(g10620) ) ;
INV     gate7047  (.A(g10553), .Z(II16298) ) ;
INV     gate7048  (.A(II16298), .Z(g10621) ) ;
INV     gate7049  (.A(g10589), .Z(II16307) ) ;
AND2    gate7050  (.A(g10518), .B(g10515), .Z(g10583) ) ;
INV     gate7051  (.A(g10583), .Z(g10629) ) ;
INV     gate7052  (.A(g10584), .Z(II16311) ) ;
INV     gate7053  (.A(II16311), .Z(g10630) ) ;
NOR2    gate7054  (.A(g10539), .B(g10322), .Z(g10563) ) ;
INV     gate7055  (.A(g10563), .Z(g10668) ) ;
INV     gate7056  (.A(g10584), .Z(g10674) ) ;
INV     gate7057  (.A(g10574), .Z(g10675) ) ;
NOR2    gate7058  (.A(g10542), .B(g10324), .Z(g10570) ) ;
INV     gate7059  (.A(g10570), .Z(g10676) ) ;
INV     gate7060  (.A(g10584), .Z(g10679) ) ;
INV     gate7061  (.A(g10612), .Z(g10683) ) ;
AND2    gate7062  (.A(g10533), .B(g4359), .Z(g10597) ) ;
INV     gate7063  (.A(g10597), .Z(II16356) ) ;
INV     gate7064  (.A(II16356), .Z(g10687) ) ;
INV     gate7065  (.A(g10590), .Z(II16360) ) ;
INV     gate7066  (.A(II16360), .Z(g10691) ) ;
AND2    gate7067  (.A(g10534), .B(g4365), .Z(g10599) ) ;
INV     gate7068  (.A(g10599), .Z(II16363) ) ;
INV     gate7069  (.A(II16363), .Z(g10692) ) ;
INV     gate7070  (.A(g10591), .Z(II16366) ) ;
INV     gate7071  (.A(II16366), .Z(g10695) ) ;
INV     gate7072  (.A(g10621), .Z(g10696) ) ;
INV     gate7073  (.A(g10592), .Z(II16370) ) ;
INV     gate7074  (.A(II16370), .Z(g10697) ) ;
INV     gate7075  (.A(g10593), .Z(II16373) ) ;
INV     gate7076  (.A(II16373), .Z(g10698) ) ;
INV     gate7077  (.A(g10596), .Z(II16376) ) ;
INV     gate7078  (.A(II16376), .Z(g10699) ) ;
INV     gate7079  (.A(g10598), .Z(II16379) ) ;
INV     gate7080  (.A(II16379), .Z(g10700) ) ;
INV     gate7081  (.A(g10629), .Z(II16387) ) ;
INV     gate7082  (.A(II16387), .Z(g10708) ) ;
INV     gate7083  (.A(g10630), .Z(g10729) ) ;
INV     gate7084  (.A(g10696), .Z(II16407) ) ;
INV     gate7085  (.A(II16407), .Z(g10730) ) ;
OR2     gate7086  (.A(g10237), .B(g10581), .Z(g10663) ) ;
INV     gate7087  (.A(g10663), .Z(II16413) ) ;
INV     gate7088  (.A(II16413), .Z(g10734) ) ;
OR2     gate7089  (.A(g10240), .B(g10582), .Z(g10664) ) ;
INV     gate7090  (.A(g10664), .Z(II16416) ) ;
INV     gate7091  (.A(II16416), .Z(g10735) ) ;
OR2     gate7092  (.A(g10562), .B(g3877), .Z(g10702) ) ;
INV     gate7093  (.A(g10702), .Z(II16432) ) ;
INV     gate7094  (.A(II16432), .Z(g10747) ) ;
INV     gate7095  (.A(g10702), .Z(II16439) ) ;
INV     gate7096  (.A(II16439), .Z(g10754) ) ;
INV     gate7097  (.A(g10734), .Z(II16458) ) ;
INV     gate7098  (.A(g10735), .Z(II16461) ) ;
OR2     gate7099  (.A(g5492), .B(g10680), .Z(g10765) ) ;
INV     gate7100  (.A(g10765), .Z(II16475) ) ;
INV     gate7101  (.A(II16475), .Z(g10781) ) ;
OR2     gate7102  (.A(g5500), .B(g10681), .Z(g10767) ) ;
INV     gate7103  (.A(g10767), .Z(II16479) ) ;
INV     gate7104  (.A(II16479), .Z(g10783) ) ;
OR2     gate7105  (.A(g5525), .B(g10682), .Z(g10770) ) ;
INV     gate7106  (.A(g10770), .Z(II16484) ) ;
INV     gate7107  (.A(II16484), .Z(g10786) ) ;
OR2     gate7108  (.A(g5533), .B(g10684), .Z(g10771) ) ;
INV     gate7109  (.A(g10771), .Z(II16487) ) ;
INV     gate7110  (.A(II16487), .Z(g10787) ) ;
OR2     gate7111  (.A(g5540), .B(g10685), .Z(g10773) ) ;
INV     gate7112  (.A(g10773), .Z(II16492) ) ;
INV     gate7113  (.A(II16492), .Z(g10792) ) ;
OR2     gate7114  (.A(g5545), .B(g10686), .Z(g10707) ) ;
INV     gate7115  (.A(g10707), .Z(II16496) ) ;
INV     gate7116  (.A(II16496), .Z(g10794) ) ;
OR2     gate7117  (.A(g5547), .B(g10690), .Z(g10711) ) ;
INV     gate7118  (.A(g10711), .Z(II16500) ) ;
INV     gate7119  (.A(II16500), .Z(g10796) ) ;
OR2     gate7120  (.A(g10662), .B(g9531), .Z(g10712) ) ;
INV     gate7121  (.A(g10712), .Z(II16507) ) ;
INV     gate7122  (.A(g10712), .Z(II16510) ) ;
INV     gate7123  (.A(II16510), .Z(g10802) ) ;
INV     gate7124  (.A(g10708), .Z(g10803) ) ;
OR2     gate7125  (.A(g6235), .B(g10705), .Z(g10717) ) ;
INV     gate7126  (.A(g10717), .Z(II16514) ) ;
INV     gate7127  (.A(II16514), .Z(g10804) ) ;
OR2     gate7128  (.A(g6238), .B(g10706), .Z(g10718) ) ;
INV     gate7129  (.A(g10718), .Z(II16518) ) ;
INV     gate7130  (.A(II16518), .Z(g10806) ) ;
OR2     gate7131  (.A(g10303), .B(g10666), .Z(g10719) ) ;
INV     gate7132  (.A(g10719), .Z(II16525) ) ;
INV     gate7133  (.A(II16525), .Z(g10819) ) ;
OR2     gate7134  (.A(g4358), .B(g10661), .Z(g10732) ) ;
INV     gate7135  (.A(g10732), .Z(II16528) ) ;
INV     gate7136  (.A(II16528), .Z(g10820) ) ;
OR2     gate7137  (.A(g10304), .B(g10667), .Z(g10720) ) ;
INV     gate7138  (.A(g10720), .Z(II16531) ) ;
INV     gate7139  (.A(II16531), .Z(g10821) ) ;
INV     gate7140  (.A(g10747), .Z(II16534) ) ;
INV     gate7141  (.A(II16534), .Z(g10822) ) ;
OR2     gate7142  (.A(g10306), .B(g10669), .Z(g10721) ) ;
INV     gate7143  (.A(g10721), .Z(II16537) ) ;
INV     gate7144  (.A(II16537), .Z(g10825) ) ;
OR2     gate7145  (.A(g10308), .B(g10671), .Z(g10722) ) ;
INV     gate7146  (.A(g10722), .Z(II16540) ) ;
INV     gate7147  (.A(II16540), .Z(g10826) ) ;
INV     gate7148  (.A(g10747), .Z(II16543) ) ;
INV     gate7149  (.A(II16543), .Z(g10827) ) ;
OR2     gate7150  (.A(g10312), .B(g10672), .Z(g10724) ) ;
INV     gate7151  (.A(g10724), .Z(II16546) ) ;
INV     gate7152  (.A(II16546), .Z(g10848) ) ;
OR2     gate7153  (.A(g10316), .B(g10673), .Z(g10726) ) ;
INV     gate7154  (.A(g10726), .Z(II16550) ) ;
INV     gate7155  (.A(II16550), .Z(g10850) ) ;
INV     gate7156  (.A(g10754), .Z(II16553) ) ;
INV     gate7157  (.A(II16553), .Z(g10851) ) ;
AND2    gate7158  (.A(g10676), .B(g3384), .Z(g10740) ) ;
INV     gate7159  (.A(g10740), .Z(g10852) ) ;
INV     gate7160  (.A(g10708), .Z(g10854) ) ;
INV     gate7161  (.A(g10819), .Z(II16571) ) ;
INV     gate7162  (.A(g10821), .Z(II16574) ) ;
INV     gate7163  (.A(g10825), .Z(II16577) ) ;
INV     gate7164  (.A(g10826), .Z(II16580) ) ;
INV     gate7165  (.A(g10848), .Z(II16583) ) ;
INV     gate7166  (.A(g10850), .Z(II16586) ) ;
INV     gate7167  (.A(g10820), .Z(II16589) ) ;
INV     gate7168  (.A(g10781), .Z(II16592) ) ;
INV     gate7169  (.A(g10783), .Z(II16595) ) ;
INV     gate7170  (.A(g10804), .Z(II16598) ) ;
INV     gate7171  (.A(g10806), .Z(II16601) ) ;
INV     gate7172  (.A(g10786), .Z(II16604) ) ;
INV     gate7173  (.A(g10787), .Z(II16607) ) ;
INV     gate7174  (.A(g10792), .Z(II16610) ) ;
INV     gate7175  (.A(g10794), .Z(II16613) ) ;
INV     gate7176  (.A(g10796), .Z(II16616) ) ;
AND2    gate7177  (.A(g4811), .B(g10754), .Z(g10809) ) ;
INV     gate7178  (.A(g10809), .Z(g10883) ) ;
INV     gate7179  (.A(g10809), .Z(g10884) ) ;
INV     gate7180  (.A(g10809), .Z(g10885) ) ;
OR2     gate7181  (.A(g5501), .B(g10741), .Z(g10858) ) ;
INV     gate7182  (.A(g10858), .Z(II16623) ) ;
INV     gate7183  (.A(II16623), .Z(g10887) ) ;
OR2     gate7184  (.A(g5512), .B(g10742), .Z(g10859) ) ;
INV     gate7185  (.A(g10859), .Z(II16626) ) ;
INV     gate7186  (.A(II16626), .Z(g10888) ) ;
OR2     gate7187  (.A(g5513), .B(g10743), .Z(g10860) ) ;
INV     gate7188  (.A(g10860), .Z(II16629) ) ;
INV     gate7189  (.A(II16629), .Z(g10889) ) ;
OR2     gate7190  (.A(g5523), .B(g10745), .Z(g10861) ) ;
INV     gate7191  (.A(g10861), .Z(II16632) ) ;
INV     gate7192  (.A(II16632), .Z(g10890) ) ;
OR2     gate7193  (.A(g5524), .B(g10746), .Z(g10862) ) ;
INV     gate7194  (.A(g10862), .Z(II16635) ) ;
INV     gate7195  (.A(II16635), .Z(g10891) ) ;
OR2     gate7196  (.A(g5531), .B(g10750), .Z(g10863) ) ;
INV     gate7197  (.A(g10863), .Z(II16638) ) ;
INV     gate7198  (.A(II16638), .Z(g10892) ) ;
OR2     gate7199  (.A(g5532), .B(g10751), .Z(g10864) ) ;
INV     gate7200  (.A(g10864), .Z(II16641) ) ;
INV     gate7201  (.A(II16641), .Z(g10893) ) ;
OR2     gate7202  (.A(g5538), .B(g10752), .Z(g10865) ) ;
INV     gate7203  (.A(g10865), .Z(II16644) ) ;
INV     gate7204  (.A(II16644), .Z(g10894) ) ;
OR2     gate7205  (.A(g5539), .B(g10753), .Z(g10866) ) ;
INV     gate7206  (.A(g10866), .Z(II16647) ) ;
INV     gate7207  (.A(II16647), .Z(g10895) ) ;
OR2     gate7208  (.A(g5544), .B(g10758), .Z(g10776) ) ;
INV     gate7209  (.A(g10776), .Z(II16650) ) ;
INV     gate7210  (.A(II16650), .Z(g10896) ) ;
INV     gate7211  (.A(g10827), .Z(g10897) ) ;
INV     gate7212  (.A(g10803), .Z(g10899) ) ;
OR2     gate7213  (.A(g6186), .B(g10762), .Z(g10791) ) ;
INV     gate7214  (.A(g10791), .Z(II16656) ) ;
INV     gate7215  (.A(II16656), .Z(g10900) ) ;
INV     gate7216  (.A(g10802), .Z(g10901) ) ;
OR2     gate7217  (.A(g6194), .B(g10763), .Z(g10793) ) ;
INV     gate7218  (.A(g10793), .Z(II16660) ) ;
INV     gate7219  (.A(II16660), .Z(g10902) ) ;
INV     gate7220  (.A(g10809), .Z(g10903) ) ;
OR2     gate7221  (.A(g6199), .B(g10764), .Z(g10795) ) ;
INV     gate7222  (.A(g10795), .Z(II16664) ) ;
INV     gate7223  (.A(II16664), .Z(g10904) ) ;
AND2    gate7224  (.A(g10723), .B(g5124), .Z(g10780) ) ;
INV     gate7225  (.A(g10780), .Z(II16667) ) ;
INV     gate7226  (.A(II16667), .Z(g10905) ) ;
OR2     gate7227  (.A(g6206), .B(g10766), .Z(g10797) ) ;
INV     gate7228  (.A(g10797), .Z(II16670) ) ;
INV     gate7229  (.A(II16670), .Z(g10906) ) ;
AND2    gate7230  (.A(g10725), .B(g5146), .Z(g10782) ) ;
INV     gate7231  (.A(g10782), .Z(II16673) ) ;
INV     gate7232  (.A(II16673), .Z(g10907) ) ;
OR2     gate7233  (.A(g6217), .B(g10768), .Z(g10798) ) ;
INV     gate7234  (.A(g10798), .Z(II16676) ) ;
INV     gate7235  (.A(II16676), .Z(g10908) ) ;
AND2    gate7236  (.A(g10727), .B(g5169), .Z(g10784) ) ;
INV     gate7237  (.A(g10784), .Z(II16679) ) ;
INV     gate7238  (.A(II16679), .Z(g10909) ) ;
OR2     gate7239  (.A(g6225), .B(g10769), .Z(g10799) ) ;
INV     gate7240  (.A(g10799), .Z(II16682) ) ;
INV     gate7241  (.A(II16682), .Z(g10910) ) ;
AND2    gate7242  (.A(g10728), .B(g5177), .Z(g10785) ) ;
INV     gate7243  (.A(g10785), .Z(II16685) ) ;
INV     gate7244  (.A(II16685), .Z(g10911) ) ;
OR2     gate7245  (.A(g6245), .B(g10772), .Z(g10800) ) ;
INV     gate7246  (.A(g10800), .Z(II16688) ) ;
INV     gate7247  (.A(II16688), .Z(g10912) ) ;
AND2    gate7248  (.A(g8303), .B(g10754), .Z(g10788) ) ;
INV     gate7249  (.A(g10788), .Z(II16691) ) ;
INV     gate7250  (.A(II16691), .Z(g10913) ) ;
INV     gate7251  (.A(g10827), .Z(g10926) ) ;
INV     gate7252  (.A(g10827), .Z(g10927) ) ;
INV     gate7253  (.A(g10827), .Z(g10928) ) ;
INV     gate7254  (.A(g10827), .Z(g10929) ) ;
INV     gate7255  (.A(g10827), .Z(g10930) ) ;
INV     gate7256  (.A(g10827), .Z(g10931) ) ;
INV     gate7257  (.A(g10827), .Z(g10932) ) ;
INV     gate7258  (.A(g10827), .Z(g10934) ) ;
INV     gate7259  (.A(g10827), .Z(g10935) ) ;
INV     gate7260  (.A(g10822), .Z(II16708) ) ;
INV     gate7261  (.A(II16708), .Z(g10947) ) ;
NAND2   gate7262  (.A(II16468), .B(II16469), .Z(g10779) ) ;
INV     gate7263  (.A(g10779), .Z(II16717) ) ;
INV     gate7264  (.A(II16717), .Z(g10972) ) ;
INV     gate7265  (.A(g10854), .Z(II16720) ) ;
INV     gate7266  (.A(II16720), .Z(g10973) ) ;
INV     gate7267  (.A(g10851), .Z(II16723) ) ;
INV     gate7268  (.A(II16723), .Z(g10974) ) ;
OR2     gate7269  (.A(g6075), .B(g10736), .Z(g10855) ) ;
INV     gate7270  (.A(g10855), .Z(II16735) ) ;
INV     gate7271  (.A(II16735), .Z(g11014) ) ;
OR2     gate7272  (.A(g6083), .B(g10737), .Z(g10856) ) ;
INV     gate7273  (.A(g10856), .Z(II16739) ) ;
INV     gate7274  (.A(II16739), .Z(g11016) ) ;
OR2     gate7275  (.A(g6090), .B(g10738), .Z(g10857) ) ;
INV     gate7276  (.A(g10857), .Z(II16742) ) ;
INV     gate7277  (.A(II16742), .Z(g11017) ) ;
INV     gate7278  (.A(g10888), .Z(II16760) ) ;
INV     gate7279  (.A(g10890), .Z(II16763) ) ;
INV     gate7280  (.A(g10892), .Z(II16766) ) ;
INV     gate7281  (.A(g10894), .Z(II16769) ) ;
INV     gate7282  (.A(g10887), .Z(II16772) ) ;
INV     gate7283  (.A(g10889), .Z(II16775) ) ;
INV     gate7284  (.A(g10891), .Z(II16778) ) ;
INV     gate7285  (.A(g10893), .Z(II16781) ) ;
INV     gate7286  (.A(g10895), .Z(II16784) ) ;
INV     gate7287  (.A(g10896), .Z(II16787) ) ;
INV     gate7288  (.A(g10900), .Z(II16790) ) ;
INV     gate7289  (.A(g11014), .Z(II16793) ) ;
INV     gate7290  (.A(g11016), .Z(II16796) ) ;
INV     gate7291  (.A(g11017), .Z(II16799) ) ;
INV     gate7292  (.A(g10902), .Z(II16802) ) ;
INV     gate7293  (.A(g10904), .Z(II16805) ) ;
INV     gate7294  (.A(g10906), .Z(II16808) ) ;
INV     gate7295  (.A(g10908), .Z(II16811) ) ;
INV     gate7296  (.A(g10910), .Z(II16814) ) ;
INV     gate7297  (.A(g10912), .Z(II16817) ) ;
AND2    gate7298  (.A(g10788), .B(g6355), .Z(g10950) ) ;
INV     gate7299  (.A(g10950), .Z(g11053) ) ;
INV     gate7300  (.A(g10950), .Z(g11054) ) ;
INV     gate7301  (.A(g10950), .Z(g11055) ) ;
INV     gate7302  (.A(g10950), .Z(g11056) ) ;
AND2    gate7303  (.A(g4822), .B(g10822), .Z(g10937) ) ;
INV     gate7304  (.A(g10937), .Z(g11057) ) ;
INV     gate7305  (.A(g10974), .Z(g11059) ) ;
INV     gate7306  (.A(g10937), .Z(g11060) ) ;
INV     gate7307  (.A(g10974), .Z(g11061) ) ;
INV     gate7308  (.A(g10937), .Z(g11062) ) ;
INV     gate7309  (.A(g10974), .Z(g11063) ) ;
INV     gate7310  (.A(g10974), .Z(g11064) ) ;
INV     gate7311  (.A(g10974), .Z(g11065) ) ;
INV     gate7312  (.A(g10974), .Z(g11066) ) ;
INV     gate7313  (.A(g10974), .Z(g11067) ) ;
INV     gate7314  (.A(g10974), .Z(g11068) ) ;
INV     gate7315  (.A(g10974), .Z(g11069) ) ;
INV     gate7316  (.A(g10913), .Z(g11071) ) ;
INV     gate7317  (.A(g10913), .Z(g11072) ) ;
INV     gate7318  (.A(g10913), .Z(g11073) ) ;
INV     gate7319  (.A(g10901), .Z(g11074) ) ;
INV     gate7320  (.A(g10937), .Z(g11075) ) ;
OR2     gate7321  (.A(g4220), .B(g10777), .Z(g10898) ) ;
INV     gate7322  (.A(g10898), .Z(II16843) ) ;
INV     gate7323  (.A(II16843), .Z(g11076) ) ;
NAND2   gate7324  (.A(g10807), .B(g10805), .Z(g10886) ) ;
INV     gate7325  (.A(g10886), .Z(II16847) ) ;
INV     gate7326  (.A(II16847), .Z(g11078) ) ;
INV     gate7327  (.A(g10905), .Z(II16850) ) ;
INV     gate7328  (.A(II16850), .Z(g11079) ) ;
INV     gate7329  (.A(g10907), .Z(II16853) ) ;
INV     gate7330  (.A(II16853), .Z(g11080) ) ;
INV     gate7331  (.A(g10909), .Z(II16856) ) ;
INV     gate7332  (.A(II16856), .Z(g11081) ) ;
INV     gate7333  (.A(g10911), .Z(II16859) ) ;
INV     gate7334  (.A(II16859), .Z(g11082) ) ;
INV     gate7335  (.A(g10913), .Z(g11083) ) ;
INV     gate7336  (.A(g10972), .Z(II16863) ) ;
INV     gate7337  (.A(II16863), .Z(g11084) ) ;
INV     gate7338  (.A(g10913), .Z(II16867) ) ;
INV     gate7339  (.A(II16867), .Z(g11086) ) ;
INV     gate7340  (.A(g10973), .Z(II16871) ) ;
INV     gate7341  (.A(II16871), .Z(g11088) ) ;
OR2     gate7342  (.A(g5170), .B(g10808), .Z(g10936) ) ;
INV     gate7343  (.A(g10936), .Z(II16879) ) ;
INV     gate7344  (.A(II16879), .Z(g11096) ) ;
INV     gate7345  (.A(g10974), .Z(g11106) ) ;
INV     gate7346  (.A(g10974), .Z(g11107) ) ;
INV     gate7347  (.A(g10974), .Z(g11108) ) ;
INV     gate7348  (.A(g10974), .Z(g11109) ) ;
INV     gate7349  (.A(g10974), .Z(g11110) ) ;
INV     gate7350  (.A(g10974), .Z(g11111) ) ;
INV     gate7351  (.A(g10947), .Z(II16897) ) ;
INV     gate7352  (.A(II16897), .Z(g11112) ) ;
INV     gate7353  (.A(g10950), .Z(g11155) ) ;
INV     gate7354  (.A(g10950), .Z(g11157) ) ;
INV     gate7355  (.A(g10950), .Z(g11159) ) ;
INV     gate7356  (.A(g10950), .Z(g11160) ) ;
INV     gate7357  (.A(g10950), .Z(g11162) ) ;
INV     gate7358  (.A(g11084), .Z(II16920) ) ;
INV     gate7359  (.A(g11086), .Z(II16938) ) ;
INV     gate7360  (.A(g11076), .Z(II16941) ) ;
INV     gate7361  (.A(g11079), .Z(II16944) ) ;
INV     gate7362  (.A(g11080), .Z(II16947) ) ;
INV     gate7363  (.A(g11081), .Z(II16950) ) ;
INV     gate7364  (.A(g11082), .Z(II16953) ) ;
INV     gate7365  (.A(g11096), .Z(II16956) ) ;
INV     gate7366  (.A(g11112), .Z(g11191) ) ;
INV     gate7367  (.A(g11112), .Z(g11193) ) ;
INV     gate7368  (.A(g11112), .Z(g11195) ) ;
INV     gate7369  (.A(g11112), .Z(g11197) ) ;
INV     gate7370  (.A(g11112), .Z(g11199) ) ;
INV     gate7371  (.A(g11112), .Z(g11200) ) ;
INV     gate7372  (.A(g11112), .Z(g11202) ) ;
INV     gate7373  (.A(g11112), .Z(g11203) ) ;
INV     gate7374  (.A(g11112), .Z(g11205) ) ;
INV     gate7375  (.A(g11088), .Z(II16979) ) ;
INV     gate7376  (.A(g11088), .Z(II16982) ) ;
INV     gate7377  (.A(II16982), .Z(g11207) ) ;
NOR2    gate7378  (.A(g10970), .B(g10971), .Z(g11077) ) ;
INV     gate7379  (.A(g11077), .Z(g11208) ) ;
INV     gate7380  (.A(g11112), .Z(g11239) ) ;
INV     gate7381  (.A(g11112), .Z(g11241) ) ;
INV     gate7382  (.A(g11112), .Z(g11242) ) ;
INV     gate7383  (.A(g11112), .Z(g11243) ) ;
INV     gate7384  (.A(g11112), .Z(g11244) ) ;
INV     gate7385  (.A(g11112), .Z(g11245) ) ;
INV     gate7386  (.A(g11208), .Z(g11284) ) ;
INV     gate7387  (.A(g11207), .Z(g11287) ) ;
OR2     gate7388  (.A(g11085), .B(g10946), .Z(g11233) ) ;
INV     gate7389  (.A(g11233), .Z(II17070) ) ;
INV     gate7390  (.A(II17070), .Z(g11289) ) ;
OR2     gate7391  (.A(g6162), .B(g11143), .Z(g11249) ) ;
INV     gate7392  (.A(g11249), .Z(II17084) ) ;
INV     gate7393  (.A(II17084), .Z(g11301) ) ;
OR2     gate7394  (.A(g11144), .B(g11005), .Z(g11217) ) ;
INV     gate7395  (.A(g11217), .Z(II17092) ) ;
INV     gate7396  (.A(II17092), .Z(g11307) ) ;
OR2     gate7397  (.A(g11145), .B(g11006), .Z(g11219) ) ;
INV     gate7398  (.A(g11219), .Z(II17096) ) ;
INV     gate7399  (.A(II17096), .Z(g11309) ) ;
OR2     gate7400  (.A(g11146), .B(g11007), .Z(g11221) ) ;
INV     gate7401  (.A(g11221), .Z(II17100) ) ;
INV     gate7402  (.A(II17100), .Z(g11311) ) ;
OR2     gate7403  (.A(g11147), .B(g11008), .Z(g11223) ) ;
INV     gate7404  (.A(g11223), .Z(II17104) ) ;
INV     gate7405  (.A(II17104), .Z(g11313) ) ;
OR2     gate7406  (.A(g11149), .B(g11009), .Z(g11225) ) ;
INV     gate7407  (.A(g11225), .Z(II17108) ) ;
INV     gate7408  (.A(II17108), .Z(g11315) ) ;
OR2     gate7409  (.A(g11151), .B(g11010), .Z(g11227) ) ;
INV     gate7410  (.A(g11227), .Z(II17112) ) ;
INV     gate7411  (.A(II17112), .Z(g11317) ) ;
OR2     gate7412  (.A(g11154), .B(g11012), .Z(g11229) ) ;
INV     gate7413  (.A(g11229), .Z(II17116) ) ;
INV     gate7414  (.A(II17116), .Z(g11319) ) ;
OR2     gate7415  (.A(g11156), .B(g11013), .Z(g11231) ) ;
INV     gate7416  (.A(g11231), .Z(II17121) ) ;
INV     gate7417  (.A(II17121), .Z(g11322) ) ;
OR2     gate7418  (.A(g11158), .B(g11015), .Z(g11232) ) ;
INV     gate7419  (.A(g11232), .Z(II17124) ) ;
INV     gate7420  (.A(II17124), .Z(g11323) ) ;
INV     gate7421  (.A(g11301), .Z(II17142) ) ;
INV     gate7422  (.A(II17142), .Z(g11339) ) ;
OR2     gate7423  (.A(g11215), .B(g11093), .Z(g11305) ) ;
INV     gate7424  (.A(g11305), .Z(II17146) ) ;
INV     gate7425  (.A(II17146), .Z(g11341) ) ;
OR2     gate7426  (.A(g11216), .B(g11095), .Z(g11306) ) ;
INV     gate7427  (.A(g11306), .Z(II17149) ) ;
INV     gate7428  (.A(II17149), .Z(g11342) ) ;
OR2     gate7429  (.A(g11218), .B(g11098), .Z(g11308) ) ;
INV     gate7430  (.A(g11308), .Z(II17152) ) ;
INV     gate7431  (.A(II17152), .Z(g11343) ) ;
OR2     gate7432  (.A(g11220), .B(g11100), .Z(g11310) ) ;
INV     gate7433  (.A(g11310), .Z(II17155) ) ;
INV     gate7434  (.A(II17155), .Z(g11344) ) ;
OR2     gate7435  (.A(g11222), .B(g11101), .Z(g11312) ) ;
INV     gate7436  (.A(g11312), .Z(II17158) ) ;
INV     gate7437  (.A(II17158), .Z(g11345) ) ;
OR2     gate7438  (.A(g11224), .B(g11102), .Z(g11314) ) ;
INV     gate7439  (.A(g11314), .Z(II17161) ) ;
INV     gate7440  (.A(II17161), .Z(g11346) ) ;
AND2    gate7441  (.A(g11201), .B(g4379), .Z(g11320) ) ;
INV     gate7442  (.A(g11320), .Z(II17164) ) ;
INV     gate7443  (.A(II17164), .Z(g11347) ) ;
NAND2   gate7444  (.A(II17052), .B(II17053), .Z(g11276) ) ;
INV     gate7445  (.A(g11276), .Z(g11348) ) ;
INV     gate7446  (.A(g11287), .Z(g11350) ) ;
OR2     gate7447  (.A(g6576), .B(g11210), .Z(g11294) ) ;
INV     gate7448  (.A(g11294), .Z(II17170) ) ;
INV     gate7449  (.A(II17170), .Z(g11351) ) ;
OR2     gate7450  (.A(g11211), .B(g10818), .Z(g11293) ) ;
INV     gate7451  (.A(g11293), .Z(II17173) ) ;
INV     gate7452  (.A(II17173), .Z(g11352) ) ;
OR2     gate7453  (.A(g10670), .B(g11209), .Z(g11286) ) ;
INV     gate7454  (.A(g11286), .Z(II17176) ) ;
INV     gate7455  (.A(II17176), .Z(g11353) ) ;
INV     gate7456  (.A(g11307), .Z(II17179) ) ;
INV     gate7457  (.A(II17179), .Z(g11354) ) ;
INV     gate7458  (.A(g11309), .Z(II17182) ) ;
INV     gate7459  (.A(II17182), .Z(g11357) ) ;
INV     gate7460  (.A(g11311), .Z(II17185) ) ;
INV     gate7461  (.A(II17185), .Z(g11360) ) ;
INV     gate7462  (.A(g11313), .Z(II17188) ) ;
INV     gate7463  (.A(II17188), .Z(g11363) ) ;
INV     gate7464  (.A(g11315), .Z(II17191) ) ;
INV     gate7465  (.A(II17191), .Z(g11366) ) ;
INV     gate7466  (.A(g11317), .Z(II17194) ) ;
INV     gate7467  (.A(II17194), .Z(g11369) ) ;
INV     gate7468  (.A(g11319), .Z(II17198) ) ;
INV     gate7469  (.A(II17198), .Z(g11373) ) ;
INV     gate7470  (.A(g11322), .Z(II17202) ) ;
INV     gate7471  (.A(II17202), .Z(g11377) ) ;
INV     gate7472  (.A(g11323), .Z(II17206) ) ;
INV     gate7473  (.A(II17206), .Z(g11381) ) ;
INV     gate7474  (.A(g11289), .Z(II17209) ) ;
INV     gate7475  (.A(II17209), .Z(g11384) ) ;
AND2    gate7476  (.A(g11246), .B(g4226), .Z(g11290) ) ;
INV     gate7477  (.A(g11290), .Z(II17213) ) ;
INV     gate7478  (.A(II17213), .Z(g11388) ) ;
AND2    gate7479  (.A(g11247), .B(g4233), .Z(g11291) ) ;
INV     gate7480  (.A(g11291), .Z(II17216) ) ;
INV     gate7481  (.A(II17216), .Z(g11389) ) ;
AND2    gate7482  (.A(g11252), .B(g4250), .Z(g11292) ) ;
INV     gate7483  (.A(g11292), .Z(II17219) ) ;
INV     gate7484  (.A(II17219), .Z(g11390) ) ;
OR2     gate7485  (.A(g11212), .B(g11087), .Z(g11298) ) ;
INV     gate7486  (.A(g11298), .Z(II17225) ) ;
INV     gate7487  (.A(II17225), .Z(g11394) ) ;
OR2     gate7488  (.A(g11213), .B(g11091), .Z(g11300) ) ;
INV     gate7489  (.A(g11300), .Z(II17228) ) ;
INV     gate7490  (.A(II17228), .Z(g11395) ) ;
OR2     gate7491  (.A(g11214), .B(g11092), .Z(g11303) ) ;
INV     gate7492  (.A(g11303), .Z(II17231) ) ;
INV     gate7493  (.A(II17231), .Z(g11396) ) ;
INV     gate7494  (.A(g11353), .Z(II17234) ) ;
INV     gate7495  (.A(g11394), .Z(II17237) ) ;
INV     gate7496  (.A(g11395), .Z(II17240) ) ;
INV     gate7497  (.A(g11396), .Z(II17243) ) ;
INV     gate7498  (.A(g11341), .Z(II17246) ) ;
INV     gate7499  (.A(g11342), .Z(II17249) ) ;
INV     gate7500  (.A(g11343), .Z(II17252) ) ;
INV     gate7501  (.A(g11344), .Z(II17255) ) ;
INV     gate7502  (.A(g11345), .Z(II17258) ) ;
INV     gate7503  (.A(g11346), .Z(II17261) ) ;
INV     gate7504  (.A(g11352), .Z(II17265) ) ;
INV     gate7505  (.A(g11351), .Z(II17268) ) ;
INV     gate7506  (.A(g11388), .Z(II17271) ) ;
INV     gate7507  (.A(II17271), .Z(g11410) ) ;
INV     gate7508  (.A(g11389), .Z(II17274) ) ;
INV     gate7509  (.A(II17274), .Z(g11411) ) ;
INV     gate7510  (.A(g11390), .Z(II17277) ) ;
INV     gate7511  (.A(II17277), .Z(g11412) ) ;
AND2    gate7512  (.A(g11275), .B(g7912), .Z(g11391) ) ;
INV     gate7513  (.A(g11391), .Z(II17302) ) ;
INV     gate7514  (.A(II17302), .Z(g11417) ) ;
AND2    gate7515  (.A(g11278), .B(g7914), .Z(g11392) ) ;
INV     gate7516  (.A(g11392), .Z(II17312) ) ;
INV     gate7517  (.A(II17312), .Z(g11419) ) ;
AND2    gate7518  (.A(g11280), .B(g7916), .Z(g11393) ) ;
INV     gate7519  (.A(g11393), .Z(II17315) ) ;
INV     gate7520  (.A(II17315), .Z(g11420) ) ;
AND2    gate7521  (.A(g11285), .B(g4424), .Z(g11340) ) ;
INV     gate7522  (.A(g11340), .Z(II17318) ) ;
INV     gate7523  (.A(II17318), .Z(g11421) ) ;
INV     gate7524  (.A(g11348), .Z(II17321) ) ;
INV     gate7525  (.A(II17321), .Z(g11422) ) ;
INV     gate7526  (.A(g11347), .Z(II17324) ) ;
INV     gate7527  (.A(II17324), .Z(g11423) ) ;
AND2    gate7528  (.A(g11288), .B(g7964), .Z(g11349) ) ;
INV     gate7529  (.A(g11349), .Z(II17327) ) ;
INV     gate7530  (.A(II17327), .Z(g11424) ) ;
INV     gate7531  (.A(g11357), .Z(II17331) ) ;
INV     gate7532  (.A(II17331), .Z(g11426) ) ;
INV     gate7533  (.A(g11360), .Z(II17334) ) ;
INV     gate7534  (.A(II17334), .Z(g11427) ) ;
INV     gate7535  (.A(g11363), .Z(II17337) ) ;
INV     gate7536  (.A(II17337), .Z(g11428) ) ;
INV     gate7537  (.A(g11366), .Z(II17340) ) ;
INV     gate7538  (.A(II17340), .Z(g11429) ) ;
INV     gate7539  (.A(g11369), .Z(II17344) ) ;
INV     gate7540  (.A(II17344), .Z(g11431) ) ;
INV     gate7541  (.A(g11373), .Z(II17347) ) ;
INV     gate7542  (.A(II17347), .Z(g11432) ) ;
INV     gate7543  (.A(g11377), .Z(II17350) ) ;
INV     gate7544  (.A(II17350), .Z(g11433) ) ;
INV     gate7545  (.A(g11381), .Z(II17353) ) ;
INV     gate7546  (.A(II17353), .Z(g11434) ) ;
INV     gate7547  (.A(g11384), .Z(II17356) ) ;
INV     gate7548  (.A(II17356), .Z(g11435) ) ;
AND2    gate7549  (.A(g11316), .B(g4266), .Z(g11372) ) ;
INV     gate7550  (.A(g11372), .Z(II17359) ) ;
INV     gate7551  (.A(II17359), .Z(g11436) ) ;
AND2    gate7552  (.A(g11318), .B(g4277), .Z(g11376) ) ;
INV     gate7553  (.A(g11376), .Z(II17362) ) ;
INV     gate7554  (.A(II17362), .Z(g11437) ) ;
AND2    gate7555  (.A(g11321), .B(g4285), .Z(g11380) ) ;
INV     gate7556  (.A(g11380), .Z(II17365) ) ;
INV     gate7557  (.A(II17365), .Z(g11438) ) ;
INV     gate7558  (.A(g11423), .Z(II17368) ) ;
INV     gate7559  (.A(g11410), .Z(II17371) ) ;
INV     gate7560  (.A(g11411), .Z(II17374) ) ;
INV     gate7561  (.A(g11412), .Z(II17377) ) ;
INV     gate7562  (.A(g11436), .Z(II17381) ) ;
INV     gate7563  (.A(II17381), .Z(g11444) ) ;
INV     gate7564  (.A(g11437), .Z(II17384) ) ;
INV     gate7565  (.A(II17384), .Z(g11445) ) ;
INV     gate7566  (.A(g11438), .Z(II17387) ) ;
INV     gate7567  (.A(II17387), .Z(g11446) ) ;
OR2     gate7568  (.A(g11387), .B(g4006), .Z(g11430) ) ;
INV     gate7569  (.A(g11430), .Z(II17390) ) ;
INV     gate7570  (.A(II17390), .Z(g11447) ) ;
INV     gate7571  (.A(g11417), .Z(II17407) ) ;
INV     gate7572  (.A(II17407), .Z(g11450) ) ;
INV     gate7573  (.A(g11419), .Z(II17410) ) ;
INV     gate7574  (.A(II17410), .Z(g11451) ) ;
AND2    gate7575  (.A(g11350), .B(g10899), .Z(g11425) ) ;
INV     gate7576  (.A(g11425), .Z(II17413) ) ;
INV     gate7577  (.A(II17413), .Z(g11452) ) ;
INV     gate7578  (.A(g11420), .Z(II17416) ) ;
INV     gate7579  (.A(II17416), .Z(g11453) ) ;
INV     gate7580  (.A(g11421), .Z(II17419) ) ;
INV     gate7581  (.A(II17419), .Z(g11454) ) ;
INV     gate7582  (.A(g11424), .Z(II17424) ) ;
INV     gate7583  (.A(II17424), .Z(g11457) ) ;
INV     gate7584  (.A(g11454), .Z(II17435) ) ;
INV     gate7585  (.A(g11444), .Z(II17438) ) ;
INV     gate7586  (.A(g11445), .Z(II17441) ) ;
INV     gate7587  (.A(g11446), .Z(II17444) ) ;
INV     gate7588  (.A(g11457), .Z(II17447) ) ;
INV     gate7589  (.A(g11450), .Z(II17450) ) ;
INV     gate7590  (.A(g11451), .Z(II17453) ) ;
INV     gate7591  (.A(g11453), .Z(II17456) ) ;
INV     gate7592  (.A(g11447), .Z(II17466) ) ;
INV     gate7593  (.A(II17466), .Z(g11475) ) ;
INV     gate7594  (.A(g11452), .Z(II17470) ) ;
INV     gate7595  (.A(II17470), .Z(g11479) ) ;
INV     gate7596  (.A(g11479), .Z(II17482) ) ;
OR2     gate7597  (.A(g6532), .B(g11455), .Z(g11478) ) ;
INV     gate7598  (.A(g11478), .Z(II17500) ) ;
INV     gate7599  (.A(II17500), .Z(g11495) ) ;
OR2     gate7600  (.A(g6624), .B(g11458), .Z(g11481) ) ;
INV     gate7601  (.A(g11481), .Z(II17510) ) ;
INV     gate7602  (.A(II17510), .Z(g11497) ) ;
OR2     gate7603  (.A(g6628), .B(g11459), .Z(g11482) ) ;
INV     gate7604  (.A(g11482), .Z(II17513) ) ;
INV     gate7605  (.A(II17513), .Z(g11498) ) ;
OR2     gate7606  (.A(g6633), .B(g11460), .Z(g11483) ) ;
INV     gate7607  (.A(g11483), .Z(II17516) ) ;
INV     gate7608  (.A(II17516), .Z(g11499) ) ;
OR2     gate7609  (.A(g6639), .B(g11461), .Z(g11484) ) ;
INV     gate7610  (.A(g11484), .Z(II17519) ) ;
INV     gate7611  (.A(II17519), .Z(g11500) ) ;
OR2     gate7612  (.A(g6646), .B(g11462), .Z(g11485) ) ;
INV     gate7613  (.A(g11485), .Z(II17522) ) ;
INV     gate7614  (.A(II17522), .Z(g11501) ) ;
OR2     gate7615  (.A(g6654), .B(g11463), .Z(g11486) ) ;
INV     gate7616  (.A(g11486), .Z(II17525) ) ;
INV     gate7617  (.A(II17525), .Z(g11502) ) ;
OR2     gate7618  (.A(g6662), .B(g11464), .Z(g11487) ) ;
INV     gate7619  (.A(g11487), .Z(II17528) ) ;
INV     gate7620  (.A(II17528), .Z(g11503) ) ;
OR2     gate7621  (.A(g6671), .B(g11465), .Z(g11488) ) ;
INV     gate7622  (.A(g11488), .Z(II17531) ) ;
INV     gate7623  (.A(II17531), .Z(g11504) ) ;
INV     gate7624  (.A(g11495), .Z(II17534) ) ;
INV     gate7625  (.A(g11497), .Z(II17537) ) ;
INV     gate7626  (.A(g11498), .Z(II17540) ) ;
INV     gate7627  (.A(g11499), .Z(II17543) ) ;
INV     gate7628  (.A(g11500), .Z(II17546) ) ;
INV     gate7629  (.A(g11501), .Z(II17549) ) ;
INV     gate7630  (.A(g11502), .Z(II17552) ) ;
INV     gate7631  (.A(g11503), .Z(II17555) ) ;
INV     gate7632  (.A(g11504), .Z(II17558) ) ;
NAND2   gate7633  (.A(II17486), .B(II17487), .Z(g11490) ) ;
INV     gate7634  (.A(g11490), .Z(g11515) ) ;
AND2    gate7635  (.A(g11480), .B(g4807), .Z(g11492) ) ;
INV     gate7636  (.A(g11492), .Z(II17563) ) ;
INV     gate7637  (.A(II17563), .Z(g11518) ) ;
AND3    gate7638  (.A(g1317), .B(g3015), .C(g11492), .Z(g11519) ) ;
INV     gate7639  (.A(g11519), .Z(g11539) ) ;
INV     gate7640  (.A(g11519), .Z(g11540) ) ;
INV     gate7641  (.A(g11519), .Z(g11541) ) ;
INV     gate7642  (.A(g11519), .Z(g11542) ) ;
INV     gate7643  (.A(g11519), .Z(g11543) ) ;
INV     gate7644  (.A(g11519), .Z(g11545) ) ;
INV     gate7645  (.A(g11519), .Z(g11546) ) ;
INV     gate7646  (.A(g11519), .Z(g11547) ) ;
INV     gate7647  (.A(g11519), .Z(g11548) ) ;
AND2    gate7648  (.A(g11491), .B(g5151), .Z(g11514) ) ;
INV     gate7649  (.A(g11514), .Z(II17591) ) ;
INV     gate7650  (.A(II17591), .Z(g11550) ) ;
AND2    gate7651  (.A(g11518), .B(g3015), .Z(g11561) ) ;
INV     gate7652  (.A(g11561), .Z(g11572) ) ;
INV     gate7653  (.A(g11561), .Z(g11573) ) ;
INV     gate7654  (.A(g11561), .Z(g11574) ) ;
INV     gate7655  (.A(g11561), .Z(g11575) ) ;
NAND2   gate7656  (.A(II17585), .B(II17586), .Z(g11549) ) ;
INV     gate7657  (.A(g11549), .Z(II17610) ) ;
INV     gate7658  (.A(II17610), .Z(g11576) ) ;
INV     gate7659  (.A(g11550), .Z(II17613) ) ;
INV     gate7660  (.A(II17613), .Z(g11577) ) ;
INV     gate7661  (.A(g11561), .Z(II17616) ) ;
INV     gate7662  (.A(II17616), .Z(g11578) ) ;
INV     gate7663  (.A(g11578), .Z(II17633) ) ;
INV     gate7664  (.A(g11577), .Z(II17636) ) ;
OR2     gate7665  (.A(g11413), .B(g11544), .Z(g11580) ) ;
INV     gate7666  (.A(g11580), .Z(g11596) ) ;
OR2     gate7667  (.A(g5123), .B(g11551), .Z(g11579) ) ;
INV     gate7668  (.A(g11579), .Z(II17642) ) ;
INV     gate7669  (.A(II17642), .Z(g11598) ) ;
INV     gate7670  (.A(g11598), .Z(II17657) ) ;
OR2     gate7671  (.A(g11581), .B(g11552), .Z(g11602) ) ;
INV     gate7672  (.A(g11602), .Z(II17662) ) ;
INV     gate7673  (.A(II17662), .Z(g11614) ) ;
OR2     gate7674  (.A(g11582), .B(g11553), .Z(g11603) ) ;
INV     gate7675  (.A(g11603), .Z(II17666) ) ;
INV     gate7676  (.A(II17666), .Z(g11616) ) ;
OR2     gate7677  (.A(g11583), .B(g11554), .Z(g11604) ) ;
INV     gate7678  (.A(g11604), .Z(II17669) ) ;
INV     gate7679  (.A(II17669), .Z(g11617) ) ;
OR2     gate7680  (.A(g11584), .B(g11555), .Z(g11605) ) ;
INV     gate7681  (.A(g11605), .Z(II17672) ) ;
INV     gate7682  (.A(II17672), .Z(g11618) ) ;
OR2     gate7683  (.A(g11585), .B(g11556), .Z(g11606) ) ;
INV     gate7684  (.A(g11606), .Z(II17675) ) ;
INV     gate7685  (.A(II17675), .Z(g11619) ) ;
OR2     gate7686  (.A(g11586), .B(g11557), .Z(g11607) ) ;
INV     gate7687  (.A(g11607), .Z(II17678) ) ;
INV     gate7688  (.A(II17678), .Z(g11620) ) ;
OR2     gate7689  (.A(g11587), .B(g11558), .Z(g11608) ) ;
INV     gate7690  (.A(g11608), .Z(II17681) ) ;
INV     gate7691  (.A(II17681), .Z(g11621) ) ;
OR2     gate7692  (.A(g11588), .B(g11559), .Z(g11609) ) ;
INV     gate7693  (.A(g11609), .Z(II17684) ) ;
INV     gate7694  (.A(II17684), .Z(g11622) ) ;
OR2     gate7695  (.A(g11589), .B(g11560), .Z(g11610) ) ;
INV     gate7696  (.A(g11610), .Z(II17687) ) ;
INV     gate7697  (.A(II17687), .Z(g11623) ) ;
INV     gate7698  (.A(g11596), .Z(II17692) ) ;
INV     gate7699  (.A(II17692), .Z(g11626) ) ;
INV     gate7700  (.A(g11614), .Z(II17695) ) ;
INV     gate7701  (.A(g11616), .Z(II17698) ) ;
INV     gate7702  (.A(g11617), .Z(II17701) ) ;
INV     gate7703  (.A(g11618), .Z(II17704) ) ;
INV     gate7704  (.A(g11619), .Z(II17707) ) ;
INV     gate7705  (.A(g11620), .Z(II17710) ) ;
INV     gate7706  (.A(g11621), .Z(II17713) ) ;
INV     gate7707  (.A(g11622), .Z(II17716) ) ;
INV     gate7708  (.A(g11623), .Z(II17719) ) ;
OR2     gate7709  (.A(g6535), .B(g11597), .Z(g11625) ) ;
INV     gate7710  (.A(g11625), .Z(II17724) ) ;
INV     gate7711  (.A(II17724), .Z(g11638) ) ;
INV     gate7712  (.A(g11638), .Z(II17730) ) ;
AND2    gate7713  (.A(g11612), .B(g7897), .Z(g11639) ) ;
INV     gate7714  (.A(g11639), .Z(II17733) ) ;
INV     gate7715  (.A(II17733), .Z(g11643) ) ;
AND2    gate7716  (.A(g11613), .B(g7900), .Z(g11640) ) ;
INV     gate7717  (.A(g11640), .Z(II17736) ) ;
INV     gate7718  (.A(II17736), .Z(g11644) ) ;
AND2    gate7719  (.A(g11615), .B(g7901), .Z(g11641) ) ;
INV     gate7720  (.A(g11641), .Z(II17739) ) ;
INV     gate7721  (.A(II17739), .Z(g11645) ) ;
AND2    gate7722  (.A(g11624), .B(g7936), .Z(g11636) ) ;
INV     gate7723  (.A(g11636), .Z(II17742) ) ;
INV     gate7724  (.A(II17742), .Z(g11646) ) ;
INV     gate7725  (.A(g11643), .Z(II17746) ) ;
INV     gate7726  (.A(II17746), .Z(g11648) ) ;
INV     gate7727  (.A(g11644), .Z(II17749) ) ;
INV     gate7728  (.A(II17749), .Z(g11649) ) ;
INV     gate7729  (.A(g11645), .Z(II17752) ) ;
INV     gate7730  (.A(II17752), .Z(g11650) ) ;
INV     gate7731  (.A(g11646), .Z(II17755) ) ;
INV     gate7732  (.A(II17755), .Z(g11651) ) ;
OR2     gate7733  (.A(g6622), .B(g11637), .Z(g11647) ) ;
INV     gate7734  (.A(g11647), .Z(II17758) ) ;
INV     gate7735  (.A(II17758), .Z(g11652) ) ;
INV     gate7736  (.A(g11652), .Z(II17761) ) ;
INV     gate7737  (.A(g11651), .Z(II17764) ) ;
INV     gate7738  (.A(g11648), .Z(II17767) ) ;
INV     gate7739  (.A(g11649), .Z(II17770) ) ;
INV     gate7740  (.A(g11650), .Z(II17773) ) ;
AND2    gate7741  (.A(g932), .B(g928), .Z(g2081) ) ;
AND2    gate7742  (.A(g976), .B(g971), .Z(g2091) ) ;
AND2    gate7743  (.A(g1872), .B(g1882), .Z(g2132) ) ;
AND2    gate7744  (.A(g745), .B(g746), .Z(g2160) ) ;
AND4    gate7745  (.A(g1462), .B(g1470), .C(g1474), .D(g1478), .Z(II5084) ) ;
AND4    gate7746  (.A(g1490), .B(g1494), .C(g1504), .D(g1508), .Z(II5085) ) ;
AND2    gate7747  (.A(g1771), .B(g1766), .Z(g2264) ) ;
AND2    gate7748  (.A(g1223), .B(g1218), .Z(g2306) ) ;
AND2    gate7749  (.A(g744), .B(g743), .Z(g2379) ) ;
AND2    gate7750  (.A(g374), .B(g369), .Z(g2496) ) ;
AND2    gate7751  (.A(g461), .B(g456), .Z(g2511) ) ;
AND2    gate7752  (.A(g762), .B(g758), .Z(g2525) ) ;
AND2    gate7753  (.A(g658), .B(g668), .Z(g2531) ) ;
AND2    gate7754  (.A(g798), .B(g794), .Z(g2534) ) ;
AND2    gate7755  (.A(g1341), .B(g1336), .Z(g2544) ) ;
AND2    gate7756  (.A(g742), .B(g741), .Z(g2561) ) ;
AND4    gate7757  (.A(g1419), .B(g1424), .C(g1428), .D(g1432), .Z(II5689) ) ;
AND4    gate7758  (.A(g1436), .B(g1440), .C(g1444), .D(g1448), .Z(II5690) ) ;
AND2    gate7759  (.A(g936), .B(g2081), .Z(g2756) ) ;
AND2    gate7760  (.A(g981), .B(g2091), .Z(g2760) ) ;
AND4    gate7761  (.A(g174), .B(g170), .C(g2249), .D(g2254), .Z(II5886) ) ;
AND4    gate7762  (.A(g2078), .B(g2083), .C(g166), .D(g2095), .Z(II5887) ) ;
AND3    gate7763  (.A(g2399), .B(g2369), .C(g591), .Z(g2800) ) ;
AND2    gate7764  (.A(g2132), .B(g1891), .Z(g2804) ) ;
AND2    gate7765  (.A(g1980), .B(g1976), .Z(g2892) ) ;
AND2    gate7766  (.A(g2411), .B(g1678), .Z(g2895) ) ;
AND2    gate7767  (.A(g2424), .B(g1660), .Z(g2910) ) ;
AND2    gate7768  (.A(g2411), .B(g1675), .Z(g2911) ) ;
AND2    gate7769  (.A(g2424), .B(g1657), .Z(g2917) ) ;
AND2    gate7770  (.A(g2411), .B(g1672), .Z(g2918) ) ;
AND2    gate7771  (.A(g2411), .B(g1687), .Z(g2939) ) ;
AND2    gate7772  (.A(g2424), .B(g1654), .Z(g2940) ) ;
AND2    gate7773  (.A(g2424), .B(g1669), .Z(g2944) ) ;
AND2    gate7774  (.A(g2411), .B(g1684), .Z(g2945) ) ;
AND2    gate7775  (.A(g2424), .B(g1666), .Z(g2950) ) ;
AND2    gate7776  (.A(g2411), .B(g1681), .Z(g2951) ) ;
AND2    gate7777  (.A(g2424), .B(g1663), .Z(g2957) ) ;
AND2    gate7778  (.A(g1776), .B(g2264), .Z(g2981) ) ;
AND3    gate7779  (.A(g2061), .B(g2557), .C(g1814), .Z(g2990) ) ;
AND2    gate7780  (.A(g1227), .B(g2306), .Z(g3047) ) ;
AND2    gate7781  (.A(g2054), .B(g2050), .Z(g3089) ) ;
AND2    gate7782  (.A(g2331), .B(g2198), .Z(g3098) ) ;
AND4    gate7783  (.A(g2446), .B(g2451), .C(g2456), .D(g2475), .Z(II6309) ) ;
AND4    gate7784  (.A(g2396), .B(g2407), .C(g2421), .D(g2435), .Z(II6310) ) ;
AND4    gate7785  (.A(g2082), .B(g2087), .C(g2381), .D(g2395), .Z(II6316) ) ;
AND4    gate7786  (.A(g2406), .B(g2420), .C(g2434), .D(g2438), .Z(II6317) ) ;
AND4    gate7787  (.A(g2549), .B(g2556), .C(g2562), .D(g2570), .Z(II6330) ) ;
AND4    gate7788  (.A(g2060), .B(g2070), .C(g2074), .D(g2077), .Z(II6331) ) ;
AND4    gate7789  (.A(g201), .B(g2421), .C(g2407), .D(g2396), .Z(II6337) ) ;
AND4    gate7790  (.A(g2475), .B(g2456), .C(g2451), .D(g2446), .Z(II6338) ) ;
AND2    gate7791  (.A(g378), .B(g2496), .Z(g3257) ) ;
AND2    gate7792  (.A(g2503), .B(g2328), .Z(g3263) ) ;
AND2    gate7793  (.A(g466), .B(g2511), .Z(g3268) ) ;
AND2    gate7794  (.A(g115), .B(g2356), .Z(g3275) ) ;
AND2    gate7795  (.A(g766), .B(g2525), .Z(g3281) ) ;
AND2    gate7796  (.A(g2531), .B(g677), .Z(g3284) ) ;
AND2    gate7797  (.A(g802), .B(g2534), .Z(g3287) ) ;
AND2    gate7798  (.A(g1346), .B(g2544), .Z(g3301) ) ;
AND2    gate7799  (.A(g186), .B(g3228), .Z(g3383) ) ;
AND2    gate7800  (.A(g207), .B(g3228), .Z(g3389) ) ;
AND2    gate7801  (.A(g213), .B(g3228), .Z(g3396) ) ;
AND2    gate7802  (.A(g115), .B(g3164), .Z(g3400) ) ;
AND2    gate7803  (.A(g219), .B(g3228), .Z(g3412) ) ;
AND2    gate7804  (.A(g225), .B(g3228), .Z(g3422) ) ;
AND4    gate7805  (.A(g2677), .B(g2683), .C(g2689), .D(g2701), .Z(II6630) ) ;
AND4    gate7806  (.A(g2707), .B(g2713), .C(g2719), .D(g2765), .Z(II6631) ) ;
AND2    gate7807  (.A(g231), .B(g3228), .Z(g3429) ) ;
AND2    gate7808  (.A(g237), .B(g3228), .Z(g3434) ) ;
AND2    gate7809  (.A(g2804), .B(g1900), .Z(g3497) ) ;
AND2    gate7810  (.A(g2050), .B(g2971), .Z(g3512) ) ;
AND2    gate7811  (.A(g1209), .B(g3015), .Z(g3516) ) ;
AND2    gate7812  (.A(g1981), .B(g2892), .Z(g3533) ) ;
AND2    gate7813  (.A(g2390), .B(g3103), .Z(g3536) ) ;
AND2    gate7814  (.A(g3275), .B(g2126), .Z(g3563) ) ;
AND2    gate7815  (.A(g1710), .B(g3015), .Z(g3684) ) ;
AND2    gate7816  (.A(g1781), .B(g2981), .Z(g3685) ) ;
AND2    gate7817  (.A(g1712), .B(g3015), .Z(g3695) ) ;
AND2    gate7818  (.A(g1713), .B(g3015), .Z(g3696) ) ;
AND2    gate7819  (.A(g1690), .B(g2991), .Z(g3714) ) ;
AND2    gate7820  (.A(g192), .B(g3164), .Z(g3718) ) ;
AND2    gate7821  (.A(g2542), .B(g3089), .Z(g3772) ) ;
AND2    gate7822  (.A(g3098), .B(g2203), .Z(g3804) ) ;
AND2    gate7823  (.A(g3003), .B(g3062), .Z(g3807) ) ;
NAND2   gate7824  (.A(II6144), .B(II6145), .Z(g2948) ) ;
AND2    gate7825  (.A(g2948), .B(g2779), .Z(g3904) ) ;
AND2    gate7826  (.A(g186), .B(g3164), .Z(g3908) ) ;
AND2    gate7827  (.A(g207), .B(g3164), .Z(g3912) ) ;
AND2    gate7828  (.A(g213), .B(g3164), .Z(g3939) ) ;
AND2    gate7829  (.A(g219), .B(g3164), .Z(g3942) ) ;
AND2    gate7830  (.A(g225), .B(g3164), .Z(g3970) ) ;
AND2    gate7831  (.A(g231), .B(g3164), .Z(g3974) ) ;
AND2    gate7832  (.A(g237), .B(g3164), .Z(g3979) ) ;
AND2    gate7833  (.A(g243), .B(g3164), .Z(g3987) ) ;
AND2    gate7834  (.A(g248), .B(g3164), .Z(g3989) ) ;
AND2    gate7835  (.A(g1738), .B(g2774), .Z(g3991) ) ;
AND2    gate7836  (.A(g2677), .B(g2276), .Z(g3998) ) ;
AND2    gate7837  (.A(g1741), .B(g2777), .Z(g3999) ) ;
AND2    gate7838  (.A(g1744), .B(g2778), .Z(g4000) ) ;
AND2    gate7839  (.A(g201), .B(g3228), .Z(g4006) ) ;
AND2    gate7840  (.A(g2683), .B(g2276), .Z(g4007) ) ;
AND2    gate7841  (.A(g2689), .B(g2276), .Z(g4008) ) ;
AND2    gate7842  (.A(g1747), .B(g2789), .Z(g4009) ) ;
AND2    gate7843  (.A(g2695), .B(g2276), .Z(g4047) ) ;
AND2    gate7844  (.A(g1750), .B(g2790), .Z(g4048) ) ;
AND2    gate7845  (.A(g2701), .B(g2276), .Z(g4053) ) ;
AND2    gate7846  (.A(g1753), .B(g2793), .Z(g4054) ) ;
AND2    gate7847  (.A(g2707), .B(g2276), .Z(g4058) ) ;
AND2    gate7848  (.A(g1756), .B(g2796), .Z(g4059) ) ;
AND2    gate7849  (.A(g2713), .B(g2276), .Z(g4063) ) ;
AND2    gate7850  (.A(g1759), .B(g2799), .Z(g4064) ) ;
AND2    gate7851  (.A(g2719), .B(g2276), .Z(g4068) ) ;
AND2    gate7852  (.A(g1762), .B(g2802), .Z(g4069) ) ;
AND2    gate7853  (.A(g3263), .B(g2330), .Z(g4070) ) ;
AND2    gate7854  (.A(g3200), .B(g3222), .Z(g4073) ) ;
AND2    gate7855  (.A(g2765), .B(g2276), .Z(g4079) ) ;
AND2    gate7856  (.A(g2677), .B(g2989), .Z(g4097) ) ;
AND2    gate7857  (.A(g770), .B(g3281), .Z(g4099) ) ;
AND2    gate7858  (.A(g2683), .B(g2997), .Z(g4103) ) ;
AND2    gate7859  (.A(g3284), .B(g686), .Z(g4106) ) ;
AND2    gate7860  (.A(g806), .B(g3287), .Z(g4109) ) ;
AND2    gate7861  (.A(g2689), .B(g3009), .Z(g4115) ) ;
AND2    gate7862  (.A(g2695), .B(g3037), .Z(g4123) ) ;
AND2    gate7863  (.A(g2701), .B(g3040), .Z(g4126) ) ;
AND2    gate7864  (.A(g1976), .B(g2779), .Z(g4128) ) ;
AND2    gate7865  (.A(g2707), .B(g3051), .Z(g4141) ) ;
AND2    gate7866  (.A(g2713), .B(g3055), .Z(g4157) ) ;
AND2    gate7867  (.A(g2719), .B(g3060), .Z(g4161) ) ;
NAND2   gate7868  (.A(II6323), .B(II6324), .Z(g3106) ) ;
AND2    gate7869  (.A(g3106), .B(g2971), .Z(g4162) ) ;
AND2    gate7870  (.A(g2765), .B(g3066), .Z(g4169) ) ;
AND2    gate7871  (.A(g105), .B(g3539), .Z(g4220) ) ;
AND2    gate7872  (.A(g1003), .B(g3914), .Z(g4223) ) ;
AND2    gate7873  (.A(g1092), .B(g3638), .Z(g4224) ) ;
AND2    gate7874  (.A(g999), .B(g3914), .Z(g4229) ) ;
AND2    gate7875  (.A(g1095), .B(g3638), .Z(g4230) ) ;
AND2    gate7876  (.A(g1011), .B(g3914), .Z(g4235) ) ;
AND2    gate7877  (.A(g1098), .B(g3638), .Z(g4236) ) ;
AND2    gate7878  (.A(g1007), .B(g3914), .Z(g4252) ) ;
AND2    gate7879  (.A(g1074), .B(g3638), .Z(g4253) ) ;
AND2    gate7880  (.A(g1019), .B(g3914), .Z(g4261) ) ;
AND2    gate7881  (.A(g1015), .B(g3914), .Z(g4269) ) ;
AND2    gate7882  (.A(g1965), .B(g3400), .Z(g4316) ) ;
AND2    gate7883  (.A(g339), .B(g3586), .Z(g4341) ) ;
AND2    gate7884  (.A(g345), .B(g3586), .Z(g4343) ) ;
AND2    gate7885  (.A(g1169), .B(g3730), .Z(g4345) ) ;
AND2    gate7886  (.A(g3497), .B(g1909), .Z(g4348) ) ;
AND2    gate7887  (.A(g1209), .B(g3747), .Z(g4358) ) ;
AND2    gate7888  (.A(g1861), .B(g3748), .Z(g4360) ) ;
AND2    gate7889  (.A(g1215), .B(g3756), .Z(g4364) ) ;
NAND2   gate7890  (.A(II5619), .B(II5620), .Z(g2517) ) ;
AND2    gate7891  (.A(g2517), .B(g3829), .Z(g4383) ) ;
NAND3   gate7892  (.A(g2310), .B(g3062), .C(g2325), .Z(g3529) ) ;
AND2    gate7893  (.A(g3529), .B(g3092), .Z(g4389) ) ;
NAND2   gate7894  (.A(II6448), .B(II6449), .Z(g3273) ) ;
AND2    gate7895  (.A(g3273), .B(g3829), .Z(g4392) ) ;
AND2    gate7896  (.A(g3475), .B(g2181), .Z(g4397) ) ;
NAND2   gate7897  (.A(II7224), .B(II7225), .Z(g4088) ) ;
AND2    gate7898  (.A(g4088), .B(g3829), .Z(g4400) ) ;
AND2    gate7899  (.A(g2971), .B(g3772), .Z(g4401) ) ;
AND2    gate7900  (.A(g2268), .B(g3533), .Z(g4431) ) ;
AND2    gate7901  (.A(g3723), .B(g1975), .Z(g4432) ) ;
AND2    gate7902  (.A(g1713), .B(g3906), .Z(g4481) ) ;
AND2    gate7903  (.A(g336), .B(g3586), .Z(g4483) ) ;
AND2    gate7904  (.A(g1711), .B(g3910), .Z(g4486) ) ;
AND2    gate7905  (.A(g1718), .B(g3911), .Z(g4487) ) ;
AND2    gate7906  (.A(g348), .B(g3586), .Z(g4489) ) ;
AND2    gate7907  (.A(g1786), .B(g3685), .Z(g4492) ) ;
AND2    gate7908  (.A(g351), .B(g3586), .Z(g4497) ) ;
AND2    gate7909  (.A(g2031), .B(g3938), .Z(g4502) ) ;
AND2    gate7910  (.A(g654), .B(g3943), .Z(g4503) ) ;
AND2    gate7911  (.A(g354), .B(g3586), .Z(g4505) ) ;
AND2    gate7912  (.A(g357), .B(g3586), .Z(g4512) ) ;
AND2    gate7913  (.A(g360), .B(g3586), .Z(g4522) ) ;
AND2    gate7914  (.A(g363), .B(g3586), .Z(g4534) ) ;
AND2    gate7915  (.A(g366), .B(g3586), .Z(g4542) ) ;
AND2    gate7916  (.A(g342), .B(g3586), .Z(g4550) ) ;
AND2    gate7917  (.A(g2034), .B(g3829), .Z(g4559) ) ;
NAND3   gate7918  (.A(g2439), .B(g3222), .C(g2493), .Z(g3766) ) ;
AND2    gate7919  (.A(g3766), .B(g3254), .Z(g4581) ) ;
AND2    gate7920  (.A(g3710), .B(g2322), .Z(g4584) ) ;
NAND2   gate7921  (.A(g611), .B(g617), .Z(g2325) ) ;
AND3    gate7922  (.A(g3056), .B(g3753), .C(g2325), .Z(g4604) ) ;
AND2    gate7923  (.A(g3804), .B(g2212), .Z(g4610) ) ;
NOR3    gate7924  (.A(g3141), .B(g2354), .C(g2353), .Z(g3879) ) ;
AND2    gate7925  (.A(g3275), .B(g3879), .Z(g4617) ) ;
AND2    gate7926  (.A(g192), .B(g3946), .Z(g4670) ) ;
AND2    gate7927  (.A(g1071), .B(g3638), .Z(g4712) ) ;
AND2    gate7928  (.A(g646), .B(g3333), .Z(g4714) ) ;
AND2    gate7929  (.A(g1077), .B(g3638), .Z(g4715) ) ;
AND2    gate7930  (.A(g650), .B(g3343), .Z(g4718) ) ;
AND2    gate7931  (.A(g1023), .B(g3914), .Z(g4720) ) ;
NAND2   gate7932  (.A(II6778), .B(II6779), .Z(g3626) ) ;
AND2    gate7933  (.A(g3626), .B(g2779), .Z(g4723) ) ;
AND2    gate7934  (.A(g1032), .B(g3914), .Z(g4725) ) ;
NAND2   gate7935  (.A(g1834), .B(g1840), .Z(g2493) ) ;
AND3    gate7936  (.A(g3215), .B(g3992), .C(g2493), .Z(g4806) ) ;
AND2    gate7937  (.A(g4070), .B(g2336), .Z(g4816) ) ;
AND2    gate7938  (.A(g186), .B(g3946), .Z(g4820) ) ;
AND2    gate7939  (.A(g207), .B(g3946), .Z(g4823) ) ;
AND2    gate7940  (.A(g774), .B(g4099), .Z(g4824) ) ;
AND2    gate7941  (.A(g213), .B(g3946), .Z(g4827) ) ;
AND2    gate7942  (.A(g4106), .B(g695), .Z(g4828) ) ;
AND2    gate7943  (.A(g810), .B(g4109), .Z(g4831) ) ;
AND2    gate7944  (.A(g219), .B(g3946), .Z(g4834) ) ;
AND2    gate7945  (.A(g643), .B(g3520), .Z(g4836) ) ;
AND2    gate7946  (.A(g1068), .B(g3638), .Z(g4837) ) ;
NOR3    gate7947  (.A(g3291), .B(g2410), .C(g2538), .Z(g4122) ) ;
AND2    gate7948  (.A(g3275), .B(g4122), .Z(g4838) ) ;
AND2    gate7949  (.A(g225), .B(g3946), .Z(g4839) ) ;
AND2    gate7950  (.A(g1080), .B(g3638), .Z(g4865) ) ;
AND2    gate7951  (.A(g231), .B(g3946), .Z(g4866) ) ;
AND2    gate7952  (.A(g1027), .B(g3914), .Z(g4868) ) ;
AND2    gate7953  (.A(g1083), .B(g3638), .Z(g4869) ) ;
AND2    gate7954  (.A(g237), .B(g3946), .Z(g4870) ) ;
AND2    gate7955  (.A(g1864), .B(g3523), .Z(g4871) ) ;
AND2    gate7956  (.A(g995), .B(g3914), .Z(g4875) ) ;
AND2    gate7957  (.A(g1086), .B(g3638), .Z(g4876) ) ;
AND2    gate7958  (.A(g243), .B(g3946), .Z(g4877) ) ;
AND2    gate7959  (.A(g1868), .B(g3531), .Z(g4878) ) ;
AND2    gate7960  (.A(g991), .B(g3914), .Z(g4881) ) ;
AND2    gate7961  (.A(g1089), .B(g3638), .Z(g4882) ) ;
AND2    gate7962  (.A(g248), .B(g3946), .Z(g4883) ) ;
NAND2   gate7963  (.A(II7034), .B(II7035), .Z(g3813) ) ;
AND2    gate7964  (.A(g3813), .B(g2971), .Z(g4884) ) ;
AND2    gate7965  (.A(g1062), .B(g4436), .Z(g4914) ) ;
AND2    gate7966  (.A(g2779), .B(g4431), .Z(g4921) ) ;
AND2    gate7967  (.A(g1065), .B(g4442), .Z(g4932) ) ;
AND2    gate7968  (.A(g1038), .B(g4451), .Z(g4941) ) ;
AND2    gate7969  (.A(g3505), .B(g4449), .Z(g4949) ) ;
AND2    gate7970  (.A(g1415), .B(g4682), .Z(g4950) ) ;
AND2    gate7971  (.A(g1648), .B(g4457), .Z(g4952) ) ;
AND2    gate7972  (.A(g1520), .B(g4682), .Z(g4959) ) ;
AND2    gate7973  (.A(g1403), .B(g4682), .Z(g4960) ) ;
AND2    gate7974  (.A(g1651), .B(g4461), .Z(g4962) ) ;
AND2    gate7975  (.A(g1515), .B(g4682), .Z(g4967) ) ;
AND2    gate7976  (.A(g1432), .B(g4682), .Z(g4968) ) ;
AND2    gate7977  (.A(g1642), .B(g4463), .Z(g4969) ) ;
AND2    gate7978  (.A(g1419), .B(g4682), .Z(g4971) ) ;
AND2    gate7979  (.A(g1436), .B(g4682), .Z(g4972) ) ;
AND2    gate7980  (.A(g1645), .B(g4467), .Z(g4973) ) ;
AND2    gate7981  (.A(g1411), .B(g4682), .Z(g4986) ) ;
AND2    gate7982  (.A(g1440), .B(g4682), .Z(g4987) ) ;
AND2    gate7983  (.A(g1424), .B(g4682), .Z(g4989) ) ;
AND2    gate7984  (.A(g1444), .B(g4682), .Z(g4990) ) ;
AND2    gate7985  (.A(g1508), .B(g4640), .Z(g4991) ) ;
AND2    gate7986  (.A(g1407), .B(g4682), .Z(g4992) ) ;
AND2    gate7987  (.A(g1448), .B(g4682), .Z(g4993) ) ;
AND2    gate7988  (.A(g1504), .B(g4640), .Z(g4994) ) ;
AND2    gate7989  (.A(g1474), .B(g4640), .Z(g4995) ) ;
AND2    gate7990  (.A(g1428), .B(g4682), .Z(g4996) ) ;
AND2    gate7991  (.A(g1499), .B(g4640), .Z(g4999) ) ;
AND2    gate7992  (.A(g1470), .B(g4640), .Z(g5000) ) ;
AND2    gate7993  (.A(g1494), .B(g4640), .Z(g5002) ) ;
AND2    gate7994  (.A(g1466), .B(g4640), .Z(g5003) ) ;
AND2    gate7995  (.A(g1490), .B(g4640), .Z(g5005) ) ;
AND2    gate7996  (.A(g1462), .B(g4640), .Z(g5006) ) ;
AND2    gate7997  (.A(g1486), .B(g4640), .Z(g5009) ) ;
AND2    gate7998  (.A(g1458), .B(g4640), .Z(g5010) ) ;
AND2    gate7999  (.A(g1071), .B(g4511), .Z(g5023) ) ;
AND2    gate8000  (.A(g1482), .B(g4640), .Z(g5025) ) ;
AND2    gate8001  (.A(g1453), .B(g4640), .Z(g5026) ) ;
AND2    gate8002  (.A(g1077), .B(g4521), .Z(g5029) ) ;
AND2    gate8003  (.A(g1478), .B(g4640), .Z(g5031) ) ;
AND2    gate8004  (.A(g3983), .B(g4401), .Z(g5041) ) ;
AND2    gate8005  (.A(g4348), .B(g1918), .Z(g5044) ) ;
AND2    gate8006  (.A(g4432), .B(g2834), .Z(g5051) ) ;
AND2    gate8007  (.A(g305), .B(g4811), .Z(g5067) ) ;
AND2    gate8008  (.A(g1771), .B(g4587), .Z(g5074) ) ;
AND2    gate8009  (.A(g1776), .B(g4591), .Z(g5084) ) ;
AND2    gate8010  (.A(g1781), .B(g4592), .Z(g5090) ) ;
AND2    gate8011  (.A(g1786), .B(g4603), .Z(g5097) ) ;
NAND2   gate8012  (.A(II8179), .B(II8180), .Z(g4821) ) ;
AND2    gate8013  (.A(g4821), .B(g3829), .Z(g5099) ) ;
AND2    gate8014  (.A(g1791), .B(g4606), .Z(g5100) ) ;
AND2    gate8015  (.A(g1796), .B(g4608), .Z(g5104) ) ;
AND2    gate8016  (.A(g1801), .B(g4614), .Z(g5108) ) ;
AND2    gate8017  (.A(g1806), .B(g4618), .Z(g5110) ) ;
NOR3    gate8018  (.A(g3419), .B(g3408), .C(g3628), .Z(g4572) ) ;
AND2    gate8019  (.A(g1394), .B(g4572), .Z(g5115) ) ;
AND2    gate8020  (.A(g1618), .B(g4669), .Z(g5123) ) ;
AND2    gate8021  (.A(g4474), .B(g2733), .Z(g5128) ) ;
AND2    gate8022  (.A(g1639), .B(g4673), .Z(g5145) ) ;
AND2    gate8023  (.A(g4478), .B(g2733), .Z(g5151) ) ;
AND2    gate8024  (.A(g1512), .B(g4679), .Z(g5168) ) ;
AND2    gate8025  (.A(g1811), .B(g4680), .Z(g5170) ) ;
AND2    gate8026  (.A(g4555), .B(g4549), .Z(g5172) ) ;
NAND4   gate8027  (.A(g3215), .B(g3247), .C(g2439), .D(g3200), .Z(g4104) ) ;
AND3    gate8028  (.A(g2047), .B(g4401), .C(g4104), .Z(g5178) ) ;
AND2    gate8029  (.A(g4541), .B(g4533), .Z(g5180) ) ;
AND2    gate8030  (.A(g4520), .B(g4510), .Z(g5181) ) ;
AND2    gate8031  (.A(g4504), .B(g4496), .Z(g5188) ) ;
AND2    gate8032  (.A(g1068), .B(g4719), .Z(g5199) ) ;
AND2    gate8033  (.A(g4838), .B(g2126), .Z(g5204) ) ;
AND2    gate8034  (.A(g1080), .B(g4724), .Z(g5211) ) ;
NOR3    gate8035  (.A(g4065), .B(g3261), .C(g2500), .Z(g4276) ) ;
AND2    gate8036  (.A(g4276), .B(g3400), .Z(g5215) ) ;
AND2    gate8037  (.A(g1083), .B(g4729), .Z(g5220) ) ;
AND2    gate8038  (.A(g1086), .B(g4734), .Z(g5228) ) ;
AND2    gate8039  (.A(g1791), .B(g4492), .Z(g5233) ) ;
AND2    gate8040  (.A(g1089), .B(g4747), .Z(g5249) ) ;
AND2    gate8041  (.A(g4335), .B(g4165), .Z(g5254) ) ;
NAND2   gate8042  (.A(II7563), .B(II7564), .Z(g4297) ) ;
AND2    gate8043  (.A(g4297), .B(g2779), .Z(g5256) ) ;
AND2    gate8044  (.A(g627), .B(g4739), .Z(g5259) ) ;
AND2    gate8045  (.A(g1092), .B(g4758), .Z(g5260) ) ;
AND2    gate8046  (.A(g1095), .B(g4763), .Z(g5264) ) ;
AND2    gate8047  (.A(g1098), .B(g4769), .Z(g5268) ) ;
AND2    gate8048  (.A(g1074), .B(g4776), .Z(g5273) ) ;
AND2    gate8049  (.A(g1766), .B(g4783), .Z(g5279) ) ;
AND2    gate8050  (.A(g4593), .B(g3052), .Z(g5280) ) ;
AND2    gate8051  (.A(g4401), .B(g1857), .Z(g5318) ) ;
AND2    gate8052  (.A(g2126), .B(g4617), .Z(g5349) ) ;
AND2    gate8053  (.A(g4610), .B(g2224), .Z(g5398) ) ;
AND2    gate8054  (.A(g1512), .B(g4344), .Z(g5418) ) ;
OR2     gate8055  (.A(g3275), .B(g9), .Z(g3819) ) ;
AND2    gate8056  (.A(g1041), .B(g4880), .Z(g5444) ) ;
OR2     gate8057  (.A(g3275), .B(g12), .Z(g3875) ) ;
AND2    gate8058  (.A(g1044), .B(g4222), .Z(g5470) ) ;
AND2    gate8059  (.A(g4268), .B(g3518), .Z(g5473) ) ;
AND2    gate8060  (.A(g1615), .B(g4237), .Z(g5476) ) ;
AND2    gate8061  (.A(g1845), .B(g4243), .Z(g5479) ) ;
AND2    gate8062  (.A(g4279), .B(g3519), .Z(g5480) ) ;
AND2    gate8063  (.A(g1621), .B(g4254), .Z(g5483) ) ;
AND2    gate8064  (.A(g4287), .B(g3521), .Z(g5489) ) ;
AND2    gate8065  (.A(g1624), .B(g4262), .Z(g5491) ) ;
AND2    gate8066  (.A(g1654), .B(g4263), .Z(g5492) ) ;
AND2    gate8067  (.A(g4296), .B(g3522), .Z(g5497) ) ;
AND2    gate8068  (.A(g1627), .B(g4270), .Z(g5499) ) ;
AND2    gate8069  (.A(g1657), .B(g4272), .Z(g5500) ) ;
AND2    gate8070  (.A(g1672), .B(g4273), .Z(g5501) ) ;
AND2    gate8071  (.A(g4310), .B(g3528), .Z(g5507) ) ;
AND2    gate8072  (.A(g1630), .B(g4280), .Z(g5510) ) ;
AND2    gate8073  (.A(g1660), .B(g4281), .Z(g5512) ) ;
AND2    gate8074  (.A(g1675), .B(g4282), .Z(g5513) ) ;
AND2    gate8075  (.A(g4317), .B(g3532), .Z(g5518) ) ;
AND2    gate8076  (.A(g1633), .B(g4289), .Z(g5522) ) ;
AND2    gate8077  (.A(g1663), .B(g4290), .Z(g5523) ) ;
AND2    gate8078  (.A(g1678), .B(g4291), .Z(g5524) ) ;
AND2    gate8079  (.A(g1721), .B(g4292), .Z(g5525) ) ;
AND2    gate8080  (.A(g4322), .B(g3537), .Z(g5528) ) ;
AND2    gate8081  (.A(g1636), .B(g4305), .Z(g5530) ) ;
AND2    gate8082  (.A(g1666), .B(g4306), .Z(g5531) ) ;
AND2    gate8083  (.A(g1681), .B(g4307), .Z(g5532) ) ;
AND2    gate8084  (.A(g1724), .B(g4308), .Z(g5533) ) ;
AND2    gate8085  (.A(g4327), .B(g3544), .Z(g5535) ) ;
AND2    gate8086  (.A(g4143), .B(g4299), .Z(g5537) ) ;
AND2    gate8087  (.A(g1669), .B(g4313), .Z(g5538) ) ;
AND2    gate8088  (.A(g1684), .B(g4314), .Z(g5539) ) ;
AND2    gate8089  (.A(g1727), .B(g4315), .Z(g5540) ) ;
AND2    gate8090  (.A(g4331), .B(g3582), .Z(g5541) ) ;
AND2    gate8091  (.A(g1687), .B(g4320), .Z(g5544) ) ;
AND2    gate8092  (.A(g1730), .B(g4321), .Z(g5545) ) ;
AND2    gate8093  (.A(g1733), .B(g4326), .Z(g5547) ) ;
AND2    gate8094  (.A(g4816), .B(g2338), .Z(g5569) ) ;
AND2    gate8095  (.A(g1618), .B(g4501), .Z(g5575) ) ;
AND2    gate8096  (.A(g1639), .B(g4508), .Z(g5588) ) ;
AND2    gate8097  (.A(g1615), .B(g4514), .Z(g5591) ) ;
AND2    gate8098  (.A(g1621), .B(g4524), .Z(g5595) ) ;
AND2    gate8099  (.A(g778), .B(g4824), .Z(g5598) ) ;
AND2    gate8100  (.A(g1035), .B(g4375), .Z(g5601) ) ;
AND2    gate8101  (.A(g1624), .B(g4535), .Z(g5602) ) ;
AND2    gate8102  (.A(g4828), .B(g704), .Z(g5605) ) ;
AND2    gate8103  (.A(g814), .B(g4831), .Z(g5608) ) ;
AND2    gate8104  (.A(g1047), .B(g4382), .Z(g5611) ) ;
AND2    gate8105  (.A(g1627), .B(g4543), .Z(g5612) ) ;
AND2    gate8106  (.A(g1050), .B(g4391), .Z(g5617) ) ;
AND2    gate8107  (.A(g1630), .B(g4551), .Z(g5618) ) ;
AND2    gate8108  (.A(g1053), .B(g4399), .Z(g5625) ) ;
AND2    gate8109  (.A(g1633), .B(g4557), .Z(g5626) ) ;
AND2    gate8110  (.A(g1056), .B(g4416), .Z(g5631) ) ;
AND2    gate8111  (.A(g1636), .B(g4563), .Z(g5632) ) ;
AND2    gate8112  (.A(g1059), .B(g4427), .Z(g5640) ) ;
AND2    gate8113  (.A(g148), .B(g5361), .Z(g5674) ) ;
AND2    gate8114  (.A(g131), .B(g5361), .Z(g5675) ) ;
AND2    gate8115  (.A(g153), .B(g5361), .Z(g5680) ) ;
AND2    gate8116  (.A(g135), .B(g5361), .Z(g5681) ) ;
AND2    gate8117  (.A(g158), .B(g5361), .Z(g5686) ) ;
AND2    gate8118  (.A(g139), .B(g5361), .Z(g5687) ) ;
AND2    gate8119  (.A(g1567), .B(g5112), .Z(g5690) ) ;
AND2    gate8120  (.A(g162), .B(g5361), .Z(g5694) ) ;
AND2    gate8121  (.A(g166), .B(g5361), .Z(g5695) ) ;
AND2    gate8122  (.A(g1571), .B(g5116), .Z(g5698) ) ;
AND2    gate8123  (.A(g1592), .B(g5117), .Z(g5699) ) ;
AND2    gate8124  (.A(g174), .B(g5361), .Z(g5703) ) ;
AND2    gate8125  (.A(g143), .B(g5361), .Z(g5704) ) ;
AND2    gate8126  (.A(g1574), .B(g5121), .Z(g5706) ) ;
AND2    gate8127  (.A(g1595), .B(g5122), .Z(g5707) ) ;
AND2    gate8128  (.A(g170), .B(g5361), .Z(g5720) ) ;
AND2    gate8129  (.A(g1577), .B(g5143), .Z(g5721) ) ;
AND2    gate8130  (.A(g1598), .B(g5144), .Z(g5722) ) ;
AND2    gate8131  (.A(g1580), .B(g5166), .Z(g5725) ) ;
AND2    gate8132  (.A(g1601), .B(g5167), .Z(g5726) ) ;
AND2    gate8133  (.A(g1583), .B(g5175), .Z(g5731) ) ;
AND2    gate8134  (.A(g1604), .B(g5176), .Z(g5732) ) ;
AND2    gate8135  (.A(g1524), .B(g5183), .Z(g5737) ) ;
AND2    gate8136  (.A(g1586), .B(g5184), .Z(g5738) ) ;
AND2    gate8137  (.A(g1607), .B(g5185), .Z(g5739) ) ;
AND2    gate8138  (.A(g1528), .B(g5191), .Z(g5744) ) ;
AND2    gate8139  (.A(g1549), .B(g5192), .Z(g5745) ) ;
AND2    gate8140  (.A(g1589), .B(g5193), .Z(g5746) ) ;
NAND2   gate8141  (.A(II8480), .B(II8481), .Z(g5103) ) ;
AND2    gate8142  (.A(g1531), .B(g5202), .Z(g5756) ) ;
AND2    gate8143  (.A(g1552), .B(g5203), .Z(g5757) ) ;
NAND4   gate8144  (.A(g3056), .B(g3071), .C(g2310), .D(g3003), .Z(g3818) ) ;
AND3    gate8145  (.A(g2112), .B(g4921), .C(g3818), .Z(g5769) ) ;
AND2    gate8146  (.A(g1534), .B(g5213), .Z(g5771) ) ;
AND2    gate8147  (.A(g1555), .B(g5214), .Z(g5772) ) ;
AND2    gate8148  (.A(g1537), .B(g5222), .Z(g5781) ) ;
AND2    gate8149  (.A(g1558), .B(g5223), .Z(g5782) ) ;
AND2    gate8150  (.A(g1540), .B(g5231), .Z(g5788) ) ;
AND2    gate8151  (.A(g1561), .B(g5232), .Z(g5789) ) ;
AND2    gate8152  (.A(g1543), .B(g5251), .Z(g5795) ) ;
AND2    gate8153  (.A(g1564), .B(g5252), .Z(g5796) ) ;
AND2    gate8154  (.A(g1546), .B(g5261), .Z(g5804) ) ;
NAND2   gate8155  (.A(g2571), .B(g2061), .Z(g3204) ) ;
AND2    gate8156  (.A(g3204), .B(g5318), .Z(g5825) ) ;
OR2     gate8157  (.A(g3107), .B(g2167), .Z(g3860) ) ;
AND2    gate8158  (.A(g3860), .B(g5519), .Z(g5848) ) ;
AND2    gate8159  (.A(g5044), .B(g1927), .Z(g5853) ) ;
AND2    gate8160  (.A(g4921), .B(g639), .Z(g5877) ) ;
NAND2   gate8161  (.A(II9007), .B(II9008), .Z(g5592) ) ;
AND2    gate8162  (.A(g5592), .B(g3829), .Z(g5882) ) ;
OR2     gate8163  (.A(g1393), .B(g1394), .Z(g2204) ) ;
AND2    gate8164  (.A(g2204), .B(g5354), .Z(g5897) ) ;
NAND2   gate8165  (.A(II5676), .B(II5677), .Z(g2555) ) ;
AND2    gate8166  (.A(g2555), .B(g4977), .Z(g5902) ) ;
NAND2   gate8167  (.A(II6488), .B(II6489), .Z(g3322) ) ;
AND2    gate8168  (.A(g3322), .B(g4977), .Z(g5911) ) ;
AND2    gate8169  (.A(g1041), .B(g5320), .Z(g5913) ) ;
NAND2   gate8170  (.A(II7322), .B(II7323), .Z(g4168) ) ;
AND2    gate8171  (.A(g4168), .B(g4977), .Z(g5915) ) ;
AND2    gate8172  (.A(g1044), .B(g5320), .Z(g5917) ) ;
OR2     gate8173  (.A(g3400), .B(g119), .Z(g4609) ) ;
AND2    gate8174  (.A(g5216), .B(g2965), .Z(g5919) ) ;
AND2    gate8175  (.A(g5215), .B(g1965), .Z(g5934) ) ;
AND2    gate8176  (.A(g1796), .B(g5233), .Z(g5944) ) ;
AND2    gate8177  (.A(g2017), .B(g4977), .Z(g6047) ) ;
AND2    gate8178  (.A(g1035), .B(g5320), .Z(g6058) ) ;
AND2    gate8179  (.A(g5398), .B(g2230), .Z(g6064) ) ;
AND2    gate8180  (.A(g1047), .B(g5320), .Z(g6067) ) ;
AND2    gate8181  (.A(g1050), .B(g5320), .Z(g6070) ) ;
AND2    gate8182  (.A(g549), .B(g5613), .Z(g6075) ) ;
AND2    gate8183  (.A(g1053), .B(g5320), .Z(g6079) ) ;
AND2    gate8184  (.A(g552), .B(g5619), .Z(g6083) ) ;
AND2    gate8185  (.A(g1056), .B(g5320), .Z(g6087) ) ;
AND2    gate8186  (.A(g553), .B(g5627), .Z(g6090) ) ;
AND2    gate8187  (.A(g1059), .B(g5320), .Z(g6092) ) ;
AND2    gate8188  (.A(g1062), .B(g5320), .Z(g6095) ) ;
AND2    gate8189  (.A(g1065), .B(g5320), .Z(g6098) ) ;
AND2    gate8190  (.A(g1038), .B(g5320), .Z(g6102) ) ;
OR2     gate8191  (.A(g2863), .B(g2516), .Z(g3584) ) ;
AND2    gate8192  (.A(g3584), .B(g5200), .Z(g6162) ) ;
AND2    gate8193  (.A(g546), .B(g5042), .Z(g6186) ) ;
AND2    gate8194  (.A(g5569), .B(g2340), .Z(g6187) ) ;
AND2    gate8195  (.A(g554), .B(g5043), .Z(g6194) ) ;
AND2    gate8196  (.A(g557), .B(g5062), .Z(g6199) ) ;
AND2    gate8197  (.A(g3738), .B(g4921), .Z(g6204) ) ;
AND2    gate8198  (.A(g560), .B(g5068), .Z(g6206) ) ;
AND2    gate8199  (.A(g563), .B(g5073), .Z(g6217) ) ;
AND2    gate8200  (.A(g782), .B(g5598), .Z(g6221) ) ;
AND2    gate8201  (.A(g566), .B(g5082), .Z(g6225) ) ;
AND2    gate8202  (.A(g5605), .B(g713), .Z(g6228) ) ;
AND2    gate8203  (.A(g818), .B(g5608), .Z(g6231) ) ;
AND2    gate8204  (.A(g569), .B(g5089), .Z(g6235) ) ;
AND2    gate8205  (.A(g572), .B(g5096), .Z(g6238) ) ;
AND2    gate8206  (.A(g182), .B(g5361), .Z(g6240) ) ;
AND2    gate8207  (.A(g575), .B(g5098), .Z(g6245) ) ;
AND2    gate8208  (.A(g178), .B(g5361), .Z(g6246) ) ;
AND2    gate8209  (.A(g127), .B(g5361), .Z(g6247) ) ;
AND2    gate8210  (.A(g1270), .B(g5949), .Z(g6316) ) ;
AND2    gate8211  (.A(g1304), .B(g5949), .Z(g6317) ) ;
AND2    gate8212  (.A(g1300), .B(g5949), .Z(g6318) ) ;
AND2    gate8213  (.A(g1296), .B(g5949), .Z(g6319) ) ;
AND2    gate8214  (.A(g1292), .B(g5949), .Z(g6320) ) ;
AND2    gate8215  (.A(g1284), .B(g5949), .Z(g6321) ) ;
AND2    gate8216  (.A(g1275), .B(g5949), .Z(g6322) ) ;
AND2    gate8217  (.A(g1235), .B(g5949), .Z(g6323) ) ;
AND2    gate8218  (.A(g1240), .B(g5949), .Z(g6324) ) ;
AND2    gate8219  (.A(g1245), .B(g5949), .Z(g6325) ) ;
AND2    gate8220  (.A(g1250), .B(g5949), .Z(g6326) ) ;
AND2    gate8221  (.A(g1255), .B(g5949), .Z(g6327) ) ;
AND2    gate8222  (.A(g1260), .B(g5949), .Z(g6328) ) ;
AND2    gate8223  (.A(g1265), .B(g5949), .Z(g6329) ) ;
AND2    gate8224  (.A(g272), .B(g5885), .Z(g6341) ) ;
AND2    gate8225  (.A(g293), .B(g5886), .Z(g6342) ) ;
OR2     gate8226  (.A(g5631), .B(g4882), .Z(g5823) ) ;
AND2    gate8227  (.A(g5823), .B(g4426), .Z(g6345) ) ;
OR2     gate8228  (.A(g4878), .B(g4884), .Z(g5038) ) ;
AND2    gate8229  (.A(g5038), .B(g5883), .Z(g6346) ) ;
AND2    gate8230  (.A(g275), .B(g5890), .Z(g6347) ) ;
AND2    gate8231  (.A(g296), .B(g5891), .Z(g6348) ) ;
OR2     gate8232  (.A(g5640), .B(g4224), .Z(g5837) ) ;
AND2    gate8233  (.A(g5837), .B(g4435), .Z(g6350) ) ;
AND2    gate8234  (.A(g278), .B(g5894), .Z(g6352) ) ;
AND2    gate8235  (.A(g299), .B(g5895), .Z(g6353) ) ;
OR2     gate8236  (.A(g4914), .B(g4230), .Z(g5841) ) ;
AND2    gate8237  (.A(g5841), .B(g4441), .Z(g6358) ) ;
AND2    gate8238  (.A(g281), .B(g5898), .Z(g6359) ) ;
AND2    gate8239  (.A(g302), .B(g5899), .Z(g6360) ) ;
OR2     gate8240  (.A(g4932), .B(g4236), .Z(g5846) ) ;
AND2    gate8241  (.A(g5846), .B(g4450), .Z(g6362) ) ;
AND2    gate8242  (.A(g284), .B(g5901), .Z(g6363) ) ;
OR2     gate8243  (.A(g4941), .B(g4253), .Z(g5851) ) ;
AND2    gate8244  (.A(g5851), .B(g4454), .Z(g6364) ) ;
AND2    gate8245  (.A(g2132), .B(g5748), .Z(g6404) ) ;
AND2    gate8246  (.A(g2804), .B(g5759), .Z(g6410) ) ;
AND2    gate8247  (.A(g3497), .B(g5774), .Z(g6416) ) ;
AND2    gate8248  (.A(g4348), .B(g5784), .Z(g6423) ) ;
AND2    gate8249  (.A(g5044), .B(g5791), .Z(g6430) ) ;
AND2    gate8250  (.A(g5853), .B(g5797), .Z(g6438) ) ;
AND2    gate8251  (.A(g5052), .B(g6210), .Z(g6463) ) ;
OR2     gate8252  (.A(g4360), .B(g3512), .Z(g5224) ) ;
AND2    gate8253  (.A(g5853), .B(g1936), .Z(g6472) ) ;
OR2     gate8254  (.A(g5074), .B(g4383), .Z(g5981) ) ;
OR2     gate8255  (.A(g5084), .B(g4392), .Z(g5983) ) ;
OR2     gate8256  (.A(g5090), .B(g4400), .Z(g5993) ) ;
OR2     gate8257  (.A(g5097), .B(g5099), .Z(g5995) ) ;
NAND2   gate8258  (.A(II9947), .B(II9948), .Z(g6207) ) ;
AND2    gate8259  (.A(g6207), .B(g3829), .Z(g6530) ) ;
AND2    gate8260  (.A(g339), .B(g6057), .Z(g6532) ) ;
AND2    gate8261  (.A(g345), .B(g6063), .Z(g6535) ) ;
AND2    gate8262  (.A(g1223), .B(g6072), .Z(g6540) ) ;
AND2    gate8263  (.A(g1227), .B(g6081), .Z(g6544) ) ;
AND2    gate8264  (.A(g5515), .B(g6175), .Z(g6549) ) ;
AND2    gate8265  (.A(g1231), .B(g6089), .Z(g6550) ) ;
AND2    gate8266  (.A(g5075), .B(g6183), .Z(g6554) ) ;
OR2     gate8267  (.A(g5178), .B(g5186), .Z(g5762) ) ;
AND2    gate8268  (.A(g5762), .B(g5503), .Z(g6576) ) ;
AND2    gate8269  (.A(g1801), .B(g5944), .Z(g6580) ) ;
OR2     gate8270  (.A(g5279), .B(g4559), .Z(g6105) ) ;
AND2    gate8271  (.A(g6105), .B(g3246), .Z(g6616) ) ;
AND2    gate8272  (.A(g658), .B(g6016), .Z(g6618) ) ;
AND2    gate8273  (.A(g49), .B(g6156), .Z(g6619) ) ;
AND2    gate8274  (.A(g336), .B(g6165), .Z(g6622) ) ;
AND2    gate8275  (.A(g55), .B(g6170), .Z(g6623) ) ;
AND2    gate8276  (.A(g348), .B(g6171), .Z(g6624) ) ;
AND2    gate8277  (.A(g1218), .B(g6178), .Z(g6625) ) ;
AND2    gate8278  (.A(g351), .B(g6182), .Z(g6628) ) ;
AND2    gate8279  (.A(g61), .B(g6190), .Z(g6632) ) ;
AND2    gate8280  (.A(g354), .B(g6191), .Z(g6633) ) ;
AND2    gate8281  (.A(g357), .B(g6196), .Z(g6639) ) ;
AND2    gate8282  (.A(g5281), .B(g5801), .Z(g6640) ) ;
AND2    gate8283  (.A(g67), .B(g6202), .Z(g6645) ) ;
AND2    gate8284  (.A(g360), .B(g6203), .Z(g6646) ) ;
AND2    gate8285  (.A(g5288), .B(g5808), .Z(g6647) ) ;
AND2    gate8286  (.A(g363), .B(g6214), .Z(g6654) ) ;
AND2    gate8287  (.A(g5296), .B(g5812), .Z(g6655) ) ;
OR2     gate8288  (.A(g5204), .B(g4), .Z(g6061) ) ;
AND2    gate8289  (.A(g73), .B(g6219), .Z(g6661) ) ;
AND2    gate8290  (.A(g366), .B(g6220), .Z(g6662) ) ;
AND2    gate8291  (.A(g6064), .B(g2237), .Z(g6663) ) ;
AND2    gate8292  (.A(g5301), .B(g5818), .Z(g6666) ) ;
AND2    gate8293  (.A(g342), .B(g6227), .Z(g6671) ) ;
AND2    gate8294  (.A(g5305), .B(g5822), .Z(g6673) ) ;
OR2     gate8295  (.A(g5349), .B(g1), .Z(g6074) ) ;
AND2    gate8296  (.A(g5314), .B(g5836), .Z(g6684) ) ;
AND2    gate8297  (.A(g5486), .B(g5840), .Z(g6687) ) ;
AND2    gate8298  (.A(g5494), .B(g5845), .Z(g6693) ) ;
AND2    gate8299  (.A(g5504), .B(g5850), .Z(g6696) ) ;
OR2     gate8300  (.A(g5444), .B(g4712), .Z(g6177) ) ;
AND2    gate8301  (.A(g6177), .B(g4221), .Z(g6699) ) ;
OR2     gate8302  (.A(g5470), .B(g4715), .Z(g6185) ) ;
AND2    gate8303  (.A(g6185), .B(g4228), .Z(g6701) ) ;
AND2    gate8304  (.A(g1872), .B(g6128), .Z(g6730) ) ;
AND2    gate8305  (.A(g2531), .B(g6137), .Z(g6738) ) ;
AND2    gate8306  (.A(g3284), .B(g6141), .Z(g6741) ) ;
AND2    gate8307  (.A(g4106), .B(g6146), .Z(g6743) ) ;
AND2    gate8308  (.A(g4828), .B(g6151), .Z(g6744) ) ;
AND2    gate8309  (.A(g5605), .B(g6158), .Z(g6745) ) ;
AND2    gate8310  (.A(g6228), .B(g6166), .Z(g6746) ) ;
AND2    gate8311  (.A(g6187), .B(g2343), .Z(g6752) ) ;
NAND2   gate8312  (.A(g2382), .B(g2399), .Z(g3010) ) ;
AND2    gate8313  (.A(g3010), .B(g5877), .Z(g6756) ) ;
AND2    gate8314  (.A(g786), .B(g6221), .Z(g6760) ) ;
OR2     gate8315  (.A(g5601), .B(g4837), .Z(g5802) ) ;
AND2    gate8316  (.A(g5802), .B(g4381), .Z(g6763) ) ;
AND2    gate8317  (.A(g263), .B(g5866), .Z(g6771) ) ;
AND2    gate8318  (.A(g6228), .B(g722), .Z(g6772) ) ;
AND2    gate8319  (.A(g822), .B(g6231), .Z(g6775) ) ;
OR2     gate8320  (.A(g5611), .B(g4865), .Z(g5809) ) ;
AND2    gate8321  (.A(g5809), .B(g4390), .Z(g6776) ) ;
AND2    gate8322  (.A(g266), .B(g5875), .Z(g6787) ) ;
AND2    gate8323  (.A(g287), .B(g5876), .Z(g6788) ) ;
OR2     gate8324  (.A(g5617), .B(g4869), .Z(g5813) ) ;
AND2    gate8325  (.A(g5813), .B(g4398), .Z(g6790) ) ;
AND2    gate8326  (.A(g269), .B(g5880), .Z(g6791) ) ;
AND2    gate8327  (.A(g290), .B(g5881), .Z(g6792) ) ;
OR2     gate8328  (.A(g5625), .B(g4876), .Z(g5819) ) ;
AND2    gate8329  (.A(g5819), .B(g4415), .Z(g6794) ) ;
OR2     gate8330  (.A(g4871), .B(g4162), .Z(g5036) ) ;
AND2    gate8331  (.A(g1964), .B(g6392), .Z(g6855) ) ;
AND2    gate8332  (.A(g1896), .B(g6389), .Z(g6872) ) ;
AND2    gate8333  (.A(g3263), .B(g6557), .Z(g6873) ) ;
AND2    gate8334  (.A(g1905), .B(g6400), .Z(g6875) ) ;
AND2    gate8335  (.A(g4070), .B(g6560), .Z(g6876) ) ;
AND2    gate8336  (.A(g1914), .B(g6407), .Z(g6879) ) ;
AND2    gate8337  (.A(g4816), .B(g6562), .Z(g6880) ) ;
AND2    gate8338  (.A(g1923), .B(g6413), .Z(g6883) ) ;
AND2    gate8339  (.A(g5569), .B(g6564), .Z(g6884) ) ;
AND2    gate8340  (.A(g1932), .B(g6420), .Z(g6886) ) ;
AND2    gate8341  (.A(g6187), .B(g6566), .Z(g6887) ) ;
AND2    gate8342  (.A(g1941), .B(g6427), .Z(g6889) ) ;
AND2    gate8343  (.A(g6752), .B(g6568), .Z(g6890) ) ;
AND2    gate8344  (.A(g1950), .B(g6435), .Z(g6891) ) ;
AND2    gate8345  (.A(g6472), .B(g5805), .Z(g6892) ) ;
AND2    gate8346  (.A(g6472), .B(g1945), .Z(g6940) ) ;
OR2     gate8347  (.A(g5100), .B(g5882), .Z(g6592) ) ;
NAND2   gate8348  (.A(II10770), .B(II10771), .Z(g6758) ) ;
AND2    gate8349  (.A(g6758), .B(g3829), .Z(g6994) ) ;
OR2     gate8350  (.A(g5934), .B(g123), .Z(g6626) ) ;
AND2    gate8351  (.A(g5892), .B(g6570), .Z(g7046) ) ;
AND2    gate8352  (.A(g5896), .B(g6575), .Z(g7050) ) ;
AND2    gate8353  (.A(g5900), .B(g6579), .Z(g7055) ) ;
OR2     gate8354  (.A(g4503), .B(g5256), .Z(g6078) ) ;
AND2    gate8355  (.A(g6078), .B(g6714), .Z(g7059) ) ;
OR2     gate8356  (.A(g5769), .B(g5780), .Z(g6739) ) ;
AND2    gate8357  (.A(g6739), .B(g5521), .Z(g7060) ) ;
AND2    gate8358  (.A(g790), .B(g6760), .Z(g7061) ) ;
AND2    gate8359  (.A(g5903), .B(g6582), .Z(g7063) ) ;
AND2    gate8360  (.A(g5912), .B(g6586), .Z(g7068) ) ;
AND2    gate8361  (.A(g5916), .B(g6590), .Z(g7071) ) ;
AND2    gate8362  (.A(g2331), .B(g6737), .Z(g7088) ) ;
AND2    gate8363  (.A(g1212), .B(g6648), .Z(g7125) ) ;
AND2    gate8364  (.A(g6663), .B(g2241), .Z(g7127) ) ;
AND2    gate8365  (.A(g6041), .B(g6697), .Z(g7130) ) ;
AND2    gate8366  (.A(g6044), .B(g6700), .Z(g7131) ) ;
AND2    gate8367  (.A(g6048), .B(g6702), .Z(g7132) ) ;
OR2     gate8368  (.A(g4714), .B(g3904), .Z(g5587) ) ;
NOR2    gate8369  (.A(g6032), .B(g6023), .Z(g6355) ) ;
AND2    gate8370  (.A(g869), .B(g6355), .Z(g7135) ) ;
AND2    gate8371  (.A(g6050), .B(g6704), .Z(g7136) ) ;
OR2     gate8372  (.A(g4718), .B(g4723), .Z(g5590) ) ;
AND2    gate8373  (.A(g6055), .B(g6707), .Z(g7138) ) ;
AND2    gate8374  (.A(g6060), .B(g6709), .Z(g7139) ) ;
AND2    gate8375  (.A(g6069), .B(g6711), .Z(g7140) ) ;
AND2    gate8376  (.A(g6073), .B(g6716), .Z(g7141) ) ;
AND2    gate8377  (.A(g6082), .B(g6718), .Z(g7145) ) ;
AND2    gate8378  (.A(g1878), .B(g6720), .Z(g7182) ) ;
AND2    gate8379  (.A(g1887), .B(g6724), .Z(g7185) ) ;
AND2    gate8380  (.A(g2503), .B(g6403), .Z(g7186) ) ;
AND2    gate8381  (.A(g3098), .B(g6418), .Z(g7200) ) ;
AND2    gate8382  (.A(g3804), .B(g6425), .Z(g7209) ) ;
AND2    gate8383  (.A(g4610), .B(g6432), .Z(g7217) ) ;
AND2    gate8384  (.A(g5398), .B(g6441), .Z(g7224) ) ;
AND2    gate8385  (.A(g6064), .B(g6444), .Z(g7230) ) ;
AND2    gate8386  (.A(g6663), .B(g6447), .Z(g7235) ) ;
AND2    gate8387  (.A(g6772), .B(g6172), .Z(g7241) ) ;
AND2    gate8388  (.A(g6752), .B(g2345), .Z(g7260) ) ;
OR2     gate8389  (.A(g4836), .B(g4128), .Z(g5028) ) ;
AND2    gate8390  (.A(g5028), .B(g6499), .Z(g7271) ) ;
AND2    gate8391  (.A(g6772), .B(g731), .Z(g7277) ) ;
AND2    gate8392  (.A(g6980), .B(g3880), .Z(g7368) ) ;
AND2    gate8393  (.A(g6990), .B(g3880), .Z(g7378) ) ;
AND2    gate8394  (.A(g7001), .B(g3880), .Z(g7389) ) ;
NAND3   gate8395  (.A(g2310), .B(g4604), .C(g3807), .Z(g4976) ) ;
NAND2   gate8396  (.A(II10931), .B(II10932), .Z(g6858) ) ;
AND3    gate8397  (.A(g4976), .B(g632), .C(g6858), .Z(g7409) ) ;
AND2    gate8398  (.A(g7260), .B(g6572), .Z(g7435) ) ;
AND2    gate8399  (.A(g7277), .B(g5827), .Z(g7444) ) ;
AND2    gate8400  (.A(g6868), .B(g4355), .Z(g7449) ) ;
AND2    gate8401  (.A(g7148), .B(g2809), .Z(g7453) ) ;
AND2    gate8402  (.A(g7148), .B(g2814), .Z(g7459) ) ;
AND2    gate8403  (.A(g7148), .B(g2821), .Z(g7466) ) ;
AND2    gate8404  (.A(g7148), .B(g2829), .Z(g7472) ) ;
AND2    gate8405  (.A(g7148), .B(g2840), .Z(g7496) ) ;
AND2    gate8406  (.A(g7148), .B(g2847), .Z(g7504) ) ;
AND2    gate8407  (.A(g7148), .B(g2855), .Z(g7515) ) ;
AND2    gate8408  (.A(g7148), .B(g2868), .Z(g7526) ) ;
AND2    gate8409  (.A(g7148), .B(g2874), .Z(g7535) ) ;
AND2    gate8410  (.A(g7148), .B(g2877), .Z(g7536) ) ;
OR2     gate8411  (.A(g5104), .B(g6530), .Z(g7075) ) ;
AND2    gate8412  (.A(g7148), .B(g2885), .Z(g7542) ) ;
NAND2   gate8413  (.A(II11509), .B(II11510), .Z(g7269) ) ;
AND2    gate8414  (.A(g7269), .B(g3829), .Z(g7549) ) ;
OR2     gate8415  (.A(g6540), .B(g5902), .Z(g7092) ) ;
OR2     gate8416  (.A(g6544), .B(g5911), .Z(g7096) ) ;
OR2     gate8417  (.A(g6550), .B(g5915), .Z(g7102) ) ;
AND2    gate8418  (.A(g6940), .B(g5984), .Z(g7613) ) ;
AND2    gate8419  (.A(g664), .B(g7079), .Z(g7623) ) ;
AND2    gate8420  (.A(g673), .B(g7085), .Z(g7625) ) ;
OR2     gate8421  (.A(g6625), .B(g6047), .Z(g7184) ) ;
AND2    gate8422  (.A(g7127), .B(g2251), .Z(g7661) ) ;
AND2    gate8423  (.A(g7004), .B(g3880), .Z(g7674) ) ;
AND2    gate8424  (.A(g1950), .B(g6863), .Z(g7679) ) ;
AND2    gate8425  (.A(g682), .B(g7197), .Z(g7704) ) ;
AND2    gate8426  (.A(g691), .B(g7206), .Z(g7707) ) ;
AND2    gate8427  (.A(g700), .B(g7214), .Z(g7710) ) ;
AND2    gate8428  (.A(g709), .B(g7221), .Z(g7718) ) ;
AND2    gate8429  (.A(g718), .B(g7227), .Z(g7719) ) ;
AND2    gate8430  (.A(g727), .B(g7232), .Z(g7720) ) ;
AND2    gate8431  (.A(g736), .B(g7237), .Z(g7721) ) ;
AND2    gate8432  (.A(g7127), .B(g6449), .Z(g7722) ) ;
AND2    gate8433  (.A(g7260), .B(g2347), .Z(g7730) ) ;
AND2    gate8434  (.A(g6935), .B(g3880), .Z(g7732) ) ;
AND2    gate8435  (.A(g6944), .B(g3880), .Z(g7734) ) ;
AND2    gate8436  (.A(g6951), .B(g3880), .Z(g7736) ) ;
AND2    gate8437  (.A(g6957), .B(g3880), .Z(g7739) ) ;
AND2    gate8438  (.A(g6961), .B(g3880), .Z(g7741) ) ;
AND2    gate8439  (.A(g6967), .B(g3880), .Z(g7743) ) ;
AND2    gate8440  (.A(g1878), .B(g7479), .Z(g7818) ) ;
AND2    gate8441  (.A(g1887), .B(g7479), .Z(g7819) ) ;
AND2    gate8442  (.A(g1896), .B(g7479), .Z(g7820) ) ;
AND2    gate8443  (.A(g1905), .B(g7479), .Z(g7821) ) ;
AND2    gate8444  (.A(g1914), .B(g7479), .Z(g7822) ) ;
AND2    gate8445  (.A(g1923), .B(g7479), .Z(g7823) ) ;
AND2    gate8446  (.A(g1932), .B(g7479), .Z(g7824) ) ;
AND2    gate8447  (.A(g1941), .B(g7479), .Z(g7825) ) ;
NAND2   gate8448  (.A(II12144), .B(II12145), .Z(g7599) ) ;
AND2    gate8449  (.A(g7609), .B(g3790), .Z(g7876) ) ;
AND2    gate8450  (.A(g7610), .B(g3798), .Z(g7879) ) ;
AND2    gate8451  (.A(g7612), .B(g3810), .Z(g7881) ) ;
OR2     gate8452  (.A(g6873), .B(g6404), .Z(g7457) ) ;
AND2    gate8453  (.A(g7457), .B(g7022), .Z(g7884) ) ;
AND2    gate8454  (.A(g7614), .B(g3812), .Z(g7885) ) ;
OR2     gate8455  (.A(g6876), .B(g6410), .Z(g7465) ) ;
AND2    gate8456  (.A(g7465), .B(g7025), .Z(g7888) ) ;
AND2    gate8457  (.A(g7615), .B(g3814), .Z(g7889) ) ;
OR2     gate8458  (.A(g6880), .B(g6416), .Z(g7471) ) ;
AND2    gate8459  (.A(g7471), .B(g7028), .Z(g7891) ) ;
AND2    gate8460  (.A(g7616), .B(g3815), .Z(g7892) ) ;
OR2     gate8461  (.A(g6884), .B(g6423), .Z(g7478) ) ;
AND2    gate8462  (.A(g7478), .B(g7031), .Z(g7893) ) ;
AND2    gate8463  (.A(g7617), .B(g3816), .Z(g7894) ) ;
OR2     gate8464  (.A(g6887), .B(g6430), .Z(g7503) ) ;
AND2    gate8465  (.A(g7503), .B(g7036), .Z(g7895) ) ;
OR2     gate8466  (.A(g6890), .B(g6438), .Z(g7511) ) ;
AND2    gate8467  (.A(g7511), .B(g7041), .Z(g7898) ) ;
AND2    gate8468  (.A(g7661), .B(g6587), .Z(g7902) ) ;
OR2     gate8469  (.A(g5108), .B(g6994), .Z(g7621) ) ;
AND2    gate8470  (.A(g2809), .B(g7446), .Z(g7931) ) ;
AND2    gate8471  (.A(g2814), .B(g7450), .Z(g7933) ) ;
AND2    gate8472  (.A(g2821), .B(g7454), .Z(g7935) ) ;
AND2    gate8473  (.A(g7606), .B(g4013), .Z(g7937) ) ;
AND2    gate8474  (.A(g2829), .B(g7460), .Z(g7939) ) ;
AND2    gate8475  (.A(g7620), .B(g4013), .Z(g7940) ) ;
AND2    gate8476  (.A(g2840), .B(g7467), .Z(g7943) ) ;
AND2    gate8477  (.A(g2847), .B(g7473), .Z(g7945) ) ;
AND2    gate8478  (.A(g2855), .B(g7497), .Z(g7948) ) ;
AND2    gate8479  (.A(g2868), .B(g7505), .Z(g7951) ) ;
AND2    gate8480  (.A(g2874), .B(g7512), .Z(g7954) ) ;
AND2    gate8481  (.A(g2877), .B(g7516), .Z(g7955) ) ;
AND2    gate8482  (.A(g2885), .B(g7527), .Z(g7957) ) ;
AND2    gate8483  (.A(g736), .B(g7697), .Z(g7958) ) ;
AND2    gate8484  (.A(g7730), .B(g6712), .Z(g7962) ) ;
OR2     gate8485  (.A(g7088), .B(g6618), .Z(g7384) ) ;
AND2    gate8486  (.A(g7384), .B(g7703), .Z(g7970) ) ;
AND2    gate8487  (.A(g1878), .B(g7379), .Z(g7988) ) ;
OR2     gate8488  (.A(g7186), .B(g6730), .Z(g7510) ) ;
AND2    gate8489  (.A(g7510), .B(g6871), .Z(g8005) ) ;
OR2     gate8490  (.A(g7200), .B(g6738), .Z(g7738) ) ;
AND2    gate8491  (.A(g7738), .B(g7413), .Z(g8010) ) ;
OR2     gate8492  (.A(g7209), .B(g6741), .Z(g7740) ) ;
AND2    gate8493  (.A(g7740), .B(g7419), .Z(g8014) ) ;
OR2     gate8494  (.A(g7217), .B(g6743), .Z(g7742) ) ;
AND2    gate8495  (.A(g7742), .B(g7425), .Z(g8018) ) ;
OR2     gate8496  (.A(g7224), .B(g6744), .Z(g7367) ) ;
AND2    gate8497  (.A(g7367), .B(g7430), .Z(g8023) ) ;
OR2     gate8498  (.A(g7230), .B(g6745), .Z(g7375) ) ;
AND2    gate8499  (.A(g7375), .B(g7436), .Z(g8028) ) ;
OR2     gate8500  (.A(g7235), .B(g6746), .Z(g7385) ) ;
AND2    gate8501  (.A(g7385), .B(g7438), .Z(g8032) ) ;
NAND2   gate8502  (.A(II12086), .B(II12087), .Z(g7587) ) ;
NAND2   gate8503  (.A(II11908), .B(II11909), .Z(g7523) ) ;
NAND2   gate8504  (.A(II11915), .B(II11916), .Z(g7524) ) ;
NAND2   gate8505  (.A(II11936), .B(II11937), .Z(g7533) ) ;
NAND2   gate8506  (.A(II12061), .B(II12062), .Z(g7582) ) ;
NAND2   gate8507  (.A(II12137), .B(II12138), .Z(g7598) ) ;
NAND2   gate8508  (.A(II11974), .B(II11975), .Z(g7547) ) ;
NAND2   gate8509  (.A(II11981), .B(II11982), .Z(g7548) ) ;
NAND2   gate8510  (.A(II11996), .B(II11997), .Z(g7557) ) ;
NAND2   gate8511  (.A(II12003), .B(II12004), .Z(g7558) ) ;
NAND2   gate8512  (.A(II12020), .B(II12021), .Z(g7567) ) ;
NAND2   gate8513  (.A(II12127), .B(II12128), .Z(g7596) ) ;
NAND2   gate8514  (.A(II12039), .B(II12040), .Z(g7572) ) ;
NAND2   gate8515  (.A(II12046), .B(II12047), .Z(g7573) ) ;
NAND2   gate8516  (.A(II12068), .B(II12069), .Z(g7583) ) ;
NAND2   gate8517  (.A(II12075), .B(II12076), .Z(g7584) ) ;
NAND2   gate8518  (.A(II12093), .B(II12094), .Z(g7588) ) ;
NAND2   gate8519  (.A(II12107), .B(II12108), .Z(g7592) ) ;
NAND2   gate8520  (.A(II12114), .B(II12115), .Z(g7593) ) ;
AND2    gate8521  (.A(g664), .B(g7826), .Z(g8068) ) ;
AND2    gate8522  (.A(g673), .B(g7826), .Z(g8069) ) ;
AND2    gate8523  (.A(g682), .B(g7826), .Z(g8070) ) ;
AND2    gate8524  (.A(g691), .B(g7826), .Z(g8071) ) ;
AND2    gate8525  (.A(g700), .B(g7826), .Z(g8072) ) ;
AND2    gate8526  (.A(g709), .B(g7826), .Z(g8073) ) ;
AND2    gate8527  (.A(g718), .B(g7826), .Z(g8074) ) ;
AND2    gate8528  (.A(g727), .B(g7826), .Z(g8075) ) ;
AND2    gate8529  (.A(g6200), .B(g7851), .Z(g8097) ) ;
AND2    gate8530  (.A(g6201), .B(g7852), .Z(g8098) ) ;
AND2    gate8531  (.A(g6208), .B(g7877), .Z(g8101) ) ;
AND2    gate8532  (.A(g6209), .B(g7878), .Z(g8102) ) ;
AND2    gate8533  (.A(g6218), .B(g7880), .Z(g8104) ) ;
AND2    gate8534  (.A(g6226), .B(g7882), .Z(g8107) ) ;
AND2    gate8535  (.A(g1891), .B(g7938), .Z(g8108) ) ;
AND2    gate8536  (.A(g6236), .B(g7886), .Z(g8117) ) ;
AND2    gate8537  (.A(g1900), .B(g7941), .Z(g8118) ) ;
AND2    gate8538  (.A(g6239), .B(g7890), .Z(g8119) ) ;
AND2    gate8539  (.A(g1909), .B(g7944), .Z(g8120) ) ;
AND2    gate8540  (.A(g1918), .B(g7946), .Z(g8123) ) ;
AND2    gate8541  (.A(g1927), .B(g7949), .Z(g8127) ) ;
AND2    gate8542  (.A(g1936), .B(g7952), .Z(g8130) ) ;
AND2    gate8543  (.A(g1945), .B(g7956), .Z(g8135) ) ;
OR2     gate8544  (.A(g7435), .B(g6892), .Z(g7926) ) ;
AND2    gate8545  (.A(g7926), .B(g7045), .Z(g8136) ) ;
NAND2   gate8546  (.A(g7409), .B(g5573), .Z(g7960) ) ;
AND2    gate8547  (.A(g7960), .B(g3737), .Z(g8163) ) ;
AND2    gate8548  (.A(g5253), .B(g7853), .Z(g8167) ) ;
AND2    gate8549  (.A(g5262), .B(g7853), .Z(g8168) ) ;
AND2    gate8550  (.A(g5265), .B(g7853), .Z(g8169) ) ;
AND2    gate8551  (.A(g5270), .B(g7853), .Z(g8170) ) ;
AND2    gate8552  (.A(g5275), .B(g7853), .Z(g8172) ) ;
OR2     gate8553  (.A(g5110), .B(g7549), .Z(g7971) ) ;
AND2    gate8554  (.A(g5284), .B(g7853), .Z(g8174) ) ;
AND2    gate8555  (.A(g5291), .B(g7853), .Z(g8175) ) ;
AND2    gate8556  (.A(g5299), .B(g7853), .Z(g8176) ) ;
AND2    gate8557  (.A(g664), .B(g7997), .Z(g8185) ) ;
AND3    gate8558  (.A(g4094), .B(g3792), .C(g7980), .Z(g8209) ) ;
AND2    gate8559  (.A(g1872), .B(g7883), .Z(g8217) ) ;
AND2    gate8560  (.A(g1882), .B(g7887), .Z(g8224) ) ;
OR2     gate8561  (.A(g7722), .B(g7241), .Z(g7846) ) ;
AND2    gate8562  (.A(g7846), .B(g7442), .Z(g8246) ) ;
OR2     gate8563  (.A(g5691), .B(g5052), .Z(g6777) ) ;
NAND2   gate8564  (.A(g5052), .B(g7853), .Z(g8109) ) ;
AND2    gate8565  (.A(g658), .B(g8235), .Z(g8364) ) ;
AND2    gate8566  (.A(g668), .B(g8240), .Z(g8365) ) ;
OR2     gate8567  (.A(g7902), .B(g7444), .Z(g8199) ) ;
OR2     gate8568  (.A(g6756), .B(g6204), .Z(g7265) ) ;
OR2     gate8569  (.A(g7988), .B(g7679), .Z(g8252) ) ;
AND2    gate8570  (.A(g8252), .B(g4240), .Z(g8380) ) ;
AND2    gate8571  (.A(g6077), .B(g8213), .Z(g8382) ) ;
NAND2   gate8572  (.A(II13090), .B(II13091), .Z(g8180) ) ;
AND2    gate8573  (.A(g6084), .B(g8218), .Z(g8385) ) ;
AND2    gate8574  (.A(g6085), .B(g8219), .Z(g8386) ) ;
AND2    gate8575  (.A(g6086), .B(g8220), .Z(g8387) ) ;
NAND2   gate8576  (.A(II13077), .B(II13078), .Z(g8177) ) ;
AND2    gate8577  (.A(g8177), .B(g7689), .Z(g8388) ) ;
AND2    gate8578  (.A(g6091), .B(g8225), .Z(g8389) ) ;
OR2     gate8579  (.A(g7962), .B(g7613), .Z(g8268) ) ;
OR2     gate8580  (.A(g5825), .B(g5041), .Z(g6465) ) ;
AND2    gate8581  (.A(g6094), .B(g8229), .Z(g8399) ) ;
AND2    gate8582  (.A(g6097), .B(g8234), .Z(g8400) ) ;
AND2    gate8583  (.A(g677), .B(g8124), .Z(g8401) ) ;
AND2    gate8584  (.A(g6101), .B(g8239), .Z(g8403) ) ;
AND2    gate8585  (.A(g686), .B(g8129), .Z(g8404) ) ;
AND2    gate8586  (.A(g695), .B(g8131), .Z(g8406) ) ;
AND2    gate8587  (.A(g704), .B(g8139), .Z(g8408) ) ;
AND2    gate8588  (.A(g713), .B(g8143), .Z(g8410) ) ;
AND2    gate8589  (.A(g722), .B(g8146), .Z(g8413) ) ;
AND2    gate8590  (.A(g731), .B(g8151), .Z(g8416) ) ;
NAND2   gate8591  (.A(II13249), .B(II13250), .Z(g8298) ) ;
AND2    gate8592  (.A(g8298), .B(g7403), .Z(g8461) ) ;
NAND2   gate8593  (.A(II13259), .B(II13260), .Z(g8300) ) ;
AND2    gate8594  (.A(g8300), .B(g7406), .Z(g8462) ) ;
NAND2   gate8595  (.A(II13266), .B(II13267), .Z(g8301) ) ;
AND2    gate8596  (.A(g8301), .B(g7410), .Z(g8463) ) ;
NAND2   gate8597  (.A(II13273), .B(II13274), .Z(g8302) ) ;
AND2    gate8598  (.A(g8302), .B(g7416), .Z(g8464) ) ;
NAND2   gate8599  (.A(II13284), .B(II13285), .Z(g8305) ) ;
AND2    gate8600  (.A(g8305), .B(g7422), .Z(g8469) ) ;
NAND2   gate8601  (.A(II13301), .B(II13302), .Z(g8308) ) ;
AND2    gate8602  (.A(g8308), .B(g7427), .Z(g8470) ) ;
OR2     gate8603  (.A(g8163), .B(g5051), .Z(g8383) ) ;
AND2    gate8604  (.A(g8383), .B(g5285), .Z(g8474) ) ;
OR2     gate8605  (.A(g8185), .B(g7958), .Z(g8377) ) ;
AND2    gate8606  (.A(g8377), .B(g4737), .Z(g8499) ) ;
NAND2   gate8607  (.A(II13308), .B(II13309), .Z(g8309) ) ;
NAND2   gate8608  (.A(II13538), .B(II13539), .Z(g8411) ) ;
AND2    gate8609  (.A(g8411), .B(g7967), .Z(g8508) ) ;
NAND2   gate8610  (.A(II13553), .B(II13554), .Z(g8414) ) ;
AND2    gate8611  (.A(g8414), .B(g7972), .Z(g8510) ) ;
NAND2   gate8612  (.A(II13294), .B(II13295), .Z(g8307) ) ;
AND2    gate8613  (.A(g8307), .B(g7693), .Z(g8547) ) ;
NAND2   gate8614  (.A(II13505), .B(II13506), .Z(g8402) ) ;
AND2    gate8615  (.A(g8402), .B(g8011), .Z(g8550) ) ;
NAND2   gate8616  (.A(II13514), .B(II13515), .Z(g8405) ) ;
AND2    gate8617  (.A(g8405), .B(g8015), .Z(g8553) ) ;
NAND2   gate8618  (.A(II13522), .B(II13523), .Z(g8407) ) ;
AND2    gate8619  (.A(g8407), .B(g8020), .Z(g8554) ) ;
NAND2   gate8620  (.A(II13530), .B(II13531), .Z(g8409) ) ;
AND2    gate8621  (.A(g8409), .B(g8025), .Z(g8555) ) ;
NAND2   gate8622  (.A(II13545), .B(II13546), .Z(g8412) ) ;
AND2    gate8623  (.A(g8412), .B(g8029), .Z(g8556) ) ;
NAND2   gate8624  (.A(II13560), .B(II13561), .Z(g8415) ) ;
AND2    gate8625  (.A(g8415), .B(g8033), .Z(g8557) ) ;
NAND2   gate8626  (.A(II13660), .B(II13661), .Z(g8471) ) ;
AND2    gate8627  (.A(g8471), .B(g7432), .Z(g8598) ) ;
NAND2   gate8628  (.A(g3440), .B(g2745), .Z(g4588) ) ;
NAND2   gate8629  (.A(g5277), .B(g8366), .Z(g8511) ) ;
AND2    gate8630  (.A(g4588), .B(g8511), .Z(g8648) ) ;
AND2    gate8631  (.A(g8520), .B(g4013), .Z(g8651) ) ;
AND2    gate8632  (.A(g8523), .B(g4013), .Z(g8652) ) ;
AND2    gate8633  (.A(g8526), .B(g4013), .Z(g8653) ) ;
AND2    gate8634  (.A(g8529), .B(g4013), .Z(g8654) ) ;
AND2    gate8635  (.A(g8532), .B(g4013), .Z(g8655) ) ;
AND2    gate8636  (.A(g8535), .B(g4013), .Z(g8659) ) ;
AND2    gate8637  (.A(g8538), .B(g4013), .Z(g8663) ) ;
NAND2   gate8638  (.A(g3664), .B(g2356), .Z(g4803) ) ;
NAND2   gate8639  (.A(g5527), .B(g8390), .Z(g8549) ) ;
AND2    gate8640  (.A(g4803), .B(g8549), .Z(g8683) ) ;
NAND2   gate8641  (.A(II13766), .B(II13767), .Z(g8558) ) ;
AND2    gate8642  (.A(g8558), .B(g8036), .Z(g8687) ) ;
AND2    gate8643  (.A(g3738), .B(g8509), .Z(g8693) ) ;
AND2    gate8644  (.A(g7591), .B(g8576), .Z(g8698) ) ;
AND2    gate8645  (.A(g7595), .B(g8579), .Z(g8699) ) ;
AND2    gate8646  (.A(g7597), .B(g8582), .Z(g8701) ) ;
AND2    gate8647  (.A(g7601), .B(g8585), .Z(g8703) ) ;
AND2    gate8648  (.A(g7602), .B(g8589), .Z(g8706) ) ;
AND2    gate8649  (.A(g7605), .B(g8592), .Z(g8708) ) ;
AND2    gate8650  (.A(g7607), .B(g8595), .Z(g8710) ) ;
AND2    gate8651  (.A(g8600), .B(g7903), .Z(g8718) ) ;
AND2    gate8652  (.A(g8601), .B(g7905), .Z(g8720) ) ;
AND2    gate8653  (.A(g8604), .B(g7908), .Z(g8722) ) ;
AND2    gate8654  (.A(g8606), .B(g7910), .Z(g8724) ) ;
AND2    gate8655  (.A(g8608), .B(g7913), .Z(g8726) ) ;
AND2    gate8656  (.A(g8610), .B(g7915), .Z(g8728) ) ;
AND2    gate8657  (.A(g8613), .B(g7917), .Z(g8730) ) ;
AND2    gate8658  (.A(g8622), .B(g7918), .Z(g8731) ) ;
AND2    gate8659  (.A(g8624), .B(g7919), .Z(g8732) ) ;
AND2    gate8660  (.A(g8625), .B(g7920), .Z(g8733) ) ;
AND2    gate8661  (.A(g8626), .B(g7923), .Z(g8734) ) ;
AND2    gate8662  (.A(g7600), .B(g8632), .Z(g8735) ) ;
AND2    gate8663  (.A(g7439), .B(g8635), .Z(g8736) ) ;
AND2    gate8664  (.A(g7670), .B(g8656), .Z(g8748) ) ;
AND2    gate8665  (.A(g7604), .B(g8660), .Z(g8749) ) ;
AND2    gate8666  (.A(g7414), .B(g8664), .Z(g8753) ) ;
AND2    gate8667  (.A(g7420), .B(g8667), .Z(g8754) ) ;
AND2    gate8668  (.A(g7426), .B(g8671), .Z(g8755) ) ;
AND2    gate8669  (.A(g7431), .B(g8674), .Z(g8756) ) ;
AND2    gate8670  (.A(g7437), .B(g8677), .Z(g8759) ) ;
AND2    gate8671  (.A(g7440), .B(g8680), .Z(g8763) ) ;
AND2    gate8672  (.A(g7443), .B(g8684), .Z(g8764) ) ;
NAND2   gate8673  (.A(II13908), .B(II13909), .Z(g8630) ) ;
NAND2   gate8674  (.A(II13858), .B(II13859), .Z(g8612) ) ;
NAND2   gate8675  (.A(II13868), .B(II13869), .Z(g8616) ) ;
NAND2   gate8676  (.A(II13877), .B(II13878), .Z(g8623) ) ;
NAND2   gate8677  (.A(II13901), .B(II13902), .Z(g8629) ) ;
NAND2   gate8678  (.A(II13887), .B(II13888), .Z(g8627) ) ;
NAND2   gate8679  (.A(II13894), .B(II13895), .Z(g8628) ) ;
AND2    gate8680  (.A(g8688), .B(g2317), .Z(g8778) ) ;
OR2     gate8681  (.A(g8108), .B(g8461), .Z(g8638) ) ;
AND2    gate8682  (.A(g8638), .B(g8716), .Z(g8786) ) ;
OR2     gate8683  (.A(g8118), .B(g8462), .Z(g8639) ) ;
AND2    gate8684  (.A(g8639), .B(g8719), .Z(g8789) ) ;
OR2     gate8685  (.A(g8120), .B(g8463), .Z(g8641) ) ;
AND2    gate8686  (.A(g8641), .B(g8721), .Z(g8791) ) ;
OR2     gate8687  (.A(g8123), .B(g8464), .Z(g8644) ) ;
AND2    gate8688  (.A(g8644), .B(g8723), .Z(g8793) ) ;
OR2     gate8689  (.A(g8127), .B(g8469), .Z(g8645) ) ;
AND2    gate8690  (.A(g8645), .B(g8725), .Z(g8796) ) ;
OR2     gate8691  (.A(g8130), .B(g8470), .Z(g8647) ) ;
AND2    gate8692  (.A(g8647), .B(g8727), .Z(g8799) ) ;
OR2     gate8693  (.A(g8135), .B(g8598), .Z(g8742) ) ;
AND2    gate8694  (.A(g8742), .B(g8729), .Z(g8801) ) ;
NAND2   gate8695  (.A(II13991), .B(II13992), .Z(g8705) ) ;
OR2     gate8696  (.A(g8364), .B(g8508), .Z(g8643) ) ;
AND2    gate8697  (.A(g8643), .B(g8751), .Z(g8821) ) ;
OR2     gate8698  (.A(g8365), .B(g8510), .Z(g8614) ) ;
AND2    gate8699  (.A(g8614), .B(g8752), .Z(g8822) ) ;
OR2     gate8700  (.A(g8217), .B(g8388), .Z(g8552) ) ;
AND2    gate8701  (.A(g8552), .B(g8696), .Z(g8827) ) ;
OR2     gate8702  (.A(g8224), .B(g8547), .Z(g8646) ) ;
AND2    gate8703  (.A(g8646), .B(g8697), .Z(g8837) ) ;
OR2     gate8704  (.A(g8401), .B(g8550), .Z(g8602) ) ;
AND2    gate8705  (.A(g8602), .B(g8702), .Z(g8838) ) ;
OR2     gate8706  (.A(g8404), .B(g8553), .Z(g8605) ) ;
AND2    gate8707  (.A(g8605), .B(g8704), .Z(g8841) ) ;
OR2     gate8708  (.A(g8406), .B(g8554), .Z(g8607) ) ;
AND2    gate8709  (.A(g8607), .B(g8707), .Z(g8842) ) ;
OR2     gate8710  (.A(g8408), .B(g8555), .Z(g8609) ) ;
AND2    gate8711  (.A(g8609), .B(g8709), .Z(g8844) ) ;
OR2     gate8712  (.A(g8410), .B(g8556), .Z(g8611) ) ;
AND2    gate8713  (.A(g8611), .B(g8711), .Z(g8845) ) ;
OR2     gate8714  (.A(g8413), .B(g8557), .Z(g8615) ) ;
AND2    gate8715  (.A(g8615), .B(g8712), .Z(g8846) ) ;
OR2     gate8716  (.A(g8416), .B(g8687), .Z(g8715) ) ;
AND2    gate8717  (.A(g8715), .B(g8713), .Z(g8848) ) ;
AND3    gate8718  (.A(g8255), .B(g6368), .C(g8858), .Z(g8875) ) ;
AND3    gate8719  (.A(g8105), .B(g6764), .C(g8858), .Z(g8876) ) ;
AND3    gate8720  (.A(g8103), .B(g6764), .C(g8858), .Z(g8877) ) ;
AND3    gate8721  (.A(g8099), .B(g6368), .C(g8858), .Z(g8878) ) ;
AND3    gate8722  (.A(g8110), .B(g6764), .C(g8858), .Z(g8879) ) ;
AND2    gate8723  (.A(g7872), .B(g8807), .Z(g8927) ) ;
AND3    gate8724  (.A(g8095), .B(g6368), .C(g8828), .Z(g8929) ) ;
AND3    gate8725  (.A(g8100), .B(g6368), .C(g8828), .Z(g8930) ) ;
AND2    gate8726  (.A(g8807), .B(g8164), .Z(g8931) ) ;
AND3    gate8727  (.A(g8106), .B(g6778), .C(g8849), .Z(g8935) ) ;
AND3    gate8728  (.A(g8115), .B(g6778), .C(g8849), .Z(g8936) ) ;
AND3    gate8729  (.A(g8056), .B(g6368), .C(g8828), .Z(g8947) ) ;
AND3    gate8730  (.A(g8255), .B(g6368), .C(g8828), .Z(g8949) ) ;
AND3    gate8731  (.A(g8110), .B(g6368), .C(g8828), .Z(g8955) ) ;
AND3    gate8732  (.A(g8081), .B(g6368), .C(g8828), .Z(g8957) ) ;
AND3    gate8733  (.A(g8085), .B(g6368), .C(g8828), .Z(g8960) ) ;
AND3    gate8734  (.A(g8089), .B(g6368), .C(g8828), .Z(g8962) ) ;
AND3    gate8735  (.A(g8056), .B(g6368), .C(g8849), .Z(g8963) ) ;
AND3    gate8736  (.A(g8255), .B(g6368), .C(g8849), .Z(g8964) ) ;
AND3    gate8737  (.A(g8110), .B(g6778), .C(g8849), .Z(g8965) ) ;
AND3    gate8738  (.A(g8081), .B(g6778), .C(g8849), .Z(g8966) ) ;
AND3    gate8739  (.A(g8085), .B(g6778), .C(g8849), .Z(g8967) ) ;
AND3    gate8740  (.A(g8089), .B(g6778), .C(g8849), .Z(g8968) ) ;
AND3    gate8741  (.A(g8081), .B(g6764), .C(g8858), .Z(g8971) ) ;
AND3    gate8742  (.A(g8085), .B(g6764), .C(g8858), .Z(g8972) ) ;
AND3    gate8743  (.A(g8094), .B(g6368), .C(g8858), .Z(g8974) ) ;
AND3    gate8744  (.A(g8089), .B(g6764), .C(g8858), .Z(g8975) ) ;
AND3    gate8745  (.A(g8110), .B(g6778), .C(g8925), .Z(g8994) ) ;
AND2    gate8746  (.A(g6454), .B(g8929), .Z(g8995) ) ;
AND2    gate8747  (.A(g6454), .B(g8930), .Z(g9010) ) ;
AND2    gate8748  (.A(g8935), .B(g7192), .Z(g9030) ) ;
NAND2   gate8749  (.A(II14203), .B(II14204), .Z(g8880) ) ;
AND2    gate8750  (.A(g8965), .B(g6674), .Z(g9111) ) ;
NAND2   gate8751  (.A(II14210), .B(II14211), .Z(g8881) ) ;
AND2    gate8752  (.A(g8966), .B(g6674), .Z(g9125) ) ;
NAND2   gate8753  (.A(II14217), .B(II14218), .Z(g8882) ) ;
AND2    gate8754  (.A(g8967), .B(g6674), .Z(g9151) ) ;
AND2    gate8755  (.A(g8968), .B(g6674), .Z(g9173) ) ;
AND2    gate8756  (.A(g6454), .B(g8955), .Z(g9192) ) ;
AND2    gate8757  (.A(g6454), .B(g8957), .Z(g9205) ) ;
AND2    gate8758  (.A(g6454), .B(g8960), .Z(g9223) ) ;
AND2    gate8759  (.A(g6454), .B(g8962), .Z(g9240) ) ;
NAND2   gate8760  (.A(II14264), .B(II14265), .Z(g8932) ) ;
NAND2   gate8761  (.A(II14271), .B(II14272), .Z(g8933) ) ;
NAND2   gate8762  (.A(II14278), .B(II14279), .Z(g8934) ) ;
AND2    gate8763  (.A(g8974), .B(g5708), .Z(g9274) ) ;
AND2    gate8764  (.A(g8878), .B(g5708), .Z(g9292) ) ;
AND2    gate8765  (.A(g8877), .B(g5708), .Z(g9316) ) ;
AND2    gate8766  (.A(g6109), .B(g8875), .Z(g9317) ) ;
AND2    gate8767  (.A(g8971), .B(g5708), .Z(g9328) ) ;
AND2    gate8768  (.A(g8975), .B(g5708), .Z(g9335) ) ;
AND2    gate8769  (.A(g962), .B(g9223), .Z(g9357) ) ;
AND2    gate8770  (.A(g1318), .B(g9151), .Z(g9358) ) ;
AND2    gate8771  (.A(g1308), .B(g9173), .Z(g9359) ) ;
AND2    gate8772  (.A(g965), .B(g9223), .Z(g9364) ) ;
AND2    gate8773  (.A(g1321), .B(g9151), .Z(g9365) ) ;
AND2    gate8774  (.A(g1311), .B(g9173), .Z(g9366) ) ;
AND2    gate8775  (.A(g968), .B(g9223), .Z(g9384) ) ;
AND2    gate8776  (.A(g1324), .B(g9151), .Z(g9385) ) ;
AND2    gate8777  (.A(g1327), .B(g9151), .Z(g9386) ) ;
AND2    gate8778  (.A(g1330), .B(g9151), .Z(g9389) ) ;
AND2    gate8779  (.A(g1333), .B(g9151), .Z(g9390) ) ;
AND2    gate8780  (.A(g1721), .B(g9052), .Z(g9409) ) ;
AND2    gate8781  (.A(g1724), .B(g9052), .Z(g9411) ) ;
AND2    gate8782  (.A(g1727), .B(g9052), .Z(g9412) ) ;
AND2    gate8783  (.A(g1730), .B(g9052), .Z(g9414) ) ;
AND2    gate8784  (.A(g1733), .B(g9052), .Z(g9415) ) ;
AND2    gate8785  (.A(g1738), .B(g9052), .Z(g9417) ) ;
AND2    gate8786  (.A(g1741), .B(g9052), .Z(g9418) ) ;
AND2    gate8787  (.A(g1744), .B(g9030), .Z(g9419) ) ;
AND2    gate8788  (.A(g1747), .B(g9030), .Z(g9420) ) ;
AND2    gate8789  (.A(g1750), .B(g9030), .Z(g9422) ) ;
AND2    gate8790  (.A(g1753), .B(g9030), .Z(g9425) ) ;
AND2    gate8791  (.A(g1756), .B(g9030), .Z(g9428) ) ;
AND2    gate8792  (.A(g1759), .B(g9030), .Z(g9430) ) ;
AND2    gate8793  (.A(g1762), .B(g9030), .Z(g9447) ) ;
NAND2   gate8794  (.A(II14443), .B(II14444), .Z(g9107) ) ;
AND2    gate8795  (.A(g2725), .B(g9173), .Z(g9582) ) ;
AND2    gate8796  (.A(g886), .B(g8995), .Z(g9583) ) ;
AND2    gate8797  (.A(g2726), .B(g9173), .Z(g9584) ) ;
AND2    gate8798  (.A(g889), .B(g8995), .Z(g9585) ) ;
AND2    gate8799  (.A(g2727), .B(g9173), .Z(g9586) ) ;
AND2    gate8800  (.A(g892), .B(g8995), .Z(g9587) ) ;
AND2    gate8801  (.A(g3272), .B(g9173), .Z(g9588) ) ;
AND2    gate8802  (.A(g895), .B(g8995), .Z(g9590) ) ;
AND2    gate8803  (.A(g4), .B(g9292), .Z(g9592) ) ;
AND2    gate8804  (.A(g898), .B(g9205), .Z(g9593) ) ;
AND2    gate8805  (.A(g1), .B(g9292), .Z(g9594) ) ;
AND2    gate8806  (.A(g901), .B(g9205), .Z(g9595) ) ;
AND2    gate8807  (.A(g2649), .B(g9010), .Z(g9596) ) ;
AND2    gate8808  (.A(g1170), .B(g9125), .Z(g9597) ) ;
AND2    gate8809  (.A(g2086), .B(g9274), .Z(g9598) ) ;
AND2    gate8810  (.A(g8), .B(g9292), .Z(g9599) ) ;
AND2    gate8811  (.A(g904), .B(g9205), .Z(g9600) ) ;
AND2    gate8812  (.A(g922), .B(g9192), .Z(g9601) ) ;
AND2    gate8813  (.A(g2650), .B(g9010), .Z(g9602) ) ;
AND2    gate8814  (.A(g1173), .B(g9125), .Z(g9603) ) ;
AND2    gate8815  (.A(g1194), .B(g9111), .Z(g9604) ) ;
AND2    gate8816  (.A(g12), .B(g9274), .Z(g9607) ) ;
AND2    gate8817  (.A(g7), .B(g9292), .Z(g9608) ) ;
AND2    gate8818  (.A(g907), .B(g9205), .Z(g9609) ) ;
AND2    gate8819  (.A(g925), .B(g9192), .Z(g9610) ) ;
AND2    gate8820  (.A(g2651), .B(g9010), .Z(g9611) ) ;
AND2    gate8821  (.A(g2652), .B(g9240), .Z(g9612) ) ;
AND2    gate8822  (.A(g1176), .B(g9125), .Z(g9613) ) ;
AND2    gate8823  (.A(g1197), .B(g9111), .Z(g9614) ) ;
AND2    gate8824  (.A(g9), .B(g9274), .Z(g9617) ) ;
AND2    gate8825  (.A(g910), .B(g9205), .Z(g9618) ) ;
AND2    gate8826  (.A(g2772), .B(g9010), .Z(g9619) ) ;
AND2    gate8827  (.A(g2653), .B(g9240), .Z(g9620) ) ;
AND2    gate8828  (.A(g1179), .B(g9125), .Z(g9621) ) ;
AND2    gate8829  (.A(g1200), .B(g9111), .Z(g9622) ) ;
AND2    gate8830  (.A(g17), .B(g9274), .Z(g9623) ) ;
AND2    gate8831  (.A(g913), .B(g9205), .Z(g9641) ) ;
AND2    gate8832  (.A(g2654), .B(g9240), .Z(g9642) ) ;
AND2    gate8833  (.A(g950), .B(g9223), .Z(g9643) ) ;
AND2    gate8834  (.A(g1182), .B(g9125), .Z(g9644) ) ;
AND2    gate8835  (.A(g1203), .B(g9111), .Z(g9645) ) ;
AND2    gate8836  (.A(g16), .B(g9274), .Z(g9648) ) ;
AND2    gate8837  (.A(g916), .B(g9205), .Z(g9649) ) ;
AND2    gate8838  (.A(g2797), .B(g9240), .Z(g9650) ) ;
AND2    gate8839  (.A(g944), .B(g9240), .Z(g9651) ) ;
AND2    gate8840  (.A(g953), .B(g9223), .Z(g9652) ) ;
AND2    gate8841  (.A(g1185), .B(g9125), .Z(g9653) ) ;
AND2    gate8842  (.A(g919), .B(g9205), .Z(g9657) ) ;
AND2    gate8843  (.A(g947), .B(g9240), .Z(g9658) ) ;
AND2    gate8844  (.A(g956), .B(g9223), .Z(g9659) ) ;
AND2    gate8845  (.A(g1188), .B(g9125), .Z(g9660) ) ;
AND2    gate8846  (.A(g2094), .B(g9292), .Z(g9662) ) ;
AND2    gate8847  (.A(g959), .B(g9223), .Z(g9663) ) ;
AND2    gate8848  (.A(g1191), .B(g9125), .Z(g9664) ) ;
AND2    gate8849  (.A(g1314), .B(g9151), .Z(g9665) ) ;
AND2    gate8850  (.A(g263), .B(g9432), .Z(g9689) ) ;
AND2    gate8851  (.A(g266), .B(g9432), .Z(g9690) ) ;
AND2    gate8852  (.A(g269), .B(g9432), .Z(g9691) ) ;
AND2    gate8853  (.A(g272), .B(g9432), .Z(g9692) ) ;
AND2    gate8854  (.A(g275), .B(g9432), .Z(g9693) ) ;
AND2    gate8855  (.A(g278), .B(g9432), .Z(g9694) ) ;
AND2    gate8856  (.A(g1567), .B(g9474), .Z(g9695) ) ;
AND2    gate8857  (.A(g1571), .B(g9474), .Z(g9698) ) ;
AND2    gate8858  (.A(g1574), .B(g9474), .Z(g9701) ) ;
AND2    gate8859  (.A(g1577), .B(g9474), .Z(g9703) ) ;
AND2    gate8860  (.A(g1580), .B(g9474), .Z(g9705) ) ;
AND2    gate8861  (.A(g1583), .B(g9474), .Z(g9707) ) ;
AND2    gate8862  (.A(g1524), .B(g9490), .Z(g9709) ) ;
AND2    gate8863  (.A(g1528), .B(g9490), .Z(g9712) ) ;
AND2    gate8864  (.A(g1531), .B(g9490), .Z(g9715) ) ;
AND2    gate8865  (.A(g1534), .B(g9490), .Z(g9716) ) ;
AND2    gate8866  (.A(g1537), .B(g9490), .Z(g9717) ) ;
AND2    gate8867  (.A(g1540), .B(g9490), .Z(g9718) ) ;
NAND2   gate8868  (.A(II14613), .B(II14614), .Z(g9413) ) ;
OR4     gate8869  (.A(g9612), .B(g9643), .C(g9410), .D(II14855), .Z(g9722) ) ;
OR4     gate8870  (.A(g9010), .B(g8995), .C(g9388), .D(g9363), .Z(g9785) ) ;
AND2    gate8871  (.A(g9722), .B(g9785), .Z(g9828) ) ;
OR4     gate8872  (.A(g9620), .B(g9652), .C(g9391), .D(II14858), .Z(g9723) ) ;
AND2    gate8873  (.A(g9723), .B(g9785), .Z(g9829) ) ;
OR4     gate8874  (.A(g9642), .B(g9659), .C(g9616), .D(II14862), .Z(g9725) ) ;
AND2    gate8875  (.A(g9725), .B(g9785), .Z(g9830) ) ;
OR4     gate8876  (.A(g9650), .B(g9663), .C(g9362), .D(II14866), .Z(g9727) ) ;
AND2    gate8877  (.A(g9727), .B(g9785), .Z(g9831) ) ;
OR3     gate8878  (.A(g9618), .B(g9357), .C(g9656), .Z(g9729) ) ;
AND2    gate8879  (.A(g9729), .B(g9785), .Z(g9833) ) ;
OR3     gate8880  (.A(g9641), .B(g9364), .C(g9387), .Z(g9731) ) ;
AND2    gate8881  (.A(g9731), .B(g9785), .Z(g9834) ) ;
OR4     gate8882  (.A(g9649), .B(g9651), .C(g9384), .D(g9361), .Z(g9735) ) ;
AND2    gate8883  (.A(g9735), .B(g9785), .Z(g9835) ) ;
OR3     gate8884  (.A(g9657), .B(g9658), .C(g9655), .Z(g9737) ) ;
AND2    gate8885  (.A(g9737), .B(g9785), .Z(g9836) ) ;
OR3     gate8886  (.A(g9665), .B(g9606), .C(II14822), .Z(g9697) ) ;
OR2     gate8887  (.A(g9515), .B(g9510), .Z(g9751) ) ;
AND2    gate8888  (.A(g9697), .B(g9751), .Z(g9837) ) ;
OR3     gate8889  (.A(g9358), .B(g9667), .C(II14827), .Z(g9700) ) ;
OR2     gate8890  (.A(g9173), .B(g9511), .Z(g9754) ) ;
AND2    gate8891  (.A(g9700), .B(g9754), .Z(g9838) ) ;
OR3     gate8892  (.A(g9365), .B(g9647), .C(II14831), .Z(g9702) ) ;
OR2     gate8893  (.A(g9173), .B(g9528), .Z(g9742) ) ;
AND2    gate8894  (.A(g9702), .B(g9742), .Z(g9839) ) ;
OR3     gate8895  (.A(g9385), .B(g9605), .C(II14835), .Z(g9704) ) ;
OR2     gate8896  (.A(g9173), .B(g9509), .Z(g9747) ) ;
AND2    gate8897  (.A(g9704), .B(g9747), .Z(g9840) ) ;
OR3     gate8898  (.A(g9644), .B(g9386), .C(g9591), .Z(g9706) ) ;
OR2     gate8899  (.A(g9151), .B(g9125), .Z(g9512) ) ;
AND2    gate8900  (.A(g9706), .B(g9512), .Z(g9841) ) ;
OR3     gate8901  (.A(g9653), .B(g9389), .C(g9646), .Z(g9708) ) ;
OR2     gate8902  (.A(g9151), .B(g9125), .Z(g9516) ) ;
AND2    gate8903  (.A(g9708), .B(g9516), .Z(g9842) ) ;
OR4     gate8904  (.A(g9660), .B(g9390), .C(g9359), .D(g9589), .Z(g9711) ) ;
OR3     gate8905  (.A(g9173), .B(g9151), .C(g9125), .Z(g9519) ) ;
AND2    gate8906  (.A(g9711), .B(g9519), .Z(g9843) ) ;
OR3     gate8907  (.A(g9664), .B(g9366), .C(g9654), .Z(g9714) ) ;
OR2     gate8908  (.A(g9173), .B(g9125), .Z(g9522) ) ;
AND2    gate8909  (.A(g9714), .B(g9522), .Z(g9844) ) ;
AND2    gate8910  (.A(g287), .B(g9764), .Z(g9846) ) ;
AND2    gate8911  (.A(g290), .B(g9766), .Z(g9847) ) ;
OR3     gate8912  (.A(g9409), .B(g9419), .C(g9615), .Z(g9724) ) ;
OR2     gate8913  (.A(g9052), .B(g9030), .Z(g9557) ) ;
AND2    gate8914  (.A(g9724), .B(g9557), .Z(g9848) ) ;
AND2    gate8915  (.A(g293), .B(g9768), .Z(g9849) ) ;
OR3     gate8916  (.A(g9411), .B(g9420), .C(g9489), .Z(g9726) ) ;
OR2     gate8917  (.A(g9052), .B(g9030), .Z(g9560) ) ;
AND2    gate8918  (.A(g9726), .B(g9560), .Z(g9850) ) ;
AND2    gate8919  (.A(g296), .B(g9770), .Z(g9851) ) ;
OR3     gate8920  (.A(g9412), .B(g9422), .C(g9426), .Z(g9728) ) ;
OR2     gate8921  (.A(g9052), .B(g9030), .Z(g9563) ) ;
AND2    gate8922  (.A(g9728), .B(g9563), .Z(g9852) ) ;
AND2    gate8923  (.A(g299), .B(g9771), .Z(g9853) ) ;
OR3     gate8924  (.A(g9414), .B(g9425), .C(g9423), .Z(g9730) ) ;
OR2     gate8925  (.A(g9052), .B(g9030), .Z(g9566) ) ;
AND2    gate8926  (.A(g9730), .B(g9566), .Z(g9854) ) ;
AND2    gate8927  (.A(g302), .B(g9772), .Z(g9855) ) ;
AND2    gate8928  (.A(g1592), .B(g9773), .Z(g9856) ) ;
OR3     gate8929  (.A(g9415), .B(g9428), .C(g9421), .Z(g9734) ) ;
OR2     gate8930  (.A(g9052), .B(g9030), .Z(g9569) ) ;
AND2    gate8931  (.A(g9734), .B(g9569), .Z(g9857) ) ;
AND2    gate8932  (.A(g1595), .B(g9774), .Z(g9858) ) ;
OR2     gate8933  (.A(g9430), .B(g9416), .Z(g9736) ) ;
OR2     gate8934  (.A(g9052), .B(g9030), .Z(g9573) ) ;
AND2    gate8935  (.A(g9736), .B(g9573), .Z(g9859) ) ;
AND2    gate8936  (.A(g1598), .B(g9775), .Z(g9860) ) ;
OR3     gate8937  (.A(g9417), .B(g9447), .C(g9506), .Z(g9738) ) ;
OR2     gate8938  (.A(g9052), .B(g9030), .Z(g9579) ) ;
AND2    gate8939  (.A(g9738), .B(g9579), .Z(g9861) ) ;
AND2    gate8940  (.A(g1601), .B(g9777), .Z(g9862) ) ;
OR2     gate8941  (.A(g9418), .B(g9505), .Z(g9740) ) ;
AND2    gate8942  (.A(g9740), .B(g9576), .Z(g9863) ) ;
AND2    gate8943  (.A(g1604), .B(g9778), .Z(g9864) ) ;
AND2    gate8944  (.A(g1607), .B(g9780), .Z(g9865) ) ;
AND2    gate8945  (.A(g1549), .B(g9802), .Z(g9866) ) ;
AND2    gate8946  (.A(g1552), .B(g9807), .Z(g9867) ) ;
AND2    gate8947  (.A(g1555), .B(g9812), .Z(g9868) ) ;
AND2    gate8948  (.A(g1558), .B(g9814), .Z(g9869) ) ;
AND2    gate8949  (.A(g1561), .B(g9816), .Z(g9870) ) ;
AND2    gate8950  (.A(g1564), .B(g9668), .Z(g9871) ) ;
OR2     gate8951  (.A(g9316), .B(g9313), .Z(g9624) ) ;
AND2    gate8952  (.A(g9883), .B(g9624), .Z(g9896) ) ;
AND2    gate8953  (.A(g9884), .B(g9624), .Z(g9897) ) ;
OR2     gate8954  (.A(g9335), .B(g9331), .Z(g9367) ) ;
AND2    gate8955  (.A(g9887), .B(g9367), .Z(g9898) ) ;
AND2    gate8956  (.A(g9889), .B(g9367), .Z(g9899) ) ;
AND2    gate8957  (.A(g9845), .B(g8327), .Z(g9900) ) ;
OR2     gate8958  (.A(g9328), .B(g9324), .Z(g9392) ) ;
AND2    gate8959  (.A(g9893), .B(g9392), .Z(g9901) ) ;
AND2    gate8960  (.A(g9894), .B(g9392), .Z(g9902) ) ;
OR4     gate8961  (.A(g9739), .B(g9598), .C(g9662), .D(g9746), .Z(g9885) ) ;
OR3     gate8962  (.A(g9454), .B(g9292), .C(g9274), .Z(g9673) ) ;
AND2    gate8963  (.A(g9885), .B(g9673), .Z(g9903) ) ;
OR3     gate8964  (.A(g9607), .B(g9592), .C(g9759), .Z(g9886) ) ;
OR3     gate8965  (.A(g9454), .B(g9292), .C(g9274), .Z(g9676) ) ;
AND2    gate8966  (.A(g9886), .B(g9676), .Z(g9904) ) ;
OR3     gate8967  (.A(g9617), .B(g9594), .C(g9750), .Z(g9872) ) ;
OR3     gate8968  (.A(g9454), .B(g9292), .C(g9274), .Z(g9680) ) ;
AND2    gate8969  (.A(g9872), .B(g9680), .Z(g9905) ) ;
OR3     gate8970  (.A(g9623), .B(g9599), .C(g9758), .Z(g9873) ) ;
OR3     gate8971  (.A(g9454), .B(g9292), .C(g9274), .Z(g9683) ) ;
AND2    gate8972  (.A(g9873), .B(g9683), .Z(g9906) ) ;
OR3     gate8973  (.A(g9648), .B(g9608), .C(g9757), .Z(g9888) ) ;
OR3     gate8974  (.A(g9454), .B(g9292), .C(g9274), .Z(g9686) ) ;
AND2    gate8975  (.A(g9888), .B(g9686), .Z(g9907) ) ;
AND2    gate8976  (.A(g9890), .B(g9782), .Z(g9908) ) ;
OR2     gate8977  (.A(g9741), .B(g9760), .Z(g9891) ) ;
AND2    gate8978  (.A(g9891), .B(g9804), .Z(g9909) ) ;
AND2    gate8979  (.A(g9892), .B(g9809), .Z(g9910) ) ;
OR2     gate8980  (.A(g9846), .B(g9689), .Z(g9911) ) ;
AND2    gate8981  (.A(g9911), .B(g9624), .Z(g9932) ) ;
OR2     gate8982  (.A(g9847), .B(g9690), .Z(g9912) ) ;
AND2    gate8983  (.A(g9912), .B(g9624), .Z(g9933) ) ;
OR2     gate8984  (.A(g9849), .B(g9691), .Z(g9913) ) ;
AND2    gate8985  (.A(g9913), .B(g9624), .Z(g9934) ) ;
OR2     gate8986  (.A(g9851), .B(g9692), .Z(g9914) ) ;
AND2    gate8987  (.A(g9914), .B(g9624), .Z(g9935) ) ;
OR2     gate8988  (.A(g9853), .B(g9693), .Z(g9915) ) ;
AND2    gate8989  (.A(g9915), .B(g9624), .Z(g9936) ) ;
OR2     gate8990  (.A(g9855), .B(g9694), .Z(g9916) ) ;
AND2    gate8991  (.A(g9916), .B(g9624), .Z(g9937) ) ;
OR2     gate8992  (.A(g9856), .B(g9695), .Z(g9917) ) ;
AND2    gate8993  (.A(g9917), .B(g9367), .Z(g9938) ) ;
OR2     gate8994  (.A(g9858), .B(g9698), .Z(g9918) ) ;
AND2    gate8995  (.A(g9918), .B(g9367), .Z(g9939) ) ;
OR2     gate8996  (.A(g9860), .B(g9701), .Z(g9920) ) ;
AND2    gate8997  (.A(g9920), .B(g9367), .Z(g9940) ) ;
OR2     gate8998  (.A(g9862), .B(g9703), .Z(g9921) ) ;
AND2    gate8999  (.A(g9921), .B(g9367), .Z(g9941) ) ;
OR2     gate9000  (.A(g9864), .B(g9705), .Z(g9922) ) ;
AND2    gate9001  (.A(g9922), .B(g9367), .Z(g9942) ) ;
OR2     gate9002  (.A(g9865), .B(g9707), .Z(g9923) ) ;
AND2    gate9003  (.A(g9923), .B(g9367), .Z(g9943) ) ;
OR2     gate9004  (.A(g9866), .B(g9709), .Z(g9924) ) ;
AND2    gate9005  (.A(g9924), .B(g9392), .Z(g9944) ) ;
OR2     gate9006  (.A(g9867), .B(g9712), .Z(g9925) ) ;
AND2    gate9007  (.A(g9925), .B(g9392), .Z(g9945) ) ;
OR2     gate9008  (.A(g9868), .B(g9715), .Z(g9926) ) ;
AND2    gate9009  (.A(g9926), .B(g9392), .Z(g9946) ) ;
OR2     gate9010  (.A(g9869), .B(g9716), .Z(g9927) ) ;
AND2    gate9011  (.A(g9927), .B(g9392), .Z(g9947) ) ;
OR2     gate9012  (.A(g9870), .B(g9717), .Z(g9928) ) ;
AND2    gate9013  (.A(g9928), .B(g9392), .Z(g9948) ) ;
OR2     gate9014  (.A(g9871), .B(g9718), .Z(g9929) ) ;
AND2    gate9015  (.A(g9929), .B(g9392), .Z(g9949) ) ;
OR3     gate9016  (.A(g9901), .B(g9898), .C(g9779), .Z(g9950) ) ;
OR4     gate9017  (.A(g9335), .B(g9331), .C(g9328), .D(g9324), .Z(g9536) ) ;
AND2    gate9018  (.A(g9950), .B(g9536), .Z(g9959) ) ;
OR3     gate9019  (.A(g9902), .B(g9899), .C(g9803), .Z(g9951) ) ;
AND2    gate9020  (.A(g9951), .B(g9536), .Z(g9960) ) ;
OR3     gate9021  (.A(g9944), .B(g9938), .C(g9817), .Z(g9952) ) ;
AND2    gate9022  (.A(g9952), .B(g9536), .Z(g9962) ) ;
OR3     gate9023  (.A(g9945), .B(g9939), .C(g9669), .Z(g9953) ) ;
AND2    gate9024  (.A(g9953), .B(g9536), .Z(g9963) ) ;
OR3     gate9025  (.A(g9946), .B(g9940), .C(g9781), .Z(g9954) ) ;
AND2    gate9026  (.A(g9954), .B(g9536), .Z(g9964) ) ;
OR3     gate9027  (.A(g9947), .B(g9941), .C(g9808), .Z(g9955) ) ;
AND2    gate9028  (.A(g9955), .B(g9536), .Z(g9965) ) ;
OR3     gate9029  (.A(g9948), .B(g9942), .C(g9815), .Z(g9956) ) ;
AND2    gate9030  (.A(g9956), .B(g9536), .Z(g9966) ) ;
OR3     gate9031  (.A(g9949), .B(g9943), .C(g9776), .Z(g9957) ) ;
AND2    gate9032  (.A(g9957), .B(g9536), .Z(g9967) ) ;
AND2    gate9033  (.A(g8892), .B(g10145), .Z(g10230) ) ;
AND2    gate9034  (.A(g8892), .B(g10150), .Z(g10232) ) ;
AND2    gate9035  (.A(g10145), .B(g9100), .Z(g10237) ) ;
AND2    gate9036  (.A(g10150), .B(g9103), .Z(g10240) ) ;
AND2    gate9037  (.A(g8892), .B(g10208), .Z(g10295) ) ;
AND2    gate9038  (.A(g8892), .B(g10211), .Z(g10297) ) ;
AND2    gate9039  (.A(g8892), .B(g10214), .Z(g10298) ) ;
AND2    gate9040  (.A(g8892), .B(g10217), .Z(g10299) ) ;
AND2    gate9041  (.A(g8892), .B(g10220), .Z(g10300) ) ;
AND2    gate9042  (.A(g8892), .B(g10223), .Z(g10301) ) ;
AND2    gate9043  (.A(g10208), .B(g9076), .Z(g10303) ) ;
AND2    gate9044  (.A(g10211), .B(g9079), .Z(g10304) ) ;
AND2    gate9045  (.A(g10214), .B(g9082), .Z(g10306) ) ;
AND2    gate9046  (.A(g10217), .B(g9085), .Z(g10308) ) ;
AND2    gate9047  (.A(g10220), .B(g9094), .Z(g10312) ) ;
AND2    gate9048  (.A(g10223), .B(g9097), .Z(g10316) ) ;
AND2    gate9049  (.A(g10319), .B(g2135), .Z(g10365) ) ;
NOR2    gate9050  (.A(g10228), .B(g3507), .Z(g10362) ) ;
AND2    gate9051  (.A(g10362), .B(g3375), .Z(g10367) ) ;
AND2    gate9052  (.A(g10311), .B(g2135), .Z(g10442) ) ;
AND2    gate9053  (.A(g10315), .B(g2135), .Z(g10445) ) ;
NOR2    gate9054  (.A(g10329), .B(g3744), .Z(g10420) ) ;
AND2    gate9055  (.A(g10420), .B(g3345), .Z(g10449) ) ;
NOR2    gate9056  (.A(g10327), .B(g3744), .Z(g10364) ) ;
AND2    gate9057  (.A(g10364), .B(g3359), .Z(g10450) ) ;
AND2    gate9058  (.A(g10444), .B(g3365), .Z(g10451) ) ;
NOR2    gate9059  (.A(g10332), .B(g3507), .Z(g10435) ) ;
NOR2    gate9060  (.A(g10330), .B(g3507), .Z(g10433) ) ;
AND2    gate9061  (.A(g10431), .B(g3971), .Z(g10495) ) ;
NOR2    gate9062  (.A(g10326), .B(g3507), .Z(g10429) ) ;
AND2    gate9063  (.A(g10388), .B(g2135), .Z(g10503) ) ;
AND2    gate9064  (.A(g10389), .B(g2135), .Z(g10504) ) ;
AND2    gate9065  (.A(g10390), .B(g2135), .Z(g10506) ) ;
AND2    gate9066  (.A(g10391), .B(g2135), .Z(g10508) ) ;
AND2    gate9067  (.A(g10393), .B(g2135), .Z(g10510) ) ;
AND2    gate9068  (.A(g10395), .B(g2135), .Z(g10512) ) ;
OR2     gate9069  (.A(g4961), .B(g10367), .Z(g10489) ) ;
AND2    gate9070  (.A(g10489), .B(g4580), .Z(g10514) ) ;
NAND2   gate9071  (.A(g10438), .B(g6032), .Z(g10511) ) ;
NAND2   gate9072  (.A(g10436), .B(g6023), .Z(g10509) ) ;
NAND2   gate9073  (.A(g10434), .B(g5859), .Z(g10507) ) ;
AND3    gate9074  (.A(g10511), .B(g10509), .C(g10507), .Z(II16142) ) ;
NAND2   gate9075  (.A(g10432), .B(g5938), .Z(g10505) ) ;
NAND2   gate9076  (.A(g10430), .B(g5999), .Z(g10469) ) ;
NAND2   gate9077  (.A(g10285), .B(g5392), .Z(g10366) ) ;
NAND2   gate9078  (.A(g10363), .B(g5360), .Z(g10447) ) ;
NAND2   gate9079  (.A(g10443), .B(g5350), .Z(g10446) ) ;
AND3    gate9080  (.A(g10366), .B(g10447), .C(g10446), .Z(II16145) ) ;
NAND2   gate9081  (.A(g10441), .B(g5345), .Z(g10513) ) ;
NAND2   gate9082  (.A(g10360), .B(g6037), .Z(g10440) ) ;
AND3    gate9083  (.A(g10513), .B(g10440), .C(II16145), .Z(g10518) ) ;
AND2    gate9084  (.A(g10487), .B(g4575), .Z(g10560) ) ;
OR2     gate9085  (.A(g4951), .B(g10451), .Z(g10549) ) ;
AND2    gate9086  (.A(g10549), .B(g4583), .Z(g10561) ) ;
AND2    gate9087  (.A(g10531), .B(g9453), .Z(g10581) ) ;
AND2    gate9088  (.A(g10532), .B(g9473), .Z(g10582) ) ;
OR2     gate9089  (.A(g4942), .B(g10450), .Z(g10550) ) ;
AND2    gate9090  (.A(g10550), .B(g4347), .Z(g10595) ) ;
OR2     gate9091  (.A(g4933), .B(g10449), .Z(g10533) ) ;
AND2    gate9092  (.A(g10543), .B(g4525), .Z(g10622) ) ;
OR2     gate9093  (.A(g5511), .B(g10495), .Z(g10544) ) ;
AND2    gate9094  (.A(g10544), .B(g4536), .Z(g10623) ) ;
AND2    gate9095  (.A(g10545), .B(g4544), .Z(g10624) ) ;
AND2    gate9096  (.A(g10546), .B(g4552), .Z(g10625) ) ;
AND2    gate9097  (.A(g10547), .B(g4558), .Z(g10626) ) ;
AND2    gate9098  (.A(g10548), .B(g4564), .Z(g10627) ) ;
AND2    gate9099  (.A(g10600), .B(g3829), .Z(g10633) ) ;
AND2    gate9100  (.A(g10604), .B(g3829), .Z(g10634) ) ;
AND2    gate9101  (.A(g10608), .B(g3829), .Z(g10638) ) ;
AND2    gate9102  (.A(g10612), .B(g3829), .Z(g10642) ) ;
NOR2    gate9103  (.A(g10480), .B(g10521), .Z(g10594) ) ;
AND2    gate9104  (.A(g10594), .B(g3015), .Z(g10661) ) ;
AND2    gate9105  (.A(g8892), .B(g10571), .Z(g10662) ) ;
AND2    gate9106  (.A(g10575), .B(g9424), .Z(g10666) ) ;
AND2    gate9107  (.A(g10576), .B(g9427), .Z(g10667) ) ;
AND2    gate9108  (.A(g10577), .B(g9429), .Z(g10669) ) ;
AND2    gate9109  (.A(g10571), .B(g9091), .Z(g10670) ) ;
AND2    gate9110  (.A(g10578), .B(g9431), .Z(g10671) ) ;
AND2    gate9111  (.A(g10579), .B(g9449), .Z(g10672) ) ;
AND2    gate9112  (.A(g10580), .B(g9450), .Z(g10673) ) ;
OR2     gate9113  (.A(g10560), .B(g7368), .Z(g10564) ) ;
AND2    gate9114  (.A(g10564), .B(g3586), .Z(g10680) ) ;
OR2     gate9115  (.A(g10514), .B(g7378), .Z(g10567) ) ;
AND2    gate9116  (.A(g10567), .B(g3586), .Z(g10681) ) ;
AND2    gate9117  (.A(g10600), .B(g3863), .Z(g10682) ) ;
AND2    gate9118  (.A(g10604), .B(g3863), .Z(g10684) ) ;
AND2    gate9119  (.A(g10608), .B(g3863), .Z(g10685) ) ;
AND2    gate9120  (.A(g10612), .B(g3863), .Z(g10686) ) ;
AND2    gate9121  (.A(g10616), .B(g3863), .Z(g10690) ) ;
AND2    gate9122  (.A(g10620), .B(g10619), .Z(g10701) ) ;
AND2    gate9123  (.A(g10564), .B(g4840), .Z(g10705) ) ;
AND2    gate9124  (.A(g10567), .B(g4840), .Z(g10706) ) ;
NAND2   gate9125  (.A(II5316), .B(II5317), .Z(g2272) ) ;
AND2    gate9126  (.A(g2272), .B(g10630), .Z(g10715) ) ;
OR2     gate9127  (.A(g5052), .B(g10396), .Z(g10497) ) ;
AND2    gate9128  (.A(g10497), .B(g10675), .Z(g10716) ) ;
NAND3   gate9129  (.A(g2439), .B(g4806), .C(g4073), .Z(g5118) ) ;
NAND2   gate9130  (.A(II16331), .B(II16332), .Z(g10665) ) ;
AND3    gate9131  (.A(g5118), .B(g1850), .C(g10665), .Z(g10731) ) ;
OR2     gate9132  (.A(g10595), .B(g7674), .Z(g10658) ) ;
AND2    gate9133  (.A(g10658), .B(g4840), .Z(g10736) ) ;
AND2    gate9134  (.A(g10687), .B(g4840), .Z(g10737) ) ;
AND2    gate9135  (.A(g10692), .B(g4840), .Z(g10738) ) ;
AND2    gate9136  (.A(g10676), .B(g3368), .Z(g10739) ) ;
OR2     gate9137  (.A(g10622), .B(g7732), .Z(g10635) ) ;
AND2    gate9138  (.A(g10635), .B(g4013), .Z(g10741) ) ;
OR2     gate9139  (.A(g10561), .B(g7389), .Z(g10655) ) ;
AND2    gate9140  (.A(g10655), .B(g3586), .Z(g10742) ) ;
OR2     gate9141  (.A(g10623), .B(g7734), .Z(g10639) ) ;
AND2    gate9142  (.A(g10639), .B(g4013), .Z(g10743) ) ;
AND2    gate9143  (.A(g10658), .B(g3586), .Z(g10745) ) ;
OR2     gate9144  (.A(g10624), .B(g7736), .Z(g10643) ) ;
AND2    gate9145  (.A(g10643), .B(g4013), .Z(g10746) ) ;
AND2    gate9146  (.A(g10687), .B(g3586), .Z(g10750) ) ;
OR2     gate9147  (.A(g10625), .B(g7739), .Z(g10646) ) ;
AND2    gate9148  (.A(g10646), .B(g4013), .Z(g10751) ) ;
AND2    gate9149  (.A(g10692), .B(g3586), .Z(g10752) ) ;
OR2     gate9150  (.A(g10626), .B(g7741), .Z(g10649) ) ;
AND2    gate9151  (.A(g10649), .B(g4013), .Z(g10753) ) ;
OR2     gate9152  (.A(g10627), .B(g7743), .Z(g10652) ) ;
AND2    gate9153  (.A(g10652), .B(g4013), .Z(g10758) ) ;
AND2    gate9154  (.A(g10698), .B(g10697), .Z(g10759) ) ;
AND2    gate9155  (.A(g10695), .B(g10691), .Z(g10760) ) ;
AND2    gate9156  (.A(g10700), .B(g10699), .Z(g10761) ) ;
AND2    gate9157  (.A(g10635), .B(g4840), .Z(g10762) ) ;
AND2    gate9158  (.A(g10639), .B(g4840), .Z(g10763) ) ;
AND2    gate9159  (.A(g10643), .B(g4840), .Z(g10764) ) ;
AND2    gate9160  (.A(g10646), .B(g4840), .Z(g10766) ) ;
AND2    gate9161  (.A(g10649), .B(g4840), .Z(g10768) ) ;
AND2    gate9162  (.A(g10652), .B(g4840), .Z(g10769) ) ;
AND2    gate9163  (.A(g10655), .B(g4840), .Z(g10772) ) ;
OR2     gate9164  (.A(g5227), .B(g10674), .Z(g10733) ) ;
AND2    gate9165  (.A(g10733), .B(g3015), .Z(g10777) ) ;
AND2    gate9166  (.A(g1027), .B(g10729), .Z(g10778) ) ;
OR2     gate9167  (.A(g4952), .B(g10633), .Z(g10723) ) ;
OR2     gate9168  (.A(g4962), .B(g10634), .Z(g10725) ) ;
OR2     gate9169  (.A(g4969), .B(g10638), .Z(g10727) ) ;
OR2     gate9170  (.A(g4973), .B(g10642), .Z(g10728) ) ;
NOR2    gate9171  (.A(g8209), .B(g4811), .Z(g8303) ) ;
OR3     gate9172  (.A(g10600), .B(g10668), .C(II16427), .Z(g10744) ) ;
AND2    gate9173  (.A(g10744), .B(g3829), .Z(g10808) ) ;
AND2    gate9174  (.A(g10730), .B(g4545), .Z(g10818) ) ;
NAND2   gate9175  (.A(g10731), .B(g5034), .Z(g10853) ) ;
AND2    gate9176  (.A(g10853), .B(g3982), .Z(g10933) ) ;
NAND2   gate9177  (.A(II8663), .B(II8664), .Z(g5225) ) ;
AND2    gate9178  (.A(g5225), .B(g10827), .Z(g10946) ) ;
NAND2   gate9179  (.A(II5203), .B(II5204), .Z(g2223) ) ;
AND2    gate9180  (.A(g2223), .B(g10809), .Z(g10948) ) ;
NAND2   gate9181  (.A(II6137), .B(II6138), .Z(g2947) ) ;
AND2    gate9182  (.A(g2947), .B(g10809), .Z(g10949) ) ;
NAND2   gate9183  (.A(II6771), .B(II6772), .Z(g3625) ) ;
AND2    gate9184  (.A(g3625), .B(g10809), .Z(g10969) ) ;
AND2    gate9185  (.A(g10852), .B(g3390), .Z(g10970) ) ;
NOR2    gate9186  (.A(g10739), .B(g3903), .Z(g10849) ) ;
AND2    gate9187  (.A(g10849), .B(g3161), .Z(g10971) ) ;
NAND2   gate9188  (.A(II8514), .B(II8515), .Z(g5119) ) ;
AND2    gate9189  (.A(g5119), .B(g10827), .Z(g11005) ) ;
NAND2   gate9190  (.A(II8528), .B(II8529), .Z(g5125) ) ;
AND2    gate9191  (.A(g5125), .B(g10827), .Z(g11006) ) ;
NAND2   gate9192  (.A(II8544), .B(II8545), .Z(g5147) ) ;
AND2    gate9193  (.A(g5147), .B(g10827), .Z(g11007) ) ;
NAND2   gate9194  (.A(II8562), .B(II8563), .Z(g5171) ) ;
AND2    gate9195  (.A(g5171), .B(g10827), .Z(g11008) ) ;
NAND2   gate9196  (.A(II8576), .B(II8577), .Z(g5179) ) ;
AND2    gate9197  (.A(g5179), .B(g10827), .Z(g11009) ) ;
NAND2   gate9198  (.A(II8590), .B(II8591), .Z(g5187) ) ;
AND2    gate9199  (.A(g5187), .B(g10827), .Z(g11010) ) ;
AND2    gate9200  (.A(g1968), .B(g10809), .Z(g11011) ) ;
NAND2   gate9201  (.A(II8605), .B(II8606), .Z(g5196) ) ;
AND2    gate9202  (.A(g5196), .B(g10827), .Z(g11012) ) ;
NAND2   gate9203  (.A(II8625), .B(II8626), .Z(g5209) ) ;
AND2    gate9204  (.A(g5209), .B(g10827), .Z(g11013) ) ;
NAND2   gate9205  (.A(II8641), .B(II8642), .Z(g5217) ) ;
AND2    gate9206  (.A(g5217), .B(g10827), .Z(g11015) ) ;
AND2    gate9207  (.A(g7286), .B(g10974), .Z(g11018) ) ;
AND2    gate9208  (.A(g421), .B(g10974), .Z(g11019) ) ;
AND2    gate9209  (.A(g452), .B(g10974), .Z(g11020) ) ;
AND2    gate9210  (.A(g448), .B(g10974), .Z(g11021) ) ;
AND2    gate9211  (.A(g444), .B(g10974), .Z(g11022) ) ;
AND2    gate9212  (.A(g440), .B(g10974), .Z(g11023) ) ;
AND2    gate9213  (.A(g435), .B(g10974), .Z(g11024) ) ;
AND2    gate9214  (.A(g426), .B(g10974), .Z(g11025) ) ;
AND2    gate9215  (.A(g386), .B(g10974), .Z(g11026) ) ;
AND2    gate9216  (.A(g391), .B(g10974), .Z(g11027) ) ;
AND2    gate9217  (.A(g396), .B(g10974), .Z(g11028) ) ;
AND2    gate9218  (.A(g401), .B(g10974), .Z(g11029) ) ;
AND2    gate9219  (.A(g406), .B(g10974), .Z(g11030) ) ;
AND2    gate9220  (.A(g411), .B(g10974), .Z(g11031) ) ;
AND2    gate9221  (.A(g416), .B(g10974), .Z(g11032) ) ;
AND2    gate9222  (.A(g2008), .B(g10913), .Z(g11070) ) ;
AND2    gate9223  (.A(g312), .B(g10897), .Z(g11085) ) ;
AND2    gate9224  (.A(g829), .B(g10950), .Z(g11087) ) ;
AND2    gate9225  (.A(g833), .B(g10950), .Z(g11091) ) ;
AND2    gate9226  (.A(g837), .B(g10950), .Z(g11092) ) ;
AND2    gate9227  (.A(g841), .B(g10950), .Z(g11093) ) ;
AND2    gate9228  (.A(g374), .B(g10883), .Z(g11094) ) ;
AND2    gate9229  (.A(g845), .B(g10950), .Z(g11095) ) ;
AND2    gate9230  (.A(g378), .B(g10884), .Z(g11097) ) ;
AND2    gate9231  (.A(g849), .B(g10950), .Z(g11098) ) ;
AND2    gate9232  (.A(g382), .B(g10885), .Z(g11099) ) ;
AND2    gate9233  (.A(g853), .B(g10950), .Z(g11100) ) ;
AND2    gate9234  (.A(g857), .B(g10950), .Z(g11101) ) ;
AND2    gate9235  (.A(g861), .B(g10950), .Z(g11102) ) ;
NAND2   gate9236  (.A(II5264), .B(II5265), .Z(g2250) ) ;
AND2    gate9237  (.A(g2250), .B(g10937), .Z(g11103) ) ;
NAND2   gate9238  (.A(II6187), .B(II6188), .Z(g2963) ) ;
AND2    gate9239  (.A(g2963), .B(g10937), .Z(g11104) ) ;
NAND2   gate9240  (.A(II6806), .B(II6807), .Z(g3634) ) ;
AND2    gate9241  (.A(g3634), .B(g10937), .Z(g11105) ) ;
OR2     gate9242  (.A(g10778), .B(g10715), .Z(g10923) ) ;
AND2    gate9243  (.A(g10923), .B(g4567), .Z(g11143) ) ;
AND2    gate9244  (.A(g305), .B(g10926), .Z(g11144) ) ;
AND2    gate9245  (.A(g315), .B(g10927), .Z(g11145) ) ;
AND2    gate9246  (.A(g318), .B(g10928), .Z(g11146) ) ;
AND2    gate9247  (.A(g321), .B(g10929), .Z(g11147) ) ;
NAND2   gate9248  (.A(II5372), .B(II5373), .Z(g2321) ) ;
AND2    gate9249  (.A(g2321), .B(g10913), .Z(g11148) ) ;
AND2    gate9250  (.A(g324), .B(g10930), .Z(g11149) ) ;
NAND2   gate9251  (.A(II6288), .B(II6289), .Z(g3087) ) ;
AND2    gate9252  (.A(g3087), .B(g10913), .Z(g11150) ) ;
AND2    gate9253  (.A(g327), .B(g10931), .Z(g11151) ) ;
AND2    gate9254  (.A(g369), .B(g10903), .Z(g11152) ) ;
NAND2   gate9255  (.A(II6989), .B(II6990), .Z(g3771) ) ;
AND2    gate9256  (.A(g3771), .B(g10913), .Z(g11153) ) ;
AND2    gate9257  (.A(g330), .B(g10932), .Z(g11154) ) ;
AND2    gate9258  (.A(g333), .B(g10934), .Z(g11156) ) ;
AND2    gate9259  (.A(g309), .B(g10935), .Z(g11158) ) ;
AND2    gate9260  (.A(g1969), .B(g10937), .Z(g11161) ) ;
AND2    gate9261  (.A(g4889), .B(g11112), .Z(g11164) ) ;
AND2    gate9262  (.A(g476), .B(g11112), .Z(g11165) ) ;
AND2    gate9263  (.A(g542), .B(g11112), .Z(g11166) ) ;
AND2    gate9264  (.A(g538), .B(g11112), .Z(g11167) ) ;
AND2    gate9265  (.A(g534), .B(g11112), .Z(g11168) ) ;
AND2    gate9266  (.A(g530), .B(g11112), .Z(g11169) ) ;
AND2    gate9267  (.A(g525), .B(g11112), .Z(g11170) ) ;
AND2    gate9268  (.A(g481), .B(g11112), .Z(g11171) ) ;
AND2    gate9269  (.A(g486), .B(g11112), .Z(g11172) ) ;
AND2    gate9270  (.A(g491), .B(g11112), .Z(g11173) ) ;
AND2    gate9271  (.A(g496), .B(g11112), .Z(g11174) ) ;
AND2    gate9272  (.A(g501), .B(g11112), .Z(g11175) ) ;
AND2    gate9273  (.A(g506), .B(g11112), .Z(g11176) ) ;
AND2    gate9274  (.A(g511), .B(g11112), .Z(g11177) ) ;
AND2    gate9275  (.A(g516), .B(g11112), .Z(g11178) ) ;
AND2    gate9276  (.A(g5594), .B(g11059), .Z(g11186) ) ;
AND2    gate9277  (.A(g5597), .B(g11061), .Z(g11187) ) ;
AND2    gate9278  (.A(g5604), .B(g11063), .Z(g11188) ) ;
AND2    gate9279  (.A(g5616), .B(g11064), .Z(g11189) ) ;
AND2    gate9280  (.A(g5623), .B(g11065), .Z(g11190) ) ;
AND2    gate9281  (.A(g5628), .B(g11066), .Z(g11192) ) ;
AND2    gate9282  (.A(g5637), .B(g11067), .Z(g11194) ) ;
AND2    gate9283  (.A(g4912), .B(g11068), .Z(g11196) ) ;
AND2    gate9284  (.A(g4919), .B(g11069), .Z(g11198) ) ;
AND2    gate9285  (.A(g971), .B(g11083), .Z(g11204) ) ;
AND2    gate9286  (.A(g11074), .B(g9448), .Z(g11209) ) ;
AND2    gate9287  (.A(g11078), .B(g4515), .Z(g11210) ) ;
OR2     gate9288  (.A(g10933), .B(g5280), .Z(g11058) ) ;
AND2    gate9289  (.A(g11058), .B(g5534), .Z(g11211) ) ;
AND2    gate9290  (.A(g944), .B(g11155), .Z(g11212) ) ;
AND2    gate9291  (.A(g947), .B(g11157), .Z(g11213) ) ;
AND2    gate9292  (.A(g950), .B(g11159), .Z(g11214) ) ;
AND2    gate9293  (.A(g953), .B(g11160), .Z(g11215) ) ;
AND2    gate9294  (.A(g956), .B(g11162), .Z(g11216) ) ;
AND2    gate9295  (.A(g959), .B(g11053), .Z(g11218) ) ;
AND2    gate9296  (.A(g962), .B(g11054), .Z(g11220) ) ;
AND2    gate9297  (.A(g965), .B(g11055), .Z(g11222) ) ;
AND2    gate9298  (.A(g968), .B(g11056), .Z(g11224) ) ;
AND2    gate9299  (.A(g461), .B(g11057), .Z(g11226) ) ;
AND2    gate9300  (.A(g466), .B(g11060), .Z(g11228) ) ;
AND2    gate9301  (.A(g471), .B(g11062), .Z(g11230) ) ;
AND2    gate9302  (.A(g5424), .B(g11106), .Z(g11234) ) ;
AND2    gate9303  (.A(g5443), .B(g11107), .Z(g11235) ) ;
AND2    gate9304  (.A(g5469), .B(g11108), .Z(g11236) ) ;
AND2    gate9305  (.A(g5472), .B(g11109), .Z(g11237) ) ;
AND2    gate9306  (.A(g5474), .B(g11110), .Z(g11238) ) ;
AND2    gate9307  (.A(g5481), .B(g11111), .Z(g11240) ) ;
AND2    gate9308  (.A(g976), .B(g11071), .Z(g11248) ) ;
AND2    gate9309  (.A(g981), .B(g11072), .Z(g11253) ) ;
AND2    gate9310  (.A(g986), .B(g11073), .Z(g11254) ) ;
AND2    gate9311  (.A(g456), .B(g11075), .Z(g11255) ) ;
AND2    gate9312  (.A(g5624), .B(g11191), .Z(g11271) ) ;
AND2    gate9313  (.A(g5629), .B(g11193), .Z(g11272) ) ;
AND2    gate9314  (.A(g5638), .B(g11195), .Z(g11273) ) ;
AND2    gate9315  (.A(g4913), .B(g11197), .Z(g11274) ) ;
AND2    gate9316  (.A(g4920), .B(g11199), .Z(g11277) ) ;
AND2    gate9317  (.A(g4939), .B(g11200), .Z(g11279) ) ;
AND2    gate9318  (.A(g4948), .B(g11202), .Z(g11281) ) ;
AND2    gate9319  (.A(g4958), .B(g11203), .Z(g11282) ) ;
AND2    gate9320  (.A(g4966), .B(g11205), .Z(g11283) ) ;
OR2     gate9321  (.A(g11094), .B(g10948), .Z(g11246) ) ;
OR2     gate9322  (.A(g11097), .B(g10949), .Z(g11247) ) ;
OR2     gate9323  (.A(g11099), .B(g10969), .Z(g11252) ) ;
AND2    gate9324  (.A(g5475), .B(g11239), .Z(g11295) ) ;
AND2    gate9325  (.A(g5482), .B(g11241), .Z(g11296) ) ;
AND2    gate9326  (.A(g5490), .B(g11242), .Z(g11297) ) ;
AND2    gate9327  (.A(g5498), .B(g11243), .Z(g11299) ) ;
AND2    gate9328  (.A(g5508), .B(g11244), .Z(g11302) ) ;
AND2    gate9329  (.A(g5520), .B(g11245), .Z(g11304) ) ;
OR2     gate9330  (.A(g11152), .B(g11011), .Z(g11201) ) ;
OR2     gate9331  (.A(g11255), .B(g11161), .Z(g11285) ) ;
OR2     gate9332  (.A(g11204), .B(g11070), .Z(g11288) ) ;
OR2     gate9333  (.A(g11226), .B(g11103), .Z(g11316) ) ;
OR2     gate9334  (.A(g11228), .B(g11104), .Z(g11318) ) ;
OR2     gate9335  (.A(g11230), .B(g11105), .Z(g11321) ) ;
AND2    gate9336  (.A(g11284), .B(g3629), .Z(g11387) ) ;
OR2     gate9337  (.A(g11248), .B(g11148), .Z(g11275) ) ;
OR2     gate9338  (.A(g11253), .B(g11150), .Z(g11278) ) ;
OR2     gate9339  (.A(g11254), .B(g11153), .Z(g11280) ) ;
AND2    gate9340  (.A(g11339), .B(g5949), .Z(g11407) ) ;
AND2    gate9341  (.A(g11354), .B(g10679), .Z(g11413) ) ;
AND2    gate9342  (.A(g11435), .B(g5446), .Z(g11455) ) ;
AND3    gate9343  (.A(g3765), .B(g3517), .C(g11422), .Z(g11456) ) ;
AND2    gate9344  (.A(g11426), .B(g5446), .Z(g11458) ) ;
AND2    gate9345  (.A(g11427), .B(g5446), .Z(g11459) ) ;
AND2    gate9346  (.A(g11428), .B(g5446), .Z(g11460) ) ;
AND2    gate9347  (.A(g11429), .B(g5446), .Z(g11461) ) ;
AND2    gate9348  (.A(g11431), .B(g5446), .Z(g11462) ) ;
AND2    gate9349  (.A(g11432), .B(g5446), .Z(g11463) ) ;
AND2    gate9350  (.A(g11433), .B(g5446), .Z(g11464) ) ;
AND2    gate9351  (.A(g11434), .B(g5446), .Z(g11465) ) ;
NOR2    gate9352  (.A(g11456), .B(g4567), .Z(g11480) ) ;
NAND2   gate9353  (.A(II17493), .B(II17494), .Z(g11491) ) ;
AND2    gate9354  (.A(g11515), .B(g10584), .Z(g11544) ) ;
NAND2   gate9355  (.A(II17568), .B(II17569), .Z(g11538) ) ;
AND2    gate9356  (.A(g11538), .B(g4013), .Z(g11551) ) ;
AND2    gate9357  (.A(g2677), .B(g11519), .Z(g11552) ) ;
AND2    gate9358  (.A(g2683), .B(g11519), .Z(g11553) ) ;
AND2    gate9359  (.A(g2689), .B(g11519), .Z(g11554) ) ;
AND2    gate9360  (.A(g2695), .B(g11519), .Z(g11555) ) ;
AND2    gate9361  (.A(g2701), .B(g11519), .Z(g11556) ) ;
AND2    gate9362  (.A(g2707), .B(g11519), .Z(g11557) ) ;
AND2    gate9363  (.A(g2713), .B(g11519), .Z(g11558) ) ;
AND2    gate9364  (.A(g2719), .B(g11519), .Z(g11559) ) ;
AND2    gate9365  (.A(g2765), .B(g11519), .Z(g11560) ) ;
AND2    gate9366  (.A(g2018), .B(g11561), .Z(g11571) ) ;
AND2    gate9367  (.A(g1308), .B(g11539), .Z(g11581) ) ;
AND2    gate9368  (.A(g1311), .B(g11540), .Z(g11582) ) ;
AND2    gate9369  (.A(g1314), .B(g11541), .Z(g11583) ) ;
AND2    gate9370  (.A(g1318), .B(g11542), .Z(g11584) ) ;
AND2    gate9371  (.A(g1321), .B(g11543), .Z(g11585) ) ;
AND2    gate9372  (.A(g1324), .B(g11545), .Z(g11586) ) ;
AND2    gate9373  (.A(g1327), .B(g11546), .Z(g11587) ) ;
AND2    gate9374  (.A(g1330), .B(g11547), .Z(g11588) ) ;
AND2    gate9375  (.A(g1333), .B(g11548), .Z(g11589) ) ;
NAND2   gate9376  (.A(II5324), .B(II5325), .Z(g2274) ) ;
AND2    gate9377  (.A(g2274), .B(g11561), .Z(g11590) ) ;
NAND2   gate9378  (.A(II6225), .B(II6226), .Z(g2988) ) ;
AND2    gate9379  (.A(g2988), .B(g11561), .Z(g11591) ) ;
NAND2   gate9380  (.A(II6880), .B(II6881), .Z(g3717) ) ;
AND2    gate9381  (.A(g3717), .B(g11561), .Z(g11592) ) ;
AND2    gate9382  (.A(g1336), .B(g11575), .Z(g11595) ) ;
AND2    gate9383  (.A(g11576), .B(g5446), .Z(g11597) ) ;
AND2    gate9384  (.A(g1341), .B(g11572), .Z(g11599) ) ;
AND2    gate9385  (.A(g1346), .B(g11573), .Z(g11600) ) ;
AND2    gate9386  (.A(g1351), .B(g11574), .Z(g11601) ) ;
OR2     gate9387  (.A(g11595), .B(g11571), .Z(g11624) ) ;
AND2    gate9388  (.A(g11626), .B(g5446), .Z(g11637) ) ;
OR2     gate9389  (.A(g11599), .B(g11590), .Z(g11612) ) ;
OR2     gate9390  (.A(g11600), .B(g11591), .Z(g11613) ) ;
OR2     gate9391  (.A(g11601), .B(g11592), .Z(g11615) ) ;
OR4     gate9392  (.A(g1145), .B(g1141), .C(g1137), .D(g1133), .Z(II5351) ) ;
OR4     gate9393  (.A(g1129), .B(g1125), .C(g1121), .D(g1117), .Z(II5352) ) ;
OR2     gate9394  (.A(II5351), .B(II5352), .Z(g2305) ) ;
OR4     gate9395  (.A(g1265), .B(g1260), .C(g1255), .D(g1250), .Z(II5357) ) ;
OR4     gate9396  (.A(g1245), .B(g1240), .C(g1235), .D(g1275), .Z(II5358) ) ;
OR2     gate9397  (.A(II5357), .B(II5358), .Z(g2309) ) ;
OR4     gate9398  (.A(g1149), .B(g1153), .C(g1157), .D(g1160), .Z(II5363) ) ;
OR4     gate9399  (.A(g1163), .B(g1166), .C(g1113), .D(II5363), .Z(g2315) ) ;
OR4     gate9400  (.A(g1280), .B(g1284), .C(g1292), .D(g1296), .Z(II5366) ) ;
OR4     gate9401  (.A(g1300), .B(g1304), .C(g1270), .D(II5366), .Z(g2316) ) ;
OR4     gate9402  (.A(g1403), .B(g1407), .C(g1411), .D(g1415), .Z(g2353) ) ;
OR4     gate9403  (.A(g416), .B(g411), .C(g406), .D(g401), .Z(II5570) ) ;
OR4     gate9404  (.A(g396), .B(g391), .C(g386), .D(g426), .Z(II5571) ) ;
OR2     gate9405  (.A(II5570), .B(II5571), .Z(g2499) ) ;
OR4     gate9406  (.A(g431), .B(g435), .C(g440), .D(g444), .Z(II5576) ) ;
OR4     gate9407  (.A(g448), .B(g452), .C(g421), .D(II5576), .Z(g2501) ) ;
OR4     gate9408  (.A(g516), .B(g511), .C(g506), .D(g501), .Z(II5599) ) ;
OR4     gate9409  (.A(g496), .B(g491), .C(g486), .D(g481), .Z(II5600) ) ;
OR2     gate9410  (.A(II5599), .B(II5600), .Z(g2514) ) ;
OR4     gate9411  (.A(g521), .B(g525), .C(g530), .D(g534), .Z(II5626) ) ;
OR4     gate9412  (.A(g538), .B(g542), .C(g476), .D(II5626), .Z(g2521) ) ;
OR3     gate9413  (.A(g845), .B(g841), .C(g837), .Z(II5629) ) ;
OR3     gate9414  (.A(g833), .B(g829), .C(II5629), .Z(g2522) ) ;
OR4     gate9415  (.A(g861), .B(g857), .C(g853), .D(g849), .Z(g2528) ) ;
OR3     gate9416  (.A(g1499), .B(g1486), .C(g1482), .Z(II5649) ) ;
OR3     gate9417  (.A(g1466), .B(g1458), .C(II5649), .Z(g2538) ) ;
NAND2   gate9418  (.A(II5006), .B(II5007), .Z(g2111) ) ;
NAND2   gate9419  (.A(II4996), .B(II4997), .Z(g2109) ) ;
NAND2   gate9420  (.A(II4979), .B(II4980), .Z(g2106) ) ;
NAND2   gate9421  (.A(II4965), .B(II4966), .Z(g2104) ) ;
OR4     gate9422  (.A(g2111), .B(g2109), .C(g2106), .D(g2104), .Z(II5804) ) ;
NAND2   gate9423  (.A(II4955), .B(II4956), .Z(g2102) ) ;
NAND2   gate9424  (.A(II4942), .B(II4943), .Z(g2099) ) ;
NAND2   gate9425  (.A(II4929), .B(II4930), .Z(g2096) ) ;
NAND2   gate9426  (.A(II4911), .B(II4912), .Z(g2088) ) ;
OR4     gate9427  (.A(g2102), .B(g2099), .C(g2096), .D(g2088), .Z(II5805) ) ;
NAND2   gate9428  (.A(II5539), .B(II5540), .Z(g2445) ) ;
NAND2   gate9429  (.A(II5529), .B(II5530), .Z(g2437) ) ;
NAND2   gate9430  (.A(II5517), .B(II5518), .Z(g2433) ) ;
NAND2   gate9431  (.A(II5501), .B(II5502), .Z(g2419) ) ;
OR4     gate9432  (.A(g2445), .B(g2437), .C(g2433), .D(g2419), .Z(II6350) ) ;
NAND2   gate9433  (.A(II5485), .B(II5486), .Z(g2405) ) ;
NAND2   gate9434  (.A(II5469), .B(II5470), .Z(g2389) ) ;
NAND2   gate9435  (.A(II5460), .B(II5461), .Z(g2380) ) ;
NAND2   gate9436  (.A(II5450), .B(II5451), .Z(g2372) ) ;
OR4     gate9437  (.A(g2405), .B(g2389), .C(g2380), .D(g2372), .Z(II6351) ) ;
NOR2    gate9438  (.A(g2521), .B(g2514), .Z(g3118) ) ;
NAND2   gate9439  (.A(II5136), .B(II5137), .Z(g2180) ) ;
NOR2    gate9440  (.A(g2316), .B(g2309), .Z(g2863) ) ;
NAND2   gate9441  (.A(II5612), .B(II5613), .Z(g2516) ) ;
NOR2    gate9442  (.A(g2501), .B(g2499), .Z(g3107) ) ;
NAND2   gate9443  (.A(II5105), .B(II5106), .Z(g2167) ) ;
NOR2    gate9444  (.A(g2315), .B(g2305), .Z(g2862) ) ;
NAND2   gate9445  (.A(II5605), .B(II5606), .Z(g2515) ) ;
OR2     gate9446  (.A(g2862), .B(g2515), .Z(g4052) ) ;
OR2     gate9447  (.A(g4581), .B(g4584), .Z(g4997) ) ;
NAND2   gate9448  (.A(g3807), .B(g3071), .Z(g4476) ) ;
OR2     gate9449  (.A(g4389), .B(g4397), .Z(g5555) ) ;
NAND2   gate9450  (.A(g4073), .B(g3247), .Z(g4675) ) ;
NOR2    gate9451  (.A(g2047), .B(g4401), .Z(g5186) ) ;
OR2     gate9452  (.A(g5172), .B(g5180), .Z(g6122) ) ;
OR2     gate9453  (.A(g5181), .B(g5188), .Z(g6124) ) ;
NOR2    gate9454  (.A(g2112), .B(g4921), .Z(g5780) ) ;
OR2     gate9455  (.A(g6463), .B(g5471), .Z(g6899) ) ;
OR2     gate9456  (.A(g7687), .B(g7182), .Z(g7963) ) ;
OR2     gate9457  (.A(g7884), .B(g6872), .Z(g8148) ) ;
OR2     gate9458  (.A(g7888), .B(g6875), .Z(g8153) ) ;
OR2     gate9459  (.A(g7891), .B(g6879), .Z(g8154) ) ;
OR2     gate9460  (.A(g7965), .B(g7623), .Z(g8157) ) ;
OR2     gate9461  (.A(g7893), .B(g6883), .Z(g8158) ) ;
OR2     gate9462  (.A(g7895), .B(g6886), .Z(g8159) ) ;
OR2     gate9463  (.A(g8005), .B(g7185), .Z(g8161) ) ;
OR2     gate9464  (.A(g7898), .B(g6889), .Z(g8162) ) ;
OR2     gate9465  (.A(g8010), .B(g7704), .Z(g8247) ) ;
OR2     gate9466  (.A(g8014), .B(g7707), .Z(g8248) ) ;
OR2     gate9467  (.A(g8018), .B(g7710), .Z(g8249) ) ;
OR2     gate9468  (.A(g8023), .B(g7718), .Z(g8253) ) ;
OR2     gate9469  (.A(g8028), .B(g7719), .Z(g8259) ) ;
OR2     gate9470  (.A(g7970), .B(g7625), .Z(g8262) ) ;
OR2     gate9471  (.A(g8032), .B(g7720), .Z(g8263) ) ;
OR2     gate9472  (.A(g8136), .B(g6891), .Z(g8322) ) ;
OR2     gate9473  (.A(g8246), .B(g7721), .Z(g8417) ) ;
OR2     gate9474  (.A(g8778), .B(g8693), .Z(g8823) ) ;
OR3     gate9475  (.A(g8995), .B(g9205), .C(g9192), .Z(II14582) ) ;
OR3     gate9476  (.A(g8995), .B(g9205), .C(g9192), .Z(II14585) ) ;
OR2     gate9477  (.A(g9205), .B(g9192), .Z(g9363) ) ;
OR3     gate9478  (.A(g8995), .B(g9205), .C(g9192), .Z(II14596) ) ;
OR2     gate9479  (.A(g9240), .B(g9223), .Z(g9388) ) ;
OR3     gate9480  (.A(g8995), .B(g9205), .C(g9192), .Z(II14602) ) ;
OR3     gate9481  (.A(g8995), .B(g9205), .C(g9192), .Z(II14607) ) ;
OR3     gate9482  (.A(g9151), .B(g9125), .C(g9111), .Z(g9509) ) ;
OR2     gate9483  (.A(g9125), .B(g9111), .Z(g9510) ) ;
OR3     gate9484  (.A(g9151), .B(g9125), .C(g9111), .Z(g9511) ) ;
OR2     gate9485  (.A(g9173), .B(g9151), .Z(g9515) ) ;
OR3     gate9486  (.A(g9151), .B(g9125), .C(g9111), .Z(g9528) ) ;
OR3     gate9487  (.A(g8995), .B(g9205), .C(g9192), .Z(II14751) ) ;
OR3     gate9488  (.A(g8995), .B(g9205), .C(g9192), .Z(II14776) ) ;
OR3     gate9489  (.A(g8995), .B(g9205), .C(g9192), .Z(II14779) ) ;
OR3     gate9490  (.A(g9597), .B(g9604), .C(g9582), .Z(II14822) ) ;
NOR4    gate9491  (.A(g9125), .B(g9111), .C(g9173), .D(g9151), .Z(g9606) ) ;
OR3     gate9492  (.A(g9603), .B(g9614), .C(g9584), .Z(II14827) ) ;
NOR4    gate9493  (.A(g9125), .B(g9111), .C(g9173), .D(g9151), .Z(g9667) ) ;
OR3     gate9494  (.A(g9613), .B(g9622), .C(g9586), .Z(II14831) ) ;
NOR4    gate9495  (.A(g9125), .B(g9111), .C(g9173), .D(g9151), .Z(g9647) ) ;
OR3     gate9496  (.A(g9621), .B(g9645), .C(g9588), .Z(II14835) ) ;
NOR4    gate9497  (.A(g9125), .B(g9111), .C(g9173), .D(g9151), .Z(g9605) ) ;
NOR2    gate9498  (.A(g9125), .B(g9151), .Z(g9591) ) ;
NOR2    gate9499  (.A(g9125), .B(g9151), .Z(g9646) ) ;
NOR3    gate9500  (.A(g9125), .B(g9173), .C(g9151), .Z(g9589) ) ;
NOR2    gate9501  (.A(g9125), .B(g9173), .Z(g9654) ) ;
OR4     gate9502  (.A(g9583), .B(g9593), .C(g9601), .D(g9596), .Z(II14855) ) ;
NOR4    gate9503  (.A(g9010), .B(g9240), .C(g9223), .D(II14607), .Z(g9410) ) ;
OR4     gate9504  (.A(g9585), .B(g9595), .C(g9610), .D(g9602), .Z(II14858) ) ;
NOR4    gate9505  (.A(g9010), .B(g9240), .C(g9223), .D(II14602), .Z(g9391) ) ;
NOR2    gate9506  (.A(g9052), .B(g9030), .Z(g9615) ) ;
OR3     gate9507  (.A(g9587), .B(g9600), .C(g9611), .Z(II14862) ) ;
NOR4    gate9508  (.A(g9010), .B(g9240), .C(g9223), .D(II14751), .Z(g9616) ) ;
NOR2    gate9509  (.A(g9052), .B(g9030), .Z(g9489) ) ;
OR3     gate9510  (.A(g9590), .B(g9609), .C(g9619), .Z(II14866) ) ;
NOR4    gate9511  (.A(g9010), .B(g9240), .C(g9223), .D(II14585), .Z(g9362) ) ;
NOR2    gate9512  (.A(g9052), .B(g9030), .Z(g9426) ) ;
NOR4    gate9513  (.A(g9010), .B(g9240), .C(g9223), .D(II14779), .Z(g9656) ) ;
NOR2    gate9514  (.A(g9052), .B(g9030), .Z(g9423) ) ;
NOR4    gate9515  (.A(g9010), .B(g9240), .C(g9223), .D(II14596), .Z(g9387) ) ;
NOR2    gate9516  (.A(g9052), .B(g9030), .Z(g9421) ) ;
NOR4    gate9517  (.A(g9010), .B(g9240), .C(g9223), .D(II14582), .Z(g9361) ) ;
NOR2    gate9518  (.A(g9052), .B(g9030), .Z(g9416) ) ;
NOR4    gate9519  (.A(g9010), .B(g9240), .C(g9223), .D(II14776), .Z(g9655) ) ;
NOR2    gate9520  (.A(g9052), .B(g9030), .Z(g9506) ) ;
NOR3    gate9521  (.A(g9454), .B(g9274), .C(g9292), .Z(g9750) ) ;
NOR3    gate9522  (.A(g9454), .B(g9274), .C(g9292), .Z(g9758) ) ;
OR4     gate9523  (.A(g7853), .B(g9804), .C(g9624), .D(g9785), .Z(II15033) ) ;
OR4     gate9524  (.A(g7853), .B(g9809), .C(g9624), .D(g9785), .Z(II15039) ) ;
OR4     gate9525  (.A(g7853), .B(g9686), .C(g9624), .D(g9785), .Z(II15042) ) ;
OR4     gate9526  (.A(g7853), .B(g9676), .C(g9624), .D(g9785), .Z(II15045) ) ;
OR4     gate9527  (.A(g7853), .B(g9683), .C(g9624), .D(g9785), .Z(II15048) ) ;
OR4     gate9528  (.A(g7853), .B(g9673), .C(g9624), .D(g9785), .Z(II15051) ) ;
OR4     gate9529  (.A(g7853), .B(g9782), .C(g9624), .D(g9785), .Z(II15054) ) ;
OR4     gate9530  (.A(g7853), .B(g9680), .C(g9624), .D(g9785), .Z(II15057) ) ;
NOR3    gate9531  (.A(g9454), .B(g9274), .C(g9292), .Z(g9746) ) ;
NOR3    gate9532  (.A(g9454), .B(g9274), .C(g9292), .Z(g9759) ) ;
NOR3    gate9533  (.A(g9454), .B(g9274), .C(g9292), .Z(g9757) ) ;
NOR2    gate9534  (.A(g9392), .B(g9367), .Z(g9779) ) ;
NOR2    gate9535  (.A(g9392), .B(g9367), .Z(g9803) ) ;
NOR2    gate9536  (.A(g9392), .B(g9367), .Z(g9817) ) ;
NOR2    gate9537  (.A(g9392), .B(g9367), .Z(g9669) ) ;
NOR2    gate9538  (.A(g9392), .B(g9367), .Z(g9781) ) ;
NOR2    gate9539  (.A(g9392), .B(g9367), .Z(g9808) ) ;
NOR2    gate9540  (.A(g9392), .B(g9367), .Z(g9815) ) ;
NOR2    gate9541  (.A(g9392), .B(g9367), .Z(g9776) ) ;
OR4     gate9542  (.A(g8175), .B(g9909), .C(g9896), .D(g9835), .Z(II15171) ) ;
NOR4    gate9543  (.A(g9519), .B(g9536), .C(g9579), .D(II15033), .Z(g9874) ) ;
OR4     gate9544  (.A(g9843), .B(g9959), .C(g9861), .D(g9874), .Z(II15172) ) ;
OR4     gate9545  (.A(g8176), .B(g9910), .C(g9897), .D(g9836), .Z(II15176) ) ;
NOR4    gate9546  (.A(g9522), .B(g9536), .C(g9576), .D(II15039), .Z(g9876) ) ;
OR4     gate9547  (.A(g9844), .B(g9960), .C(g9863), .D(g9876), .Z(II15177) ) ;
OR4     gate9548  (.A(g8167), .B(g9903), .C(g9932), .D(g9828), .Z(II15199) ) ;
NOR4    gate9549  (.A(g9751), .B(g9536), .C(g9557), .D(II15051), .Z(g9880) ) ;
OR4     gate9550  (.A(g9837), .B(g9962), .C(g9848), .D(g9880), .Z(II15200) ) ;
OR4     gate9551  (.A(g8168), .B(g9904), .C(g9933), .D(g9829), .Z(II15204) ) ;
NOR4    gate9552  (.A(g9754), .B(g9536), .C(g9560), .D(II15045), .Z(g9878) ) ;
OR4     gate9553  (.A(g9838), .B(g9963), .C(g9850), .D(g9878), .Z(II15205) ) ;
OR4     gate9554  (.A(g8169), .B(g9905), .C(g9934), .D(g9830), .Z(II15209) ) ;
NOR4    gate9555  (.A(g9742), .B(g9536), .C(g9563), .D(II15057), .Z(g9882) ) ;
OR4     gate9556  (.A(g9839), .B(g9964), .C(g9852), .D(g9882), .Z(II15210) ) ;
OR4     gate9557  (.A(g8170), .B(g9906), .C(g9935), .D(g9831), .Z(II15214) ) ;
NOR4    gate9558  (.A(g9747), .B(g9536), .C(g9566), .D(II15048), .Z(g9879) ) ;
OR4     gate9559  (.A(g9840), .B(g9965), .C(g9854), .D(g9879), .Z(II15215) ) ;
OR4     gate9560  (.A(g8172), .B(g9907), .C(g9936), .D(g9833), .Z(II15219) ) ;
NOR4    gate9561  (.A(g9512), .B(g9536), .C(g9569), .D(II15042), .Z(g9877) ) ;
OR4     gate9562  (.A(g9841), .B(g9966), .C(g9857), .D(g9877), .Z(II15220) ) ;
OR4     gate9563  (.A(g8174), .B(g9908), .C(g9937), .D(g9834), .Z(II15224) ) ;
NOR4    gate9564  (.A(g9516), .B(g9536), .C(g9573), .D(II15054), .Z(g9881) ) ;
OR4     gate9565  (.A(g9842), .B(g9967), .C(g9859), .D(g9881), .Z(II15225) ) ;
NOR2    gate9566  (.A(g10247), .B(g3113), .Z(g10291) ) ;
NOR2    gate9567  (.A(g10323), .B(g3113), .Z(g10376) ) ;
NAND2   gate9568  (.A(II15879), .B(II15880), .Z(g10386) ) ;
NAND2   gate9569  (.A(II15871), .B(II15872), .Z(g10384) ) ;
NAND2   gate9570  (.A(II16038), .B(II16039), .Z(g10476) ) ;
NAND2   gate9571  (.A(II16024), .B(II16025), .Z(g10474) ) ;
OR4     gate9572  (.A(g10386), .B(g10384), .C(g10476), .D(g10474), .Z(II16148) ) ;
NAND2   gate9573  (.A(II16016), .B(II16017), .Z(g10472) ) ;
NAND2   gate9574  (.A(II16008), .B(II16009), .Z(g10470) ) ;
NAND2   gate9575  (.A(II16000), .B(II16001), .Z(g10468) ) ;
NAND2   gate9576  (.A(II15993), .B(II15994), .Z(g10467) ) ;
OR4     gate9577  (.A(g10472), .B(g10470), .C(g10468), .D(g10467), .Z(II16149) ) ;
OR2     gate9578  (.A(II16148), .B(II16149), .Z(g10521) ) ;
NAND2   gate9579  (.A(II15899), .B(II15900), .Z(g10394) ) ;
NAND2   gate9580  (.A(II15891), .B(II15892), .Z(g10392) ) ;
NAND2   gate9581  (.A(II16080), .B(II16081), .Z(g10482) ) ;
NAND2   gate9582  (.A(II16073), .B(II16074), .Z(g10481) ) ;
OR4     gate9583  (.A(g10394), .B(g10392), .C(g10482), .D(g10481), .Z(II16160) ) ;
NAND2   gate9584  (.A(II16059), .B(II16060), .Z(g10479) ) ;
NAND2   gate9585  (.A(II16052), .B(II16053), .Z(g10478) ) ;
NAND2   gate9586  (.A(II16045), .B(II16046), .Z(g10477) ) ;
NAND2   gate9587  (.A(II16031), .B(II16032), .Z(g10475) ) ;
OR4     gate9588  (.A(g10479), .B(g10478), .C(g10477), .D(g10475), .Z(II16161) ) ;
OR2     gate9589  (.A(II16160), .B(II16161), .Z(g10529) ) ;
NOR2    gate9590  (.A(g10483), .B(g10529), .Z(g10562) ) ;
NAND2   gate9591  (.A(II8677), .B(II8678), .Z(g5227) ) ;
OR3     gate9592  (.A(g10683), .B(g10608), .C(g10604), .Z(II16427) ) ;
OR2     gate9593  (.A(g10759), .B(g10760), .Z(g10805) ) ;
OR2     gate9594  (.A(g10701), .B(g10761), .Z(g10807) ) ;
NAND2   gate9595  (.A(g386), .B(g318), .Z(II4910) ) ;
NAND2   gate9596  (.A(g386), .B(II4910), .Z(II4911) ) ;
NAND2   gate9597  (.A(g318), .B(II4910), .Z(II4912) ) ;
NAND2   gate9598  (.A(g391), .B(g321), .Z(II4928) ) ;
NAND2   gate9599  (.A(g391), .B(II4928), .Z(II4929) ) ;
NAND2   gate9600  (.A(g321), .B(II4928), .Z(II4930) ) ;
NAND2   gate9601  (.A(g396), .B(g324), .Z(II4941) ) ;
NAND2   gate9602  (.A(g396), .B(II4941), .Z(II4942) ) ;
NAND2   gate9603  (.A(g324), .B(II4941), .Z(II4943) ) ;
NAND2   gate9604  (.A(g401), .B(g327), .Z(II4954) ) ;
NAND2   gate9605  (.A(g401), .B(II4954), .Z(II4955) ) ;
NAND2   gate9606  (.A(g327), .B(II4954), .Z(II4956) ) ;
NAND2   gate9607  (.A(g406), .B(g330), .Z(II4964) ) ;
NAND2   gate9608  (.A(g406), .B(II4964), .Z(II4965) ) ;
NAND2   gate9609  (.A(g330), .B(II4964), .Z(II4966) ) ;
NAND2   gate9610  (.A(g991), .B(g995), .Z(II4971) ) ;
NAND2   gate9611  (.A(g991), .B(II4971), .Z(II4972) ) ;
NAND2   gate9612  (.A(g995), .B(II4971), .Z(II4973) ) ;
NAND2   gate9613  (.A(II4972), .B(II4973), .Z(g2105) ) ;
NAND2   gate9614  (.A(g411), .B(g333), .Z(II4978) ) ;
NAND2   gate9615  (.A(g411), .B(II4978), .Z(II4979) ) ;
NAND2   gate9616  (.A(g333), .B(II4978), .Z(II4980) ) ;
NAND2   gate9617  (.A(g999), .B(g1003), .Z(II4985) ) ;
NAND2   gate9618  (.A(g999), .B(II4985), .Z(II4986) ) ;
NAND2   gate9619  (.A(g1003), .B(II4985), .Z(II4987) ) ;
NAND2   gate9620  (.A(II4986), .B(II4987), .Z(g2107) ) ;
NAND2   gate9621  (.A(g416), .B(g309), .Z(II4995) ) ;
NAND2   gate9622  (.A(g416), .B(II4995), .Z(II4996) ) ;
NAND2   gate9623  (.A(g309), .B(II4995), .Z(II4997) ) ;
NAND2   gate9624  (.A(g421), .B(g312), .Z(II5005) ) ;
NAND2   gate9625  (.A(g421), .B(II5005), .Z(II5006) ) ;
NAND2   gate9626  (.A(g312), .B(II5005), .Z(II5007) ) ;
NAND2   gate9627  (.A(g1007), .B(g1011), .Z(II5013) ) ;
NAND2   gate9628  (.A(g1007), .B(II5013), .Z(II5014) ) ;
NAND2   gate9629  (.A(g1011), .B(II5013), .Z(II5015) ) ;
NAND2   gate9630  (.A(II5014), .B(II5015), .Z(g2115) ) ;
NAND2   gate9631  (.A(g995), .B(g1275), .Z(II5023) ) ;
NAND2   gate9632  (.A(g995), .B(II5023), .Z(II5024) ) ;
NAND2   gate9633  (.A(g1275), .B(II5023), .Z(II5025) ) ;
NAND2   gate9634  (.A(g1015), .B(g1019), .Z(II5034) ) ;
NAND2   gate9635  (.A(g1015), .B(II5034), .Z(II5035) ) ;
NAND2   gate9636  (.A(g1019), .B(II5034), .Z(II5036) ) ;
NAND2   gate9637  (.A(II5035), .B(II5036), .Z(g2120) ) ;
NAND2   gate9638  (.A(g431), .B(g435), .Z(II5104) ) ;
NAND2   gate9639  (.A(g431), .B(II5104), .Z(II5105) ) ;
NAND2   gate9640  (.A(g435), .B(II5104), .Z(II5106) ) ;
NAND2   gate9641  (.A(g1386), .B(g1389), .Z(II5126) ) ;
NAND2   gate9642  (.A(g1386), .B(II5126), .Z(II5127) ) ;
NAND2   gate9643  (.A(g1389), .B(II5126), .Z(II5128) ) ;
NAND2   gate9644  (.A(II5127), .B(II5128), .Z(g2177) ) ;
NAND2   gate9645  (.A(g521), .B(g525), .Z(II5135) ) ;
NAND2   gate9646  (.A(g521), .B(II5135), .Z(II5136) ) ;
NAND2   gate9647  (.A(g525), .B(II5135), .Z(II5137) ) ;
NAND2   gate9648  (.A(g1508), .B(g1499), .Z(II5164) ) ;
NAND2   gate9649  (.A(g1508), .B(II5164), .Z(II5165) ) ;
NAND2   gate9650  (.A(g1499), .B(II5164), .Z(II5166) ) ;
NAND2   gate9651  (.A(II5165), .B(II5166), .Z(g2205) ) ;
NAND2   gate9652  (.A(g1415), .B(g1515), .Z(II5184) ) ;
NAND2   gate9653  (.A(g1415), .B(II5184), .Z(II5185) ) ;
NAND2   gate9654  (.A(g1515), .B(II5184), .Z(II5186) ) ;
NAND2   gate9655  (.A(II5185), .B(II5186), .Z(g2215) ) ;
NAND2   gate9656  (.A(g369), .B(g374), .Z(II5202) ) ;
NAND2   gate9657  (.A(g369), .B(II5202), .Z(II5203) ) ;
NAND2   gate9658  (.A(g374), .B(II5202), .Z(II5204) ) ;
NAND2   gate9659  (.A(g182), .B(g148), .Z(II5229) ) ;
NAND2   gate9660  (.A(g182), .B(II5229), .Z(II5230) ) ;
NAND2   gate9661  (.A(g148), .B(II5229), .Z(II5231) ) ;
NAND2   gate9662  (.A(II5230), .B(II5231), .Z(g2236) ) ;
NAND2   gate9663  (.A(g456), .B(g461), .Z(II5263) ) ;
NAND2   gate9664  (.A(g456), .B(II5263), .Z(II5264) ) ;
NAND2   gate9665  (.A(g461), .B(II5263), .Z(II5265) ) ;
NAND2   gate9666  (.A(g758), .B(g762), .Z(II5282) ) ;
NAND2   gate9667  (.A(g758), .B(II5282), .Z(II5283) ) ;
NAND2   gate9668  (.A(g762), .B(II5282), .Z(II5284) ) ;
NAND2   gate9669  (.A(g794), .B(g798), .Z(II5295) ) ;
NAND2   gate9670  (.A(g794), .B(II5295), .Z(II5296) ) ;
NAND2   gate9671  (.A(g798), .B(II5295), .Z(II5297) ) ;
NAND2   gate9672  (.A(g1032), .B(g1027), .Z(II5315) ) ;
NAND2   gate9673  (.A(g1032), .B(II5315), .Z(II5316) ) ;
NAND2   gate9674  (.A(g1027), .B(II5315), .Z(II5317) ) ;
NAND2   gate9675  (.A(g1336), .B(g1341), .Z(II5323) ) ;
NAND2   gate9676  (.A(g1336), .B(II5323), .Z(II5324) ) ;
NAND2   gate9677  (.A(g1341), .B(II5323), .Z(II5325) ) ;
NAND2   gate9678  (.A(g315), .B(g426), .Z(II5341) ) ;
NAND2   gate9679  (.A(g315), .B(II5341), .Z(II5342) ) ;
NAND2   gate9680  (.A(g426), .B(II5341), .Z(II5343) ) ;
NAND2   gate9681  (.A(g971), .B(g976), .Z(II5371) ) ;
NAND2   gate9682  (.A(g971), .B(II5371), .Z(II5372) ) ;
NAND2   gate9683  (.A(g976), .B(II5371), .Z(II5373) ) ;
NAND2   gate9684  (.A(g1515), .B(g1520), .Z(g2354) ) ;
NAND2   gate9685  (.A(g1235), .B(g991), .Z(II5449) ) ;
NAND2   gate9686  (.A(g1235), .B(II5449), .Z(II5450) ) ;
NAND2   gate9687  (.A(g991), .B(II5449), .Z(II5451) ) ;
NAND2   gate9688  (.A(g1240), .B(g1003), .Z(II5459) ) ;
NAND2   gate9689  (.A(g1240), .B(II5459), .Z(II5460) ) ;
NAND2   gate9690  (.A(g1003), .B(II5459), .Z(II5461) ) ;
NAND2   gate9691  (.A(g1245), .B(g999), .Z(II5468) ) ;
NAND2   gate9692  (.A(g1245), .B(II5468), .Z(II5469) ) ;
NAND2   gate9693  (.A(g999), .B(II5468), .Z(II5470) ) ;
NAND2   gate9694  (.A(g1250), .B(g1011), .Z(II5484) ) ;
NAND2   gate9695  (.A(g1250), .B(II5484), .Z(II5485) ) ;
NAND2   gate9696  (.A(g1011), .B(II5484), .Z(II5486) ) ;
NAND2   gate9697  (.A(g1255), .B(g1007), .Z(II5500) ) ;
NAND2   gate9698  (.A(g1255), .B(II5500), .Z(II5501) ) ;
NAND2   gate9699  (.A(g1007), .B(II5500), .Z(II5502) ) ;
NAND2   gate9700  (.A(g1260), .B(g1019), .Z(II5516) ) ;
NAND2   gate9701  (.A(g1260), .B(II5516), .Z(II5517) ) ;
NAND2   gate9702  (.A(g1019), .B(II5516), .Z(II5518) ) ;
NAND2   gate9703  (.A(g1265), .B(g1015), .Z(II5528) ) ;
NAND2   gate9704  (.A(g1265), .B(II5528), .Z(II5529) ) ;
NAND2   gate9705  (.A(g1015), .B(II5528), .Z(II5530) ) ;
NAND2   gate9706  (.A(g1270), .B(g1023), .Z(II5538) ) ;
NAND2   gate9707  (.A(g1270), .B(II5538), .Z(II5539) ) ;
NAND2   gate9708  (.A(g1023), .B(II5538), .Z(II5540) ) ;
NAND2   gate9709  (.A(g178), .B(g182), .Z(g2500) ) ;
NAND2   gate9710  (.A(g1696), .B(g1703), .Z(II5591) ) ;
NAND2   gate9711  (.A(g1696), .B(II5591), .Z(II5592) ) ;
NAND2   gate9712  (.A(g1703), .B(II5591), .Z(II5593) ) ;
NAND2   gate9713  (.A(g1149), .B(g1153), .Z(II5604) ) ;
NAND2   gate9714  (.A(g1149), .B(II5604), .Z(II5605) ) ;
NAND2   gate9715  (.A(g1153), .B(II5604), .Z(II5606) ) ;
NAND2   gate9716  (.A(g1280), .B(g1284), .Z(II5611) ) ;
NAND2   gate9717  (.A(g1280), .B(II5611), .Z(II5612) ) ;
NAND2   gate9718  (.A(g1284), .B(II5611), .Z(II5613) ) ;
NAND2   gate9719  (.A(g1766), .B(g1771), .Z(II5618) ) ;
NAND2   gate9720  (.A(g1766), .B(II5618), .Z(II5619) ) ;
NAND2   gate9721  (.A(g1771), .B(II5618), .Z(II5620) ) ;
NAND2   gate9722  (.A(g1218), .B(g1223), .Z(II5675) ) ;
NAND2   gate9723  (.A(g1218), .B(II5675), .Z(II5676) ) ;
NAND2   gate9724  (.A(g1223), .B(II5675), .Z(II5677) ) ;
NAND2   gate9725  (.A(g2107), .B(g2105), .Z(II5865) ) ;
NAND2   gate9726  (.A(g2107), .B(II5865), .Z(II5866) ) ;
NAND2   gate9727  (.A(g2105), .B(II5865), .Z(II5867) ) ;
NAND2   gate9728  (.A(II5866), .B(II5867), .Z(g2776) ) ;
NAND2   gate9729  (.A(g2120), .B(g2115), .Z(II5878) ) ;
NAND2   gate9730  (.A(g2120), .B(II5878), .Z(II5879) ) ;
NAND2   gate9731  (.A(g2115), .B(II5878), .Z(II5880) ) ;
NAND2   gate9732  (.A(II5879), .B(II5880), .Z(g2792) ) ;
NAND2   gate9733  (.A(g750), .B(g2057), .Z(II5891) ) ;
NAND2   gate9734  (.A(g750), .B(II5891), .Z(II5892) ) ;
NAND2   gate9735  (.A(g2057), .B(II5891), .Z(II5893) ) ;
NAND2   gate9736  (.A(II5892), .B(II5893), .Z(g2795) ) ;
NAND2   gate9737  (.A(g2205), .B(g1494), .Z(II6109) ) ;
NAND2   gate9738  (.A(g2205), .B(II6109), .Z(II6110) ) ;
NAND2   gate9739  (.A(g1494), .B(II6109), .Z(II6111) ) ;
NAND2   gate9740  (.A(II6110), .B(II6111), .Z(g2938) ) ;
NAND2   gate9741  (.A(g2215), .B(g1419), .Z(II6124) ) ;
NAND2   gate9742  (.A(g2215), .B(II6124), .Z(II6125) ) ;
NAND2   gate9743  (.A(g1419), .B(II6124), .Z(II6126) ) ;
NAND2   gate9744  (.A(II6125), .B(II6126), .Z(g2943) ) ;
NAND2   gate9745  (.A(g2496), .B(g378), .Z(II6136) ) ;
NAND2   gate9746  (.A(g2496), .B(II6136), .Z(II6137) ) ;
NAND2   gate9747  (.A(g378), .B(II6136), .Z(II6138) ) ;
NAND2   gate9748  (.A(g1976), .B(g646), .Z(II6143) ) ;
NAND2   gate9749  (.A(g1976), .B(II6143), .Z(II6144) ) ;
NAND2   gate9750  (.A(g646), .B(II6143), .Z(II6145) ) ;
NAND2   gate9751  (.A(g2236), .B(g153), .Z(II6166) ) ;
NAND2   gate9752  (.A(g2236), .B(II6166), .Z(II6167) ) ;
NAND2   gate9753  (.A(g153), .B(II6166), .Z(II6168) ) ;
NAND2   gate9754  (.A(II6167), .B(II6168), .Z(g2959) ) ;
NAND2   gate9755  (.A(g2177), .B(g197), .Z(II6176) ) ;
NAND2   gate9756  (.A(g2177), .B(II6176), .Z(II6177) ) ;
NAND2   gate9757  (.A(g197), .B(II6176), .Z(II6178) ) ;
NAND2   gate9758  (.A(II6177), .B(II6178), .Z(g2961) ) ;
NAND2   gate9759  (.A(g2511), .B(g466), .Z(II6186) ) ;
NAND2   gate9760  (.A(g2511), .B(II6186), .Z(II6187) ) ;
NAND2   gate9761  (.A(g466), .B(II6186), .Z(II6188) ) ;
NAND2   gate9762  (.A(g2525), .B(g766), .Z(II6199) ) ;
NAND2   gate9763  (.A(g2525), .B(II6199), .Z(II6200) ) ;
NAND2   gate9764  (.A(g766), .B(II6199), .Z(II6201) ) ;
NAND2   gate9765  (.A(g2534), .B(g802), .Z(II6207) ) ;
NAND2   gate9766  (.A(g2534), .B(II6207), .Z(II6208) ) ;
NAND2   gate9767  (.A(g802), .B(II6207), .Z(II6209) ) ;
NAND2   gate9768  (.A(g2544), .B(g1346), .Z(II6224) ) ;
NAND2   gate9769  (.A(g2544), .B(II6224), .Z(II6225) ) ;
NAND2   gate9770  (.A(g1346), .B(II6224), .Z(II6226) ) ;
NAND2   gate9771  (.A(g591), .B(g2382), .Z(g3011) ) ;
NAND2   gate9772  (.A(g611), .B(g2374), .Z(g3061) ) ;
NAND2   gate9773  (.A(g2091), .B(g981), .Z(II6287) ) ;
NAND2   gate9774  (.A(g2091), .B(II6287), .Z(II6288) ) ;
NAND2   gate9775  (.A(g981), .B(II6287), .Z(II6289) ) ;
NAND2   gate9776  (.A(g2050), .B(g1864), .Z(II6322) ) ;
NAND2   gate9777  (.A(g2050), .B(II6322), .Z(II6323) ) ;
NAND2   gate9778  (.A(g1864), .B(II6322), .Z(II6324) ) ;
NAND2   gate9779  (.A(g1814), .B(g2571), .Z(g3205) ) ;
NAND2   gate9780  (.A(g1834), .B(g2564), .Z(g3221) ) ;
NAND4   gate9781  (.A(g2229), .B(g2222), .C(g2211), .D(g2202), .Z(g3261) ) ;
NAND2   gate9782  (.A(g2264), .B(g1776), .Z(II6447) ) ;
NAND2   gate9783  (.A(g2264), .B(II6447), .Z(II6448) ) ;
NAND2   gate9784  (.A(g1776), .B(II6447), .Z(II6449) ) ;
NAND2   gate9785  (.A(g23), .B(g2479), .Z(II6467) ) ;
NAND2   gate9786  (.A(g23), .B(II6467), .Z(II6468) ) ;
NAND2   gate9787  (.A(g2479), .B(II6467), .Z(II6469) ) ;
NAND2   gate9788  (.A(g2306), .B(g1227), .Z(II6487) ) ;
NAND2   gate9789  (.A(g2306), .B(II6487), .Z(II6488) ) ;
NAND2   gate9790  (.A(g1227), .B(II6487), .Z(II6489) ) ;
NAND2   gate9791  (.A(g2792), .B(g2776), .Z(II6664) ) ;
NAND2   gate9792  (.A(g2792), .B(II6664), .Z(II6665) ) ;
NAND2   gate9793  (.A(g2776), .B(II6664), .Z(II6666) ) ;
NAND2   gate9794  (.A(II6665), .B(II6666), .Z(g3460) ) ;
NAND2   gate9795  (.A(g2961), .B(g201), .Z(II6714) ) ;
NAND2   gate9796  (.A(g2961), .B(II6714), .Z(II6715) ) ;
NAND2   gate9797  (.A(g201), .B(II6714), .Z(II6716) ) ;
NAND2   gate9798  (.A(II6715), .B(II6716), .Z(g3530) ) ;
NAND2   gate9799  (.A(g2938), .B(g1453), .Z(II6746) ) ;
NAND2   gate9800  (.A(g2938), .B(II6746), .Z(II6747) ) ;
NAND2   gate9801  (.A(g1453), .B(II6746), .Z(II6748) ) ;
NAND2   gate9802  (.A(g2943), .B(g1448), .Z(II6760) ) ;
NAND2   gate9803  (.A(g2943), .B(II6760), .Z(II6761) ) ;
NAND2   gate9804  (.A(g1448), .B(II6760), .Z(II6762) ) ;
NAND2   gate9805  (.A(II6761), .B(II6762), .Z(g3623) ) ;
NAND2   gate9806  (.A(g3257), .B(g382), .Z(II6770) ) ;
NAND2   gate9807  (.A(g3257), .B(II6770), .Z(II6771) ) ;
NAND2   gate9808  (.A(g382), .B(II6770), .Z(II6772) ) ;
NAND2   gate9809  (.A(g2892), .B(g650), .Z(II6777) ) ;
NAND2   gate9810  (.A(g2892), .B(II6777), .Z(II6778) ) ;
NAND2   gate9811  (.A(g650), .B(II6777), .Z(II6779) ) ;
NAND2   gate9812  (.A(g2959), .B(g143), .Z(II6792) ) ;
NAND2   gate9813  (.A(g2959), .B(II6792), .Z(II6793) ) ;
NAND2   gate9814  (.A(g143), .B(II6792), .Z(II6794) ) ;
NAND2   gate9815  (.A(g3268), .B(g471), .Z(II6805) ) ;
NAND2   gate9816  (.A(g3268), .B(II6805), .Z(II6806) ) ;
NAND2   gate9817  (.A(g471), .B(II6805), .Z(II6807) ) ;
NAND2   gate9818  (.A(g3281), .B(g770), .Z(II6825) ) ;
NAND2   gate9819  (.A(g3281), .B(II6825), .Z(II6826) ) ;
NAND2   gate9820  (.A(g770), .B(II6825), .Z(II6827) ) ;
NAND2   gate9821  (.A(g3287), .B(g806), .Z(II6836) ) ;
NAND2   gate9822  (.A(g3287), .B(II6836), .Z(II6837) ) ;
NAND2   gate9823  (.A(g806), .B(II6836), .Z(II6838) ) ;
NAND2   gate9824  (.A(g3301), .B(g1351), .Z(II6879) ) ;
NAND2   gate9825  (.A(g3301), .B(II6879), .Z(II6880) ) ;
NAND2   gate9826  (.A(g1351), .B(II6879), .Z(II6881) ) ;
NAND2   gate9827  (.A(g3039), .B(g599), .Z(g3734) ) ;
NAND2   gate9828  (.A(g2760), .B(g986), .Z(II6988) ) ;
NAND2   gate9829  (.A(g2760), .B(II6988), .Z(II6989) ) ;
NAND2   gate9830  (.A(g986), .B(II6988), .Z(II6990) ) ;
NAND2   gate9831  (.A(g3089), .B(g1868), .Z(II7033) ) ;
NAND2   gate9832  (.A(g3089), .B(II7033), .Z(II7034) ) ;
NAND2   gate9833  (.A(g1868), .B(II7033), .Z(II7035) ) ;
NAND2   gate9834  (.A(g3207), .B(g1822), .Z(g3978) ) ;
NAND2   gate9835  (.A(g2981), .B(g1781), .Z(II7223) ) ;
NAND2   gate9836  (.A(g2981), .B(II7223), .Z(II7224) ) ;
NAND2   gate9837  (.A(g1781), .B(II7223), .Z(II7225) ) ;
NAND2   gate9838  (.A(g3047), .B(g1231), .Z(II7321) ) ;
NAND2   gate9839  (.A(g3047), .B(II7321), .Z(II7322) ) ;
NAND2   gate9840  (.A(g1231), .B(II7321), .Z(II7323) ) ;
NAND2   gate9841  (.A(g3533), .B(g654), .Z(II7562) ) ;
NAND2   gate9842  (.A(g3533), .B(II7562), .Z(II7563) ) ;
NAND2   gate9843  (.A(g654), .B(II7562), .Z(II7564) ) ;
NAND2   gate9844  (.A(g1023), .B(g3460), .Z(II7683) ) ;
NAND2   gate9845  (.A(g1023), .B(II7683), .Z(II7684) ) ;
NAND2   gate9846  (.A(g3460), .B(II7683), .Z(II7685) ) ;
NAND2   gate9847  (.A(II7684), .B(II7685), .Z(g4374) ) ;
NAND2   gate9848  (.A(g4099), .B(g774), .Z(II7863) ) ;
NAND2   gate9849  (.A(g4099), .B(II7863), .Z(II7864) ) ;
NAND2   gate9850  (.A(g774), .B(II7863), .Z(II7865) ) ;
NAND2   gate9851  (.A(g4109), .B(g810), .Z(II7875) ) ;
NAND2   gate9852  (.A(g4109), .B(II7875), .Z(II7876) ) ;
NAND2   gate9853  (.A(g810), .B(II7875), .Z(II7877) ) ;
NAND2   gate9854  (.A(g3475), .B(g2399), .Z(g4538) ) ;
NAND2   gate9855  (.A(g3710), .B(g2061), .Z(g4749) ) ;
NAND2   gate9856  (.A(g3685), .B(g1786), .Z(II8178) ) ;
NAND2   gate9857  (.A(g3685), .B(II8178), .Z(II8179) ) ;
NAND2   gate9858  (.A(g1786), .B(II8178), .Z(II8180) ) ;
NOR3    gate9859  (.A(g3543), .B(g3419), .C(g3408), .Z(g4455) ) ;
NAND2   gate9860  (.A(g4455), .B(g3530), .Z(II8479) ) ;
NAND2   gate9861  (.A(g4455), .B(II8479), .Z(II8480) ) ;
NAND2   gate9862  (.A(g3530), .B(II8479), .Z(II8481) ) ;
NOR4    gate9863  (.A(g3292), .B(g2593), .C(g2586), .D(g3776), .Z(g4873) ) ;
NAND2   gate9864  (.A(g4873), .B(g3513), .Z(II8513) ) ;
NAND2   gate9865  (.A(g4873), .B(II8513), .Z(II8514) ) ;
NAND2   gate9866  (.A(g3513), .B(II8513), .Z(II8515) ) ;
NOR4    gate9867  (.A(g3292), .B(g2593), .C(g3784), .D(g2579), .Z(g4879) ) ;
NAND2   gate9868  (.A(g4879), .B(g481), .Z(II8527) ) ;
NAND2   gate9869  (.A(g4879), .B(II8527), .Z(II8528) ) ;
NAND2   gate9870  (.A(g481), .B(II8527), .Z(II8529) ) ;
NOR4    gate9871  (.A(g3292), .B(g2593), .C(g3784), .D(g3776), .Z(g4218) ) ;
NAND2   gate9872  (.A(g4218), .B(g486), .Z(II8543) ) ;
NAND2   gate9873  (.A(g4218), .B(II8543), .Z(II8544) ) ;
NAND2   gate9874  (.A(g486), .B(II8543), .Z(II8545) ) ;
NOR4    gate9875  (.A(g3292), .B(g3793), .C(g2586), .D(g2579), .Z(g4227) ) ;
NAND2   gate9876  (.A(g4227), .B(g491), .Z(II8561) ) ;
NAND2   gate9877  (.A(g4227), .B(II8561), .Z(II8562) ) ;
NAND2   gate9878  (.A(g491), .B(II8561), .Z(II8563) ) ;
NOR4    gate9879  (.A(g3292), .B(g3793), .C(g2586), .D(g3776), .Z(g4234) ) ;
NAND2   gate9880  (.A(g4234), .B(g496), .Z(II8575) ) ;
NAND2   gate9881  (.A(g4234), .B(II8575), .Z(II8576) ) ;
NAND2   gate9882  (.A(g496), .B(II8575), .Z(II8577) ) ;
NOR4    gate9883  (.A(g3292), .B(g3793), .C(g3784), .D(g2579), .Z(g4251) ) ;
NAND2   gate9884  (.A(g4251), .B(g501), .Z(II8589) ) ;
NAND2   gate9885  (.A(g4251), .B(II8589), .Z(II8590) ) ;
NAND2   gate9886  (.A(g501), .B(II8589), .Z(II8591) ) ;
NOR4    gate9887  (.A(g3292), .B(g3793), .C(g3784), .D(g3776), .Z(g4259) ) ;
NAND2   gate9888  (.A(g4259), .B(g506), .Z(II8604) ) ;
NAND2   gate9889  (.A(g4259), .B(II8604), .Z(II8605) ) ;
NAND2   gate9890  (.A(g506), .B(II8604), .Z(II8606) ) ;
NOR4    gate9891  (.A(g3800), .B(g2593), .C(g2586), .D(g2579), .Z(g4267) ) ;
NAND2   gate9892  (.A(g4267), .B(g511), .Z(II8624) ) ;
NAND2   gate9893  (.A(g4267), .B(II8624), .Z(II8625) ) ;
NAND2   gate9894  (.A(g511), .B(II8624), .Z(II8626) ) ;
NOR4    gate9895  (.A(g3800), .B(g2593), .C(g2586), .D(g3776), .Z(g4278) ) ;
NAND2   gate9896  (.A(g4278), .B(g516), .Z(II8640) ) ;
NAND2   gate9897  (.A(g4278), .B(II8640), .Z(II8641) ) ;
NAND2   gate9898  (.A(g516), .B(II8640), .Z(II8642) ) ;
NAND2   gate9899  (.A(g4824), .B(g778), .Z(II8650) ) ;
NAND2   gate9900  (.A(g4824), .B(II8650), .Z(II8651) ) ;
NAND2   gate9901  (.A(g778), .B(II8650), .Z(II8652) ) ;
NOR4    gate9902  (.A(g3800), .B(g2593), .C(g3784), .D(g2579), .Z(g4286) ) ;
NAND2   gate9903  (.A(g4286), .B(g476), .Z(II8662) ) ;
NAND2   gate9904  (.A(g4286), .B(II8662), .Z(II8663) ) ;
NAND2   gate9905  (.A(g476), .B(II8662), .Z(II8664) ) ;
NAND2   gate9906  (.A(g4831), .B(g814), .Z(II8669) ) ;
NAND2   gate9907  (.A(g4831), .B(II8669), .Z(II8670) ) ;
NAND2   gate9908  (.A(g814), .B(II8669), .Z(II8671) ) ;
NAND2   gate9909  (.A(g4374), .B(g1027), .Z(II8676) ) ;
NAND2   gate9910  (.A(g4374), .B(II8676), .Z(II8677) ) ;
NAND2   gate9911  (.A(g1027), .B(II8676), .Z(II8678) ) ;
NOR4    gate9912  (.A(g3077), .B(g2669), .C(g2662), .D(g3479), .Z(g4601) ) ;
NAND2   gate9913  (.A(g4601), .B(g4052), .Z(II8715) ) ;
NAND2   gate9914  (.A(g4601), .B(II8715), .Z(II8716) ) ;
NAND2   gate9915  (.A(g4052), .B(II8715), .Z(II8717) ) ;
NOR4    gate9916  (.A(g3077), .B(g2669), .C(g3485), .D(g2655), .Z(g4605) ) ;
NAND2   gate9917  (.A(g4605), .B(g1117), .Z(II8728) ) ;
NAND2   gate9918  (.A(g4605), .B(II8728), .Z(II8729) ) ;
NAND2   gate9919  (.A(g1117), .B(II8728), .Z(II8730) ) ;
NAND2   gate9920  (.A(g3734), .B(g4538), .Z(g5277) ) ;
NOR4    gate9921  (.A(g3077), .B(g2669), .C(g3485), .D(g3479), .Z(g4607) ) ;
NAND2   gate9922  (.A(g4607), .B(g1121), .Z(II8738) ) ;
NAND2   gate9923  (.A(g4607), .B(II8738), .Z(II8739) ) ;
NAND2   gate9924  (.A(g1121), .B(II8738), .Z(II8740) ) ;
NOR4    gate9925  (.A(g3077), .B(g3491), .C(g2662), .D(g2655), .Z(g4613) ) ;
NAND2   gate9926  (.A(g4613), .B(g1125), .Z(II8750) ) ;
NAND2   gate9927  (.A(g4613), .B(II8750), .Z(II8751) ) ;
NAND2   gate9928  (.A(g1125), .B(II8750), .Z(II8752) ) ;
NOR4    gate9929  (.A(g3077), .B(g3491), .C(g2662), .D(g3479), .Z(g4616) ) ;
NAND2   gate9930  (.A(g4616), .B(g1129), .Z(II8761) ) ;
NAND2   gate9931  (.A(g4616), .B(II8761), .Z(II8762) ) ;
NAND2   gate9932  (.A(g1129), .B(II8761), .Z(II8763) ) ;
NOR4    gate9933  (.A(g3077), .B(g3491), .C(g3485), .D(g2655), .Z(g4619) ) ;
NAND2   gate9934  (.A(g4619), .B(g1133), .Z(II8770) ) ;
NAND2   gate9935  (.A(g4619), .B(II8770), .Z(II8771) ) ;
NAND2   gate9936  (.A(g1133), .B(II8770), .Z(II8772) ) ;
NOR4    gate9937  (.A(g3077), .B(g3491), .C(g3485), .D(g3479), .Z(g4630) ) ;
NAND2   gate9938  (.A(g4630), .B(g1137), .Z(II8778) ) ;
NAND2   gate9939  (.A(g4630), .B(II8778), .Z(II8779) ) ;
NAND2   gate9940  (.A(g1137), .B(II8778), .Z(II8780) ) ;
NOR4    gate9941  (.A(g3501), .B(g2669), .C(g2662), .D(g2655), .Z(g4639) ) ;
NAND2   gate9942  (.A(g4639), .B(g1141), .Z(II8786) ) ;
NAND2   gate9943  (.A(g4639), .B(II8786), .Z(II8787) ) ;
NAND2   gate9944  (.A(g1141), .B(II8786), .Z(II8788) ) ;
NOR4    gate9945  (.A(g3501), .B(g2669), .C(g2662), .D(g3479), .Z(g4672) ) ;
NAND2   gate9946  (.A(g4672), .B(g1145), .Z(II8795) ) ;
NAND2   gate9947  (.A(g4672), .B(II8795), .Z(II8796) ) ;
NAND2   gate9948  (.A(g1145), .B(II8795), .Z(II8797) ) ;
NOR4    gate9949  (.A(g3501), .B(g2669), .C(g3485), .D(g2655), .Z(g4677) ) ;
NAND2   gate9950  (.A(g4677), .B(g1113), .Z(II8803) ) ;
NAND2   gate9951  (.A(g4677), .B(II8803), .Z(II8804) ) ;
NAND2   gate9952  (.A(g1113), .B(II8803), .Z(II8805) ) ;
NAND2   gate9953  (.A(g3978), .B(g4749), .Z(g5527) ) ;
NAND2   gate9954  (.A(g4777), .B(g4401), .Z(g5552) ) ;
NAND2   gate9955  (.A(g4492), .B(g1791), .Z(II9006) ) ;
NAND2   gate9956  (.A(g4492), .B(II9006), .Z(II9007) ) ;
NAND2   gate9957  (.A(g1791), .B(II9006), .Z(II9008) ) ;
NAND2   gate9958  (.A(g5598), .B(g782), .Z(II9557) ) ;
NAND2   gate9959  (.A(g5598), .B(II9557), .Z(II9558) ) ;
NAND2   gate9960  (.A(g782), .B(II9557), .Z(II9559) ) ;
NAND2   gate9961  (.A(g5608), .B(g818), .Z(II9574) ) ;
NAND2   gate9962  (.A(g5608), .B(II9574), .Z(II9575) ) ;
NAND2   gate9963  (.A(g818), .B(II9574), .Z(II9576) ) ;
NAND2   gate9964  (.A(g4566), .B(g4921), .Z(g6027) ) ;
NAND2   gate9965  (.A(g5233), .B(g1796), .Z(II9946) ) ;
NAND2   gate9966  (.A(g5233), .B(II9946), .Z(II9947) ) ;
NAND2   gate9967  (.A(g1796), .B(II9946), .Z(II9948) ) ;
NAND2   gate9968  (.A(g6221), .B(g786), .Z(II10507) ) ;
NAND2   gate9969  (.A(g6221), .B(II10507), .Z(II10508) ) ;
NAND2   gate9970  (.A(g786), .B(II10507), .Z(II10509) ) ;
NAND2   gate9971  (.A(g6231), .B(g822), .Z(II10519) ) ;
NAND2   gate9972  (.A(g6231), .B(II10519), .Z(II10520) ) ;
NAND2   gate9973  (.A(g822), .B(II10519), .Z(II10521) ) ;
NAND2   gate9974  (.A(g5944), .B(g1801), .Z(II10769) ) ;
NAND2   gate9975  (.A(g5944), .B(II10769), .Z(II10770) ) ;
NAND2   gate9976  (.A(g1801), .B(II10769), .Z(II10771) ) ;
NAND2   gate9977  (.A(g6395), .B(g5555), .Z(II10930) ) ;
NAND2   gate9978  (.A(g6395), .B(II10930), .Z(II10931) ) ;
NAND2   gate9979  (.A(g5555), .B(II10930), .Z(II10932) ) ;
NAND2   gate9980  (.A(g6760), .B(g790), .Z(II11241) ) ;
NAND2   gate9981  (.A(g6760), .B(II11241), .Z(II11242) ) ;
NAND2   gate9982  (.A(g790), .B(II11241), .Z(II11243) ) ;
NAND2   gate9983  (.A(g6775), .B(g826), .Z(II11261) ) ;
NAND2   gate9984  (.A(g6775), .B(II11261), .Z(II11262) ) ;
NAND2   gate9985  (.A(g826), .B(II11261), .Z(II11263) ) ;
NAND2   gate9986  (.A(g305), .B(g6485), .Z(II11278) ) ;
NAND2   gate9987  (.A(g305), .B(II11278), .Z(II11279) ) ;
NAND2   gate9988  (.A(g6485), .B(II11278), .Z(II11280) ) ;
NAND2   gate9989  (.A(g6580), .B(g1806), .Z(II11508) ) ;
NAND2   gate9990  (.A(g6580), .B(II11508), .Z(II11509) ) ;
NAND2   gate9991  (.A(g1806), .B(II11508), .Z(II11510) ) ;
NAND2   gate9992  (.A(g6967), .B(g1474), .Z(II11907) ) ;
NAND2   gate9993  (.A(g6967), .B(II11907), .Z(II11908) ) ;
NAND2   gate9994  (.A(g1474), .B(II11907), .Z(II11909) ) ;
NAND2   gate9995  (.A(g6935), .B(g1494), .Z(II11914) ) ;
NAND2   gate9996  (.A(g6935), .B(II11914), .Z(II11915) ) ;
NAND2   gate9997  (.A(g1494), .B(II11914), .Z(II11916) ) ;
NAND2   gate9998  (.A(g7004), .B(g1458), .Z(II11935) ) ;
NAND2   gate9999  (.A(g7004), .B(II11935), .Z(II11936) ) ;
NAND2   gate10000  (.A(g1458), .B(II11935), .Z(II11937) ) ;
NAND2   gate10001  (.A(g7001), .B(g1462), .Z(II11973) ) ;
NAND2   gate10002  (.A(g7001), .B(II11973), .Z(II11974) ) ;
NAND2   gate10003  (.A(g1462), .B(II11973), .Z(II11975) ) ;
NAND2   gate10004  (.A(g6957), .B(g1482), .Z(II11980) ) ;
NAND2   gate10005  (.A(g6957), .B(II11980), .Z(II11981) ) ;
NAND2   gate10006  (.A(g1482), .B(II11980), .Z(II11982) ) ;
NAND2   gate10007  (.A(g7107), .B(g127), .Z(II11995) ) ;
NAND2   gate10008  (.A(g7107), .B(II11995), .Z(II11996) ) ;
NAND2   gate10009  (.A(g127), .B(II11995), .Z(II11997) ) ;
NAND2   gate10010  (.A(g7082), .B(g153), .Z(II12002) ) ;
NAND2   gate10011  (.A(g7082), .B(II12002), .Z(II12003) ) ;
NAND2   gate10012  (.A(g153), .B(II12002), .Z(II12004) ) ;
NAND2   gate10013  (.A(g7119), .B(g166), .Z(II12019) ) ;
NAND2   gate10014  (.A(g7119), .B(II12019), .Z(II12020) ) ;
NAND2   gate10015  (.A(g166), .B(II12019), .Z(II12021) ) ;
NAND2   gate10016  (.A(g6990), .B(g1466), .Z(II12038) ) ;
NAND2   gate10017  (.A(g6990), .B(II12038), .Z(II12039) ) ;
NAND2   gate10018  (.A(g1466), .B(II12038), .Z(II12040) ) ;
NAND2   gate10019  (.A(g6951), .B(g1486), .Z(II12045) ) ;
NAND2   gate10020  (.A(g6951), .B(II12045), .Z(II12046) ) ;
NAND2   gate10021  (.A(g1486), .B(II12045), .Z(II12047) ) ;
NAND2   gate10022  (.A(g6961), .B(g1478), .Z(II12060) ) ;
NAND2   gate10023  (.A(g6961), .B(II12060), .Z(II12061) ) ;
NAND2   gate10024  (.A(g1478), .B(II12060), .Z(II12062) ) ;
NAND2   gate10025  (.A(g7116), .B(g139), .Z(II12067) ) ;
NAND2   gate10026  (.A(g7116), .B(II12067), .Z(II12068) ) ;
NAND2   gate10027  (.A(g139), .B(II12067), .Z(II12069) ) ;
NAND2   gate10028  (.A(g7098), .B(g174), .Z(II12074) ) ;
NAND2   gate10029  (.A(g7098), .B(II12074), .Z(II12075) ) ;
NAND2   gate10030  (.A(g174), .B(II12074), .Z(II12076) ) ;
NAND2   gate10031  (.A(g6980), .B(g1470), .Z(II12085) ) ;
NAND2   gate10032  (.A(g6980), .B(II12085), .Z(II12086) ) ;
NAND2   gate10033  (.A(g1470), .B(II12085), .Z(II12087) ) ;
NAND2   gate10034  (.A(g6944), .B(g1490), .Z(II12092) ) ;
NAND2   gate10035  (.A(g6944), .B(II12092), .Z(II12093) ) ;
NAND2   gate10036  (.A(g1490), .B(II12092), .Z(II12094) ) ;
NAND2   gate10037  (.A(g7113), .B(g135), .Z(II12106) ) ;
NAND2   gate10038  (.A(g7113), .B(II12106), .Z(II12107) ) ;
NAND2   gate10039  (.A(g135), .B(II12106), .Z(II12108) ) ;
NAND2   gate10040  (.A(g7093), .B(g162), .Z(II12113) ) ;
NAND2   gate10041  (.A(g7093), .B(II12113), .Z(II12114) ) ;
NAND2   gate10042  (.A(g162), .B(II12113), .Z(II12115) ) ;
NAND2   gate10043  (.A(g7103), .B(g170), .Z(II12126) ) ;
NAND2   gate10044  (.A(g7103), .B(II12126), .Z(II12127) ) ;
NAND2   gate10045  (.A(g170), .B(II12126), .Z(II12128) ) ;
NAND2   gate10046  (.A(g7110), .B(g131), .Z(II12136) ) ;
NAND2   gate10047  (.A(g7110), .B(II12136), .Z(II12137) ) ;
NAND2   gate10048  (.A(g131), .B(II12136), .Z(II12138) ) ;
NAND2   gate10049  (.A(g7089), .B(g158), .Z(II12143) ) ;
NAND2   gate10050  (.A(g7089), .B(II12143), .Z(II12144) ) ;
NAND2   gate10051  (.A(g158), .B(II12143), .Z(II12145) ) ;
NAND2   gate10052  (.A(g7061), .B(g2518), .Z(II12214) ) ;
NAND2   gate10053  (.A(g7061), .B(II12214), .Z(II12215) ) ;
NAND2   gate10054  (.A(g2518), .B(II12214), .Z(II12216) ) ;
NAND2   gate10055  (.A(g6863), .B(g3206), .Z(g7717) ) ;
NOR2    gate10056  (.A(g4117), .B(g4432), .Z(g5573) ) ;
NAND2   gate10057  (.A(g7697), .B(g3038), .Z(g7978) ) ;
NAND2   gate10058  (.A(g5552), .B(g7717), .Z(g8006) ) ;
NAND2   gate10059  (.A(g1872), .B(g7963), .Z(II13076) ) ;
NAND2   gate10060  (.A(g1872), .B(II13076), .Z(II13077) ) ;
NAND2   gate10061  (.A(g7963), .B(II13076), .Z(II13078) ) ;
NAND2   gate10062  (.A(g8006), .B(g1840), .Z(II13089) ) ;
NAND2   gate10063  (.A(g8006), .B(II13089), .Z(II13090) ) ;
NAND2   gate10064  (.A(g1840), .B(II13089), .Z(II13091) ) ;
NAND2   gate10065  (.A(g6027), .B(g7978), .Z(g8190) ) ;
NAND2   gate10066  (.A(g1891), .B(g8148), .Z(II13248) ) ;
NAND2   gate10067  (.A(g1891), .B(II13248), .Z(II13249) ) ;
NAND2   gate10068  (.A(g8148), .B(II13248), .Z(II13250) ) ;
NAND2   gate10069  (.A(g1900), .B(g8153), .Z(II13258) ) ;
NAND2   gate10070  (.A(g1900), .B(II13258), .Z(II13259) ) ;
NAND2   gate10071  (.A(g8153), .B(II13258), .Z(II13260) ) ;
NAND2   gate10072  (.A(g1909), .B(g8154), .Z(II13265) ) ;
NAND2   gate10073  (.A(g1909), .B(II13265), .Z(II13266) ) ;
NAND2   gate10074  (.A(g8154), .B(II13265), .Z(II13267) ) ;
NAND2   gate10075  (.A(g1918), .B(g8158), .Z(II13272) ) ;
NAND2   gate10076  (.A(g1918), .B(II13272), .Z(II13273) ) ;
NAND2   gate10077  (.A(g8158), .B(II13272), .Z(II13274) ) ;
NAND2   gate10078  (.A(g1927), .B(g8159), .Z(II13283) ) ;
NAND2   gate10079  (.A(g1927), .B(II13283), .Z(II13284) ) ;
NAND2   gate10080  (.A(g8159), .B(II13283), .Z(II13285) ) ;
NAND2   gate10081  (.A(g1882), .B(g8161), .Z(II13293) ) ;
NAND2   gate10082  (.A(g1882), .B(II13293), .Z(II13294) ) ;
NAND2   gate10083  (.A(g8161), .B(II13293), .Z(II13295) ) ;
NAND2   gate10084  (.A(g1936), .B(g8162), .Z(II13300) ) ;
NAND2   gate10085  (.A(g1936), .B(II13300), .Z(II13301) ) ;
NAND2   gate10086  (.A(g8162), .B(II13300), .Z(II13302) ) ;
NAND2   gate10087  (.A(g8190), .B(g617), .Z(II13307) ) ;
NAND2   gate10088  (.A(g8190), .B(II13307), .Z(II13308) ) ;
NAND2   gate10089  (.A(g617), .B(II13307), .Z(II13309) ) ;
NAND2   gate10090  (.A(g677), .B(g8247), .Z(II13504) ) ;
NAND2   gate10091  (.A(g677), .B(II13504), .Z(II13505) ) ;
NAND2   gate10092  (.A(g8247), .B(II13504), .Z(II13506) ) ;
NAND2   gate10093  (.A(g686), .B(g8248), .Z(II13513) ) ;
NAND2   gate10094  (.A(g686), .B(II13513), .Z(II13514) ) ;
NAND2   gate10095  (.A(g8248), .B(II13513), .Z(II13515) ) ;
NAND2   gate10096  (.A(g695), .B(g8249), .Z(II13521) ) ;
NAND2   gate10097  (.A(g695), .B(II13521), .Z(II13522) ) ;
NAND2   gate10098  (.A(g8249), .B(II13521), .Z(II13523) ) ;
NAND2   gate10099  (.A(g704), .B(g8253), .Z(II13529) ) ;
NAND2   gate10100  (.A(g704), .B(II13529), .Z(II13530) ) ;
NAND2   gate10101  (.A(g8253), .B(II13529), .Z(II13531) ) ;
NAND2   gate10102  (.A(g658), .B(g8157), .Z(II13537) ) ;
NAND2   gate10103  (.A(g658), .B(II13537), .Z(II13538) ) ;
NAND2   gate10104  (.A(g8157), .B(II13537), .Z(II13539) ) ;
NAND2   gate10105  (.A(g713), .B(g8259), .Z(II13544) ) ;
NAND2   gate10106  (.A(g713), .B(II13544), .Z(II13545) ) ;
NAND2   gate10107  (.A(g8259), .B(II13544), .Z(II13546) ) ;
NAND2   gate10108  (.A(g668), .B(g8262), .Z(II13552) ) ;
NAND2   gate10109  (.A(g668), .B(II13552), .Z(II13553) ) ;
NAND2   gate10110  (.A(g8262), .B(II13552), .Z(II13554) ) ;
NAND2   gate10111  (.A(g722), .B(g8263), .Z(II13559) ) ;
NAND2   gate10112  (.A(g722), .B(II13559), .Z(II13560) ) ;
NAND2   gate10113  (.A(g8263), .B(II13559), .Z(II13561) ) ;
NAND2   gate10114  (.A(g1945), .B(g8322), .Z(II13659) ) ;
NAND2   gate10115  (.A(g1945), .B(II13659), .Z(II13660) ) ;
NAND2   gate10116  (.A(g8322), .B(II13659), .Z(II13661) ) ;
NAND2   gate10117  (.A(g3760), .B(g8366), .Z(g8501) ) ;
NAND4   gate10118  (.A(g2382), .B(g605), .C(g591), .D(g8366), .Z(g8502) ) ;
NAND2   gate10119  (.A(g3475), .B(g8366), .Z(g8506) ) ;
NAND2   gate10120  (.A(g4001), .B(g8390), .Z(g8541) ) ;
NAND4   gate10121  (.A(g2571), .B(g1828), .C(g1814), .D(g8390), .Z(g8542) ) ;
NAND2   gate10122  (.A(g3710), .B(g8390), .Z(g8545) ) ;
NAND2   gate10123  (.A(g731), .B(g8417), .Z(II13765) ) ;
NAND2   gate10124  (.A(g731), .B(II13765), .Z(II13766) ) ;
NAND2   gate10125  (.A(g8417), .B(II13765), .Z(II13767) ) ;
NAND2   gate10126  (.A(g8538), .B(g1448), .Z(II13857) ) ;
NAND2   gate10127  (.A(g8538), .B(II13857), .Z(II13858) ) ;
NAND2   gate10128  (.A(g1448), .B(II13857), .Z(II13859) ) ;
NAND2   gate10129  (.A(g8523), .B(g1403), .Z(II13867) ) ;
NAND2   gate10130  (.A(g8523), .B(II13867), .Z(II13868) ) ;
NAND2   gate10131  (.A(g1403), .B(II13867), .Z(II13869) ) ;
NAND2   gate10132  (.A(g8535), .B(g1444), .Z(II13876) ) ;
NAND2   gate10133  (.A(g8535), .B(II13876), .Z(II13877) ) ;
NAND2   gate10134  (.A(g1444), .B(II13876), .Z(II13878) ) ;
NAND2   gate10135  (.A(g8532), .B(g1440), .Z(II13886) ) ;
NAND2   gate10136  (.A(g8532), .B(II13886), .Z(II13887) ) ;
NAND2   gate10137  (.A(g1440), .B(II13886), .Z(II13888) ) ;
NAND2   gate10138  (.A(g8529), .B(g1436), .Z(II13893) ) ;
NAND2   gate10139  (.A(g8529), .B(II13893), .Z(II13894) ) ;
NAND2   gate10140  (.A(g1436), .B(II13893), .Z(II13895) ) ;
NAND2   gate10141  (.A(g8520), .B(g1428), .Z(II13900) ) ;
NAND2   gate10142  (.A(g8520), .B(II13900), .Z(II13901) ) ;
NAND2   gate10143  (.A(g1428), .B(II13900), .Z(II13902) ) ;
NAND2   gate10144  (.A(g8526), .B(g1432), .Z(II13907) ) ;
NAND2   gate10145  (.A(g8526), .B(II13907), .Z(II13908) ) ;
NAND2   gate10146  (.A(g1432), .B(II13907), .Z(II13909) ) ;
NAND2   gate10147  (.A(g622), .B(g8688), .Z(II13990) ) ;
NAND2   gate10148  (.A(g622), .B(II13990), .Z(II13991) ) ;
NAND2   gate10149  (.A(g8688), .B(II13990), .Z(II13992) ) ;
NAND3   gate10150  (.A(g2317), .B(g4921), .C(g8688), .Z(g8737) ) ;
NAND2   gate10151  (.A(g8688), .B(g4921), .Z(g8738) ) ;
NAND2   gate10152  (.A(g8599), .B(g4401), .Z(g8757) ) ;
NAND3   gate10153  (.A(g8502), .B(g8501), .C(g8739), .Z(g8824) ) ;
NAND3   gate10154  (.A(g8502), .B(g8738), .C(g8506), .Z(g8825) ) ;
NAND3   gate10155  (.A(g8739), .B(g8737), .C(g8648), .Z(g8826) ) ;
NAND2   gate10156  (.A(g8750), .B(g4401), .Z(g8839) ) ;
NAND3   gate10157  (.A(g8542), .B(g8541), .C(g8760), .Z(g8840) ) ;
NAND3   gate10158  (.A(g8542), .B(g8757), .C(g8545), .Z(g8843) ) ;
NAND2   gate10159  (.A(g8760), .B(g8683), .Z(g8847) ) ;
NAND2   gate10160  (.A(g8825), .B(g591), .Z(II14202) ) ;
NAND2   gate10161  (.A(g8825), .B(II14202), .Z(II14203) ) ;
NAND2   gate10162  (.A(g591), .B(II14202), .Z(II14204) ) ;
NAND2   gate10163  (.A(g8824), .B(g599), .Z(II14209) ) ;
NAND2   gate10164  (.A(g8824), .B(II14209), .Z(II14210) ) ;
NAND2   gate10165  (.A(g599), .B(II14209), .Z(II14211) ) ;
NAND2   gate10166  (.A(g8826), .B(g605), .Z(II14216) ) ;
NAND2   gate10167  (.A(g8826), .B(II14216), .Z(II14217) ) ;
NAND2   gate10168  (.A(g605), .B(II14216), .Z(II14218) ) ;
NAND2   gate10169  (.A(g8843), .B(g1814), .Z(II14263) ) ;
NAND2   gate10170  (.A(g8843), .B(II14263), .Z(II14264) ) ;
NAND2   gate10171  (.A(g1814), .B(II14263), .Z(II14265) ) ;
NAND2   gate10172  (.A(g8840), .B(g1822), .Z(II14270) ) ;
NAND2   gate10173  (.A(g8840), .B(II14270), .Z(II14271) ) ;
NAND2   gate10174  (.A(g1822), .B(II14270), .Z(II14272) ) ;
NAND2   gate10175  (.A(g8847), .B(g1828), .Z(II14277) ) ;
NAND2   gate10176  (.A(g8847), .B(II14277), .Z(II14278) ) ;
NAND2   gate10177  (.A(g1828), .B(II14277), .Z(II14279) ) ;
NAND2   gate10178  (.A(g8823), .B(g4921), .Z(g8942) ) ;
NAND2   gate10179  (.A(g5548), .B(g8839), .Z(g8970) ) ;
NAND2   gate10180  (.A(g8970), .B(g1834), .Z(II14442) ) ;
NAND2   gate10181  (.A(g8970), .B(II14442), .Z(II14443) ) ;
NAND2   gate10182  (.A(g1834), .B(II14442), .Z(II14444) ) ;
NAND2   gate10183  (.A(g6019), .B(g8942), .Z(g9204) ) ;
NAND2   gate10184  (.A(g9204), .B(g611), .Z(II14612) ) ;
NAND2   gate10185  (.A(g9204), .B(II14612), .Z(II14613) ) ;
NAND2   gate10186  (.A(g611), .B(II14612), .Z(II14614) ) ;
NAND2   gate10187  (.A(g9984), .B(g9980), .Z(II15256) ) ;
NAND2   gate10188  (.A(g9984), .B(II15256), .Z(II15257) ) ;
NAND2   gate10189  (.A(g9980), .B(II15256), .Z(II15258) ) ;
NAND2   gate10190  (.A(II15257), .B(II15258), .Z(g10043) ) ;
NAND2   gate10191  (.A(g10047), .B(g10044), .Z(II15430) ) ;
NAND2   gate10192  (.A(g10047), .B(II15430), .Z(II15431) ) ;
NAND2   gate10193  (.A(g10044), .B(II15430), .Z(II15432) ) ;
NAND2   gate10194  (.A(II15431), .B(II15432), .Z(g10144) ) ;
NAND2   gate10195  (.A(g10035), .B(g10122), .Z(II15441) ) ;
NAND2   gate10196  (.A(g10035), .B(II15441), .Z(II15442) ) ;
NAND2   gate10197  (.A(g10122), .B(II15441), .Z(II15443) ) ;
NAND2   gate10198  (.A(II15442), .B(II15443), .Z(g10149) ) ;
NAND2   gate10199  (.A(g10058), .B(g10051), .Z(II15451) ) ;
NAND2   gate10200  (.A(g10058), .B(II15451), .Z(II15452) ) ;
NAND2   gate10201  (.A(g10051), .B(II15451), .Z(II15453) ) ;
NAND2   gate10202  (.A(II15452), .B(II15453), .Z(g10153) ) ;
NAND2   gate10203  (.A(g10149), .B(g10144), .Z(II15607) ) ;
NAND2   gate10204  (.A(g10149), .B(II15607), .Z(II15608) ) ;
NAND2   gate10205  (.A(g10144), .B(II15607), .Z(II15609) ) ;
NAND2   gate10206  (.A(II15608), .B(II15609), .Z(g10229) ) ;
NAND2   gate10207  (.A(g10043), .B(g10153), .Z(II15615) ) ;
NAND2   gate10208  (.A(g10043), .B(II15615), .Z(II15616) ) ;
NAND2   gate10209  (.A(g10153), .B(II15615), .Z(II15617) ) ;
NAND2   gate10210  (.A(II15616), .B(II15617), .Z(g10231) ) ;
NAND2   gate10211  (.A(g10231), .B(g10229), .Z(II15716) ) ;
NAND2   gate10212  (.A(g10231), .B(II15716), .Z(II15717) ) ;
NAND2   gate10213  (.A(g10229), .B(II15716), .Z(II15718) ) ;
NAND2   gate10214  (.A(II15717), .B(II15718), .Z(g10302) ) ;
NOR2    gate10215  (.A(g10276), .B(g3566), .Z(g10285) ) ;
NOR2    gate10216  (.A(g10226), .B(g4620), .Z(g10358) ) ;
NAND2   gate10217  (.A(g10358), .B(g2713), .Z(II15870) ) ;
NAND2   gate10218  (.A(g10358), .B(II15870), .Z(II15871) ) ;
NAND2   gate10219  (.A(g2713), .B(II15870), .Z(II15872) ) ;
NOR2    gate10220  (.A(g10227), .B(g4620), .Z(g10359) ) ;
NAND2   gate10221  (.A(g10359), .B(g2719), .Z(II15878) ) ;
NAND2   gate10222  (.A(g10359), .B(II15878), .Z(II15879) ) ;
NAND2   gate10223  (.A(g2719), .B(II15878), .Z(II15880) ) ;
NOR2    gate10224  (.A(g10271), .B(g3463), .Z(g10286) ) ;
NAND2   gate10225  (.A(g853), .B(g10286), .Z(II15890) ) ;
NAND2   gate10226  (.A(g853), .B(II15890), .Z(II15891) ) ;
NAND2   gate10227  (.A(g10286), .B(II15890), .Z(II15892) ) ;
NOR2    gate10228  (.A(g10275), .B(g3463), .Z(g10287) ) ;
NAND2   gate10229  (.A(g857), .B(g10287), .Z(II15898) ) ;
NAND2   gate10230  (.A(g857), .B(II15898), .Z(II15899) ) ;
NAND2   gate10231  (.A(g10287), .B(II15898), .Z(II15900) ) ;
NAND2   gate10232  (.A(g6899), .B(g10302), .Z(II15906) ) ;
NAND2   gate10233  (.A(g6899), .B(II15906), .Z(II15907) ) ;
NAND2   gate10234  (.A(g10302), .B(II15906), .Z(II15908) ) ;
NOR2    gate10235  (.A(g10277), .B(g3566), .Z(g10360) ) ;
NOR2    gate10236  (.A(g3305), .B(g5614), .Z(g6037) ) ;
NOR2    gate10237  (.A(g10353), .B(g3566), .Z(g10443) ) ;
NOR2    gate10238  (.A(g4163), .B(g4872), .Z(g5350) ) ;
NOR2    gate10239  (.A(g10355), .B(g3566), .Z(g10363) ) ;
NOR2    gate10240  (.A(g2071), .B(g4225), .Z(g5360) ) ;
NOR2    gate10241  (.A(g10289), .B(g4620), .Z(g10422) ) ;
NAND2   gate10242  (.A(g10422), .B(g2677), .Z(II15992) ) ;
NAND2   gate10243  (.A(g10422), .B(II15992), .Z(II15993) ) ;
NAND2   gate10244  (.A(g2677), .B(II15992), .Z(II15994) ) ;
NOR2    gate10245  (.A(g10290), .B(g4620), .Z(g10423) ) ;
NAND2   gate10246  (.A(g10423), .B(g2683), .Z(II15999) ) ;
NAND2   gate10247  (.A(g10423), .B(II15999), .Z(II16000) ) ;
NAND2   gate10248  (.A(g2683), .B(II15999), .Z(II16001) ) ;
NOR2    gate10249  (.A(g10349), .B(g3566), .Z(g10430) ) ;
NOR2    gate10250  (.A(g2753), .B(g4953), .Z(g5999) ) ;
NOR2    gate10251  (.A(g10292), .B(g4620), .Z(g10424) ) ;
NAND2   gate10252  (.A(g10424), .B(g2689), .Z(II16007) ) ;
NAND2   gate10253  (.A(g10424), .B(II16007), .Z(II16008) ) ;
NAND2   gate10254  (.A(g2689), .B(II16007), .Z(II16009) ) ;
NOR2    gate10255  (.A(g10293), .B(g4620), .Z(g10425) ) ;
NAND2   gate10256  (.A(g10425), .B(g2695), .Z(II16015) ) ;
NAND2   gate10257  (.A(g10425), .B(II16015), .Z(II16016) ) ;
NAND2   gate10258  (.A(g2695), .B(II16015), .Z(II16017) ) ;
NOR2    gate10259  (.A(g10294), .B(g4620), .Z(g10426) ) ;
NAND2   gate10260  (.A(g10426), .B(g2701), .Z(II16023) ) ;
NAND2   gate10261  (.A(g10426), .B(II16023), .Z(II16024) ) ;
NAND2   gate10262  (.A(g2701), .B(II16023), .Z(II16025) ) ;
NOR2    gate10263  (.A(g10342), .B(g3463), .Z(g10368) ) ;
NAND2   gate10264  (.A(g829), .B(g10368), .Z(II16030) ) ;
NAND2   gate10265  (.A(g829), .B(II16030), .Z(II16031) ) ;
NAND2   gate10266  (.A(g10368), .B(II16030), .Z(II16032) ) ;
NOR2    gate10267  (.A(g10296), .B(g4620), .Z(g10427) ) ;
NAND2   gate10268  (.A(g10427), .B(g2707), .Z(II16037) ) ;
NAND2   gate10269  (.A(g10427), .B(II16037), .Z(II16038) ) ;
NAND2   gate10270  (.A(g2707), .B(II16037), .Z(II16039) ) ;
NOR2    gate10271  (.A(g10343), .B(g3463), .Z(g10370) ) ;
NAND2   gate10272  (.A(g833), .B(g10370), .Z(II16044) ) ;
NAND2   gate10273  (.A(g833), .B(II16044), .Z(II16045) ) ;
NAND2   gate10274  (.A(g10370), .B(II16044), .Z(II16046) ) ;
NOR2    gate10275  (.A(g10344), .B(g3463), .Z(g10371) ) ;
NAND2   gate10276  (.A(g837), .B(g10371), .Z(II16051) ) ;
NAND2   gate10277  (.A(g837), .B(II16051), .Z(II16052) ) ;
NAND2   gate10278  (.A(g10371), .B(II16051), .Z(II16053) ) ;
NOR2    gate10279  (.A(g10345), .B(g3463), .Z(g10372) ) ;
NAND2   gate10280  (.A(g841), .B(g10372), .Z(II16058) ) ;
NAND2   gate10281  (.A(g841), .B(II16058), .Z(II16059) ) ;
NAND2   gate10282  (.A(g10372), .B(II16058), .Z(II16060) ) ;
NOR2    gate10283  (.A(g10335), .B(g4620), .Z(g10428) ) ;
NAND2   gate10284  (.A(g10428), .B(g2765), .Z(II16065) ) ;
NAND2   gate10285  (.A(g10428), .B(II16065), .Z(II16066) ) ;
NAND2   gate10286  (.A(g2765), .B(II16065), .Z(II16067) ) ;
NAND2   gate10287  (.A(II16066), .B(II16067), .Z(g10480) ) ;
NOR2    gate10288  (.A(g10346), .B(g3463), .Z(g10373) ) ;
NAND2   gate10289  (.A(g845), .B(g10373), .Z(II16072) ) ;
NAND2   gate10290  (.A(g845), .B(II16072), .Z(II16073) ) ;
NAND2   gate10291  (.A(g10373), .B(II16072), .Z(II16074) ) ;
NOR2    gate10292  (.A(g10347), .B(g3463), .Z(g10374) ) ;
NAND2   gate10293  (.A(g849), .B(g10374), .Z(II16079) ) ;
NAND2   gate10294  (.A(g849), .B(II16079), .Z(II16080) ) ;
NAND2   gate10295  (.A(g10374), .B(II16079), .Z(II16081) ) ;
NOR2    gate10296  (.A(g10288), .B(g3463), .Z(g10375) ) ;
NAND2   gate10297  (.A(g861), .B(g10375), .Z(II16086) ) ;
NAND2   gate10298  (.A(g861), .B(II16086), .Z(II16087) ) ;
NAND2   gate10299  (.A(g10375), .B(II16086), .Z(II16088) ) ;
NAND2   gate10300  (.A(II16087), .B(II16088), .Z(g10483) ) ;
NOR2    gate10301  (.A(g10350), .B(g3566), .Z(g10432) ) ;
NOR2    gate10302  (.A(g2764), .B(g4988), .Z(g5938) ) ;
NOR2    gate10303  (.A(g10352), .B(g3566), .Z(g10434) ) ;
NOR2    gate10304  (.A(g3362), .B(g4943), .Z(g5859) ) ;
NOR2    gate10305  (.A(g10354), .B(g3566), .Z(g10436) ) ;
NOR2    gate10306  (.A(g2763), .B(g4975), .Z(g6023) ) ;
NOR2    gate10307  (.A(g10356), .B(g3566), .Z(g10438) ) ;
NOR2    gate10308  (.A(g3430), .B(g5039), .Z(g6032) ) ;
NOR2    gate10309  (.A(g10351), .B(g3566), .Z(g10441) ) ;
NOR2    gate10310  (.A(g2754), .B(g4835), .Z(g5345) ) ;
NAND2   gate10311  (.A(g10616), .B(g4997), .Z(II16330) ) ;
NAND2   gate10312  (.A(g10616), .B(II16330), .Z(II16331) ) ;
NAND2   gate10313  (.A(g4997), .B(II16330), .Z(II16332) ) ;
NAND2   gate10314  (.A(g10716), .B(g10518), .Z(II16467) ) ;
NAND2   gate10315  (.A(g10716), .B(II16467), .Z(II16468) ) ;
NAND2   gate10316  (.A(g10518), .B(II16467), .Z(II16469) ) ;
NOR2    gate10317  (.A(g3524), .B(g4593), .Z(g5034) ) ;
NAND2   gate10318  (.A(g10923), .B(g11249), .Z(II17051) ) ;
NAND2   gate10319  (.A(g10923), .B(II17051), .Z(II17052) ) ;
NAND2   gate10320  (.A(g11249), .B(II17051), .Z(II17053) ) ;
NAND2   gate10321  (.A(g11360), .B(g11357), .Z(II17281) ) ;
NAND2   gate10322  (.A(g11360), .B(II17281), .Z(II17282) ) ;
NAND2   gate10323  (.A(g11357), .B(II17281), .Z(II17283) ) ;
NAND2   gate10324  (.A(II17282), .B(II17283), .Z(g11414) ) ;
NAND2   gate10325  (.A(g11366), .B(g11363), .Z(II17288) ) ;
NAND2   gate10326  (.A(g11366), .B(II17288), .Z(II17289) ) ;
NAND2   gate10327  (.A(g11363), .B(II17288), .Z(II17290) ) ;
NAND2   gate10328  (.A(II17289), .B(II17290), .Z(g11415) ) ;
NAND2   gate10329  (.A(g11373), .B(g11369), .Z(II17295) ) ;
NAND2   gate10330  (.A(g11373), .B(II17295), .Z(II17296) ) ;
NAND2   gate10331  (.A(g11369), .B(II17295), .Z(II17297) ) ;
NAND2   gate10332  (.A(II17296), .B(II17297), .Z(g11416) ) ;
NAND2   gate10333  (.A(g11381), .B(g11377), .Z(II17305) ) ;
NAND2   gate10334  (.A(g11381), .B(II17305), .Z(II17306) ) ;
NAND2   gate10335  (.A(g11377), .B(II17305), .Z(II17307) ) ;
NAND2   gate10336  (.A(II17306), .B(II17307), .Z(g11418) ) ;
NAND2   gate10337  (.A(g11415), .B(g11414), .Z(II17393) ) ;
NAND2   gate10338  (.A(g11415), .B(II17393), .Z(II17394) ) ;
NAND2   gate10339  (.A(g11414), .B(II17393), .Z(II17395) ) ;
NAND2   gate10340  (.A(II17394), .B(II17395), .Z(g11448) ) ;
NAND2   gate10341  (.A(g11418), .B(g11416), .Z(II17400) ) ;
NAND2   gate10342  (.A(g11418), .B(II17400), .Z(II17401) ) ;
NAND2   gate10343  (.A(g11416), .B(II17400), .Z(II17402) ) ;
NAND2   gate10344  (.A(II17401), .B(II17402), .Z(g11449) ) ;
NAND2   gate10345  (.A(g11449), .B(g11448), .Z(II17459) ) ;
NAND2   gate10346  (.A(g11449), .B(II17459), .Z(II17460) ) ;
NAND2   gate10347  (.A(g11448), .B(II17459), .Z(II17461) ) ;
NAND2   gate10348  (.A(II17460), .B(II17461), .Z(g11474) ) ;
NAND2   gate10349  (.A(g11384), .B(g11474), .Z(II17485) ) ;
NAND2   gate10350  (.A(g11384), .B(II17485), .Z(II17486) ) ;
NAND2   gate10351  (.A(g11474), .B(II17485), .Z(II17487) ) ;
NAND2   gate10352  (.A(g11475), .B(g3623), .Z(II17492) ) ;
NAND2   gate10353  (.A(g11475), .B(II17492), .Z(II17493) ) ;
NAND2   gate10354  (.A(g3623), .B(II17492), .Z(II17494) ) ;
NAND2   gate10355  (.A(g11475), .B(g7603), .Z(II17503) ) ;
NAND2   gate10356  (.A(g11475), .B(II17503), .Z(II17504) ) ;
NAND2   gate10357  (.A(g7603), .B(II17503), .Z(II17505) ) ;
NAND2   gate10358  (.A(II17504), .B(II17505), .Z(g11496) ) ;
NAND2   gate10359  (.A(g11496), .B(g1610), .Z(II17567) ) ;
NAND2   gate10360  (.A(g11496), .B(II17567), .Z(II17568) ) ;
NAND2   gate10361  (.A(g1610), .B(II17567), .Z(II17569) ) ;
NAND2   gate10362  (.A(g11354), .B(g11515), .Z(II17584) ) ;
NAND2   gate10363  (.A(g11354), .B(II17584), .Z(II17585) ) ;
NAND2   gate10364  (.A(g11515), .B(II17584), .Z(II17586) ) ;
NOR2    gate10365  (.A(g4502), .B(g3714), .Z(g4974) ) ;
NOR2    gate10366  (.A(g9317), .B(g10179), .Z(g10239) ) ;
NOR2    gate10367  (.A(g9317), .B(g10272), .Z(g10322) ) ;
NOR2    gate10368  (.A(g9317), .B(g10244), .Z(g10324) ) ;

endmodule
