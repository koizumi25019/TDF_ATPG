module s35932 (DATA_0_31, DATA_0_30, DATA_0_29, DATA_0_28, DATA_0_27
    , DATA_0_26, DATA_0_25, DATA_0_24, DATA_0_23, DATA_0_22
    , DATA_0_21, DATA_0_20, DATA_0_19, DATA_0_18, DATA_0_17
    , DATA_0_16, DATA_0_15, DATA_0_14, DATA_0_13, DATA_0_12
    , DATA_0_11, DATA_0_10, DATA_0_9, DATA_0_8, DATA_0_7
    , DATA_0_6, DATA_0_5, DATA_0_4, DATA_0_3, DATA_0_2
    , DATA_0_1, DATA_0_0, RESET, TM1, TM0
    , CLK
    , DATA_9_31, DATA_9_30, DATA_9_29, DATA_9_28, DATA_9_27
    , DATA_9_26, DATA_9_25, DATA_9_24, DATA_9_23, DATA_9_22
    , DATA_9_21, DATA_9_20, DATA_9_19, DATA_9_18, DATA_9_17
    , DATA_9_16, DATA_9_15, DATA_9_14, DATA_9_13, DATA_9_12
    , DATA_9_11, DATA_9_10, DATA_9_9, DATA_9_8, DATA_9_7
    , DATA_9_6, DATA_9_5, DATA_9_4, DATA_9_3, DATA_9_2
    , DATA_9_1, DATA_9_0, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_2
    , CRC_OUT_9_3, CRC_OUT_9_4, CRC_OUT_9_5, CRC_OUT_9_6, CRC_OUT_9_7
    , CRC_OUT_9_8, CRC_OUT_9_9, CRC_OUT_9_10, CRC_OUT_9_11, CRC_OUT_9_12
    , CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, CRC_OUT_9_16, CRC_OUT_9_17
    , CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_20, CRC_OUT_9_21, CRC_OUT_9_22
    , CRC_OUT_9_23, CRC_OUT_9_24, CRC_OUT_9_25, CRC_OUT_9_26, CRC_OUT_9_27
    , CRC_OUT_9_28, CRC_OUT_9_29, CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_8_0
    , CRC_OUT_8_1, CRC_OUT_8_2, CRC_OUT_8_3, CRC_OUT_8_4, CRC_OUT_8_5
    , CRC_OUT_8_6, CRC_OUT_8_7, CRC_OUT_8_8, CRC_OUT_8_9, CRC_OUT_8_10
    , CRC_OUT_8_11, CRC_OUT_8_12, CRC_OUT_8_13, CRC_OUT_8_14, CRC_OUT_8_15
    , CRC_OUT_8_16, CRC_OUT_8_17, CRC_OUT_8_18, CRC_OUT_8_19, CRC_OUT_8_20
    , CRC_OUT_8_21, CRC_OUT_8_22, CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25
    , CRC_OUT_8_26, CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_30
    , CRC_OUT_8_31, CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_2, CRC_OUT_7_3
    , CRC_OUT_7_4, CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8
    , CRC_OUT_7_9, CRC_OUT_7_10, CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13
    , CRC_OUT_7_14, CRC_OUT_7_15, CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18
    , CRC_OUT_7_19, CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23
    , CRC_OUT_7_24, CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28
    , CRC_OUT_7_29, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_6_0, CRC_OUT_6_1
    , CRC_OUT_6_2, CRC_OUT_6_3, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6
    , CRC_OUT_6_7, CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_6_10, CRC_OUT_6_11
    , CRC_OUT_6_12, CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16
    , CRC_OUT_6_17, CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_20, CRC_OUT_6_21
    , CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, CRC_OUT_6_26
    , CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_30, CRC_OUT_6_31
    , CRC_OUT_5_0, CRC_OUT_5_1, CRC_OUT_5_2, CRC_OUT_5_3, CRC_OUT_5_4
    , CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, CRC_OUT_5_9
    , CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, CRC_OUT_5_14
    , CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, CRC_OUT_5_19
    , CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, CRC_OUT_5_23, CRC_OUT_5_24
    , CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, CRC_OUT_5_28, CRC_OUT_5_29
    , CRC_OUT_5_30, CRC_OUT_5_31, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_2
    , CRC_OUT_4_3, CRC_OUT_4_4, CRC_OUT_4_5, CRC_OUT_4_6, CRC_OUT_4_7
    , CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_4_10, CRC_OUT_4_11, CRC_OUT_4_12
    , CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, CRC_OUT_4_16, CRC_OUT_4_17
    , CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_20, CRC_OUT_4_21, CRC_OUT_4_22
    , CRC_OUT_4_23, CRC_OUT_4_24, CRC_OUT_4_25, CRC_OUT_4_26, CRC_OUT_4_27
    , CRC_OUT_4_28, CRC_OUT_4_29, CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_3_0
    , CRC_OUT_3_1, CRC_OUT_3_2, CRC_OUT_3_3, CRC_OUT_3_4, CRC_OUT_3_5
    , CRC_OUT_3_6, CRC_OUT_3_7, CRC_OUT_3_8, CRC_OUT_3_9, CRC_OUT_3_10
    , CRC_OUT_3_11, CRC_OUT_3_12, CRC_OUT_3_13, CRC_OUT_3_14, CRC_OUT_3_15
    , CRC_OUT_3_16, CRC_OUT_3_17, CRC_OUT_3_18, CRC_OUT_3_19, CRC_OUT_3_20
    , CRC_OUT_3_21, CRC_OUT_3_22, CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25
    , CRC_OUT_3_26, CRC_OUT_3_27, CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_30
    , CRC_OUT_3_31, CRC_OUT_2_0, CRC_OUT_2_1, CRC_OUT_2_2, CRC_OUT_2_3
    , CRC_OUT_2_4, CRC_OUT_2_5, CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8
    , CRC_OUT_2_9, CRC_OUT_2_10, CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13
    , CRC_OUT_2_14, CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18
    , CRC_OUT_2_19, CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23
    , CRC_OUT_2_24, CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28
    , CRC_OUT_2_29, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_1_0, CRC_OUT_1_1
    , CRC_OUT_1_2, CRC_OUT_1_3, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6
    , CRC_OUT_1_7, CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_1_10, CRC_OUT_1_11
    , CRC_OUT_1_12, CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16
    , CRC_OUT_1_17, CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_20, CRC_OUT_1_21
    , CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, CRC_OUT_1_26
    , CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_30, CRC_OUT_1_31
    ) ;

input   DATA_0_31, DATA_0_30, DATA_0_29, DATA_0_28, DATA_0_27
    , DATA_0_26, DATA_0_25, DATA_0_24, DATA_0_23, DATA_0_22
    , DATA_0_21, DATA_0_20, DATA_0_19, DATA_0_18, DATA_0_17
    , DATA_0_16, DATA_0_15, DATA_0_14, DATA_0_13, DATA_0_12
    , DATA_0_11, DATA_0_10, DATA_0_9, DATA_0_8, DATA_0_7
    , DATA_0_6, DATA_0_5, DATA_0_4, DATA_0_3, DATA_0_2
    , DATA_0_1, DATA_0_0, RESET, TM1, TM0
    , CLK ;

output  DATA_9_31, DATA_9_30, DATA_9_29, DATA_9_28, DATA_9_27
    , DATA_9_26, DATA_9_25, DATA_9_24, DATA_9_23, DATA_9_22
    , DATA_9_21, DATA_9_20, DATA_9_19, DATA_9_18, DATA_9_17
    , DATA_9_16, DATA_9_15, DATA_9_14, DATA_9_13, DATA_9_12
    , DATA_9_11, DATA_9_10, DATA_9_9, DATA_9_8, DATA_9_7
    , DATA_9_6, DATA_9_5, DATA_9_4, DATA_9_3, DATA_9_2
    , DATA_9_1, DATA_9_0, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_2
    , CRC_OUT_9_3, CRC_OUT_9_4, CRC_OUT_9_5, CRC_OUT_9_6, CRC_OUT_9_7
    , CRC_OUT_9_8, CRC_OUT_9_9, CRC_OUT_9_10, CRC_OUT_9_11, CRC_OUT_9_12
    , CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, CRC_OUT_9_16, CRC_OUT_9_17
    , CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_20, CRC_OUT_9_21, CRC_OUT_9_22
    , CRC_OUT_9_23, CRC_OUT_9_24, CRC_OUT_9_25, CRC_OUT_9_26, CRC_OUT_9_27
    , CRC_OUT_9_28, CRC_OUT_9_29, CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_8_0
    , CRC_OUT_8_1, CRC_OUT_8_2, CRC_OUT_8_3, CRC_OUT_8_4, CRC_OUT_8_5
    , CRC_OUT_8_6, CRC_OUT_8_7, CRC_OUT_8_8, CRC_OUT_8_9, CRC_OUT_8_10
    , CRC_OUT_8_11, CRC_OUT_8_12, CRC_OUT_8_13, CRC_OUT_8_14, CRC_OUT_8_15
    , CRC_OUT_8_16, CRC_OUT_8_17, CRC_OUT_8_18, CRC_OUT_8_19, CRC_OUT_8_20
    , CRC_OUT_8_21, CRC_OUT_8_22, CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25
    , CRC_OUT_8_26, CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_30
    , CRC_OUT_8_31, CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_2, CRC_OUT_7_3
    , CRC_OUT_7_4, CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8
    , CRC_OUT_7_9, CRC_OUT_7_10, CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13
    , CRC_OUT_7_14, CRC_OUT_7_15, CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18
    , CRC_OUT_7_19, CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23
    , CRC_OUT_7_24, CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28
    , CRC_OUT_7_29, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_6_0, CRC_OUT_6_1
    , CRC_OUT_6_2, CRC_OUT_6_3, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6
    , CRC_OUT_6_7, CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_6_10, CRC_OUT_6_11
    , CRC_OUT_6_12, CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16
    , CRC_OUT_6_17, CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_20, CRC_OUT_6_21
    , CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, CRC_OUT_6_26
    , CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_30, CRC_OUT_6_31
    , CRC_OUT_5_0, CRC_OUT_5_1, CRC_OUT_5_2, CRC_OUT_5_3, CRC_OUT_5_4
    , CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, CRC_OUT_5_9
    , CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, CRC_OUT_5_14
    , CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, CRC_OUT_5_19
    , CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, CRC_OUT_5_23, CRC_OUT_5_24
    , CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, CRC_OUT_5_28, CRC_OUT_5_29
    , CRC_OUT_5_30, CRC_OUT_5_31, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_2
    , CRC_OUT_4_3, CRC_OUT_4_4, CRC_OUT_4_5, CRC_OUT_4_6, CRC_OUT_4_7
    , CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_4_10, CRC_OUT_4_11, CRC_OUT_4_12
    , CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, CRC_OUT_4_16, CRC_OUT_4_17
    , CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_20, CRC_OUT_4_21, CRC_OUT_4_22
    , CRC_OUT_4_23, CRC_OUT_4_24, CRC_OUT_4_25, CRC_OUT_4_26, CRC_OUT_4_27
    , CRC_OUT_4_28, CRC_OUT_4_29, CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_3_0
    , CRC_OUT_3_1, CRC_OUT_3_2, CRC_OUT_3_3, CRC_OUT_3_4, CRC_OUT_3_5
    , CRC_OUT_3_6, CRC_OUT_3_7, CRC_OUT_3_8, CRC_OUT_3_9, CRC_OUT_3_10
    , CRC_OUT_3_11, CRC_OUT_3_12, CRC_OUT_3_13, CRC_OUT_3_14, CRC_OUT_3_15
    , CRC_OUT_3_16, CRC_OUT_3_17, CRC_OUT_3_18, CRC_OUT_3_19, CRC_OUT_3_20
    , CRC_OUT_3_21, CRC_OUT_3_22, CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25
    , CRC_OUT_3_26, CRC_OUT_3_27, CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_30
    , CRC_OUT_3_31, CRC_OUT_2_0, CRC_OUT_2_1, CRC_OUT_2_2, CRC_OUT_2_3
    , CRC_OUT_2_4, CRC_OUT_2_5, CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8
    , CRC_OUT_2_9, CRC_OUT_2_10, CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13
    , CRC_OUT_2_14, CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18
    , CRC_OUT_2_19, CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23
    , CRC_OUT_2_24, CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28
    , CRC_OUT_2_29, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_1_0, CRC_OUT_1_1
    , CRC_OUT_1_2, CRC_OUT_1_3, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6
    , CRC_OUT_1_7, CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_1_10, CRC_OUT_1_11
    , CRC_OUT_1_12, CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16
    , CRC_OUT_1_17, CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_20, CRC_OUT_1_21
    , CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, CRC_OUT_1_26
    , CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_30, CRC_OUT_1_31
     ;

INV     gate0  (.A(WX1011), .Z(DATA_9_31) ) ;
INV     gate1  (.A(WX1018), .Z(DATA_9_30) ) ;
INV     gate2  (.A(WX1025), .Z(DATA_9_29) ) ;
INV     gate3  (.A(WX1032), .Z(DATA_9_28) ) ;
INV     gate4  (.A(WX1039), .Z(DATA_9_27) ) ;
INV     gate5  (.A(WX1046), .Z(DATA_9_26) ) ;
INV     gate6  (.A(WX1053), .Z(DATA_9_25) ) ;
INV     gate7  (.A(WX1060), .Z(DATA_9_24) ) ;
INV     gate8  (.A(WX1067), .Z(DATA_9_23) ) ;
INV     gate9  (.A(WX1074), .Z(DATA_9_22) ) ;
INV     gate10  (.A(WX1081), .Z(DATA_9_21) ) ;
INV     gate11  (.A(WX1088), .Z(DATA_9_20) ) ;
INV     gate12  (.A(WX1095), .Z(DATA_9_19) ) ;
INV     gate13  (.A(WX1102), .Z(DATA_9_18) ) ;
INV     gate14  (.A(WX1109), .Z(DATA_9_17) ) ;
INV     gate15  (.A(WX1116), .Z(DATA_9_16) ) ;
INV     gate16  (.A(WX1123), .Z(DATA_9_15) ) ;
INV     gate17  (.A(WX1130), .Z(DATA_9_14) ) ;
INV     gate18  (.A(WX1137), .Z(DATA_9_13) ) ;
INV     gate19  (.A(WX1144), .Z(DATA_9_12) ) ;
INV     gate20  (.A(WX1151), .Z(DATA_9_11) ) ;
INV     gate21  (.A(WX1158), .Z(DATA_9_10) ) ;
INV     gate22  (.A(WX1165), .Z(DATA_9_9) ) ;
INV     gate23  (.A(WX1172), .Z(DATA_9_8) ) ;
INV     gate24  (.A(WX1179), .Z(DATA_9_7) ) ;
INV     gate25  (.A(WX1186), .Z(DATA_9_6) ) ;
INV     gate26  (.A(WX1193), .Z(DATA_9_5) ) ;
INV     gate27  (.A(WX1200), .Z(DATA_9_4) ) ;
INV     gate28  (.A(WX1207), .Z(DATA_9_3) ) ;
INV     gate29  (.A(WX1214), .Z(DATA_9_2) ) ;
INV     gate30  (.A(WX1221), .Z(DATA_9_1) ) ;
INV     gate31  (.A(WX1228), .Z(DATA_9_0) ) ;
DFF     gate32  (.D(WX1264), .CP(CLK), .Q(CRC_OUT_9_0) ) ;
DFF     gate33  (.D(WX1266), .CP(CLK), .Q(CRC_OUT_9_1) ) ;
DFF     gate34  (.D(WX1268), .CP(CLK), .Q(CRC_OUT_9_2) ) ;
DFF     gate35  (.D(WX1270), .CP(CLK), .Q(CRC_OUT_9_3) ) ;
DFF     gate36  (.D(WX1272), .CP(CLK), .Q(CRC_OUT_9_4) ) ;
DFF     gate37  (.D(WX1274), .CP(CLK), .Q(CRC_OUT_9_5) ) ;
DFF     gate38  (.D(WX1276), .CP(CLK), .Q(CRC_OUT_9_6) ) ;
DFF     gate39  (.D(WX1278), .CP(CLK), .Q(CRC_OUT_9_7) ) ;
DFF     gate40  (.D(WX1280), .CP(CLK), .Q(CRC_OUT_9_8) ) ;
DFF     gate41  (.D(WX1282), .CP(CLK), .Q(CRC_OUT_9_9) ) ;
DFF     gate42  (.D(WX1284), .CP(CLK), .Q(CRC_OUT_9_10) ) ;
DFF     gate43  (.D(WX1286), .CP(CLK), .Q(CRC_OUT_9_11) ) ;
DFF     gate44  (.D(WX1288), .CP(CLK), .Q(CRC_OUT_9_12) ) ;
DFF     gate45  (.D(WX1290), .CP(CLK), .Q(CRC_OUT_9_13) ) ;
DFF     gate46  (.D(WX1292), .CP(CLK), .Q(CRC_OUT_9_14) ) ;
DFF     gate47  (.D(WX1294), .CP(CLK), .Q(CRC_OUT_9_15) ) ;
DFF     gate48  (.D(WX1296), .CP(CLK), .Q(CRC_OUT_9_16) ) ;
DFF     gate49  (.D(WX1298), .CP(CLK), .Q(CRC_OUT_9_17) ) ;
DFF     gate50  (.D(WX1300), .CP(CLK), .Q(CRC_OUT_9_18) ) ;
DFF     gate51  (.D(WX1302), .CP(CLK), .Q(CRC_OUT_9_19) ) ;
DFF     gate52  (.D(WX1304), .CP(CLK), .Q(CRC_OUT_9_20) ) ;
DFF     gate53  (.D(WX1306), .CP(CLK), .Q(CRC_OUT_9_21) ) ;
DFF     gate54  (.D(WX1308), .CP(CLK), .Q(CRC_OUT_9_22) ) ;
DFF     gate55  (.D(WX1310), .CP(CLK), .Q(CRC_OUT_9_23) ) ;
DFF     gate56  (.D(WX1312), .CP(CLK), .Q(CRC_OUT_9_24) ) ;
DFF     gate57  (.D(WX1314), .CP(CLK), .Q(CRC_OUT_9_25) ) ;
DFF     gate58  (.D(WX1316), .CP(CLK), .Q(CRC_OUT_9_26) ) ;
DFF     gate59  (.D(WX1318), .CP(CLK), .Q(CRC_OUT_9_27) ) ;
DFF     gate60  (.D(WX1320), .CP(CLK), .Q(CRC_OUT_9_28) ) ;
DFF     gate61  (.D(WX1322), .CP(CLK), .Q(CRC_OUT_9_29) ) ;
DFF     gate62  (.D(WX1324), .CP(CLK), .Q(CRC_OUT_9_30) ) ;
DFF     gate63  (.D(WX1326), .CP(CLK), .Q(CRC_OUT_9_31) ) ;
DFF     gate64  (.D(WX2557), .CP(CLK), .Q(CRC_OUT_8_0) ) ;
DFF     gate65  (.D(WX2559), .CP(CLK), .Q(CRC_OUT_8_1) ) ;
DFF     gate66  (.D(WX2561), .CP(CLK), .Q(CRC_OUT_8_2) ) ;
DFF     gate67  (.D(WX2563), .CP(CLK), .Q(CRC_OUT_8_3) ) ;
DFF     gate68  (.D(WX2565), .CP(CLK), .Q(CRC_OUT_8_4) ) ;
DFF     gate69  (.D(WX2567), .CP(CLK), .Q(CRC_OUT_8_5) ) ;
DFF     gate70  (.D(WX2569), .CP(CLK), .Q(CRC_OUT_8_6) ) ;
DFF     gate71  (.D(WX2571), .CP(CLK), .Q(CRC_OUT_8_7) ) ;
DFF     gate72  (.D(WX2573), .CP(CLK), .Q(CRC_OUT_8_8) ) ;
DFF     gate73  (.D(WX2575), .CP(CLK), .Q(CRC_OUT_8_9) ) ;
DFF     gate74  (.D(WX2577), .CP(CLK), .Q(CRC_OUT_8_10) ) ;
DFF     gate75  (.D(WX2579), .CP(CLK), .Q(CRC_OUT_8_11) ) ;
DFF     gate76  (.D(WX2581), .CP(CLK), .Q(CRC_OUT_8_12) ) ;
DFF     gate77  (.D(WX2583), .CP(CLK), .Q(CRC_OUT_8_13) ) ;
DFF     gate78  (.D(WX2585), .CP(CLK), .Q(CRC_OUT_8_14) ) ;
DFF     gate79  (.D(WX2587), .CP(CLK), .Q(CRC_OUT_8_15) ) ;
DFF     gate80  (.D(WX2589), .CP(CLK), .Q(CRC_OUT_8_16) ) ;
DFF     gate81  (.D(WX2591), .CP(CLK), .Q(CRC_OUT_8_17) ) ;
DFF     gate82  (.D(WX2593), .CP(CLK), .Q(CRC_OUT_8_18) ) ;
DFF     gate83  (.D(WX2595), .CP(CLK), .Q(CRC_OUT_8_19) ) ;
DFF     gate84  (.D(WX2597), .CP(CLK), .Q(CRC_OUT_8_20) ) ;
DFF     gate85  (.D(WX2599), .CP(CLK), .Q(CRC_OUT_8_21) ) ;
DFF     gate86  (.D(WX2601), .CP(CLK), .Q(CRC_OUT_8_22) ) ;
DFF     gate87  (.D(WX2603), .CP(CLK), .Q(CRC_OUT_8_23) ) ;
DFF     gate88  (.D(WX2605), .CP(CLK), .Q(CRC_OUT_8_24) ) ;
DFF     gate89  (.D(WX2607), .CP(CLK), .Q(CRC_OUT_8_25) ) ;
DFF     gate90  (.D(WX2609), .CP(CLK), .Q(CRC_OUT_8_26) ) ;
DFF     gate91  (.D(WX2611), .CP(CLK), .Q(CRC_OUT_8_27) ) ;
DFF     gate92  (.D(WX2613), .CP(CLK), .Q(CRC_OUT_8_28) ) ;
DFF     gate93  (.D(WX2615), .CP(CLK), .Q(CRC_OUT_8_29) ) ;
DFF     gate94  (.D(WX2617), .CP(CLK), .Q(CRC_OUT_8_30) ) ;
DFF     gate95  (.D(WX2619), .CP(CLK), .Q(CRC_OUT_8_31) ) ;
DFF     gate96  (.D(WX3850), .CP(CLK), .Q(CRC_OUT_7_0) ) ;
DFF     gate97  (.D(WX3852), .CP(CLK), .Q(CRC_OUT_7_1) ) ;
DFF     gate98  (.D(WX3854), .CP(CLK), .Q(CRC_OUT_7_2) ) ;
DFF     gate99  (.D(WX3856), .CP(CLK), .Q(CRC_OUT_7_3) ) ;
DFF     gate100  (.D(WX3858), .CP(CLK), .Q(CRC_OUT_7_4) ) ;
DFF     gate101  (.D(WX3860), .CP(CLK), .Q(CRC_OUT_7_5) ) ;
DFF     gate102  (.D(WX3862), .CP(CLK), .Q(CRC_OUT_7_6) ) ;
DFF     gate103  (.D(WX3864), .CP(CLK), .Q(CRC_OUT_7_7) ) ;
DFF     gate104  (.D(WX3866), .CP(CLK), .Q(CRC_OUT_7_8) ) ;
DFF     gate105  (.D(WX3868), .CP(CLK), .Q(CRC_OUT_7_9) ) ;
DFF     gate106  (.D(WX3870), .CP(CLK), .Q(CRC_OUT_7_10) ) ;
DFF     gate107  (.D(WX3872), .CP(CLK), .Q(CRC_OUT_7_11) ) ;
DFF     gate108  (.D(WX3874), .CP(CLK), .Q(CRC_OUT_7_12) ) ;
DFF     gate109  (.D(WX3876), .CP(CLK), .Q(CRC_OUT_7_13) ) ;
DFF     gate110  (.D(WX3878), .CP(CLK), .Q(CRC_OUT_7_14) ) ;
DFF     gate111  (.D(WX3880), .CP(CLK), .Q(CRC_OUT_7_15) ) ;
DFF     gate112  (.D(WX3882), .CP(CLK), .Q(CRC_OUT_7_16) ) ;
DFF     gate113  (.D(WX3884), .CP(CLK), .Q(CRC_OUT_7_17) ) ;
DFF     gate114  (.D(WX3886), .CP(CLK), .Q(CRC_OUT_7_18) ) ;
DFF     gate115  (.D(WX3888), .CP(CLK), .Q(CRC_OUT_7_19) ) ;
DFF     gate116  (.D(WX3890), .CP(CLK), .Q(CRC_OUT_7_20) ) ;
DFF     gate117  (.D(WX3892), .CP(CLK), .Q(CRC_OUT_7_21) ) ;
DFF     gate118  (.D(WX3894), .CP(CLK), .Q(CRC_OUT_7_22) ) ;
DFF     gate119  (.D(WX3896), .CP(CLK), .Q(CRC_OUT_7_23) ) ;
DFF     gate120  (.D(WX3898), .CP(CLK), .Q(CRC_OUT_7_24) ) ;
DFF     gate121  (.D(WX3900), .CP(CLK), .Q(CRC_OUT_7_25) ) ;
DFF     gate122  (.D(WX3902), .CP(CLK), .Q(CRC_OUT_7_26) ) ;
DFF     gate123  (.D(WX3904), .CP(CLK), .Q(CRC_OUT_7_27) ) ;
DFF     gate124  (.D(WX3906), .CP(CLK), .Q(CRC_OUT_7_28) ) ;
DFF     gate125  (.D(WX3908), .CP(CLK), .Q(CRC_OUT_7_29) ) ;
DFF     gate126  (.D(WX3910), .CP(CLK), .Q(CRC_OUT_7_30) ) ;
DFF     gate127  (.D(WX3912), .CP(CLK), .Q(CRC_OUT_7_31) ) ;
DFF     gate128  (.D(WX5143), .CP(CLK), .Q(CRC_OUT_6_0) ) ;
DFF     gate129  (.D(WX5145), .CP(CLK), .Q(CRC_OUT_6_1) ) ;
DFF     gate130  (.D(WX5147), .CP(CLK), .Q(CRC_OUT_6_2) ) ;
DFF     gate131  (.D(WX5149), .CP(CLK), .Q(CRC_OUT_6_3) ) ;
DFF     gate132  (.D(WX5151), .CP(CLK), .Q(CRC_OUT_6_4) ) ;
DFF     gate133  (.D(WX5153), .CP(CLK), .Q(CRC_OUT_6_5) ) ;
DFF     gate134  (.D(WX5155), .CP(CLK), .Q(CRC_OUT_6_6) ) ;
DFF     gate135  (.D(WX5157), .CP(CLK), .Q(CRC_OUT_6_7) ) ;
DFF     gate136  (.D(WX5159), .CP(CLK), .Q(CRC_OUT_6_8) ) ;
DFF     gate137  (.D(WX5161), .CP(CLK), .Q(CRC_OUT_6_9) ) ;
DFF     gate138  (.D(WX5163), .CP(CLK), .Q(CRC_OUT_6_10) ) ;
DFF     gate139  (.D(WX5165), .CP(CLK), .Q(CRC_OUT_6_11) ) ;
DFF     gate140  (.D(WX5167), .CP(CLK), .Q(CRC_OUT_6_12) ) ;
DFF     gate141  (.D(WX5169), .CP(CLK), .Q(CRC_OUT_6_13) ) ;
DFF     gate142  (.D(WX5171), .CP(CLK), .Q(CRC_OUT_6_14) ) ;
DFF     gate143  (.D(WX5173), .CP(CLK), .Q(CRC_OUT_6_15) ) ;
DFF     gate144  (.D(WX5175), .CP(CLK), .Q(CRC_OUT_6_16) ) ;
DFF     gate145  (.D(WX5177), .CP(CLK), .Q(CRC_OUT_6_17) ) ;
DFF     gate146  (.D(WX5179), .CP(CLK), .Q(CRC_OUT_6_18) ) ;
DFF     gate147  (.D(WX5181), .CP(CLK), .Q(CRC_OUT_6_19) ) ;
DFF     gate148  (.D(WX5183), .CP(CLK), .Q(CRC_OUT_6_20) ) ;
DFF     gate149  (.D(WX5185), .CP(CLK), .Q(CRC_OUT_6_21) ) ;
DFF     gate150  (.D(WX5187), .CP(CLK), .Q(CRC_OUT_6_22) ) ;
DFF     gate151  (.D(WX5189), .CP(CLK), .Q(CRC_OUT_6_23) ) ;
DFF     gate152  (.D(WX5191), .CP(CLK), .Q(CRC_OUT_6_24) ) ;
DFF     gate153  (.D(WX5193), .CP(CLK), .Q(CRC_OUT_6_25) ) ;
DFF     gate154  (.D(WX5195), .CP(CLK), .Q(CRC_OUT_6_26) ) ;
DFF     gate155  (.D(WX5197), .CP(CLK), .Q(CRC_OUT_6_27) ) ;
DFF     gate156  (.D(WX5199), .CP(CLK), .Q(CRC_OUT_6_28) ) ;
DFF     gate157  (.D(WX5201), .CP(CLK), .Q(CRC_OUT_6_29) ) ;
DFF     gate158  (.D(WX5203), .CP(CLK), .Q(CRC_OUT_6_30) ) ;
DFF     gate159  (.D(WX5205), .CP(CLK), .Q(CRC_OUT_6_31) ) ;
DFF     gate160  (.D(WX6436), .CP(CLK), .Q(CRC_OUT_5_0) ) ;
DFF     gate161  (.D(WX6438), .CP(CLK), .Q(CRC_OUT_5_1) ) ;
DFF     gate162  (.D(WX6440), .CP(CLK), .Q(CRC_OUT_5_2) ) ;
DFF     gate163  (.D(WX6442), .CP(CLK), .Q(CRC_OUT_5_3) ) ;
DFF     gate164  (.D(WX6444), .CP(CLK), .Q(CRC_OUT_5_4) ) ;
DFF     gate165  (.D(WX6446), .CP(CLK), .Q(CRC_OUT_5_5) ) ;
DFF     gate166  (.D(WX6448), .CP(CLK), .Q(CRC_OUT_5_6) ) ;
DFF     gate167  (.D(WX6450), .CP(CLK), .Q(CRC_OUT_5_7) ) ;
DFF     gate168  (.D(WX6452), .CP(CLK), .Q(CRC_OUT_5_8) ) ;
DFF     gate169  (.D(WX6454), .CP(CLK), .Q(CRC_OUT_5_9) ) ;
DFF     gate170  (.D(WX6456), .CP(CLK), .Q(CRC_OUT_5_10) ) ;
DFF     gate171  (.D(WX6458), .CP(CLK), .Q(CRC_OUT_5_11) ) ;
DFF     gate172  (.D(WX6460), .CP(CLK), .Q(CRC_OUT_5_12) ) ;
DFF     gate173  (.D(WX6462), .CP(CLK), .Q(CRC_OUT_5_13) ) ;
DFF     gate174  (.D(WX6464), .CP(CLK), .Q(CRC_OUT_5_14) ) ;
DFF     gate175  (.D(WX6466), .CP(CLK), .Q(CRC_OUT_5_15) ) ;
DFF     gate176  (.D(WX6468), .CP(CLK), .Q(CRC_OUT_5_16) ) ;
DFF     gate177  (.D(WX6470), .CP(CLK), .Q(CRC_OUT_5_17) ) ;
DFF     gate178  (.D(WX6472), .CP(CLK), .Q(CRC_OUT_5_18) ) ;
DFF     gate179  (.D(WX6474), .CP(CLK), .Q(CRC_OUT_5_19) ) ;
DFF     gate180  (.D(WX6476), .CP(CLK), .Q(CRC_OUT_5_20) ) ;
DFF     gate181  (.D(WX6478), .CP(CLK), .Q(CRC_OUT_5_21) ) ;
DFF     gate182  (.D(WX6480), .CP(CLK), .Q(CRC_OUT_5_22) ) ;
DFF     gate183  (.D(WX6482), .CP(CLK), .Q(CRC_OUT_5_23) ) ;
DFF     gate184  (.D(WX6484), .CP(CLK), .Q(CRC_OUT_5_24) ) ;
DFF     gate185  (.D(WX6486), .CP(CLK), .Q(CRC_OUT_5_25) ) ;
DFF     gate186  (.D(WX6488), .CP(CLK), .Q(CRC_OUT_5_26) ) ;
DFF     gate187  (.D(WX6490), .CP(CLK), .Q(CRC_OUT_5_27) ) ;
DFF     gate188  (.D(WX6492), .CP(CLK), .Q(CRC_OUT_5_28) ) ;
DFF     gate189  (.D(WX6494), .CP(CLK), .Q(CRC_OUT_5_29) ) ;
DFF     gate190  (.D(WX6496), .CP(CLK), .Q(CRC_OUT_5_30) ) ;
DFF     gate191  (.D(WX6498), .CP(CLK), .Q(CRC_OUT_5_31) ) ;
DFF     gate192  (.D(WX7729), .CP(CLK), .Q(CRC_OUT_4_0) ) ;
DFF     gate193  (.D(WX7731), .CP(CLK), .Q(CRC_OUT_4_1) ) ;
DFF     gate194  (.D(WX7733), .CP(CLK), .Q(CRC_OUT_4_2) ) ;
DFF     gate195  (.D(WX7735), .CP(CLK), .Q(CRC_OUT_4_3) ) ;
DFF     gate196  (.D(WX7737), .CP(CLK), .Q(CRC_OUT_4_4) ) ;
DFF     gate197  (.D(WX7739), .CP(CLK), .Q(CRC_OUT_4_5) ) ;
DFF     gate198  (.D(WX7741), .CP(CLK), .Q(CRC_OUT_4_6) ) ;
DFF     gate199  (.D(WX7743), .CP(CLK), .Q(CRC_OUT_4_7) ) ;
DFF     gate200  (.D(WX7745), .CP(CLK), .Q(CRC_OUT_4_8) ) ;
DFF     gate201  (.D(WX7747), .CP(CLK), .Q(CRC_OUT_4_9) ) ;
DFF     gate202  (.D(WX7749), .CP(CLK), .Q(CRC_OUT_4_10) ) ;
DFF     gate203  (.D(WX7751), .CP(CLK), .Q(CRC_OUT_4_11) ) ;
DFF     gate204  (.D(WX7753), .CP(CLK), .Q(CRC_OUT_4_12) ) ;
DFF     gate205  (.D(WX7755), .CP(CLK), .Q(CRC_OUT_4_13) ) ;
DFF     gate206  (.D(WX7757), .CP(CLK), .Q(CRC_OUT_4_14) ) ;
DFF     gate207  (.D(WX7759), .CP(CLK), .Q(CRC_OUT_4_15) ) ;
DFF     gate208  (.D(WX7761), .CP(CLK), .Q(CRC_OUT_4_16) ) ;
DFF     gate209  (.D(WX7763), .CP(CLK), .Q(CRC_OUT_4_17) ) ;
DFF     gate210  (.D(WX7765), .CP(CLK), .Q(CRC_OUT_4_18) ) ;
DFF     gate211  (.D(WX7767), .CP(CLK), .Q(CRC_OUT_4_19) ) ;
DFF     gate212  (.D(WX7769), .CP(CLK), .Q(CRC_OUT_4_20) ) ;
DFF     gate213  (.D(WX7771), .CP(CLK), .Q(CRC_OUT_4_21) ) ;
DFF     gate214  (.D(WX7773), .CP(CLK), .Q(CRC_OUT_4_22) ) ;
DFF     gate215  (.D(WX7775), .CP(CLK), .Q(CRC_OUT_4_23) ) ;
DFF     gate216  (.D(WX7777), .CP(CLK), .Q(CRC_OUT_4_24) ) ;
DFF     gate217  (.D(WX7779), .CP(CLK), .Q(CRC_OUT_4_25) ) ;
DFF     gate218  (.D(WX7781), .CP(CLK), .Q(CRC_OUT_4_26) ) ;
DFF     gate219  (.D(WX7783), .CP(CLK), .Q(CRC_OUT_4_27) ) ;
DFF     gate220  (.D(WX7785), .CP(CLK), .Q(CRC_OUT_4_28) ) ;
DFF     gate221  (.D(WX7787), .CP(CLK), .Q(CRC_OUT_4_29) ) ;
DFF     gate222  (.D(WX7789), .CP(CLK), .Q(CRC_OUT_4_30) ) ;
DFF     gate223  (.D(WX7791), .CP(CLK), .Q(CRC_OUT_4_31) ) ;
DFF     gate224  (.D(WX9022), .CP(CLK), .Q(CRC_OUT_3_0) ) ;
DFF     gate225  (.D(WX9024), .CP(CLK), .Q(CRC_OUT_3_1) ) ;
DFF     gate226  (.D(WX9026), .CP(CLK), .Q(CRC_OUT_3_2) ) ;
DFF     gate227  (.D(WX9028), .CP(CLK), .Q(CRC_OUT_3_3) ) ;
DFF     gate228  (.D(WX9030), .CP(CLK), .Q(CRC_OUT_3_4) ) ;
DFF     gate229  (.D(WX9032), .CP(CLK), .Q(CRC_OUT_3_5) ) ;
DFF     gate230  (.D(WX9034), .CP(CLK), .Q(CRC_OUT_3_6) ) ;
DFF     gate231  (.D(WX9036), .CP(CLK), .Q(CRC_OUT_3_7) ) ;
DFF     gate232  (.D(WX9038), .CP(CLK), .Q(CRC_OUT_3_8) ) ;
DFF     gate233  (.D(WX9040), .CP(CLK), .Q(CRC_OUT_3_9) ) ;
DFF     gate234  (.D(WX9042), .CP(CLK), .Q(CRC_OUT_3_10) ) ;
DFF     gate235  (.D(WX9044), .CP(CLK), .Q(CRC_OUT_3_11) ) ;
DFF     gate236  (.D(WX9046), .CP(CLK), .Q(CRC_OUT_3_12) ) ;
DFF     gate237  (.D(WX9048), .CP(CLK), .Q(CRC_OUT_3_13) ) ;
DFF     gate238  (.D(WX9050), .CP(CLK), .Q(CRC_OUT_3_14) ) ;
DFF     gate239  (.D(WX9052), .CP(CLK), .Q(CRC_OUT_3_15) ) ;
DFF     gate240  (.D(WX9054), .CP(CLK), .Q(CRC_OUT_3_16) ) ;
DFF     gate241  (.D(WX9056), .CP(CLK), .Q(CRC_OUT_3_17) ) ;
DFF     gate242  (.D(WX9058), .CP(CLK), .Q(CRC_OUT_3_18) ) ;
DFF     gate243  (.D(WX9060), .CP(CLK), .Q(CRC_OUT_3_19) ) ;
DFF     gate244  (.D(WX9062), .CP(CLK), .Q(CRC_OUT_3_20) ) ;
DFF     gate245  (.D(WX9064), .CP(CLK), .Q(CRC_OUT_3_21) ) ;
DFF     gate246  (.D(WX9066), .CP(CLK), .Q(CRC_OUT_3_22) ) ;
DFF     gate247  (.D(WX9068), .CP(CLK), .Q(CRC_OUT_3_23) ) ;
DFF     gate248  (.D(WX9070), .CP(CLK), .Q(CRC_OUT_3_24) ) ;
DFF     gate249  (.D(WX9072), .CP(CLK), .Q(CRC_OUT_3_25) ) ;
DFF     gate250  (.D(WX9074), .CP(CLK), .Q(CRC_OUT_3_26) ) ;
DFF     gate251  (.D(WX9076), .CP(CLK), .Q(CRC_OUT_3_27) ) ;
DFF     gate252  (.D(WX9078), .CP(CLK), .Q(CRC_OUT_3_28) ) ;
DFF     gate253  (.D(WX9080), .CP(CLK), .Q(CRC_OUT_3_29) ) ;
DFF     gate254  (.D(WX9082), .CP(CLK), .Q(CRC_OUT_3_30) ) ;
DFF     gate255  (.D(WX9084), .CP(CLK), .Q(CRC_OUT_3_31) ) ;
DFF     gate256  (.D(WX10315), .CP(CLK), .Q(CRC_OUT_2_0) ) ;
DFF     gate257  (.D(WX10317), .CP(CLK), .Q(CRC_OUT_2_1) ) ;
DFF     gate258  (.D(WX10319), .CP(CLK), .Q(CRC_OUT_2_2) ) ;
DFF     gate259  (.D(WX10321), .CP(CLK), .Q(CRC_OUT_2_3) ) ;
DFF     gate260  (.D(WX10323), .CP(CLK), .Q(CRC_OUT_2_4) ) ;
DFF     gate261  (.D(WX10325), .CP(CLK), .Q(CRC_OUT_2_5) ) ;
DFF     gate262  (.D(WX10327), .CP(CLK), .Q(CRC_OUT_2_6) ) ;
DFF     gate263  (.D(WX10329), .CP(CLK), .Q(CRC_OUT_2_7) ) ;
DFF     gate264  (.D(WX10331), .CP(CLK), .Q(CRC_OUT_2_8) ) ;
DFF     gate265  (.D(WX10333), .CP(CLK), .Q(CRC_OUT_2_9) ) ;
DFF     gate266  (.D(WX10335), .CP(CLK), .Q(CRC_OUT_2_10) ) ;
DFF     gate267  (.D(WX10337), .CP(CLK), .Q(CRC_OUT_2_11) ) ;
DFF     gate268  (.D(WX10339), .CP(CLK), .Q(CRC_OUT_2_12) ) ;
DFF     gate269  (.D(WX10341), .CP(CLK), .Q(CRC_OUT_2_13) ) ;
DFF     gate270  (.D(WX10343), .CP(CLK), .Q(CRC_OUT_2_14) ) ;
DFF     gate271  (.D(WX10345), .CP(CLK), .Q(CRC_OUT_2_15) ) ;
DFF     gate272  (.D(WX10347), .CP(CLK), .Q(CRC_OUT_2_16) ) ;
DFF     gate273  (.D(WX10349), .CP(CLK), .Q(CRC_OUT_2_17) ) ;
DFF     gate274  (.D(WX10351), .CP(CLK), .Q(CRC_OUT_2_18) ) ;
DFF     gate275  (.D(WX10353), .CP(CLK), .Q(CRC_OUT_2_19) ) ;
DFF     gate276  (.D(WX10355), .CP(CLK), .Q(CRC_OUT_2_20) ) ;
DFF     gate277  (.D(WX10357), .CP(CLK), .Q(CRC_OUT_2_21) ) ;
DFF     gate278  (.D(WX10359), .CP(CLK), .Q(CRC_OUT_2_22) ) ;
DFF     gate279  (.D(WX10361), .CP(CLK), .Q(CRC_OUT_2_23) ) ;
DFF     gate280  (.D(WX10363), .CP(CLK), .Q(CRC_OUT_2_24) ) ;
DFF     gate281  (.D(WX10365), .CP(CLK), .Q(CRC_OUT_2_25) ) ;
DFF     gate282  (.D(WX10367), .CP(CLK), .Q(CRC_OUT_2_26) ) ;
DFF     gate283  (.D(WX10369), .CP(CLK), .Q(CRC_OUT_2_27) ) ;
DFF     gate284  (.D(WX10371), .CP(CLK), .Q(CRC_OUT_2_28) ) ;
DFF     gate285  (.D(WX10373), .CP(CLK), .Q(CRC_OUT_2_29) ) ;
DFF     gate286  (.D(WX10375), .CP(CLK), .Q(CRC_OUT_2_30) ) ;
DFF     gate287  (.D(WX10377), .CP(CLK), .Q(CRC_OUT_2_31) ) ;
DFF     gate288  (.D(WX11608), .CP(CLK), .Q(CRC_OUT_1_0) ) ;
DFF     gate289  (.D(WX11610), .CP(CLK), .Q(CRC_OUT_1_1) ) ;
DFF     gate290  (.D(WX11612), .CP(CLK), .Q(CRC_OUT_1_2) ) ;
DFF     gate291  (.D(WX11614), .CP(CLK), .Q(CRC_OUT_1_3) ) ;
DFF     gate292  (.D(WX11616), .CP(CLK), .Q(CRC_OUT_1_4) ) ;
DFF     gate293  (.D(WX11618), .CP(CLK), .Q(CRC_OUT_1_5) ) ;
DFF     gate294  (.D(WX11620), .CP(CLK), .Q(CRC_OUT_1_6) ) ;
DFF     gate295  (.D(WX11622), .CP(CLK), .Q(CRC_OUT_1_7) ) ;
DFF     gate296  (.D(WX11624), .CP(CLK), .Q(CRC_OUT_1_8) ) ;
DFF     gate297  (.D(WX11626), .CP(CLK), .Q(CRC_OUT_1_9) ) ;
DFF     gate298  (.D(WX11628), .CP(CLK), .Q(CRC_OUT_1_10) ) ;
DFF     gate299  (.D(WX11630), .CP(CLK), .Q(CRC_OUT_1_11) ) ;
DFF     gate300  (.D(WX11632), .CP(CLK), .Q(CRC_OUT_1_12) ) ;
DFF     gate301  (.D(WX11634), .CP(CLK), .Q(CRC_OUT_1_13) ) ;
DFF     gate302  (.D(WX11636), .CP(CLK), .Q(CRC_OUT_1_14) ) ;
DFF     gate303  (.D(WX11638), .CP(CLK), .Q(CRC_OUT_1_15) ) ;
DFF     gate304  (.D(WX11640), .CP(CLK), .Q(CRC_OUT_1_16) ) ;
DFF     gate305  (.D(WX11642), .CP(CLK), .Q(CRC_OUT_1_17) ) ;
DFF     gate306  (.D(WX11644), .CP(CLK), .Q(CRC_OUT_1_18) ) ;
DFF     gate307  (.D(WX11646), .CP(CLK), .Q(CRC_OUT_1_19) ) ;
DFF     gate308  (.D(WX11648), .CP(CLK), .Q(CRC_OUT_1_20) ) ;
DFF     gate309  (.D(WX11650), .CP(CLK), .Q(CRC_OUT_1_21) ) ;
DFF     gate310  (.D(WX11652), .CP(CLK), .Q(CRC_OUT_1_22) ) ;
DFF     gate311  (.D(WX11654), .CP(CLK), .Q(CRC_OUT_1_23) ) ;
DFF     gate312  (.D(WX11656), .CP(CLK), .Q(CRC_OUT_1_24) ) ;
DFF     gate313  (.D(WX11658), .CP(CLK), .Q(CRC_OUT_1_25) ) ;
DFF     gate314  (.D(WX11660), .CP(CLK), .Q(CRC_OUT_1_26) ) ;
DFF     gate315  (.D(WX11662), .CP(CLK), .Q(CRC_OUT_1_27) ) ;
DFF     gate316  (.D(WX11664), .CP(CLK), .Q(CRC_OUT_1_28) ) ;
DFF     gate317  (.D(WX11666), .CP(CLK), .Q(CRC_OUT_1_29) ) ;
DFF     gate318  (.D(WX11668), .CP(CLK), .Q(CRC_OUT_1_30) ) ;
DFF     gate319  (.D(WX11670), .CP(CLK), .Q(CRC_OUT_1_31) ) ;
AND2    gate320  (.A(WX487), .B(RESET), .Z(WX484) ) ;
DFF     gate321  (.D(WX484), .CP(CLK), .Q(WX485) ) ;
AND2    gate322  (.A(WX489), .B(RESET), .Z(WX486) ) ;
DFF     gate323  (.D(WX486), .CP(CLK), .Q(WX487) ) ;
AND2    gate324  (.A(WX491), .B(RESET), .Z(WX488) ) ;
DFF     gate325  (.D(WX488), .CP(CLK), .Q(WX489) ) ;
AND2    gate326  (.A(WX493), .B(RESET), .Z(WX490) ) ;
DFF     gate327  (.D(WX490), .CP(CLK), .Q(WX491) ) ;
AND2    gate328  (.A(WX495), .B(RESET), .Z(WX492) ) ;
DFF     gate329  (.D(WX492), .CP(CLK), .Q(WX493) ) ;
AND2    gate330  (.A(WX497), .B(RESET), .Z(WX494) ) ;
DFF     gate331  (.D(WX494), .CP(CLK), .Q(WX495) ) ;
AND2    gate332  (.A(WX499), .B(RESET), .Z(WX496) ) ;
DFF     gate333  (.D(WX496), .CP(CLK), .Q(WX497) ) ;
AND2    gate334  (.A(WX501), .B(RESET), .Z(WX498) ) ;
DFF     gate335  (.D(WX498), .CP(CLK), .Q(WX499) ) ;
AND2    gate336  (.A(WX503), .B(RESET), .Z(WX500) ) ;
DFF     gate337  (.D(WX500), .CP(CLK), .Q(WX501) ) ;
AND2    gate338  (.A(WX505), .B(RESET), .Z(WX502) ) ;
DFF     gate339  (.D(WX502), .CP(CLK), .Q(WX503) ) ;
AND2    gate340  (.A(WX507), .B(RESET), .Z(WX504) ) ;
DFF     gate341  (.D(WX504), .CP(CLK), .Q(WX505) ) ;
AND2    gate342  (.A(WX509), .B(RESET), .Z(WX506) ) ;
DFF     gate343  (.D(WX506), .CP(CLK), .Q(WX507) ) ;
AND2    gate344  (.A(WX511), .B(RESET), .Z(WX508) ) ;
DFF     gate345  (.D(WX508), .CP(CLK), .Q(WX509) ) ;
AND2    gate346  (.A(WX513), .B(RESET), .Z(WX510) ) ;
DFF     gate347  (.D(WX510), .CP(CLK), .Q(WX511) ) ;
AND2    gate348  (.A(WX515), .B(RESET), .Z(WX512) ) ;
DFF     gate349  (.D(WX512), .CP(CLK), .Q(WX513) ) ;
AND2    gate350  (.A(WX517), .B(RESET), .Z(WX514) ) ;
DFF     gate351  (.D(WX514), .CP(CLK), .Q(WX515) ) ;
AND2    gate352  (.A(WX519), .B(RESET), .Z(WX516) ) ;
DFF     gate353  (.D(WX516), .CP(CLK), .Q(WX517) ) ;
AND2    gate354  (.A(WX521), .B(RESET), .Z(WX518) ) ;
DFF     gate355  (.D(WX518), .CP(CLK), .Q(WX519) ) ;
AND2    gate356  (.A(WX523), .B(RESET), .Z(WX520) ) ;
DFF     gate357  (.D(WX520), .CP(CLK), .Q(WX521) ) ;
AND2    gate358  (.A(WX525), .B(RESET), .Z(WX522) ) ;
DFF     gate359  (.D(WX522), .CP(CLK), .Q(WX523) ) ;
AND2    gate360  (.A(WX527), .B(RESET), .Z(WX524) ) ;
DFF     gate361  (.D(WX524), .CP(CLK), .Q(WX525) ) ;
AND2    gate362  (.A(WX529), .B(RESET), .Z(WX526) ) ;
DFF     gate363  (.D(WX526), .CP(CLK), .Q(WX527) ) ;
AND2    gate364  (.A(WX531), .B(RESET), .Z(WX528) ) ;
DFF     gate365  (.D(WX528), .CP(CLK), .Q(WX529) ) ;
AND2    gate366  (.A(WX533), .B(RESET), .Z(WX530) ) ;
DFF     gate367  (.D(WX530), .CP(CLK), .Q(WX531) ) ;
AND2    gate368  (.A(WX535), .B(RESET), .Z(WX532) ) ;
DFF     gate369  (.D(WX532), .CP(CLK), .Q(WX533) ) ;
AND2    gate370  (.A(WX537), .B(RESET), .Z(WX534) ) ;
DFF     gate371  (.D(WX534), .CP(CLK), .Q(WX535) ) ;
AND2    gate372  (.A(WX539), .B(RESET), .Z(WX536) ) ;
DFF     gate373  (.D(WX536), .CP(CLK), .Q(WX537) ) ;
AND2    gate374  (.A(WX541), .B(RESET), .Z(WX538) ) ;
DFF     gate375  (.D(WX538), .CP(CLK), .Q(WX539) ) ;
AND2    gate376  (.A(WX543), .B(RESET), .Z(WX540) ) ;
DFF     gate377  (.D(WX540), .CP(CLK), .Q(WX541) ) ;
AND2    gate378  (.A(WX545), .B(RESET), .Z(WX542) ) ;
DFF     gate379  (.D(WX542), .CP(CLK), .Q(WX543) ) ;
AND2    gate380  (.A(WX547), .B(RESET), .Z(WX544) ) ;
DFF     gate381  (.D(WX544), .CP(CLK), .Q(WX545) ) ;
AND2    gate382  (.A(WX483), .B(RESET), .Z(WX546) ) ;
DFF     gate383  (.D(WX546), .CP(CLK), .Q(WX547) ) ;
AND2    gate384  (.A(WX48), .B(RESET), .Z(WX644) ) ;
DFF     gate385  (.D(WX644), .CP(CLK), .Q(WX645) ) ;
AND2    gate386  (.A(WX62), .B(RESET), .Z(WX646) ) ;
DFF     gate387  (.D(WX646), .CP(CLK), .Q(WX647) ) ;
AND2    gate388  (.A(WX76), .B(RESET), .Z(WX648) ) ;
DFF     gate389  (.D(WX648), .CP(CLK), .Q(WX649) ) ;
AND2    gate390  (.A(WX90), .B(RESET), .Z(WX650) ) ;
DFF     gate391  (.D(WX650), .CP(CLK), .Q(WX651) ) ;
AND2    gate392  (.A(WX104), .B(RESET), .Z(WX652) ) ;
DFF     gate393  (.D(WX652), .CP(CLK), .Q(WX653) ) ;
AND2    gate394  (.A(WX118), .B(RESET), .Z(WX654) ) ;
DFF     gate395  (.D(WX654), .CP(CLK), .Q(WX655) ) ;
AND2    gate396  (.A(WX132), .B(RESET), .Z(WX656) ) ;
DFF     gate397  (.D(WX656), .CP(CLK), .Q(WX657) ) ;
AND2    gate398  (.A(WX146), .B(RESET), .Z(WX658) ) ;
DFF     gate399  (.D(WX658), .CP(CLK), .Q(WX659) ) ;
AND2    gate400  (.A(WX160), .B(RESET), .Z(WX660) ) ;
DFF     gate401  (.D(WX660), .CP(CLK), .Q(WX661) ) ;
AND2    gate402  (.A(WX174), .B(RESET), .Z(WX662) ) ;
DFF     gate403  (.D(WX662), .CP(CLK), .Q(WX663) ) ;
AND2    gate404  (.A(WX188), .B(RESET), .Z(WX664) ) ;
DFF     gate405  (.D(WX664), .CP(CLK), .Q(WX665) ) ;
AND2    gate406  (.A(WX202), .B(RESET), .Z(WX666) ) ;
DFF     gate407  (.D(WX666), .CP(CLK), .Q(WX667) ) ;
AND2    gate408  (.A(WX216), .B(RESET), .Z(WX668) ) ;
DFF     gate409  (.D(WX668), .CP(CLK), .Q(WX669) ) ;
AND2    gate410  (.A(WX230), .B(RESET), .Z(WX670) ) ;
DFF     gate411  (.D(WX670), .CP(CLK), .Q(WX671) ) ;
AND2    gate412  (.A(WX244), .B(RESET), .Z(WX672) ) ;
DFF     gate413  (.D(WX672), .CP(CLK), .Q(WX673) ) ;
AND2    gate414  (.A(WX258), .B(RESET), .Z(WX674) ) ;
DFF     gate415  (.D(WX674), .CP(CLK), .Q(WX675) ) ;
AND2    gate416  (.A(WX272), .B(RESET), .Z(WX676) ) ;
DFF     gate417  (.D(WX676), .CP(CLK), .Q(WX677) ) ;
AND2    gate418  (.A(WX286), .B(RESET), .Z(WX678) ) ;
DFF     gate419  (.D(WX678), .CP(CLK), .Q(WX679) ) ;
AND2    gate420  (.A(WX300), .B(RESET), .Z(WX680) ) ;
DFF     gate421  (.D(WX680), .CP(CLK), .Q(WX681) ) ;
AND2    gate422  (.A(WX314), .B(RESET), .Z(WX682) ) ;
DFF     gate423  (.D(WX682), .CP(CLK), .Q(WX683) ) ;
AND2    gate424  (.A(WX328), .B(RESET), .Z(WX684) ) ;
DFF     gate425  (.D(WX684), .CP(CLK), .Q(WX685) ) ;
AND2    gate426  (.A(WX342), .B(RESET), .Z(WX686) ) ;
DFF     gate427  (.D(WX686), .CP(CLK), .Q(WX687) ) ;
AND2    gate428  (.A(WX356), .B(RESET), .Z(WX688) ) ;
DFF     gate429  (.D(WX688), .CP(CLK), .Q(WX689) ) ;
AND2    gate430  (.A(WX370), .B(RESET), .Z(WX690) ) ;
DFF     gate431  (.D(WX690), .CP(CLK), .Q(WX691) ) ;
AND2    gate432  (.A(WX384), .B(RESET), .Z(WX692) ) ;
DFF     gate433  (.D(WX692), .CP(CLK), .Q(WX693) ) ;
AND2    gate434  (.A(WX398), .B(RESET), .Z(WX694) ) ;
DFF     gate435  (.D(WX694), .CP(CLK), .Q(WX695) ) ;
AND2    gate436  (.A(WX412), .B(RESET), .Z(WX696) ) ;
DFF     gate437  (.D(WX696), .CP(CLK), .Q(WX697) ) ;
AND2    gate438  (.A(WX426), .B(RESET), .Z(WX698) ) ;
DFF     gate439  (.D(WX698), .CP(CLK), .Q(WX699) ) ;
AND2    gate440  (.A(WX440), .B(RESET), .Z(WX700) ) ;
DFF     gate441  (.D(WX700), .CP(CLK), .Q(WX701) ) ;
AND2    gate442  (.A(WX454), .B(RESET), .Z(WX702) ) ;
DFF     gate443  (.D(WX702), .CP(CLK), .Q(WX703) ) ;
AND2    gate444  (.A(WX468), .B(RESET), .Z(WX704) ) ;
DFF     gate445  (.D(WX704), .CP(CLK), .Q(WX705) ) ;
AND2    gate446  (.A(WX482), .B(RESET), .Z(WX706) ) ;
DFF     gate447  (.D(WX706), .CP(CLK), .Q(WX707) ) ;
AND2    gate448  (.A(WX645), .B(RESET), .Z(WX708) ) ;
DFF     gate449  (.D(WX708), .CP(CLK), .Q(WX709) ) ;
AND2    gate450  (.A(WX647), .B(RESET), .Z(WX710) ) ;
DFF     gate451  (.D(WX710), .CP(CLK), .Q(WX711) ) ;
AND2    gate452  (.A(WX649), .B(RESET), .Z(WX712) ) ;
DFF     gate453  (.D(WX712), .CP(CLK), .Q(WX713) ) ;
AND2    gate454  (.A(WX651), .B(RESET), .Z(WX714) ) ;
DFF     gate455  (.D(WX714), .CP(CLK), .Q(WX715) ) ;
AND2    gate456  (.A(WX653), .B(RESET), .Z(WX716) ) ;
DFF     gate457  (.D(WX716), .CP(CLK), .Q(WX717) ) ;
AND2    gate458  (.A(WX655), .B(RESET), .Z(WX718) ) ;
DFF     gate459  (.D(WX718), .CP(CLK), .Q(WX719) ) ;
AND2    gate460  (.A(WX657), .B(RESET), .Z(WX720) ) ;
DFF     gate461  (.D(WX720), .CP(CLK), .Q(WX721) ) ;
AND2    gate462  (.A(WX659), .B(RESET), .Z(WX722) ) ;
DFF     gate463  (.D(WX722), .CP(CLK), .Q(WX723) ) ;
AND2    gate464  (.A(WX661), .B(RESET), .Z(WX724) ) ;
DFF     gate465  (.D(WX724), .CP(CLK), .Q(WX725) ) ;
AND2    gate466  (.A(WX663), .B(RESET), .Z(WX726) ) ;
DFF     gate467  (.D(WX726), .CP(CLK), .Q(WX727) ) ;
AND2    gate468  (.A(WX665), .B(RESET), .Z(WX728) ) ;
DFF     gate469  (.D(WX728), .CP(CLK), .Q(WX729) ) ;
AND2    gate470  (.A(WX667), .B(RESET), .Z(WX730) ) ;
DFF     gate471  (.D(WX730), .CP(CLK), .Q(WX731) ) ;
AND2    gate472  (.A(WX669), .B(RESET), .Z(WX732) ) ;
DFF     gate473  (.D(WX732), .CP(CLK), .Q(WX733) ) ;
AND2    gate474  (.A(WX671), .B(RESET), .Z(WX734) ) ;
DFF     gate475  (.D(WX734), .CP(CLK), .Q(WX735) ) ;
AND2    gate476  (.A(WX673), .B(RESET), .Z(WX736) ) ;
DFF     gate477  (.D(WX736), .CP(CLK), .Q(WX737) ) ;
AND2    gate478  (.A(WX675), .B(RESET), .Z(WX738) ) ;
DFF     gate479  (.D(WX738), .CP(CLK), .Q(WX739) ) ;
AND2    gate480  (.A(WX677), .B(RESET), .Z(WX740) ) ;
DFF     gate481  (.D(WX740), .CP(CLK), .Q(WX741) ) ;
AND2    gate482  (.A(WX679), .B(RESET), .Z(WX742) ) ;
DFF     gate483  (.D(WX742), .CP(CLK), .Q(WX743) ) ;
AND2    gate484  (.A(WX681), .B(RESET), .Z(WX744) ) ;
DFF     gate485  (.D(WX744), .CP(CLK), .Q(WX745) ) ;
AND2    gate486  (.A(WX683), .B(RESET), .Z(WX746) ) ;
DFF     gate487  (.D(WX746), .CP(CLK), .Q(WX747) ) ;
AND2    gate488  (.A(WX685), .B(RESET), .Z(WX748) ) ;
DFF     gate489  (.D(WX748), .CP(CLK), .Q(WX749) ) ;
AND2    gate490  (.A(WX687), .B(RESET), .Z(WX750) ) ;
DFF     gate491  (.D(WX750), .CP(CLK), .Q(WX751) ) ;
AND2    gate492  (.A(WX689), .B(RESET), .Z(WX752) ) ;
DFF     gate493  (.D(WX752), .CP(CLK), .Q(WX753) ) ;
AND2    gate494  (.A(WX691), .B(RESET), .Z(WX754) ) ;
DFF     gate495  (.D(WX754), .CP(CLK), .Q(WX755) ) ;
AND2    gate496  (.A(WX693), .B(RESET), .Z(WX756) ) ;
DFF     gate497  (.D(WX756), .CP(CLK), .Q(WX757) ) ;
AND2    gate498  (.A(WX695), .B(RESET), .Z(WX758) ) ;
DFF     gate499  (.D(WX758), .CP(CLK), .Q(WX759) ) ;
AND2    gate500  (.A(WX697), .B(RESET), .Z(WX760) ) ;
DFF     gate501  (.D(WX760), .CP(CLK), .Q(WX761) ) ;
AND2    gate502  (.A(WX699), .B(RESET), .Z(WX762) ) ;
DFF     gate503  (.D(WX762), .CP(CLK), .Q(WX763) ) ;
AND2    gate504  (.A(WX701), .B(RESET), .Z(WX764) ) ;
DFF     gate505  (.D(WX764), .CP(CLK), .Q(WX765) ) ;
AND2    gate506  (.A(WX703), .B(RESET), .Z(WX766) ) ;
DFF     gate507  (.D(WX766), .CP(CLK), .Q(WX767) ) ;
AND2    gate508  (.A(WX705), .B(RESET), .Z(WX768) ) ;
DFF     gate509  (.D(WX768), .CP(CLK), .Q(WX769) ) ;
AND2    gate510  (.A(WX707), .B(RESET), .Z(WX770) ) ;
DFF     gate511  (.D(WX770), .CP(CLK), .Q(WX771) ) ;
AND2    gate512  (.A(WX709), .B(RESET), .Z(WX772) ) ;
DFF     gate513  (.D(WX772), .CP(CLK), .Q(WX773) ) ;
AND2    gate514  (.A(WX711), .B(RESET), .Z(WX774) ) ;
DFF     gate515  (.D(WX774), .CP(CLK), .Q(WX775) ) ;
AND2    gate516  (.A(WX713), .B(RESET), .Z(WX776) ) ;
DFF     gate517  (.D(WX776), .CP(CLK), .Q(WX777) ) ;
AND2    gate518  (.A(WX715), .B(RESET), .Z(WX778) ) ;
DFF     gate519  (.D(WX778), .CP(CLK), .Q(WX779) ) ;
AND2    gate520  (.A(WX717), .B(RESET), .Z(WX780) ) ;
DFF     gate521  (.D(WX780), .CP(CLK), .Q(WX781) ) ;
AND2    gate522  (.A(WX719), .B(RESET), .Z(WX782) ) ;
DFF     gate523  (.D(WX782), .CP(CLK), .Q(WX783) ) ;
AND2    gate524  (.A(WX721), .B(RESET), .Z(WX784) ) ;
DFF     gate525  (.D(WX784), .CP(CLK), .Q(WX785) ) ;
AND2    gate526  (.A(WX723), .B(RESET), .Z(WX786) ) ;
DFF     gate527  (.D(WX786), .CP(CLK), .Q(WX787) ) ;
AND2    gate528  (.A(WX725), .B(RESET), .Z(WX788) ) ;
DFF     gate529  (.D(WX788), .CP(CLK), .Q(WX789) ) ;
AND2    gate530  (.A(WX727), .B(RESET), .Z(WX790) ) ;
DFF     gate531  (.D(WX790), .CP(CLK), .Q(WX791) ) ;
AND2    gate532  (.A(WX729), .B(RESET), .Z(WX792) ) ;
DFF     gate533  (.D(WX792), .CP(CLK), .Q(WX793) ) ;
AND2    gate534  (.A(WX731), .B(RESET), .Z(WX794) ) ;
DFF     gate535  (.D(WX794), .CP(CLK), .Q(WX795) ) ;
AND2    gate536  (.A(WX733), .B(RESET), .Z(WX796) ) ;
DFF     gate537  (.D(WX796), .CP(CLK), .Q(WX797) ) ;
AND2    gate538  (.A(WX735), .B(RESET), .Z(WX798) ) ;
DFF     gate539  (.D(WX798), .CP(CLK), .Q(WX799) ) ;
AND2    gate540  (.A(WX737), .B(RESET), .Z(WX800) ) ;
DFF     gate541  (.D(WX800), .CP(CLK), .Q(WX801) ) ;
AND2    gate542  (.A(WX739), .B(RESET), .Z(WX802) ) ;
DFF     gate543  (.D(WX802), .CP(CLK), .Q(WX803) ) ;
AND2    gate544  (.A(WX741), .B(RESET), .Z(WX804) ) ;
DFF     gate545  (.D(WX804), .CP(CLK), .Q(WX805) ) ;
AND2    gate546  (.A(WX743), .B(RESET), .Z(WX806) ) ;
DFF     gate547  (.D(WX806), .CP(CLK), .Q(WX807) ) ;
AND2    gate548  (.A(WX745), .B(RESET), .Z(WX808) ) ;
DFF     gate549  (.D(WX808), .CP(CLK), .Q(WX809) ) ;
AND2    gate550  (.A(WX747), .B(RESET), .Z(WX810) ) ;
DFF     gate551  (.D(WX810), .CP(CLK), .Q(WX811) ) ;
AND2    gate552  (.A(WX749), .B(RESET), .Z(WX812) ) ;
DFF     gate553  (.D(WX812), .CP(CLK), .Q(WX813) ) ;
AND2    gate554  (.A(WX751), .B(RESET), .Z(WX814) ) ;
DFF     gate555  (.D(WX814), .CP(CLK), .Q(WX815) ) ;
AND2    gate556  (.A(WX753), .B(RESET), .Z(WX816) ) ;
DFF     gate557  (.D(WX816), .CP(CLK), .Q(WX817) ) ;
AND2    gate558  (.A(WX755), .B(RESET), .Z(WX818) ) ;
DFF     gate559  (.D(WX818), .CP(CLK), .Q(WX819) ) ;
AND2    gate560  (.A(WX757), .B(RESET), .Z(WX820) ) ;
DFF     gate561  (.D(WX820), .CP(CLK), .Q(WX821) ) ;
AND2    gate562  (.A(WX759), .B(RESET), .Z(WX822) ) ;
DFF     gate563  (.D(WX822), .CP(CLK), .Q(WX823) ) ;
AND2    gate564  (.A(WX761), .B(RESET), .Z(WX824) ) ;
DFF     gate565  (.D(WX824), .CP(CLK), .Q(WX825) ) ;
AND2    gate566  (.A(WX763), .B(RESET), .Z(WX826) ) ;
DFF     gate567  (.D(WX826), .CP(CLK), .Q(WX827) ) ;
AND2    gate568  (.A(WX765), .B(RESET), .Z(WX828) ) ;
DFF     gate569  (.D(WX828), .CP(CLK), .Q(WX829) ) ;
AND2    gate570  (.A(WX767), .B(RESET), .Z(WX830) ) ;
DFF     gate571  (.D(WX830), .CP(CLK), .Q(WX831) ) ;
AND2    gate572  (.A(WX769), .B(RESET), .Z(WX832) ) ;
DFF     gate573  (.D(WX832), .CP(CLK), .Q(WX833) ) ;
AND2    gate574  (.A(WX771), .B(RESET), .Z(WX834) ) ;
DFF     gate575  (.D(WX834), .CP(CLK), .Q(WX835) ) ;
AND2    gate576  (.A(WX773), .B(RESET), .Z(WX836) ) ;
DFF     gate577  (.D(WX836), .CP(CLK), .Q(WX837) ) ;
AND2    gate578  (.A(WX775), .B(RESET), .Z(WX838) ) ;
DFF     gate579  (.D(WX838), .CP(CLK), .Q(WX839) ) ;
AND2    gate580  (.A(WX777), .B(RESET), .Z(WX840) ) ;
DFF     gate581  (.D(WX840), .CP(CLK), .Q(WX841) ) ;
AND2    gate582  (.A(WX779), .B(RESET), .Z(WX842) ) ;
DFF     gate583  (.D(WX842), .CP(CLK), .Q(WX843) ) ;
AND2    gate584  (.A(WX781), .B(RESET), .Z(WX844) ) ;
DFF     gate585  (.D(WX844), .CP(CLK), .Q(WX845) ) ;
AND2    gate586  (.A(WX783), .B(RESET), .Z(WX846) ) ;
DFF     gate587  (.D(WX846), .CP(CLK), .Q(WX847) ) ;
AND2    gate588  (.A(WX785), .B(RESET), .Z(WX848) ) ;
DFF     gate589  (.D(WX848), .CP(CLK), .Q(WX849) ) ;
AND2    gate590  (.A(WX787), .B(RESET), .Z(WX850) ) ;
DFF     gate591  (.D(WX850), .CP(CLK), .Q(WX851) ) ;
AND2    gate592  (.A(WX789), .B(RESET), .Z(WX852) ) ;
DFF     gate593  (.D(WX852), .CP(CLK), .Q(WX853) ) ;
AND2    gate594  (.A(WX791), .B(RESET), .Z(WX854) ) ;
DFF     gate595  (.D(WX854), .CP(CLK), .Q(WX855) ) ;
AND2    gate596  (.A(WX793), .B(RESET), .Z(WX856) ) ;
DFF     gate597  (.D(WX856), .CP(CLK), .Q(WX857) ) ;
AND2    gate598  (.A(WX795), .B(RESET), .Z(WX858) ) ;
DFF     gate599  (.D(WX858), .CP(CLK), .Q(WX859) ) ;
AND2    gate600  (.A(WX797), .B(RESET), .Z(WX860) ) ;
DFF     gate601  (.D(WX860), .CP(CLK), .Q(WX861) ) ;
AND2    gate602  (.A(WX799), .B(RESET), .Z(WX862) ) ;
DFF     gate603  (.D(WX862), .CP(CLK), .Q(WX863) ) ;
AND2    gate604  (.A(WX801), .B(RESET), .Z(WX864) ) ;
DFF     gate605  (.D(WX864), .CP(CLK), .Q(WX865) ) ;
AND2    gate606  (.A(WX803), .B(RESET), .Z(WX866) ) ;
DFF     gate607  (.D(WX866), .CP(CLK), .Q(WX867) ) ;
AND2    gate608  (.A(WX805), .B(RESET), .Z(WX868) ) ;
DFF     gate609  (.D(WX868), .CP(CLK), .Q(WX869) ) ;
AND2    gate610  (.A(WX807), .B(RESET), .Z(WX870) ) ;
DFF     gate611  (.D(WX870), .CP(CLK), .Q(WX871) ) ;
AND2    gate612  (.A(WX809), .B(RESET), .Z(WX872) ) ;
DFF     gate613  (.D(WX872), .CP(CLK), .Q(WX873) ) ;
AND2    gate614  (.A(WX811), .B(RESET), .Z(WX874) ) ;
DFF     gate615  (.D(WX874), .CP(CLK), .Q(WX875) ) ;
AND2    gate616  (.A(WX813), .B(RESET), .Z(WX876) ) ;
DFF     gate617  (.D(WX876), .CP(CLK), .Q(WX877) ) ;
AND2    gate618  (.A(WX815), .B(RESET), .Z(WX878) ) ;
DFF     gate619  (.D(WX878), .CP(CLK), .Q(WX879) ) ;
AND2    gate620  (.A(WX817), .B(RESET), .Z(WX880) ) ;
DFF     gate621  (.D(WX880), .CP(CLK), .Q(WX881) ) ;
AND2    gate622  (.A(WX819), .B(RESET), .Z(WX882) ) ;
DFF     gate623  (.D(WX882), .CP(CLK), .Q(WX883) ) ;
AND2    gate624  (.A(WX821), .B(RESET), .Z(WX884) ) ;
DFF     gate625  (.D(WX884), .CP(CLK), .Q(WX885) ) ;
AND2    gate626  (.A(WX823), .B(RESET), .Z(WX886) ) ;
DFF     gate627  (.D(WX886), .CP(CLK), .Q(WX887) ) ;
AND2    gate628  (.A(WX825), .B(RESET), .Z(WX888) ) ;
DFF     gate629  (.D(WX888), .CP(CLK), .Q(WX889) ) ;
AND2    gate630  (.A(WX827), .B(RESET), .Z(WX890) ) ;
DFF     gate631  (.D(WX890), .CP(CLK), .Q(WX891) ) ;
AND2    gate632  (.A(WX829), .B(RESET), .Z(WX892) ) ;
DFF     gate633  (.D(WX892), .CP(CLK), .Q(WX893) ) ;
AND2    gate634  (.A(WX831), .B(RESET), .Z(WX894) ) ;
DFF     gate635  (.D(WX894), .CP(CLK), .Q(WX895) ) ;
AND2    gate636  (.A(WX833), .B(RESET), .Z(WX896) ) ;
DFF     gate637  (.D(WX896), .CP(CLK), .Q(WX897) ) ;
AND2    gate638  (.A(WX835), .B(RESET), .Z(WX898) ) ;
DFF     gate639  (.D(WX898), .CP(CLK), .Q(WX899) ) ;
AND2    gate640  (.A(WX1234), .B(WX1263), .Z(WX1264) ) ;
AND2    gate641  (.A(WX1262), .B(WX1263), .Z(WX1266) ) ;
AND2    gate642  (.A(WX1261), .B(WX1263), .Z(WX1268) ) ;
AND2    gate643  (.A(WX1260), .B(WX1263), .Z(WX1270) ) ;
AND2    gate644  (.A(WX1233), .B(WX1263), .Z(WX1272) ) ;
AND2    gate645  (.A(WX1259), .B(WX1263), .Z(WX1274) ) ;
AND2    gate646  (.A(WX1258), .B(WX1263), .Z(WX1276) ) ;
AND2    gate647  (.A(WX1257), .B(WX1263), .Z(WX1278) ) ;
AND2    gate648  (.A(WX1256), .B(WX1263), .Z(WX1280) ) ;
AND2    gate649  (.A(WX1255), .B(WX1263), .Z(WX1282) ) ;
AND2    gate650  (.A(WX1254), .B(WX1263), .Z(WX1284) ) ;
AND2    gate651  (.A(WX1232), .B(WX1263), .Z(WX1286) ) ;
AND2    gate652  (.A(WX1253), .B(WX1263), .Z(WX1288) ) ;
AND2    gate653  (.A(WX1252), .B(WX1263), .Z(WX1290) ) ;
AND2    gate654  (.A(WX1251), .B(WX1263), .Z(WX1292) ) ;
AND2    gate655  (.A(WX1250), .B(WX1263), .Z(WX1294) ) ;
AND2    gate656  (.A(WX1231), .B(WX1263), .Z(WX1296) ) ;
AND2    gate657  (.A(WX1249), .B(WX1263), .Z(WX1298) ) ;
AND2    gate658  (.A(WX1248), .B(WX1263), .Z(WX1300) ) ;
AND2    gate659  (.A(WX1247), .B(WX1263), .Z(WX1302) ) ;
AND2    gate660  (.A(WX1246), .B(WX1263), .Z(WX1304) ) ;
AND2    gate661  (.A(WX1245), .B(WX1263), .Z(WX1306) ) ;
AND2    gate662  (.A(WX1244), .B(WX1263), .Z(WX1308) ) ;
AND2    gate663  (.A(WX1243), .B(WX1263), .Z(WX1310) ) ;
AND2    gate664  (.A(WX1242), .B(WX1263), .Z(WX1312) ) ;
AND2    gate665  (.A(WX1241), .B(WX1263), .Z(WX1314) ) ;
AND2    gate666  (.A(WX1240), .B(WX1263), .Z(WX1316) ) ;
AND2    gate667  (.A(WX1239), .B(WX1263), .Z(WX1318) ) ;
AND2    gate668  (.A(WX1238), .B(WX1263), .Z(WX1320) ) ;
AND2    gate669  (.A(WX1237), .B(WX1263), .Z(WX1322) ) ;
AND2    gate670  (.A(WX1236), .B(WX1263), .Z(WX1324) ) ;
AND2    gate671  (.A(WX1235), .B(WX1263), .Z(WX1326) ) ;
AND2    gate672  (.A(WX1780), .B(RESET), .Z(WX1777) ) ;
DFF     gate673  (.D(WX1777), .CP(CLK), .Q(WX1778) ) ;
AND2    gate674  (.A(WX1782), .B(RESET), .Z(WX1779) ) ;
DFF     gate675  (.D(WX1779), .CP(CLK), .Q(WX1780) ) ;
AND2    gate676  (.A(WX1784), .B(RESET), .Z(WX1781) ) ;
DFF     gate677  (.D(WX1781), .CP(CLK), .Q(WX1782) ) ;
AND2    gate678  (.A(WX1786), .B(RESET), .Z(WX1783) ) ;
DFF     gate679  (.D(WX1783), .CP(CLK), .Q(WX1784) ) ;
AND2    gate680  (.A(WX1788), .B(RESET), .Z(WX1785) ) ;
DFF     gate681  (.D(WX1785), .CP(CLK), .Q(WX1786) ) ;
AND2    gate682  (.A(WX1790), .B(RESET), .Z(WX1787) ) ;
DFF     gate683  (.D(WX1787), .CP(CLK), .Q(WX1788) ) ;
AND2    gate684  (.A(WX1792), .B(RESET), .Z(WX1789) ) ;
DFF     gate685  (.D(WX1789), .CP(CLK), .Q(WX1790) ) ;
AND2    gate686  (.A(WX1794), .B(RESET), .Z(WX1791) ) ;
DFF     gate687  (.D(WX1791), .CP(CLK), .Q(WX1792) ) ;
AND2    gate688  (.A(WX1796), .B(RESET), .Z(WX1793) ) ;
DFF     gate689  (.D(WX1793), .CP(CLK), .Q(WX1794) ) ;
AND2    gate690  (.A(WX1798), .B(RESET), .Z(WX1795) ) ;
DFF     gate691  (.D(WX1795), .CP(CLK), .Q(WX1796) ) ;
AND2    gate692  (.A(WX1800), .B(RESET), .Z(WX1797) ) ;
DFF     gate693  (.D(WX1797), .CP(CLK), .Q(WX1798) ) ;
AND2    gate694  (.A(WX1802), .B(RESET), .Z(WX1799) ) ;
DFF     gate695  (.D(WX1799), .CP(CLK), .Q(WX1800) ) ;
AND2    gate696  (.A(WX1804), .B(RESET), .Z(WX1801) ) ;
DFF     gate697  (.D(WX1801), .CP(CLK), .Q(WX1802) ) ;
AND2    gate698  (.A(WX1806), .B(RESET), .Z(WX1803) ) ;
DFF     gate699  (.D(WX1803), .CP(CLK), .Q(WX1804) ) ;
AND2    gate700  (.A(WX1808), .B(RESET), .Z(WX1805) ) ;
DFF     gate701  (.D(WX1805), .CP(CLK), .Q(WX1806) ) ;
AND2    gate702  (.A(WX1810), .B(RESET), .Z(WX1807) ) ;
DFF     gate703  (.D(WX1807), .CP(CLK), .Q(WX1808) ) ;
AND2    gate704  (.A(WX1812), .B(RESET), .Z(WX1809) ) ;
DFF     gate705  (.D(WX1809), .CP(CLK), .Q(WX1810) ) ;
AND2    gate706  (.A(WX1814), .B(RESET), .Z(WX1811) ) ;
DFF     gate707  (.D(WX1811), .CP(CLK), .Q(WX1812) ) ;
AND2    gate708  (.A(WX1816), .B(RESET), .Z(WX1813) ) ;
DFF     gate709  (.D(WX1813), .CP(CLK), .Q(WX1814) ) ;
AND2    gate710  (.A(WX1818), .B(RESET), .Z(WX1815) ) ;
DFF     gate711  (.D(WX1815), .CP(CLK), .Q(WX1816) ) ;
AND2    gate712  (.A(WX1820), .B(RESET), .Z(WX1817) ) ;
DFF     gate713  (.D(WX1817), .CP(CLK), .Q(WX1818) ) ;
AND2    gate714  (.A(WX1822), .B(RESET), .Z(WX1819) ) ;
DFF     gate715  (.D(WX1819), .CP(CLK), .Q(WX1820) ) ;
AND2    gate716  (.A(WX1824), .B(RESET), .Z(WX1821) ) ;
DFF     gate717  (.D(WX1821), .CP(CLK), .Q(WX1822) ) ;
AND2    gate718  (.A(WX1826), .B(RESET), .Z(WX1823) ) ;
DFF     gate719  (.D(WX1823), .CP(CLK), .Q(WX1824) ) ;
AND2    gate720  (.A(WX1828), .B(RESET), .Z(WX1825) ) ;
DFF     gate721  (.D(WX1825), .CP(CLK), .Q(WX1826) ) ;
AND2    gate722  (.A(WX1830), .B(RESET), .Z(WX1827) ) ;
DFF     gate723  (.D(WX1827), .CP(CLK), .Q(WX1828) ) ;
AND2    gate724  (.A(WX1832), .B(RESET), .Z(WX1829) ) ;
DFF     gate725  (.D(WX1829), .CP(CLK), .Q(WX1830) ) ;
AND2    gate726  (.A(WX1834), .B(RESET), .Z(WX1831) ) ;
DFF     gate727  (.D(WX1831), .CP(CLK), .Q(WX1832) ) ;
AND2    gate728  (.A(WX1836), .B(RESET), .Z(WX1833) ) ;
DFF     gate729  (.D(WX1833), .CP(CLK), .Q(WX1834) ) ;
AND2    gate730  (.A(WX1838), .B(RESET), .Z(WX1835) ) ;
DFF     gate731  (.D(WX1835), .CP(CLK), .Q(WX1836) ) ;
AND2    gate732  (.A(WX1840), .B(RESET), .Z(WX1837) ) ;
DFF     gate733  (.D(WX1837), .CP(CLK), .Q(WX1838) ) ;
AND2    gate734  (.A(WX1776), .B(RESET), .Z(WX1839) ) ;
DFF     gate735  (.D(WX1839), .CP(CLK), .Q(WX1840) ) ;
AND2    gate736  (.A(WX1341), .B(RESET), .Z(WX1937) ) ;
DFF     gate737  (.D(WX1937), .CP(CLK), .Q(WX1938) ) ;
AND2    gate738  (.A(WX1355), .B(RESET), .Z(WX1939) ) ;
DFF     gate739  (.D(WX1939), .CP(CLK), .Q(WX1940) ) ;
AND2    gate740  (.A(WX1369), .B(RESET), .Z(WX1941) ) ;
DFF     gate741  (.D(WX1941), .CP(CLK), .Q(WX1942) ) ;
AND2    gate742  (.A(WX1383), .B(RESET), .Z(WX1943) ) ;
DFF     gate743  (.D(WX1943), .CP(CLK), .Q(WX1944) ) ;
AND2    gate744  (.A(WX1397), .B(RESET), .Z(WX1945) ) ;
DFF     gate745  (.D(WX1945), .CP(CLK), .Q(WX1946) ) ;
AND2    gate746  (.A(WX1411), .B(RESET), .Z(WX1947) ) ;
DFF     gate747  (.D(WX1947), .CP(CLK), .Q(WX1948) ) ;
AND2    gate748  (.A(WX1425), .B(RESET), .Z(WX1949) ) ;
DFF     gate749  (.D(WX1949), .CP(CLK), .Q(WX1950) ) ;
AND2    gate750  (.A(WX1439), .B(RESET), .Z(WX1951) ) ;
DFF     gate751  (.D(WX1951), .CP(CLK), .Q(WX1952) ) ;
AND2    gate752  (.A(WX1453), .B(RESET), .Z(WX1953) ) ;
DFF     gate753  (.D(WX1953), .CP(CLK), .Q(WX1954) ) ;
AND2    gate754  (.A(WX1467), .B(RESET), .Z(WX1955) ) ;
DFF     gate755  (.D(WX1955), .CP(CLK), .Q(WX1956) ) ;
AND2    gate756  (.A(WX1481), .B(RESET), .Z(WX1957) ) ;
DFF     gate757  (.D(WX1957), .CP(CLK), .Q(WX1958) ) ;
AND2    gate758  (.A(WX1495), .B(RESET), .Z(WX1959) ) ;
DFF     gate759  (.D(WX1959), .CP(CLK), .Q(WX1960) ) ;
AND2    gate760  (.A(WX1509), .B(RESET), .Z(WX1961) ) ;
DFF     gate761  (.D(WX1961), .CP(CLK), .Q(WX1962) ) ;
AND2    gate762  (.A(WX1523), .B(RESET), .Z(WX1963) ) ;
DFF     gate763  (.D(WX1963), .CP(CLK), .Q(WX1964) ) ;
AND2    gate764  (.A(WX1537), .B(RESET), .Z(WX1965) ) ;
DFF     gate765  (.D(WX1965), .CP(CLK), .Q(WX1966) ) ;
AND2    gate766  (.A(WX1551), .B(RESET), .Z(WX1967) ) ;
DFF     gate767  (.D(WX1967), .CP(CLK), .Q(WX1968) ) ;
AND2    gate768  (.A(WX1565), .B(RESET), .Z(WX1969) ) ;
DFF     gate769  (.D(WX1969), .CP(CLK), .Q(WX1970) ) ;
AND2    gate770  (.A(WX1579), .B(RESET), .Z(WX1971) ) ;
DFF     gate771  (.D(WX1971), .CP(CLK), .Q(WX1972) ) ;
AND2    gate772  (.A(WX1593), .B(RESET), .Z(WX1973) ) ;
DFF     gate773  (.D(WX1973), .CP(CLK), .Q(WX1974) ) ;
AND2    gate774  (.A(WX1607), .B(RESET), .Z(WX1975) ) ;
DFF     gate775  (.D(WX1975), .CP(CLK), .Q(WX1976) ) ;
AND2    gate776  (.A(WX1621), .B(RESET), .Z(WX1977) ) ;
DFF     gate777  (.D(WX1977), .CP(CLK), .Q(WX1978) ) ;
AND2    gate778  (.A(WX1635), .B(RESET), .Z(WX1979) ) ;
DFF     gate779  (.D(WX1979), .CP(CLK), .Q(WX1980) ) ;
AND2    gate780  (.A(WX1649), .B(RESET), .Z(WX1981) ) ;
DFF     gate781  (.D(WX1981), .CP(CLK), .Q(WX1982) ) ;
AND2    gate782  (.A(WX1663), .B(RESET), .Z(WX1983) ) ;
DFF     gate783  (.D(WX1983), .CP(CLK), .Q(WX1984) ) ;
AND2    gate784  (.A(WX1677), .B(RESET), .Z(WX1985) ) ;
DFF     gate785  (.D(WX1985), .CP(CLK), .Q(WX1986) ) ;
AND2    gate786  (.A(WX1691), .B(RESET), .Z(WX1987) ) ;
DFF     gate787  (.D(WX1987), .CP(CLK), .Q(WX1988) ) ;
AND2    gate788  (.A(WX1705), .B(RESET), .Z(WX1989) ) ;
DFF     gate789  (.D(WX1989), .CP(CLK), .Q(WX1990) ) ;
AND2    gate790  (.A(WX1719), .B(RESET), .Z(WX1991) ) ;
DFF     gate791  (.D(WX1991), .CP(CLK), .Q(WX1992) ) ;
AND2    gate792  (.A(WX1733), .B(RESET), .Z(WX1993) ) ;
DFF     gate793  (.D(WX1993), .CP(CLK), .Q(WX1994) ) ;
AND2    gate794  (.A(WX1747), .B(RESET), .Z(WX1995) ) ;
DFF     gate795  (.D(WX1995), .CP(CLK), .Q(WX1996) ) ;
AND2    gate796  (.A(WX1761), .B(RESET), .Z(WX1997) ) ;
DFF     gate797  (.D(WX1997), .CP(CLK), .Q(WX1998) ) ;
AND2    gate798  (.A(WX1775), .B(RESET), .Z(WX1999) ) ;
DFF     gate799  (.D(WX1999), .CP(CLK), .Q(WX2000) ) ;
AND2    gate800  (.A(WX1938), .B(RESET), .Z(WX2001) ) ;
DFF     gate801  (.D(WX2001), .CP(CLK), .Q(WX2002) ) ;
AND2    gate802  (.A(WX1940), .B(RESET), .Z(WX2003) ) ;
DFF     gate803  (.D(WX2003), .CP(CLK), .Q(WX2004) ) ;
AND2    gate804  (.A(WX1942), .B(RESET), .Z(WX2005) ) ;
DFF     gate805  (.D(WX2005), .CP(CLK), .Q(WX2006) ) ;
AND2    gate806  (.A(WX1944), .B(RESET), .Z(WX2007) ) ;
DFF     gate807  (.D(WX2007), .CP(CLK), .Q(WX2008) ) ;
AND2    gate808  (.A(WX1946), .B(RESET), .Z(WX2009) ) ;
DFF     gate809  (.D(WX2009), .CP(CLK), .Q(WX2010) ) ;
AND2    gate810  (.A(WX1948), .B(RESET), .Z(WX2011) ) ;
DFF     gate811  (.D(WX2011), .CP(CLK), .Q(WX2012) ) ;
AND2    gate812  (.A(WX1950), .B(RESET), .Z(WX2013) ) ;
DFF     gate813  (.D(WX2013), .CP(CLK), .Q(WX2014) ) ;
AND2    gate814  (.A(WX1952), .B(RESET), .Z(WX2015) ) ;
DFF     gate815  (.D(WX2015), .CP(CLK), .Q(WX2016) ) ;
AND2    gate816  (.A(WX1954), .B(RESET), .Z(WX2017) ) ;
DFF     gate817  (.D(WX2017), .CP(CLK), .Q(WX2018) ) ;
AND2    gate818  (.A(WX1956), .B(RESET), .Z(WX2019) ) ;
DFF     gate819  (.D(WX2019), .CP(CLK), .Q(WX2020) ) ;
AND2    gate820  (.A(WX1958), .B(RESET), .Z(WX2021) ) ;
DFF     gate821  (.D(WX2021), .CP(CLK), .Q(WX2022) ) ;
AND2    gate822  (.A(WX1960), .B(RESET), .Z(WX2023) ) ;
DFF     gate823  (.D(WX2023), .CP(CLK), .Q(WX2024) ) ;
AND2    gate824  (.A(WX1962), .B(RESET), .Z(WX2025) ) ;
DFF     gate825  (.D(WX2025), .CP(CLK), .Q(WX2026) ) ;
AND2    gate826  (.A(WX1964), .B(RESET), .Z(WX2027) ) ;
DFF     gate827  (.D(WX2027), .CP(CLK), .Q(WX2028) ) ;
AND2    gate828  (.A(WX1966), .B(RESET), .Z(WX2029) ) ;
DFF     gate829  (.D(WX2029), .CP(CLK), .Q(WX2030) ) ;
AND2    gate830  (.A(WX1968), .B(RESET), .Z(WX2031) ) ;
DFF     gate831  (.D(WX2031), .CP(CLK), .Q(WX2032) ) ;
AND2    gate832  (.A(WX1970), .B(RESET), .Z(WX2033) ) ;
DFF     gate833  (.D(WX2033), .CP(CLK), .Q(WX2034) ) ;
AND2    gate834  (.A(WX1972), .B(RESET), .Z(WX2035) ) ;
DFF     gate835  (.D(WX2035), .CP(CLK), .Q(WX2036) ) ;
AND2    gate836  (.A(WX1974), .B(RESET), .Z(WX2037) ) ;
DFF     gate837  (.D(WX2037), .CP(CLK), .Q(WX2038) ) ;
AND2    gate838  (.A(WX1976), .B(RESET), .Z(WX2039) ) ;
DFF     gate839  (.D(WX2039), .CP(CLK), .Q(WX2040) ) ;
AND2    gate840  (.A(WX1978), .B(RESET), .Z(WX2041) ) ;
DFF     gate841  (.D(WX2041), .CP(CLK), .Q(WX2042) ) ;
AND2    gate842  (.A(WX1980), .B(RESET), .Z(WX2043) ) ;
DFF     gate843  (.D(WX2043), .CP(CLK), .Q(WX2044) ) ;
AND2    gate844  (.A(WX1982), .B(RESET), .Z(WX2045) ) ;
DFF     gate845  (.D(WX2045), .CP(CLK), .Q(WX2046) ) ;
AND2    gate846  (.A(WX1984), .B(RESET), .Z(WX2047) ) ;
DFF     gate847  (.D(WX2047), .CP(CLK), .Q(WX2048) ) ;
AND2    gate848  (.A(WX1986), .B(RESET), .Z(WX2049) ) ;
DFF     gate849  (.D(WX2049), .CP(CLK), .Q(WX2050) ) ;
AND2    gate850  (.A(WX1988), .B(RESET), .Z(WX2051) ) ;
DFF     gate851  (.D(WX2051), .CP(CLK), .Q(WX2052) ) ;
AND2    gate852  (.A(WX1990), .B(RESET), .Z(WX2053) ) ;
DFF     gate853  (.D(WX2053), .CP(CLK), .Q(WX2054) ) ;
AND2    gate854  (.A(WX1992), .B(RESET), .Z(WX2055) ) ;
DFF     gate855  (.D(WX2055), .CP(CLK), .Q(WX2056) ) ;
AND2    gate856  (.A(WX1994), .B(RESET), .Z(WX2057) ) ;
DFF     gate857  (.D(WX2057), .CP(CLK), .Q(WX2058) ) ;
AND2    gate858  (.A(WX1996), .B(RESET), .Z(WX2059) ) ;
DFF     gate859  (.D(WX2059), .CP(CLK), .Q(WX2060) ) ;
AND2    gate860  (.A(WX1998), .B(RESET), .Z(WX2061) ) ;
DFF     gate861  (.D(WX2061), .CP(CLK), .Q(WX2062) ) ;
AND2    gate862  (.A(WX2000), .B(RESET), .Z(WX2063) ) ;
DFF     gate863  (.D(WX2063), .CP(CLK), .Q(WX2064) ) ;
AND2    gate864  (.A(WX2002), .B(RESET), .Z(WX2065) ) ;
DFF     gate865  (.D(WX2065), .CP(CLK), .Q(WX2066) ) ;
AND2    gate866  (.A(WX2004), .B(RESET), .Z(WX2067) ) ;
DFF     gate867  (.D(WX2067), .CP(CLK), .Q(WX2068) ) ;
AND2    gate868  (.A(WX2006), .B(RESET), .Z(WX2069) ) ;
DFF     gate869  (.D(WX2069), .CP(CLK), .Q(WX2070) ) ;
AND2    gate870  (.A(WX2008), .B(RESET), .Z(WX2071) ) ;
DFF     gate871  (.D(WX2071), .CP(CLK), .Q(WX2072) ) ;
AND2    gate872  (.A(WX2010), .B(RESET), .Z(WX2073) ) ;
DFF     gate873  (.D(WX2073), .CP(CLK), .Q(WX2074) ) ;
AND2    gate874  (.A(WX2012), .B(RESET), .Z(WX2075) ) ;
DFF     gate875  (.D(WX2075), .CP(CLK), .Q(WX2076) ) ;
AND2    gate876  (.A(WX2014), .B(RESET), .Z(WX2077) ) ;
DFF     gate877  (.D(WX2077), .CP(CLK), .Q(WX2078) ) ;
AND2    gate878  (.A(WX2016), .B(RESET), .Z(WX2079) ) ;
DFF     gate879  (.D(WX2079), .CP(CLK), .Q(WX2080) ) ;
AND2    gate880  (.A(WX2018), .B(RESET), .Z(WX2081) ) ;
DFF     gate881  (.D(WX2081), .CP(CLK), .Q(WX2082) ) ;
AND2    gate882  (.A(WX2020), .B(RESET), .Z(WX2083) ) ;
DFF     gate883  (.D(WX2083), .CP(CLK), .Q(WX2084) ) ;
AND2    gate884  (.A(WX2022), .B(RESET), .Z(WX2085) ) ;
DFF     gate885  (.D(WX2085), .CP(CLK), .Q(WX2086) ) ;
AND2    gate886  (.A(WX2024), .B(RESET), .Z(WX2087) ) ;
DFF     gate887  (.D(WX2087), .CP(CLK), .Q(WX2088) ) ;
AND2    gate888  (.A(WX2026), .B(RESET), .Z(WX2089) ) ;
DFF     gate889  (.D(WX2089), .CP(CLK), .Q(WX2090) ) ;
AND2    gate890  (.A(WX2028), .B(RESET), .Z(WX2091) ) ;
DFF     gate891  (.D(WX2091), .CP(CLK), .Q(WX2092) ) ;
AND2    gate892  (.A(WX2030), .B(RESET), .Z(WX2093) ) ;
DFF     gate893  (.D(WX2093), .CP(CLK), .Q(WX2094) ) ;
AND2    gate894  (.A(WX2032), .B(RESET), .Z(WX2095) ) ;
DFF     gate895  (.D(WX2095), .CP(CLK), .Q(WX2096) ) ;
AND2    gate896  (.A(WX2034), .B(RESET), .Z(WX2097) ) ;
DFF     gate897  (.D(WX2097), .CP(CLK), .Q(WX2098) ) ;
AND2    gate898  (.A(WX2036), .B(RESET), .Z(WX2099) ) ;
DFF     gate899  (.D(WX2099), .CP(CLK), .Q(WX2100) ) ;
AND2    gate900  (.A(WX2038), .B(RESET), .Z(WX2101) ) ;
DFF     gate901  (.D(WX2101), .CP(CLK), .Q(WX2102) ) ;
AND2    gate902  (.A(WX2040), .B(RESET), .Z(WX2103) ) ;
DFF     gate903  (.D(WX2103), .CP(CLK), .Q(WX2104) ) ;
AND2    gate904  (.A(WX2042), .B(RESET), .Z(WX2105) ) ;
DFF     gate905  (.D(WX2105), .CP(CLK), .Q(WX2106) ) ;
AND2    gate906  (.A(WX2044), .B(RESET), .Z(WX2107) ) ;
DFF     gate907  (.D(WX2107), .CP(CLK), .Q(WX2108) ) ;
AND2    gate908  (.A(WX2046), .B(RESET), .Z(WX2109) ) ;
DFF     gate909  (.D(WX2109), .CP(CLK), .Q(WX2110) ) ;
AND2    gate910  (.A(WX2048), .B(RESET), .Z(WX2111) ) ;
DFF     gate911  (.D(WX2111), .CP(CLK), .Q(WX2112) ) ;
AND2    gate912  (.A(WX2050), .B(RESET), .Z(WX2113) ) ;
DFF     gate913  (.D(WX2113), .CP(CLK), .Q(WX2114) ) ;
AND2    gate914  (.A(WX2052), .B(RESET), .Z(WX2115) ) ;
DFF     gate915  (.D(WX2115), .CP(CLK), .Q(WX2116) ) ;
AND2    gate916  (.A(WX2054), .B(RESET), .Z(WX2117) ) ;
DFF     gate917  (.D(WX2117), .CP(CLK), .Q(WX2118) ) ;
AND2    gate918  (.A(WX2056), .B(RESET), .Z(WX2119) ) ;
DFF     gate919  (.D(WX2119), .CP(CLK), .Q(WX2120) ) ;
AND2    gate920  (.A(WX2058), .B(RESET), .Z(WX2121) ) ;
DFF     gate921  (.D(WX2121), .CP(CLK), .Q(WX2122) ) ;
AND2    gate922  (.A(WX2060), .B(RESET), .Z(WX2123) ) ;
DFF     gate923  (.D(WX2123), .CP(CLK), .Q(WX2124) ) ;
AND2    gate924  (.A(WX2062), .B(RESET), .Z(WX2125) ) ;
DFF     gate925  (.D(WX2125), .CP(CLK), .Q(WX2126) ) ;
AND2    gate926  (.A(WX2064), .B(RESET), .Z(WX2127) ) ;
DFF     gate927  (.D(WX2127), .CP(CLK), .Q(WX2128) ) ;
AND2    gate928  (.A(WX2066), .B(RESET), .Z(WX2129) ) ;
DFF     gate929  (.D(WX2129), .CP(CLK), .Q(WX2130) ) ;
AND2    gate930  (.A(WX2068), .B(RESET), .Z(WX2131) ) ;
DFF     gate931  (.D(WX2131), .CP(CLK), .Q(WX2132) ) ;
AND2    gate932  (.A(WX2070), .B(RESET), .Z(WX2133) ) ;
DFF     gate933  (.D(WX2133), .CP(CLK), .Q(WX2134) ) ;
AND2    gate934  (.A(WX2072), .B(RESET), .Z(WX2135) ) ;
DFF     gate935  (.D(WX2135), .CP(CLK), .Q(WX2136) ) ;
AND2    gate936  (.A(WX2074), .B(RESET), .Z(WX2137) ) ;
DFF     gate937  (.D(WX2137), .CP(CLK), .Q(WX2138) ) ;
AND2    gate938  (.A(WX2076), .B(RESET), .Z(WX2139) ) ;
DFF     gate939  (.D(WX2139), .CP(CLK), .Q(WX2140) ) ;
AND2    gate940  (.A(WX2078), .B(RESET), .Z(WX2141) ) ;
DFF     gate941  (.D(WX2141), .CP(CLK), .Q(WX2142) ) ;
AND2    gate942  (.A(WX2080), .B(RESET), .Z(WX2143) ) ;
DFF     gate943  (.D(WX2143), .CP(CLK), .Q(WX2144) ) ;
AND2    gate944  (.A(WX2082), .B(RESET), .Z(WX2145) ) ;
DFF     gate945  (.D(WX2145), .CP(CLK), .Q(WX2146) ) ;
AND2    gate946  (.A(WX2084), .B(RESET), .Z(WX2147) ) ;
DFF     gate947  (.D(WX2147), .CP(CLK), .Q(WX2148) ) ;
AND2    gate948  (.A(WX2086), .B(RESET), .Z(WX2149) ) ;
DFF     gate949  (.D(WX2149), .CP(CLK), .Q(WX2150) ) ;
AND2    gate950  (.A(WX2088), .B(RESET), .Z(WX2151) ) ;
DFF     gate951  (.D(WX2151), .CP(CLK), .Q(WX2152) ) ;
AND2    gate952  (.A(WX2090), .B(RESET), .Z(WX2153) ) ;
DFF     gate953  (.D(WX2153), .CP(CLK), .Q(WX2154) ) ;
AND2    gate954  (.A(WX2092), .B(RESET), .Z(WX2155) ) ;
DFF     gate955  (.D(WX2155), .CP(CLK), .Q(WX2156) ) ;
AND2    gate956  (.A(WX2094), .B(RESET), .Z(WX2157) ) ;
DFF     gate957  (.D(WX2157), .CP(CLK), .Q(WX2158) ) ;
AND2    gate958  (.A(WX2096), .B(RESET), .Z(WX2159) ) ;
DFF     gate959  (.D(WX2159), .CP(CLK), .Q(WX2160) ) ;
AND2    gate960  (.A(WX2098), .B(RESET), .Z(WX2161) ) ;
DFF     gate961  (.D(WX2161), .CP(CLK), .Q(WX2162) ) ;
AND2    gate962  (.A(WX2100), .B(RESET), .Z(WX2163) ) ;
DFF     gate963  (.D(WX2163), .CP(CLK), .Q(WX2164) ) ;
AND2    gate964  (.A(WX2102), .B(RESET), .Z(WX2165) ) ;
DFF     gate965  (.D(WX2165), .CP(CLK), .Q(WX2166) ) ;
AND2    gate966  (.A(WX2104), .B(RESET), .Z(WX2167) ) ;
DFF     gate967  (.D(WX2167), .CP(CLK), .Q(WX2168) ) ;
AND2    gate968  (.A(WX2106), .B(RESET), .Z(WX2169) ) ;
DFF     gate969  (.D(WX2169), .CP(CLK), .Q(WX2170) ) ;
AND2    gate970  (.A(WX2108), .B(RESET), .Z(WX2171) ) ;
DFF     gate971  (.D(WX2171), .CP(CLK), .Q(WX2172) ) ;
AND2    gate972  (.A(WX2110), .B(RESET), .Z(WX2173) ) ;
DFF     gate973  (.D(WX2173), .CP(CLK), .Q(WX2174) ) ;
AND2    gate974  (.A(WX2112), .B(RESET), .Z(WX2175) ) ;
DFF     gate975  (.D(WX2175), .CP(CLK), .Q(WX2176) ) ;
AND2    gate976  (.A(WX2114), .B(RESET), .Z(WX2177) ) ;
DFF     gate977  (.D(WX2177), .CP(CLK), .Q(WX2178) ) ;
AND2    gate978  (.A(WX2116), .B(RESET), .Z(WX2179) ) ;
DFF     gate979  (.D(WX2179), .CP(CLK), .Q(WX2180) ) ;
AND2    gate980  (.A(WX2118), .B(RESET), .Z(WX2181) ) ;
DFF     gate981  (.D(WX2181), .CP(CLK), .Q(WX2182) ) ;
AND2    gate982  (.A(WX2120), .B(RESET), .Z(WX2183) ) ;
DFF     gate983  (.D(WX2183), .CP(CLK), .Q(WX2184) ) ;
AND2    gate984  (.A(WX2122), .B(RESET), .Z(WX2185) ) ;
DFF     gate985  (.D(WX2185), .CP(CLK), .Q(WX2186) ) ;
AND2    gate986  (.A(WX2124), .B(RESET), .Z(WX2187) ) ;
DFF     gate987  (.D(WX2187), .CP(CLK), .Q(WX2188) ) ;
AND2    gate988  (.A(WX2126), .B(RESET), .Z(WX2189) ) ;
DFF     gate989  (.D(WX2189), .CP(CLK), .Q(WX2190) ) ;
AND2    gate990  (.A(WX2128), .B(RESET), .Z(WX2191) ) ;
DFF     gate991  (.D(WX2191), .CP(CLK), .Q(WX2192) ) ;
AND2    gate992  (.A(WX2527), .B(WX2556), .Z(WX2557) ) ;
AND2    gate993  (.A(WX2555), .B(WX2556), .Z(WX2559) ) ;
AND2    gate994  (.A(WX2554), .B(WX2556), .Z(WX2561) ) ;
AND2    gate995  (.A(WX2553), .B(WX2556), .Z(WX2563) ) ;
AND2    gate996  (.A(WX2526), .B(WX2556), .Z(WX2565) ) ;
AND2    gate997  (.A(WX2552), .B(WX2556), .Z(WX2567) ) ;
AND2    gate998  (.A(WX2551), .B(WX2556), .Z(WX2569) ) ;
AND2    gate999  (.A(WX2550), .B(WX2556), .Z(WX2571) ) ;
AND2    gate1000  (.A(WX2549), .B(WX2556), .Z(WX2573) ) ;
AND2    gate1001  (.A(WX2548), .B(WX2556), .Z(WX2575) ) ;
AND2    gate1002  (.A(WX2547), .B(WX2556), .Z(WX2577) ) ;
AND2    gate1003  (.A(WX2525), .B(WX2556), .Z(WX2579) ) ;
AND2    gate1004  (.A(WX2546), .B(WX2556), .Z(WX2581) ) ;
AND2    gate1005  (.A(WX2545), .B(WX2556), .Z(WX2583) ) ;
AND2    gate1006  (.A(WX2544), .B(WX2556), .Z(WX2585) ) ;
AND2    gate1007  (.A(WX2543), .B(WX2556), .Z(WX2587) ) ;
AND2    gate1008  (.A(WX2524), .B(WX2556), .Z(WX2589) ) ;
AND2    gate1009  (.A(WX2542), .B(WX2556), .Z(WX2591) ) ;
AND2    gate1010  (.A(WX2541), .B(WX2556), .Z(WX2593) ) ;
AND2    gate1011  (.A(WX2540), .B(WX2556), .Z(WX2595) ) ;
AND2    gate1012  (.A(WX2539), .B(WX2556), .Z(WX2597) ) ;
AND2    gate1013  (.A(WX2538), .B(WX2556), .Z(WX2599) ) ;
AND2    gate1014  (.A(WX2537), .B(WX2556), .Z(WX2601) ) ;
AND2    gate1015  (.A(WX2536), .B(WX2556), .Z(WX2603) ) ;
AND2    gate1016  (.A(WX2535), .B(WX2556), .Z(WX2605) ) ;
AND2    gate1017  (.A(WX2534), .B(WX2556), .Z(WX2607) ) ;
AND2    gate1018  (.A(WX2533), .B(WX2556), .Z(WX2609) ) ;
AND2    gate1019  (.A(WX2532), .B(WX2556), .Z(WX2611) ) ;
AND2    gate1020  (.A(WX2531), .B(WX2556), .Z(WX2613) ) ;
AND2    gate1021  (.A(WX2530), .B(WX2556), .Z(WX2615) ) ;
AND2    gate1022  (.A(WX2529), .B(WX2556), .Z(WX2617) ) ;
AND2    gate1023  (.A(WX2528), .B(WX2556), .Z(WX2619) ) ;
AND2    gate1024  (.A(WX3073), .B(RESET), .Z(WX3070) ) ;
DFF     gate1025  (.D(WX3070), .CP(CLK), .Q(WX3071) ) ;
AND2    gate1026  (.A(WX3075), .B(RESET), .Z(WX3072) ) ;
DFF     gate1027  (.D(WX3072), .CP(CLK), .Q(WX3073) ) ;
AND2    gate1028  (.A(WX3077), .B(RESET), .Z(WX3074) ) ;
DFF     gate1029  (.D(WX3074), .CP(CLK), .Q(WX3075) ) ;
AND2    gate1030  (.A(WX3079), .B(RESET), .Z(WX3076) ) ;
DFF     gate1031  (.D(WX3076), .CP(CLK), .Q(WX3077) ) ;
AND2    gate1032  (.A(WX3081), .B(RESET), .Z(WX3078) ) ;
DFF     gate1033  (.D(WX3078), .CP(CLK), .Q(WX3079) ) ;
AND2    gate1034  (.A(WX3083), .B(RESET), .Z(WX3080) ) ;
DFF     gate1035  (.D(WX3080), .CP(CLK), .Q(WX3081) ) ;
AND2    gate1036  (.A(WX3085), .B(RESET), .Z(WX3082) ) ;
DFF     gate1037  (.D(WX3082), .CP(CLK), .Q(WX3083) ) ;
AND2    gate1038  (.A(WX3087), .B(RESET), .Z(WX3084) ) ;
DFF     gate1039  (.D(WX3084), .CP(CLK), .Q(WX3085) ) ;
AND2    gate1040  (.A(WX3089), .B(RESET), .Z(WX3086) ) ;
DFF     gate1041  (.D(WX3086), .CP(CLK), .Q(WX3087) ) ;
AND2    gate1042  (.A(WX3091), .B(RESET), .Z(WX3088) ) ;
DFF     gate1043  (.D(WX3088), .CP(CLK), .Q(WX3089) ) ;
AND2    gate1044  (.A(WX3093), .B(RESET), .Z(WX3090) ) ;
DFF     gate1045  (.D(WX3090), .CP(CLK), .Q(WX3091) ) ;
AND2    gate1046  (.A(WX3095), .B(RESET), .Z(WX3092) ) ;
DFF     gate1047  (.D(WX3092), .CP(CLK), .Q(WX3093) ) ;
AND2    gate1048  (.A(WX3097), .B(RESET), .Z(WX3094) ) ;
DFF     gate1049  (.D(WX3094), .CP(CLK), .Q(WX3095) ) ;
AND2    gate1050  (.A(WX3099), .B(RESET), .Z(WX3096) ) ;
DFF     gate1051  (.D(WX3096), .CP(CLK), .Q(WX3097) ) ;
AND2    gate1052  (.A(WX3101), .B(RESET), .Z(WX3098) ) ;
DFF     gate1053  (.D(WX3098), .CP(CLK), .Q(WX3099) ) ;
AND2    gate1054  (.A(WX3103), .B(RESET), .Z(WX3100) ) ;
DFF     gate1055  (.D(WX3100), .CP(CLK), .Q(WX3101) ) ;
AND2    gate1056  (.A(WX3105), .B(RESET), .Z(WX3102) ) ;
DFF     gate1057  (.D(WX3102), .CP(CLK), .Q(WX3103) ) ;
AND2    gate1058  (.A(WX3107), .B(RESET), .Z(WX3104) ) ;
DFF     gate1059  (.D(WX3104), .CP(CLK), .Q(WX3105) ) ;
AND2    gate1060  (.A(WX3109), .B(RESET), .Z(WX3106) ) ;
DFF     gate1061  (.D(WX3106), .CP(CLK), .Q(WX3107) ) ;
AND2    gate1062  (.A(WX3111), .B(RESET), .Z(WX3108) ) ;
DFF     gate1063  (.D(WX3108), .CP(CLK), .Q(WX3109) ) ;
AND2    gate1064  (.A(WX3113), .B(RESET), .Z(WX3110) ) ;
DFF     gate1065  (.D(WX3110), .CP(CLK), .Q(WX3111) ) ;
AND2    gate1066  (.A(WX3115), .B(RESET), .Z(WX3112) ) ;
DFF     gate1067  (.D(WX3112), .CP(CLK), .Q(WX3113) ) ;
AND2    gate1068  (.A(WX3117), .B(RESET), .Z(WX3114) ) ;
DFF     gate1069  (.D(WX3114), .CP(CLK), .Q(WX3115) ) ;
AND2    gate1070  (.A(WX3119), .B(RESET), .Z(WX3116) ) ;
DFF     gate1071  (.D(WX3116), .CP(CLK), .Q(WX3117) ) ;
AND2    gate1072  (.A(WX3121), .B(RESET), .Z(WX3118) ) ;
DFF     gate1073  (.D(WX3118), .CP(CLK), .Q(WX3119) ) ;
AND2    gate1074  (.A(WX3123), .B(RESET), .Z(WX3120) ) ;
DFF     gate1075  (.D(WX3120), .CP(CLK), .Q(WX3121) ) ;
AND2    gate1076  (.A(WX3125), .B(RESET), .Z(WX3122) ) ;
DFF     gate1077  (.D(WX3122), .CP(CLK), .Q(WX3123) ) ;
AND2    gate1078  (.A(WX3127), .B(RESET), .Z(WX3124) ) ;
DFF     gate1079  (.D(WX3124), .CP(CLK), .Q(WX3125) ) ;
AND2    gate1080  (.A(WX3129), .B(RESET), .Z(WX3126) ) ;
DFF     gate1081  (.D(WX3126), .CP(CLK), .Q(WX3127) ) ;
AND2    gate1082  (.A(WX3131), .B(RESET), .Z(WX3128) ) ;
DFF     gate1083  (.D(WX3128), .CP(CLK), .Q(WX3129) ) ;
AND2    gate1084  (.A(WX3133), .B(RESET), .Z(WX3130) ) ;
DFF     gate1085  (.D(WX3130), .CP(CLK), .Q(WX3131) ) ;
AND2    gate1086  (.A(WX3069), .B(RESET), .Z(WX3132) ) ;
DFF     gate1087  (.D(WX3132), .CP(CLK), .Q(WX3133) ) ;
AND2    gate1088  (.A(WX2634), .B(RESET), .Z(WX3230) ) ;
DFF     gate1089  (.D(WX3230), .CP(CLK), .Q(WX3231) ) ;
AND2    gate1090  (.A(WX2648), .B(RESET), .Z(WX3232) ) ;
DFF     gate1091  (.D(WX3232), .CP(CLK), .Q(WX3233) ) ;
AND2    gate1092  (.A(WX2662), .B(RESET), .Z(WX3234) ) ;
DFF     gate1093  (.D(WX3234), .CP(CLK), .Q(WX3235) ) ;
AND2    gate1094  (.A(WX2676), .B(RESET), .Z(WX3236) ) ;
DFF     gate1095  (.D(WX3236), .CP(CLK), .Q(WX3237) ) ;
AND2    gate1096  (.A(WX2690), .B(RESET), .Z(WX3238) ) ;
DFF     gate1097  (.D(WX3238), .CP(CLK), .Q(WX3239) ) ;
AND2    gate1098  (.A(WX2704), .B(RESET), .Z(WX3240) ) ;
DFF     gate1099  (.D(WX3240), .CP(CLK), .Q(WX3241) ) ;
AND2    gate1100  (.A(WX2718), .B(RESET), .Z(WX3242) ) ;
DFF     gate1101  (.D(WX3242), .CP(CLK), .Q(WX3243) ) ;
AND2    gate1102  (.A(WX2732), .B(RESET), .Z(WX3244) ) ;
DFF     gate1103  (.D(WX3244), .CP(CLK), .Q(WX3245) ) ;
AND2    gate1104  (.A(WX2746), .B(RESET), .Z(WX3246) ) ;
DFF     gate1105  (.D(WX3246), .CP(CLK), .Q(WX3247) ) ;
AND2    gate1106  (.A(WX2760), .B(RESET), .Z(WX3248) ) ;
DFF     gate1107  (.D(WX3248), .CP(CLK), .Q(WX3249) ) ;
AND2    gate1108  (.A(WX2774), .B(RESET), .Z(WX3250) ) ;
DFF     gate1109  (.D(WX3250), .CP(CLK), .Q(WX3251) ) ;
AND2    gate1110  (.A(WX2788), .B(RESET), .Z(WX3252) ) ;
DFF     gate1111  (.D(WX3252), .CP(CLK), .Q(WX3253) ) ;
AND2    gate1112  (.A(WX2802), .B(RESET), .Z(WX3254) ) ;
DFF     gate1113  (.D(WX3254), .CP(CLK), .Q(WX3255) ) ;
AND2    gate1114  (.A(WX2816), .B(RESET), .Z(WX3256) ) ;
DFF     gate1115  (.D(WX3256), .CP(CLK), .Q(WX3257) ) ;
AND2    gate1116  (.A(WX2830), .B(RESET), .Z(WX3258) ) ;
DFF     gate1117  (.D(WX3258), .CP(CLK), .Q(WX3259) ) ;
AND2    gate1118  (.A(WX2844), .B(RESET), .Z(WX3260) ) ;
DFF     gate1119  (.D(WX3260), .CP(CLK), .Q(WX3261) ) ;
AND2    gate1120  (.A(WX2858), .B(RESET), .Z(WX3262) ) ;
DFF     gate1121  (.D(WX3262), .CP(CLK), .Q(WX3263) ) ;
AND2    gate1122  (.A(WX2872), .B(RESET), .Z(WX3264) ) ;
DFF     gate1123  (.D(WX3264), .CP(CLK), .Q(WX3265) ) ;
AND2    gate1124  (.A(WX2886), .B(RESET), .Z(WX3266) ) ;
DFF     gate1125  (.D(WX3266), .CP(CLK), .Q(WX3267) ) ;
AND2    gate1126  (.A(WX2900), .B(RESET), .Z(WX3268) ) ;
DFF     gate1127  (.D(WX3268), .CP(CLK), .Q(WX3269) ) ;
AND2    gate1128  (.A(WX2914), .B(RESET), .Z(WX3270) ) ;
DFF     gate1129  (.D(WX3270), .CP(CLK), .Q(WX3271) ) ;
AND2    gate1130  (.A(WX2928), .B(RESET), .Z(WX3272) ) ;
DFF     gate1131  (.D(WX3272), .CP(CLK), .Q(WX3273) ) ;
AND2    gate1132  (.A(WX2942), .B(RESET), .Z(WX3274) ) ;
DFF     gate1133  (.D(WX3274), .CP(CLK), .Q(WX3275) ) ;
AND2    gate1134  (.A(WX2956), .B(RESET), .Z(WX3276) ) ;
DFF     gate1135  (.D(WX3276), .CP(CLK), .Q(WX3277) ) ;
AND2    gate1136  (.A(WX2970), .B(RESET), .Z(WX3278) ) ;
DFF     gate1137  (.D(WX3278), .CP(CLK), .Q(WX3279) ) ;
AND2    gate1138  (.A(WX2984), .B(RESET), .Z(WX3280) ) ;
DFF     gate1139  (.D(WX3280), .CP(CLK), .Q(WX3281) ) ;
AND2    gate1140  (.A(WX2998), .B(RESET), .Z(WX3282) ) ;
DFF     gate1141  (.D(WX3282), .CP(CLK), .Q(WX3283) ) ;
AND2    gate1142  (.A(WX3012), .B(RESET), .Z(WX3284) ) ;
DFF     gate1143  (.D(WX3284), .CP(CLK), .Q(WX3285) ) ;
AND2    gate1144  (.A(WX3026), .B(RESET), .Z(WX3286) ) ;
DFF     gate1145  (.D(WX3286), .CP(CLK), .Q(WX3287) ) ;
AND2    gate1146  (.A(WX3040), .B(RESET), .Z(WX3288) ) ;
DFF     gate1147  (.D(WX3288), .CP(CLK), .Q(WX3289) ) ;
AND2    gate1148  (.A(WX3054), .B(RESET), .Z(WX3290) ) ;
DFF     gate1149  (.D(WX3290), .CP(CLK), .Q(WX3291) ) ;
AND2    gate1150  (.A(WX3068), .B(RESET), .Z(WX3292) ) ;
DFF     gate1151  (.D(WX3292), .CP(CLK), .Q(WX3293) ) ;
AND2    gate1152  (.A(WX3231), .B(RESET), .Z(WX3294) ) ;
DFF     gate1153  (.D(WX3294), .CP(CLK), .Q(WX3295) ) ;
AND2    gate1154  (.A(WX3233), .B(RESET), .Z(WX3296) ) ;
DFF     gate1155  (.D(WX3296), .CP(CLK), .Q(WX3297) ) ;
AND2    gate1156  (.A(WX3235), .B(RESET), .Z(WX3298) ) ;
DFF     gate1157  (.D(WX3298), .CP(CLK), .Q(WX3299) ) ;
AND2    gate1158  (.A(WX3237), .B(RESET), .Z(WX3300) ) ;
DFF     gate1159  (.D(WX3300), .CP(CLK), .Q(WX3301) ) ;
AND2    gate1160  (.A(WX3239), .B(RESET), .Z(WX3302) ) ;
DFF     gate1161  (.D(WX3302), .CP(CLK), .Q(WX3303) ) ;
AND2    gate1162  (.A(WX3241), .B(RESET), .Z(WX3304) ) ;
DFF     gate1163  (.D(WX3304), .CP(CLK), .Q(WX3305) ) ;
AND2    gate1164  (.A(WX3243), .B(RESET), .Z(WX3306) ) ;
DFF     gate1165  (.D(WX3306), .CP(CLK), .Q(WX3307) ) ;
AND2    gate1166  (.A(WX3245), .B(RESET), .Z(WX3308) ) ;
DFF     gate1167  (.D(WX3308), .CP(CLK), .Q(WX3309) ) ;
AND2    gate1168  (.A(WX3247), .B(RESET), .Z(WX3310) ) ;
DFF     gate1169  (.D(WX3310), .CP(CLK), .Q(WX3311) ) ;
AND2    gate1170  (.A(WX3249), .B(RESET), .Z(WX3312) ) ;
DFF     gate1171  (.D(WX3312), .CP(CLK), .Q(WX3313) ) ;
AND2    gate1172  (.A(WX3251), .B(RESET), .Z(WX3314) ) ;
DFF     gate1173  (.D(WX3314), .CP(CLK), .Q(WX3315) ) ;
AND2    gate1174  (.A(WX3253), .B(RESET), .Z(WX3316) ) ;
DFF     gate1175  (.D(WX3316), .CP(CLK), .Q(WX3317) ) ;
AND2    gate1176  (.A(WX3255), .B(RESET), .Z(WX3318) ) ;
DFF     gate1177  (.D(WX3318), .CP(CLK), .Q(WX3319) ) ;
AND2    gate1178  (.A(WX3257), .B(RESET), .Z(WX3320) ) ;
DFF     gate1179  (.D(WX3320), .CP(CLK), .Q(WX3321) ) ;
AND2    gate1180  (.A(WX3259), .B(RESET), .Z(WX3322) ) ;
DFF     gate1181  (.D(WX3322), .CP(CLK), .Q(WX3323) ) ;
AND2    gate1182  (.A(WX3261), .B(RESET), .Z(WX3324) ) ;
DFF     gate1183  (.D(WX3324), .CP(CLK), .Q(WX3325) ) ;
AND2    gate1184  (.A(WX3263), .B(RESET), .Z(WX3326) ) ;
DFF     gate1185  (.D(WX3326), .CP(CLK), .Q(WX3327) ) ;
AND2    gate1186  (.A(WX3265), .B(RESET), .Z(WX3328) ) ;
DFF     gate1187  (.D(WX3328), .CP(CLK), .Q(WX3329) ) ;
AND2    gate1188  (.A(WX3267), .B(RESET), .Z(WX3330) ) ;
DFF     gate1189  (.D(WX3330), .CP(CLK), .Q(WX3331) ) ;
AND2    gate1190  (.A(WX3269), .B(RESET), .Z(WX3332) ) ;
DFF     gate1191  (.D(WX3332), .CP(CLK), .Q(WX3333) ) ;
AND2    gate1192  (.A(WX3271), .B(RESET), .Z(WX3334) ) ;
DFF     gate1193  (.D(WX3334), .CP(CLK), .Q(WX3335) ) ;
AND2    gate1194  (.A(WX3273), .B(RESET), .Z(WX3336) ) ;
DFF     gate1195  (.D(WX3336), .CP(CLK), .Q(WX3337) ) ;
AND2    gate1196  (.A(WX3275), .B(RESET), .Z(WX3338) ) ;
DFF     gate1197  (.D(WX3338), .CP(CLK), .Q(WX3339) ) ;
AND2    gate1198  (.A(WX3277), .B(RESET), .Z(WX3340) ) ;
DFF     gate1199  (.D(WX3340), .CP(CLK), .Q(WX3341) ) ;
AND2    gate1200  (.A(WX3279), .B(RESET), .Z(WX3342) ) ;
DFF     gate1201  (.D(WX3342), .CP(CLK), .Q(WX3343) ) ;
AND2    gate1202  (.A(WX3281), .B(RESET), .Z(WX3344) ) ;
DFF     gate1203  (.D(WX3344), .CP(CLK), .Q(WX3345) ) ;
AND2    gate1204  (.A(WX3283), .B(RESET), .Z(WX3346) ) ;
DFF     gate1205  (.D(WX3346), .CP(CLK), .Q(WX3347) ) ;
AND2    gate1206  (.A(WX3285), .B(RESET), .Z(WX3348) ) ;
DFF     gate1207  (.D(WX3348), .CP(CLK), .Q(WX3349) ) ;
AND2    gate1208  (.A(WX3287), .B(RESET), .Z(WX3350) ) ;
DFF     gate1209  (.D(WX3350), .CP(CLK), .Q(WX3351) ) ;
AND2    gate1210  (.A(WX3289), .B(RESET), .Z(WX3352) ) ;
DFF     gate1211  (.D(WX3352), .CP(CLK), .Q(WX3353) ) ;
AND2    gate1212  (.A(WX3291), .B(RESET), .Z(WX3354) ) ;
DFF     gate1213  (.D(WX3354), .CP(CLK), .Q(WX3355) ) ;
AND2    gate1214  (.A(WX3293), .B(RESET), .Z(WX3356) ) ;
DFF     gate1215  (.D(WX3356), .CP(CLK), .Q(WX3357) ) ;
AND2    gate1216  (.A(WX3295), .B(RESET), .Z(WX3358) ) ;
DFF     gate1217  (.D(WX3358), .CP(CLK), .Q(WX3359) ) ;
AND2    gate1218  (.A(WX3297), .B(RESET), .Z(WX3360) ) ;
DFF     gate1219  (.D(WX3360), .CP(CLK), .Q(WX3361) ) ;
AND2    gate1220  (.A(WX3299), .B(RESET), .Z(WX3362) ) ;
DFF     gate1221  (.D(WX3362), .CP(CLK), .Q(WX3363) ) ;
AND2    gate1222  (.A(WX3301), .B(RESET), .Z(WX3364) ) ;
DFF     gate1223  (.D(WX3364), .CP(CLK), .Q(WX3365) ) ;
AND2    gate1224  (.A(WX3303), .B(RESET), .Z(WX3366) ) ;
DFF     gate1225  (.D(WX3366), .CP(CLK), .Q(WX3367) ) ;
AND2    gate1226  (.A(WX3305), .B(RESET), .Z(WX3368) ) ;
DFF     gate1227  (.D(WX3368), .CP(CLK), .Q(WX3369) ) ;
AND2    gate1228  (.A(WX3307), .B(RESET), .Z(WX3370) ) ;
DFF     gate1229  (.D(WX3370), .CP(CLK), .Q(WX3371) ) ;
AND2    gate1230  (.A(WX3309), .B(RESET), .Z(WX3372) ) ;
DFF     gate1231  (.D(WX3372), .CP(CLK), .Q(WX3373) ) ;
AND2    gate1232  (.A(WX3311), .B(RESET), .Z(WX3374) ) ;
DFF     gate1233  (.D(WX3374), .CP(CLK), .Q(WX3375) ) ;
AND2    gate1234  (.A(WX3313), .B(RESET), .Z(WX3376) ) ;
DFF     gate1235  (.D(WX3376), .CP(CLK), .Q(WX3377) ) ;
AND2    gate1236  (.A(WX3315), .B(RESET), .Z(WX3378) ) ;
DFF     gate1237  (.D(WX3378), .CP(CLK), .Q(WX3379) ) ;
AND2    gate1238  (.A(WX3317), .B(RESET), .Z(WX3380) ) ;
DFF     gate1239  (.D(WX3380), .CP(CLK), .Q(WX3381) ) ;
AND2    gate1240  (.A(WX3319), .B(RESET), .Z(WX3382) ) ;
DFF     gate1241  (.D(WX3382), .CP(CLK), .Q(WX3383) ) ;
AND2    gate1242  (.A(WX3321), .B(RESET), .Z(WX3384) ) ;
DFF     gate1243  (.D(WX3384), .CP(CLK), .Q(WX3385) ) ;
AND2    gate1244  (.A(WX3323), .B(RESET), .Z(WX3386) ) ;
DFF     gate1245  (.D(WX3386), .CP(CLK), .Q(WX3387) ) ;
AND2    gate1246  (.A(WX3325), .B(RESET), .Z(WX3388) ) ;
DFF     gate1247  (.D(WX3388), .CP(CLK), .Q(WX3389) ) ;
AND2    gate1248  (.A(WX3327), .B(RESET), .Z(WX3390) ) ;
DFF     gate1249  (.D(WX3390), .CP(CLK), .Q(WX3391) ) ;
AND2    gate1250  (.A(WX3329), .B(RESET), .Z(WX3392) ) ;
DFF     gate1251  (.D(WX3392), .CP(CLK), .Q(WX3393) ) ;
AND2    gate1252  (.A(WX3331), .B(RESET), .Z(WX3394) ) ;
DFF     gate1253  (.D(WX3394), .CP(CLK), .Q(WX3395) ) ;
AND2    gate1254  (.A(WX3333), .B(RESET), .Z(WX3396) ) ;
DFF     gate1255  (.D(WX3396), .CP(CLK), .Q(WX3397) ) ;
AND2    gate1256  (.A(WX3335), .B(RESET), .Z(WX3398) ) ;
DFF     gate1257  (.D(WX3398), .CP(CLK), .Q(WX3399) ) ;
AND2    gate1258  (.A(WX3337), .B(RESET), .Z(WX3400) ) ;
DFF     gate1259  (.D(WX3400), .CP(CLK), .Q(WX3401) ) ;
AND2    gate1260  (.A(WX3339), .B(RESET), .Z(WX3402) ) ;
DFF     gate1261  (.D(WX3402), .CP(CLK), .Q(WX3403) ) ;
AND2    gate1262  (.A(WX3341), .B(RESET), .Z(WX3404) ) ;
DFF     gate1263  (.D(WX3404), .CP(CLK), .Q(WX3405) ) ;
AND2    gate1264  (.A(WX3343), .B(RESET), .Z(WX3406) ) ;
DFF     gate1265  (.D(WX3406), .CP(CLK), .Q(WX3407) ) ;
AND2    gate1266  (.A(WX3345), .B(RESET), .Z(WX3408) ) ;
DFF     gate1267  (.D(WX3408), .CP(CLK), .Q(WX3409) ) ;
AND2    gate1268  (.A(WX3347), .B(RESET), .Z(WX3410) ) ;
DFF     gate1269  (.D(WX3410), .CP(CLK), .Q(WX3411) ) ;
AND2    gate1270  (.A(WX3349), .B(RESET), .Z(WX3412) ) ;
DFF     gate1271  (.D(WX3412), .CP(CLK), .Q(WX3413) ) ;
AND2    gate1272  (.A(WX3351), .B(RESET), .Z(WX3414) ) ;
DFF     gate1273  (.D(WX3414), .CP(CLK), .Q(WX3415) ) ;
AND2    gate1274  (.A(WX3353), .B(RESET), .Z(WX3416) ) ;
DFF     gate1275  (.D(WX3416), .CP(CLK), .Q(WX3417) ) ;
AND2    gate1276  (.A(WX3355), .B(RESET), .Z(WX3418) ) ;
DFF     gate1277  (.D(WX3418), .CP(CLK), .Q(WX3419) ) ;
AND2    gate1278  (.A(WX3357), .B(RESET), .Z(WX3420) ) ;
DFF     gate1279  (.D(WX3420), .CP(CLK), .Q(WX3421) ) ;
AND2    gate1280  (.A(WX3359), .B(RESET), .Z(WX3422) ) ;
DFF     gate1281  (.D(WX3422), .CP(CLK), .Q(WX3423) ) ;
AND2    gate1282  (.A(WX3361), .B(RESET), .Z(WX3424) ) ;
DFF     gate1283  (.D(WX3424), .CP(CLK), .Q(WX3425) ) ;
AND2    gate1284  (.A(WX3363), .B(RESET), .Z(WX3426) ) ;
DFF     gate1285  (.D(WX3426), .CP(CLK), .Q(WX3427) ) ;
AND2    gate1286  (.A(WX3365), .B(RESET), .Z(WX3428) ) ;
DFF     gate1287  (.D(WX3428), .CP(CLK), .Q(WX3429) ) ;
AND2    gate1288  (.A(WX3367), .B(RESET), .Z(WX3430) ) ;
DFF     gate1289  (.D(WX3430), .CP(CLK), .Q(WX3431) ) ;
AND2    gate1290  (.A(WX3369), .B(RESET), .Z(WX3432) ) ;
DFF     gate1291  (.D(WX3432), .CP(CLK), .Q(WX3433) ) ;
AND2    gate1292  (.A(WX3371), .B(RESET), .Z(WX3434) ) ;
DFF     gate1293  (.D(WX3434), .CP(CLK), .Q(WX3435) ) ;
AND2    gate1294  (.A(WX3373), .B(RESET), .Z(WX3436) ) ;
DFF     gate1295  (.D(WX3436), .CP(CLK), .Q(WX3437) ) ;
AND2    gate1296  (.A(WX3375), .B(RESET), .Z(WX3438) ) ;
DFF     gate1297  (.D(WX3438), .CP(CLK), .Q(WX3439) ) ;
AND2    gate1298  (.A(WX3377), .B(RESET), .Z(WX3440) ) ;
DFF     gate1299  (.D(WX3440), .CP(CLK), .Q(WX3441) ) ;
AND2    gate1300  (.A(WX3379), .B(RESET), .Z(WX3442) ) ;
DFF     gate1301  (.D(WX3442), .CP(CLK), .Q(WX3443) ) ;
AND2    gate1302  (.A(WX3381), .B(RESET), .Z(WX3444) ) ;
DFF     gate1303  (.D(WX3444), .CP(CLK), .Q(WX3445) ) ;
AND2    gate1304  (.A(WX3383), .B(RESET), .Z(WX3446) ) ;
DFF     gate1305  (.D(WX3446), .CP(CLK), .Q(WX3447) ) ;
AND2    gate1306  (.A(WX3385), .B(RESET), .Z(WX3448) ) ;
DFF     gate1307  (.D(WX3448), .CP(CLK), .Q(WX3449) ) ;
AND2    gate1308  (.A(WX3387), .B(RESET), .Z(WX3450) ) ;
DFF     gate1309  (.D(WX3450), .CP(CLK), .Q(WX3451) ) ;
AND2    gate1310  (.A(WX3389), .B(RESET), .Z(WX3452) ) ;
DFF     gate1311  (.D(WX3452), .CP(CLK), .Q(WX3453) ) ;
AND2    gate1312  (.A(WX3391), .B(RESET), .Z(WX3454) ) ;
DFF     gate1313  (.D(WX3454), .CP(CLK), .Q(WX3455) ) ;
AND2    gate1314  (.A(WX3393), .B(RESET), .Z(WX3456) ) ;
DFF     gate1315  (.D(WX3456), .CP(CLK), .Q(WX3457) ) ;
AND2    gate1316  (.A(WX3395), .B(RESET), .Z(WX3458) ) ;
DFF     gate1317  (.D(WX3458), .CP(CLK), .Q(WX3459) ) ;
AND2    gate1318  (.A(WX3397), .B(RESET), .Z(WX3460) ) ;
DFF     gate1319  (.D(WX3460), .CP(CLK), .Q(WX3461) ) ;
AND2    gate1320  (.A(WX3399), .B(RESET), .Z(WX3462) ) ;
DFF     gate1321  (.D(WX3462), .CP(CLK), .Q(WX3463) ) ;
AND2    gate1322  (.A(WX3401), .B(RESET), .Z(WX3464) ) ;
DFF     gate1323  (.D(WX3464), .CP(CLK), .Q(WX3465) ) ;
AND2    gate1324  (.A(WX3403), .B(RESET), .Z(WX3466) ) ;
DFF     gate1325  (.D(WX3466), .CP(CLK), .Q(WX3467) ) ;
AND2    gate1326  (.A(WX3405), .B(RESET), .Z(WX3468) ) ;
DFF     gate1327  (.D(WX3468), .CP(CLK), .Q(WX3469) ) ;
AND2    gate1328  (.A(WX3407), .B(RESET), .Z(WX3470) ) ;
DFF     gate1329  (.D(WX3470), .CP(CLK), .Q(WX3471) ) ;
AND2    gate1330  (.A(WX3409), .B(RESET), .Z(WX3472) ) ;
DFF     gate1331  (.D(WX3472), .CP(CLK), .Q(WX3473) ) ;
AND2    gate1332  (.A(WX3411), .B(RESET), .Z(WX3474) ) ;
DFF     gate1333  (.D(WX3474), .CP(CLK), .Q(WX3475) ) ;
AND2    gate1334  (.A(WX3413), .B(RESET), .Z(WX3476) ) ;
DFF     gate1335  (.D(WX3476), .CP(CLK), .Q(WX3477) ) ;
AND2    gate1336  (.A(WX3415), .B(RESET), .Z(WX3478) ) ;
DFF     gate1337  (.D(WX3478), .CP(CLK), .Q(WX3479) ) ;
AND2    gate1338  (.A(WX3417), .B(RESET), .Z(WX3480) ) ;
DFF     gate1339  (.D(WX3480), .CP(CLK), .Q(WX3481) ) ;
AND2    gate1340  (.A(WX3419), .B(RESET), .Z(WX3482) ) ;
DFF     gate1341  (.D(WX3482), .CP(CLK), .Q(WX3483) ) ;
AND2    gate1342  (.A(WX3421), .B(RESET), .Z(WX3484) ) ;
DFF     gate1343  (.D(WX3484), .CP(CLK), .Q(WX3485) ) ;
AND2    gate1344  (.A(WX3820), .B(WX3849), .Z(WX3850) ) ;
AND2    gate1345  (.A(WX3848), .B(WX3849), .Z(WX3852) ) ;
AND2    gate1346  (.A(WX3847), .B(WX3849), .Z(WX3854) ) ;
AND2    gate1347  (.A(WX3846), .B(WX3849), .Z(WX3856) ) ;
AND2    gate1348  (.A(WX3819), .B(WX3849), .Z(WX3858) ) ;
AND2    gate1349  (.A(WX3845), .B(WX3849), .Z(WX3860) ) ;
AND2    gate1350  (.A(WX3844), .B(WX3849), .Z(WX3862) ) ;
AND2    gate1351  (.A(WX3843), .B(WX3849), .Z(WX3864) ) ;
AND2    gate1352  (.A(WX3842), .B(WX3849), .Z(WX3866) ) ;
AND2    gate1353  (.A(WX3841), .B(WX3849), .Z(WX3868) ) ;
AND2    gate1354  (.A(WX3840), .B(WX3849), .Z(WX3870) ) ;
AND2    gate1355  (.A(WX3818), .B(WX3849), .Z(WX3872) ) ;
AND2    gate1356  (.A(WX3839), .B(WX3849), .Z(WX3874) ) ;
AND2    gate1357  (.A(WX3838), .B(WX3849), .Z(WX3876) ) ;
AND2    gate1358  (.A(WX3837), .B(WX3849), .Z(WX3878) ) ;
AND2    gate1359  (.A(WX3836), .B(WX3849), .Z(WX3880) ) ;
AND2    gate1360  (.A(WX3817), .B(WX3849), .Z(WX3882) ) ;
AND2    gate1361  (.A(WX3835), .B(WX3849), .Z(WX3884) ) ;
AND2    gate1362  (.A(WX3834), .B(WX3849), .Z(WX3886) ) ;
AND2    gate1363  (.A(WX3833), .B(WX3849), .Z(WX3888) ) ;
AND2    gate1364  (.A(WX3832), .B(WX3849), .Z(WX3890) ) ;
AND2    gate1365  (.A(WX3831), .B(WX3849), .Z(WX3892) ) ;
AND2    gate1366  (.A(WX3830), .B(WX3849), .Z(WX3894) ) ;
AND2    gate1367  (.A(WX3829), .B(WX3849), .Z(WX3896) ) ;
AND2    gate1368  (.A(WX3828), .B(WX3849), .Z(WX3898) ) ;
AND2    gate1369  (.A(WX3827), .B(WX3849), .Z(WX3900) ) ;
AND2    gate1370  (.A(WX3826), .B(WX3849), .Z(WX3902) ) ;
AND2    gate1371  (.A(WX3825), .B(WX3849), .Z(WX3904) ) ;
AND2    gate1372  (.A(WX3824), .B(WX3849), .Z(WX3906) ) ;
AND2    gate1373  (.A(WX3823), .B(WX3849), .Z(WX3908) ) ;
AND2    gate1374  (.A(WX3822), .B(WX3849), .Z(WX3910) ) ;
AND2    gate1375  (.A(WX3821), .B(WX3849), .Z(WX3912) ) ;
AND2    gate1376  (.A(WX4366), .B(RESET), .Z(WX4363) ) ;
DFF     gate1377  (.D(WX4363), .CP(CLK), .Q(WX4364) ) ;
AND2    gate1378  (.A(WX4368), .B(RESET), .Z(WX4365) ) ;
DFF     gate1379  (.D(WX4365), .CP(CLK), .Q(WX4366) ) ;
AND2    gate1380  (.A(WX4370), .B(RESET), .Z(WX4367) ) ;
DFF     gate1381  (.D(WX4367), .CP(CLK), .Q(WX4368) ) ;
AND2    gate1382  (.A(WX4372), .B(RESET), .Z(WX4369) ) ;
DFF     gate1383  (.D(WX4369), .CP(CLK), .Q(WX4370) ) ;
AND2    gate1384  (.A(WX4374), .B(RESET), .Z(WX4371) ) ;
DFF     gate1385  (.D(WX4371), .CP(CLK), .Q(WX4372) ) ;
AND2    gate1386  (.A(WX4376), .B(RESET), .Z(WX4373) ) ;
DFF     gate1387  (.D(WX4373), .CP(CLK), .Q(WX4374) ) ;
AND2    gate1388  (.A(WX4378), .B(RESET), .Z(WX4375) ) ;
DFF     gate1389  (.D(WX4375), .CP(CLK), .Q(WX4376) ) ;
AND2    gate1390  (.A(WX4380), .B(RESET), .Z(WX4377) ) ;
DFF     gate1391  (.D(WX4377), .CP(CLK), .Q(WX4378) ) ;
AND2    gate1392  (.A(WX4382), .B(RESET), .Z(WX4379) ) ;
DFF     gate1393  (.D(WX4379), .CP(CLK), .Q(WX4380) ) ;
AND2    gate1394  (.A(WX4384), .B(RESET), .Z(WX4381) ) ;
DFF     gate1395  (.D(WX4381), .CP(CLK), .Q(WX4382) ) ;
AND2    gate1396  (.A(WX4386), .B(RESET), .Z(WX4383) ) ;
DFF     gate1397  (.D(WX4383), .CP(CLK), .Q(WX4384) ) ;
AND2    gate1398  (.A(WX4388), .B(RESET), .Z(WX4385) ) ;
DFF     gate1399  (.D(WX4385), .CP(CLK), .Q(WX4386) ) ;
AND2    gate1400  (.A(WX4390), .B(RESET), .Z(WX4387) ) ;
DFF     gate1401  (.D(WX4387), .CP(CLK), .Q(WX4388) ) ;
AND2    gate1402  (.A(WX4392), .B(RESET), .Z(WX4389) ) ;
DFF     gate1403  (.D(WX4389), .CP(CLK), .Q(WX4390) ) ;
AND2    gate1404  (.A(WX4394), .B(RESET), .Z(WX4391) ) ;
DFF     gate1405  (.D(WX4391), .CP(CLK), .Q(WX4392) ) ;
AND2    gate1406  (.A(WX4396), .B(RESET), .Z(WX4393) ) ;
DFF     gate1407  (.D(WX4393), .CP(CLK), .Q(WX4394) ) ;
AND2    gate1408  (.A(WX4398), .B(RESET), .Z(WX4395) ) ;
DFF     gate1409  (.D(WX4395), .CP(CLK), .Q(WX4396) ) ;
AND2    gate1410  (.A(WX4400), .B(RESET), .Z(WX4397) ) ;
DFF     gate1411  (.D(WX4397), .CP(CLK), .Q(WX4398) ) ;
AND2    gate1412  (.A(WX4402), .B(RESET), .Z(WX4399) ) ;
DFF     gate1413  (.D(WX4399), .CP(CLK), .Q(WX4400) ) ;
AND2    gate1414  (.A(WX4404), .B(RESET), .Z(WX4401) ) ;
DFF     gate1415  (.D(WX4401), .CP(CLK), .Q(WX4402) ) ;
AND2    gate1416  (.A(WX4406), .B(RESET), .Z(WX4403) ) ;
DFF     gate1417  (.D(WX4403), .CP(CLK), .Q(WX4404) ) ;
AND2    gate1418  (.A(WX4408), .B(RESET), .Z(WX4405) ) ;
DFF     gate1419  (.D(WX4405), .CP(CLK), .Q(WX4406) ) ;
AND2    gate1420  (.A(WX4410), .B(RESET), .Z(WX4407) ) ;
DFF     gate1421  (.D(WX4407), .CP(CLK), .Q(WX4408) ) ;
AND2    gate1422  (.A(WX4412), .B(RESET), .Z(WX4409) ) ;
DFF     gate1423  (.D(WX4409), .CP(CLK), .Q(WX4410) ) ;
AND2    gate1424  (.A(WX4414), .B(RESET), .Z(WX4411) ) ;
DFF     gate1425  (.D(WX4411), .CP(CLK), .Q(WX4412) ) ;
AND2    gate1426  (.A(WX4416), .B(RESET), .Z(WX4413) ) ;
DFF     gate1427  (.D(WX4413), .CP(CLK), .Q(WX4414) ) ;
AND2    gate1428  (.A(WX4418), .B(RESET), .Z(WX4415) ) ;
DFF     gate1429  (.D(WX4415), .CP(CLK), .Q(WX4416) ) ;
AND2    gate1430  (.A(WX4420), .B(RESET), .Z(WX4417) ) ;
DFF     gate1431  (.D(WX4417), .CP(CLK), .Q(WX4418) ) ;
AND2    gate1432  (.A(WX4422), .B(RESET), .Z(WX4419) ) ;
DFF     gate1433  (.D(WX4419), .CP(CLK), .Q(WX4420) ) ;
AND2    gate1434  (.A(WX4424), .B(RESET), .Z(WX4421) ) ;
DFF     gate1435  (.D(WX4421), .CP(CLK), .Q(WX4422) ) ;
AND2    gate1436  (.A(WX4426), .B(RESET), .Z(WX4423) ) ;
DFF     gate1437  (.D(WX4423), .CP(CLK), .Q(WX4424) ) ;
AND2    gate1438  (.A(WX4362), .B(RESET), .Z(WX4425) ) ;
DFF     gate1439  (.D(WX4425), .CP(CLK), .Q(WX4426) ) ;
AND2    gate1440  (.A(WX3927), .B(RESET), .Z(WX4523) ) ;
DFF     gate1441  (.D(WX4523), .CP(CLK), .Q(WX4524) ) ;
AND2    gate1442  (.A(WX3941), .B(RESET), .Z(WX4525) ) ;
DFF     gate1443  (.D(WX4525), .CP(CLK), .Q(WX4526) ) ;
AND2    gate1444  (.A(WX3955), .B(RESET), .Z(WX4527) ) ;
DFF     gate1445  (.D(WX4527), .CP(CLK), .Q(WX4528) ) ;
AND2    gate1446  (.A(WX3969), .B(RESET), .Z(WX4529) ) ;
DFF     gate1447  (.D(WX4529), .CP(CLK), .Q(WX4530) ) ;
AND2    gate1448  (.A(WX3983), .B(RESET), .Z(WX4531) ) ;
DFF     gate1449  (.D(WX4531), .CP(CLK), .Q(WX4532) ) ;
AND2    gate1450  (.A(WX3997), .B(RESET), .Z(WX4533) ) ;
DFF     gate1451  (.D(WX4533), .CP(CLK), .Q(WX4534) ) ;
AND2    gate1452  (.A(WX4011), .B(RESET), .Z(WX4535) ) ;
DFF     gate1453  (.D(WX4535), .CP(CLK), .Q(WX4536) ) ;
AND2    gate1454  (.A(WX4025), .B(RESET), .Z(WX4537) ) ;
DFF     gate1455  (.D(WX4537), .CP(CLK), .Q(WX4538) ) ;
AND2    gate1456  (.A(WX4039), .B(RESET), .Z(WX4539) ) ;
DFF     gate1457  (.D(WX4539), .CP(CLK), .Q(WX4540) ) ;
AND2    gate1458  (.A(WX4053), .B(RESET), .Z(WX4541) ) ;
DFF     gate1459  (.D(WX4541), .CP(CLK), .Q(WX4542) ) ;
AND2    gate1460  (.A(WX4067), .B(RESET), .Z(WX4543) ) ;
DFF     gate1461  (.D(WX4543), .CP(CLK), .Q(WX4544) ) ;
AND2    gate1462  (.A(WX4081), .B(RESET), .Z(WX4545) ) ;
DFF     gate1463  (.D(WX4545), .CP(CLK), .Q(WX4546) ) ;
AND2    gate1464  (.A(WX4095), .B(RESET), .Z(WX4547) ) ;
DFF     gate1465  (.D(WX4547), .CP(CLK), .Q(WX4548) ) ;
AND2    gate1466  (.A(WX4109), .B(RESET), .Z(WX4549) ) ;
DFF     gate1467  (.D(WX4549), .CP(CLK), .Q(WX4550) ) ;
AND2    gate1468  (.A(WX4123), .B(RESET), .Z(WX4551) ) ;
DFF     gate1469  (.D(WX4551), .CP(CLK), .Q(WX4552) ) ;
AND2    gate1470  (.A(WX4137), .B(RESET), .Z(WX4553) ) ;
DFF     gate1471  (.D(WX4553), .CP(CLK), .Q(WX4554) ) ;
AND2    gate1472  (.A(WX4151), .B(RESET), .Z(WX4555) ) ;
DFF     gate1473  (.D(WX4555), .CP(CLK), .Q(WX4556) ) ;
AND2    gate1474  (.A(WX4165), .B(RESET), .Z(WX4557) ) ;
DFF     gate1475  (.D(WX4557), .CP(CLK), .Q(WX4558) ) ;
AND2    gate1476  (.A(WX4179), .B(RESET), .Z(WX4559) ) ;
DFF     gate1477  (.D(WX4559), .CP(CLK), .Q(WX4560) ) ;
AND2    gate1478  (.A(WX4193), .B(RESET), .Z(WX4561) ) ;
DFF     gate1479  (.D(WX4561), .CP(CLK), .Q(WX4562) ) ;
AND2    gate1480  (.A(WX4207), .B(RESET), .Z(WX4563) ) ;
DFF     gate1481  (.D(WX4563), .CP(CLK), .Q(WX4564) ) ;
AND2    gate1482  (.A(WX4221), .B(RESET), .Z(WX4565) ) ;
DFF     gate1483  (.D(WX4565), .CP(CLK), .Q(WX4566) ) ;
AND2    gate1484  (.A(WX4235), .B(RESET), .Z(WX4567) ) ;
DFF     gate1485  (.D(WX4567), .CP(CLK), .Q(WX4568) ) ;
AND2    gate1486  (.A(WX4249), .B(RESET), .Z(WX4569) ) ;
DFF     gate1487  (.D(WX4569), .CP(CLK), .Q(WX4570) ) ;
AND2    gate1488  (.A(WX4263), .B(RESET), .Z(WX4571) ) ;
DFF     gate1489  (.D(WX4571), .CP(CLK), .Q(WX4572) ) ;
AND2    gate1490  (.A(WX4277), .B(RESET), .Z(WX4573) ) ;
DFF     gate1491  (.D(WX4573), .CP(CLK), .Q(WX4574) ) ;
AND2    gate1492  (.A(WX4291), .B(RESET), .Z(WX4575) ) ;
DFF     gate1493  (.D(WX4575), .CP(CLK), .Q(WX4576) ) ;
AND2    gate1494  (.A(WX4305), .B(RESET), .Z(WX4577) ) ;
DFF     gate1495  (.D(WX4577), .CP(CLK), .Q(WX4578) ) ;
AND2    gate1496  (.A(WX4319), .B(RESET), .Z(WX4579) ) ;
DFF     gate1497  (.D(WX4579), .CP(CLK), .Q(WX4580) ) ;
AND2    gate1498  (.A(WX4333), .B(RESET), .Z(WX4581) ) ;
DFF     gate1499  (.D(WX4581), .CP(CLK), .Q(WX4582) ) ;
AND2    gate1500  (.A(WX4347), .B(RESET), .Z(WX4583) ) ;
DFF     gate1501  (.D(WX4583), .CP(CLK), .Q(WX4584) ) ;
AND2    gate1502  (.A(WX4361), .B(RESET), .Z(WX4585) ) ;
DFF     gate1503  (.D(WX4585), .CP(CLK), .Q(WX4586) ) ;
AND2    gate1504  (.A(WX4524), .B(RESET), .Z(WX4587) ) ;
DFF     gate1505  (.D(WX4587), .CP(CLK), .Q(WX4588) ) ;
AND2    gate1506  (.A(WX4526), .B(RESET), .Z(WX4589) ) ;
DFF     gate1507  (.D(WX4589), .CP(CLK), .Q(WX4590) ) ;
AND2    gate1508  (.A(WX4528), .B(RESET), .Z(WX4591) ) ;
DFF     gate1509  (.D(WX4591), .CP(CLK), .Q(WX4592) ) ;
AND2    gate1510  (.A(WX4530), .B(RESET), .Z(WX4593) ) ;
DFF     gate1511  (.D(WX4593), .CP(CLK), .Q(WX4594) ) ;
AND2    gate1512  (.A(WX4532), .B(RESET), .Z(WX4595) ) ;
DFF     gate1513  (.D(WX4595), .CP(CLK), .Q(WX4596) ) ;
AND2    gate1514  (.A(WX4534), .B(RESET), .Z(WX4597) ) ;
DFF     gate1515  (.D(WX4597), .CP(CLK), .Q(WX4598) ) ;
AND2    gate1516  (.A(WX4536), .B(RESET), .Z(WX4599) ) ;
DFF     gate1517  (.D(WX4599), .CP(CLK), .Q(WX4600) ) ;
AND2    gate1518  (.A(WX4538), .B(RESET), .Z(WX4601) ) ;
DFF     gate1519  (.D(WX4601), .CP(CLK), .Q(WX4602) ) ;
AND2    gate1520  (.A(WX4540), .B(RESET), .Z(WX4603) ) ;
DFF     gate1521  (.D(WX4603), .CP(CLK), .Q(WX4604) ) ;
AND2    gate1522  (.A(WX4542), .B(RESET), .Z(WX4605) ) ;
DFF     gate1523  (.D(WX4605), .CP(CLK), .Q(WX4606) ) ;
AND2    gate1524  (.A(WX4544), .B(RESET), .Z(WX4607) ) ;
DFF     gate1525  (.D(WX4607), .CP(CLK), .Q(WX4608) ) ;
AND2    gate1526  (.A(WX4546), .B(RESET), .Z(WX4609) ) ;
DFF     gate1527  (.D(WX4609), .CP(CLK), .Q(WX4610) ) ;
AND2    gate1528  (.A(WX4548), .B(RESET), .Z(WX4611) ) ;
DFF     gate1529  (.D(WX4611), .CP(CLK), .Q(WX4612) ) ;
AND2    gate1530  (.A(WX4550), .B(RESET), .Z(WX4613) ) ;
DFF     gate1531  (.D(WX4613), .CP(CLK), .Q(WX4614) ) ;
AND2    gate1532  (.A(WX4552), .B(RESET), .Z(WX4615) ) ;
DFF     gate1533  (.D(WX4615), .CP(CLK), .Q(WX4616) ) ;
AND2    gate1534  (.A(WX4554), .B(RESET), .Z(WX4617) ) ;
DFF     gate1535  (.D(WX4617), .CP(CLK), .Q(WX4618) ) ;
AND2    gate1536  (.A(WX4556), .B(RESET), .Z(WX4619) ) ;
DFF     gate1537  (.D(WX4619), .CP(CLK), .Q(WX4620) ) ;
AND2    gate1538  (.A(WX4558), .B(RESET), .Z(WX4621) ) ;
DFF     gate1539  (.D(WX4621), .CP(CLK), .Q(WX4622) ) ;
AND2    gate1540  (.A(WX4560), .B(RESET), .Z(WX4623) ) ;
DFF     gate1541  (.D(WX4623), .CP(CLK), .Q(WX4624) ) ;
AND2    gate1542  (.A(WX4562), .B(RESET), .Z(WX4625) ) ;
DFF     gate1543  (.D(WX4625), .CP(CLK), .Q(WX4626) ) ;
AND2    gate1544  (.A(WX4564), .B(RESET), .Z(WX4627) ) ;
DFF     gate1545  (.D(WX4627), .CP(CLK), .Q(WX4628) ) ;
AND2    gate1546  (.A(WX4566), .B(RESET), .Z(WX4629) ) ;
DFF     gate1547  (.D(WX4629), .CP(CLK), .Q(WX4630) ) ;
AND2    gate1548  (.A(WX4568), .B(RESET), .Z(WX4631) ) ;
DFF     gate1549  (.D(WX4631), .CP(CLK), .Q(WX4632) ) ;
AND2    gate1550  (.A(WX4570), .B(RESET), .Z(WX4633) ) ;
DFF     gate1551  (.D(WX4633), .CP(CLK), .Q(WX4634) ) ;
AND2    gate1552  (.A(WX4572), .B(RESET), .Z(WX4635) ) ;
DFF     gate1553  (.D(WX4635), .CP(CLK), .Q(WX4636) ) ;
AND2    gate1554  (.A(WX4574), .B(RESET), .Z(WX4637) ) ;
DFF     gate1555  (.D(WX4637), .CP(CLK), .Q(WX4638) ) ;
AND2    gate1556  (.A(WX4576), .B(RESET), .Z(WX4639) ) ;
DFF     gate1557  (.D(WX4639), .CP(CLK), .Q(WX4640) ) ;
AND2    gate1558  (.A(WX4578), .B(RESET), .Z(WX4641) ) ;
DFF     gate1559  (.D(WX4641), .CP(CLK), .Q(WX4642) ) ;
AND2    gate1560  (.A(WX4580), .B(RESET), .Z(WX4643) ) ;
DFF     gate1561  (.D(WX4643), .CP(CLK), .Q(WX4644) ) ;
AND2    gate1562  (.A(WX4582), .B(RESET), .Z(WX4645) ) ;
DFF     gate1563  (.D(WX4645), .CP(CLK), .Q(WX4646) ) ;
AND2    gate1564  (.A(WX4584), .B(RESET), .Z(WX4647) ) ;
DFF     gate1565  (.D(WX4647), .CP(CLK), .Q(WX4648) ) ;
AND2    gate1566  (.A(WX4586), .B(RESET), .Z(WX4649) ) ;
DFF     gate1567  (.D(WX4649), .CP(CLK), .Q(WX4650) ) ;
AND2    gate1568  (.A(WX4588), .B(RESET), .Z(WX4651) ) ;
DFF     gate1569  (.D(WX4651), .CP(CLK), .Q(WX4652) ) ;
AND2    gate1570  (.A(WX4590), .B(RESET), .Z(WX4653) ) ;
DFF     gate1571  (.D(WX4653), .CP(CLK), .Q(WX4654) ) ;
AND2    gate1572  (.A(WX4592), .B(RESET), .Z(WX4655) ) ;
DFF     gate1573  (.D(WX4655), .CP(CLK), .Q(WX4656) ) ;
AND2    gate1574  (.A(WX4594), .B(RESET), .Z(WX4657) ) ;
DFF     gate1575  (.D(WX4657), .CP(CLK), .Q(WX4658) ) ;
AND2    gate1576  (.A(WX4596), .B(RESET), .Z(WX4659) ) ;
DFF     gate1577  (.D(WX4659), .CP(CLK), .Q(WX4660) ) ;
AND2    gate1578  (.A(WX4598), .B(RESET), .Z(WX4661) ) ;
DFF     gate1579  (.D(WX4661), .CP(CLK), .Q(WX4662) ) ;
AND2    gate1580  (.A(WX4600), .B(RESET), .Z(WX4663) ) ;
DFF     gate1581  (.D(WX4663), .CP(CLK), .Q(WX4664) ) ;
AND2    gate1582  (.A(WX4602), .B(RESET), .Z(WX4665) ) ;
DFF     gate1583  (.D(WX4665), .CP(CLK), .Q(WX4666) ) ;
AND2    gate1584  (.A(WX4604), .B(RESET), .Z(WX4667) ) ;
DFF     gate1585  (.D(WX4667), .CP(CLK), .Q(WX4668) ) ;
AND2    gate1586  (.A(WX4606), .B(RESET), .Z(WX4669) ) ;
DFF     gate1587  (.D(WX4669), .CP(CLK), .Q(WX4670) ) ;
AND2    gate1588  (.A(WX4608), .B(RESET), .Z(WX4671) ) ;
DFF     gate1589  (.D(WX4671), .CP(CLK), .Q(WX4672) ) ;
AND2    gate1590  (.A(WX4610), .B(RESET), .Z(WX4673) ) ;
DFF     gate1591  (.D(WX4673), .CP(CLK), .Q(WX4674) ) ;
AND2    gate1592  (.A(WX4612), .B(RESET), .Z(WX4675) ) ;
DFF     gate1593  (.D(WX4675), .CP(CLK), .Q(WX4676) ) ;
AND2    gate1594  (.A(WX4614), .B(RESET), .Z(WX4677) ) ;
DFF     gate1595  (.D(WX4677), .CP(CLK), .Q(WX4678) ) ;
AND2    gate1596  (.A(WX4616), .B(RESET), .Z(WX4679) ) ;
DFF     gate1597  (.D(WX4679), .CP(CLK), .Q(WX4680) ) ;
AND2    gate1598  (.A(WX4618), .B(RESET), .Z(WX4681) ) ;
DFF     gate1599  (.D(WX4681), .CP(CLK), .Q(WX4682) ) ;
AND2    gate1600  (.A(WX4620), .B(RESET), .Z(WX4683) ) ;
DFF     gate1601  (.D(WX4683), .CP(CLK), .Q(WX4684) ) ;
AND2    gate1602  (.A(WX4622), .B(RESET), .Z(WX4685) ) ;
DFF     gate1603  (.D(WX4685), .CP(CLK), .Q(WX4686) ) ;
AND2    gate1604  (.A(WX4624), .B(RESET), .Z(WX4687) ) ;
DFF     gate1605  (.D(WX4687), .CP(CLK), .Q(WX4688) ) ;
AND2    gate1606  (.A(WX4626), .B(RESET), .Z(WX4689) ) ;
DFF     gate1607  (.D(WX4689), .CP(CLK), .Q(WX4690) ) ;
AND2    gate1608  (.A(WX4628), .B(RESET), .Z(WX4691) ) ;
DFF     gate1609  (.D(WX4691), .CP(CLK), .Q(WX4692) ) ;
AND2    gate1610  (.A(WX4630), .B(RESET), .Z(WX4693) ) ;
DFF     gate1611  (.D(WX4693), .CP(CLK), .Q(WX4694) ) ;
AND2    gate1612  (.A(WX4632), .B(RESET), .Z(WX4695) ) ;
DFF     gate1613  (.D(WX4695), .CP(CLK), .Q(WX4696) ) ;
AND2    gate1614  (.A(WX4634), .B(RESET), .Z(WX4697) ) ;
DFF     gate1615  (.D(WX4697), .CP(CLK), .Q(WX4698) ) ;
AND2    gate1616  (.A(WX4636), .B(RESET), .Z(WX4699) ) ;
DFF     gate1617  (.D(WX4699), .CP(CLK), .Q(WX4700) ) ;
AND2    gate1618  (.A(WX4638), .B(RESET), .Z(WX4701) ) ;
DFF     gate1619  (.D(WX4701), .CP(CLK), .Q(WX4702) ) ;
AND2    gate1620  (.A(WX4640), .B(RESET), .Z(WX4703) ) ;
DFF     gate1621  (.D(WX4703), .CP(CLK), .Q(WX4704) ) ;
AND2    gate1622  (.A(WX4642), .B(RESET), .Z(WX4705) ) ;
DFF     gate1623  (.D(WX4705), .CP(CLK), .Q(WX4706) ) ;
AND2    gate1624  (.A(WX4644), .B(RESET), .Z(WX4707) ) ;
DFF     gate1625  (.D(WX4707), .CP(CLK), .Q(WX4708) ) ;
AND2    gate1626  (.A(WX4646), .B(RESET), .Z(WX4709) ) ;
DFF     gate1627  (.D(WX4709), .CP(CLK), .Q(WX4710) ) ;
AND2    gate1628  (.A(WX4648), .B(RESET), .Z(WX4711) ) ;
DFF     gate1629  (.D(WX4711), .CP(CLK), .Q(WX4712) ) ;
AND2    gate1630  (.A(WX4650), .B(RESET), .Z(WX4713) ) ;
DFF     gate1631  (.D(WX4713), .CP(CLK), .Q(WX4714) ) ;
AND2    gate1632  (.A(WX4652), .B(RESET), .Z(WX4715) ) ;
DFF     gate1633  (.D(WX4715), .CP(CLK), .Q(WX4716) ) ;
AND2    gate1634  (.A(WX4654), .B(RESET), .Z(WX4717) ) ;
DFF     gate1635  (.D(WX4717), .CP(CLK), .Q(WX4718) ) ;
AND2    gate1636  (.A(WX4656), .B(RESET), .Z(WX4719) ) ;
DFF     gate1637  (.D(WX4719), .CP(CLK), .Q(WX4720) ) ;
AND2    gate1638  (.A(WX4658), .B(RESET), .Z(WX4721) ) ;
DFF     gate1639  (.D(WX4721), .CP(CLK), .Q(WX4722) ) ;
AND2    gate1640  (.A(WX4660), .B(RESET), .Z(WX4723) ) ;
DFF     gate1641  (.D(WX4723), .CP(CLK), .Q(WX4724) ) ;
AND2    gate1642  (.A(WX4662), .B(RESET), .Z(WX4725) ) ;
DFF     gate1643  (.D(WX4725), .CP(CLK), .Q(WX4726) ) ;
AND2    gate1644  (.A(WX4664), .B(RESET), .Z(WX4727) ) ;
DFF     gate1645  (.D(WX4727), .CP(CLK), .Q(WX4728) ) ;
AND2    gate1646  (.A(WX4666), .B(RESET), .Z(WX4729) ) ;
DFF     gate1647  (.D(WX4729), .CP(CLK), .Q(WX4730) ) ;
AND2    gate1648  (.A(WX4668), .B(RESET), .Z(WX4731) ) ;
DFF     gate1649  (.D(WX4731), .CP(CLK), .Q(WX4732) ) ;
AND2    gate1650  (.A(WX4670), .B(RESET), .Z(WX4733) ) ;
DFF     gate1651  (.D(WX4733), .CP(CLK), .Q(WX4734) ) ;
AND2    gate1652  (.A(WX4672), .B(RESET), .Z(WX4735) ) ;
DFF     gate1653  (.D(WX4735), .CP(CLK), .Q(WX4736) ) ;
AND2    gate1654  (.A(WX4674), .B(RESET), .Z(WX4737) ) ;
DFF     gate1655  (.D(WX4737), .CP(CLK), .Q(WX4738) ) ;
AND2    gate1656  (.A(WX4676), .B(RESET), .Z(WX4739) ) ;
DFF     gate1657  (.D(WX4739), .CP(CLK), .Q(WX4740) ) ;
AND2    gate1658  (.A(WX4678), .B(RESET), .Z(WX4741) ) ;
DFF     gate1659  (.D(WX4741), .CP(CLK), .Q(WX4742) ) ;
AND2    gate1660  (.A(WX4680), .B(RESET), .Z(WX4743) ) ;
DFF     gate1661  (.D(WX4743), .CP(CLK), .Q(WX4744) ) ;
AND2    gate1662  (.A(WX4682), .B(RESET), .Z(WX4745) ) ;
DFF     gate1663  (.D(WX4745), .CP(CLK), .Q(WX4746) ) ;
AND2    gate1664  (.A(WX4684), .B(RESET), .Z(WX4747) ) ;
DFF     gate1665  (.D(WX4747), .CP(CLK), .Q(WX4748) ) ;
AND2    gate1666  (.A(WX4686), .B(RESET), .Z(WX4749) ) ;
DFF     gate1667  (.D(WX4749), .CP(CLK), .Q(WX4750) ) ;
AND2    gate1668  (.A(WX4688), .B(RESET), .Z(WX4751) ) ;
DFF     gate1669  (.D(WX4751), .CP(CLK), .Q(WX4752) ) ;
AND2    gate1670  (.A(WX4690), .B(RESET), .Z(WX4753) ) ;
DFF     gate1671  (.D(WX4753), .CP(CLK), .Q(WX4754) ) ;
AND2    gate1672  (.A(WX4692), .B(RESET), .Z(WX4755) ) ;
DFF     gate1673  (.D(WX4755), .CP(CLK), .Q(WX4756) ) ;
AND2    gate1674  (.A(WX4694), .B(RESET), .Z(WX4757) ) ;
DFF     gate1675  (.D(WX4757), .CP(CLK), .Q(WX4758) ) ;
AND2    gate1676  (.A(WX4696), .B(RESET), .Z(WX4759) ) ;
DFF     gate1677  (.D(WX4759), .CP(CLK), .Q(WX4760) ) ;
AND2    gate1678  (.A(WX4698), .B(RESET), .Z(WX4761) ) ;
DFF     gate1679  (.D(WX4761), .CP(CLK), .Q(WX4762) ) ;
AND2    gate1680  (.A(WX4700), .B(RESET), .Z(WX4763) ) ;
DFF     gate1681  (.D(WX4763), .CP(CLK), .Q(WX4764) ) ;
AND2    gate1682  (.A(WX4702), .B(RESET), .Z(WX4765) ) ;
DFF     gate1683  (.D(WX4765), .CP(CLK), .Q(WX4766) ) ;
AND2    gate1684  (.A(WX4704), .B(RESET), .Z(WX4767) ) ;
DFF     gate1685  (.D(WX4767), .CP(CLK), .Q(WX4768) ) ;
AND2    gate1686  (.A(WX4706), .B(RESET), .Z(WX4769) ) ;
DFF     gate1687  (.D(WX4769), .CP(CLK), .Q(WX4770) ) ;
AND2    gate1688  (.A(WX4708), .B(RESET), .Z(WX4771) ) ;
DFF     gate1689  (.D(WX4771), .CP(CLK), .Q(WX4772) ) ;
AND2    gate1690  (.A(WX4710), .B(RESET), .Z(WX4773) ) ;
DFF     gate1691  (.D(WX4773), .CP(CLK), .Q(WX4774) ) ;
AND2    gate1692  (.A(WX4712), .B(RESET), .Z(WX4775) ) ;
DFF     gate1693  (.D(WX4775), .CP(CLK), .Q(WX4776) ) ;
AND2    gate1694  (.A(WX4714), .B(RESET), .Z(WX4777) ) ;
DFF     gate1695  (.D(WX4777), .CP(CLK), .Q(WX4778) ) ;
AND2    gate1696  (.A(WX5113), .B(WX5142), .Z(WX5143) ) ;
AND2    gate1697  (.A(WX5141), .B(WX5142), .Z(WX5145) ) ;
AND2    gate1698  (.A(WX5140), .B(WX5142), .Z(WX5147) ) ;
AND2    gate1699  (.A(WX5139), .B(WX5142), .Z(WX5149) ) ;
AND2    gate1700  (.A(WX5112), .B(WX5142), .Z(WX5151) ) ;
AND2    gate1701  (.A(WX5138), .B(WX5142), .Z(WX5153) ) ;
AND2    gate1702  (.A(WX5137), .B(WX5142), .Z(WX5155) ) ;
AND2    gate1703  (.A(WX5136), .B(WX5142), .Z(WX5157) ) ;
AND2    gate1704  (.A(WX5135), .B(WX5142), .Z(WX5159) ) ;
AND2    gate1705  (.A(WX5134), .B(WX5142), .Z(WX5161) ) ;
AND2    gate1706  (.A(WX5133), .B(WX5142), .Z(WX5163) ) ;
AND2    gate1707  (.A(WX5111), .B(WX5142), .Z(WX5165) ) ;
AND2    gate1708  (.A(WX5132), .B(WX5142), .Z(WX5167) ) ;
AND2    gate1709  (.A(WX5131), .B(WX5142), .Z(WX5169) ) ;
AND2    gate1710  (.A(WX5130), .B(WX5142), .Z(WX5171) ) ;
AND2    gate1711  (.A(WX5129), .B(WX5142), .Z(WX5173) ) ;
AND2    gate1712  (.A(WX5110), .B(WX5142), .Z(WX5175) ) ;
AND2    gate1713  (.A(WX5128), .B(WX5142), .Z(WX5177) ) ;
AND2    gate1714  (.A(WX5127), .B(WX5142), .Z(WX5179) ) ;
AND2    gate1715  (.A(WX5126), .B(WX5142), .Z(WX5181) ) ;
AND2    gate1716  (.A(WX5125), .B(WX5142), .Z(WX5183) ) ;
AND2    gate1717  (.A(WX5124), .B(WX5142), .Z(WX5185) ) ;
AND2    gate1718  (.A(WX5123), .B(WX5142), .Z(WX5187) ) ;
AND2    gate1719  (.A(WX5122), .B(WX5142), .Z(WX5189) ) ;
AND2    gate1720  (.A(WX5121), .B(WX5142), .Z(WX5191) ) ;
AND2    gate1721  (.A(WX5120), .B(WX5142), .Z(WX5193) ) ;
AND2    gate1722  (.A(WX5119), .B(WX5142), .Z(WX5195) ) ;
AND2    gate1723  (.A(WX5118), .B(WX5142), .Z(WX5197) ) ;
AND2    gate1724  (.A(WX5117), .B(WX5142), .Z(WX5199) ) ;
AND2    gate1725  (.A(WX5116), .B(WX5142), .Z(WX5201) ) ;
AND2    gate1726  (.A(WX5115), .B(WX5142), .Z(WX5203) ) ;
AND2    gate1727  (.A(WX5114), .B(WX5142), .Z(WX5205) ) ;
AND2    gate1728  (.A(WX5659), .B(RESET), .Z(WX5656) ) ;
DFF     gate1729  (.D(WX5656), .CP(CLK), .Q(WX5657) ) ;
AND2    gate1730  (.A(WX5661), .B(RESET), .Z(WX5658) ) ;
DFF     gate1731  (.D(WX5658), .CP(CLK), .Q(WX5659) ) ;
AND2    gate1732  (.A(WX5663), .B(RESET), .Z(WX5660) ) ;
DFF     gate1733  (.D(WX5660), .CP(CLK), .Q(WX5661) ) ;
AND2    gate1734  (.A(WX5665), .B(RESET), .Z(WX5662) ) ;
DFF     gate1735  (.D(WX5662), .CP(CLK), .Q(WX5663) ) ;
AND2    gate1736  (.A(WX5667), .B(RESET), .Z(WX5664) ) ;
DFF     gate1737  (.D(WX5664), .CP(CLK), .Q(WX5665) ) ;
AND2    gate1738  (.A(WX5669), .B(RESET), .Z(WX5666) ) ;
DFF     gate1739  (.D(WX5666), .CP(CLK), .Q(WX5667) ) ;
AND2    gate1740  (.A(WX5671), .B(RESET), .Z(WX5668) ) ;
DFF     gate1741  (.D(WX5668), .CP(CLK), .Q(WX5669) ) ;
AND2    gate1742  (.A(WX5673), .B(RESET), .Z(WX5670) ) ;
DFF     gate1743  (.D(WX5670), .CP(CLK), .Q(WX5671) ) ;
AND2    gate1744  (.A(WX5675), .B(RESET), .Z(WX5672) ) ;
DFF     gate1745  (.D(WX5672), .CP(CLK), .Q(WX5673) ) ;
AND2    gate1746  (.A(WX5677), .B(RESET), .Z(WX5674) ) ;
DFF     gate1747  (.D(WX5674), .CP(CLK), .Q(WX5675) ) ;
AND2    gate1748  (.A(WX5679), .B(RESET), .Z(WX5676) ) ;
DFF     gate1749  (.D(WX5676), .CP(CLK), .Q(WX5677) ) ;
AND2    gate1750  (.A(WX5681), .B(RESET), .Z(WX5678) ) ;
DFF     gate1751  (.D(WX5678), .CP(CLK), .Q(WX5679) ) ;
AND2    gate1752  (.A(WX5683), .B(RESET), .Z(WX5680) ) ;
DFF     gate1753  (.D(WX5680), .CP(CLK), .Q(WX5681) ) ;
AND2    gate1754  (.A(WX5685), .B(RESET), .Z(WX5682) ) ;
DFF     gate1755  (.D(WX5682), .CP(CLK), .Q(WX5683) ) ;
AND2    gate1756  (.A(WX5687), .B(RESET), .Z(WX5684) ) ;
DFF     gate1757  (.D(WX5684), .CP(CLK), .Q(WX5685) ) ;
AND2    gate1758  (.A(WX5689), .B(RESET), .Z(WX5686) ) ;
DFF     gate1759  (.D(WX5686), .CP(CLK), .Q(WX5687) ) ;
AND2    gate1760  (.A(WX5691), .B(RESET), .Z(WX5688) ) ;
DFF     gate1761  (.D(WX5688), .CP(CLK), .Q(WX5689) ) ;
AND2    gate1762  (.A(WX5693), .B(RESET), .Z(WX5690) ) ;
DFF     gate1763  (.D(WX5690), .CP(CLK), .Q(WX5691) ) ;
AND2    gate1764  (.A(WX5695), .B(RESET), .Z(WX5692) ) ;
DFF     gate1765  (.D(WX5692), .CP(CLK), .Q(WX5693) ) ;
AND2    gate1766  (.A(WX5697), .B(RESET), .Z(WX5694) ) ;
DFF     gate1767  (.D(WX5694), .CP(CLK), .Q(WX5695) ) ;
AND2    gate1768  (.A(WX5699), .B(RESET), .Z(WX5696) ) ;
DFF     gate1769  (.D(WX5696), .CP(CLK), .Q(WX5697) ) ;
AND2    gate1770  (.A(WX5701), .B(RESET), .Z(WX5698) ) ;
DFF     gate1771  (.D(WX5698), .CP(CLK), .Q(WX5699) ) ;
AND2    gate1772  (.A(WX5703), .B(RESET), .Z(WX5700) ) ;
DFF     gate1773  (.D(WX5700), .CP(CLK), .Q(WX5701) ) ;
AND2    gate1774  (.A(WX5705), .B(RESET), .Z(WX5702) ) ;
DFF     gate1775  (.D(WX5702), .CP(CLK), .Q(WX5703) ) ;
AND2    gate1776  (.A(WX5707), .B(RESET), .Z(WX5704) ) ;
DFF     gate1777  (.D(WX5704), .CP(CLK), .Q(WX5705) ) ;
AND2    gate1778  (.A(WX5709), .B(RESET), .Z(WX5706) ) ;
DFF     gate1779  (.D(WX5706), .CP(CLK), .Q(WX5707) ) ;
AND2    gate1780  (.A(WX5711), .B(RESET), .Z(WX5708) ) ;
DFF     gate1781  (.D(WX5708), .CP(CLK), .Q(WX5709) ) ;
AND2    gate1782  (.A(WX5713), .B(RESET), .Z(WX5710) ) ;
DFF     gate1783  (.D(WX5710), .CP(CLK), .Q(WX5711) ) ;
AND2    gate1784  (.A(WX5715), .B(RESET), .Z(WX5712) ) ;
DFF     gate1785  (.D(WX5712), .CP(CLK), .Q(WX5713) ) ;
AND2    gate1786  (.A(WX5717), .B(RESET), .Z(WX5714) ) ;
DFF     gate1787  (.D(WX5714), .CP(CLK), .Q(WX5715) ) ;
AND2    gate1788  (.A(WX5719), .B(RESET), .Z(WX5716) ) ;
DFF     gate1789  (.D(WX5716), .CP(CLK), .Q(WX5717) ) ;
AND2    gate1790  (.A(WX5655), .B(RESET), .Z(WX5718) ) ;
DFF     gate1791  (.D(WX5718), .CP(CLK), .Q(WX5719) ) ;
AND2    gate1792  (.A(WX5220), .B(RESET), .Z(WX5816) ) ;
DFF     gate1793  (.D(WX5816), .CP(CLK), .Q(WX5817) ) ;
AND2    gate1794  (.A(WX5234), .B(RESET), .Z(WX5818) ) ;
DFF     gate1795  (.D(WX5818), .CP(CLK), .Q(WX5819) ) ;
AND2    gate1796  (.A(WX5248), .B(RESET), .Z(WX5820) ) ;
DFF     gate1797  (.D(WX5820), .CP(CLK), .Q(WX5821) ) ;
AND2    gate1798  (.A(WX5262), .B(RESET), .Z(WX5822) ) ;
DFF     gate1799  (.D(WX5822), .CP(CLK), .Q(WX5823) ) ;
AND2    gate1800  (.A(WX5276), .B(RESET), .Z(WX5824) ) ;
DFF     gate1801  (.D(WX5824), .CP(CLK), .Q(WX5825) ) ;
AND2    gate1802  (.A(WX5290), .B(RESET), .Z(WX5826) ) ;
DFF     gate1803  (.D(WX5826), .CP(CLK), .Q(WX5827) ) ;
AND2    gate1804  (.A(WX5304), .B(RESET), .Z(WX5828) ) ;
DFF     gate1805  (.D(WX5828), .CP(CLK), .Q(WX5829) ) ;
AND2    gate1806  (.A(WX5318), .B(RESET), .Z(WX5830) ) ;
DFF     gate1807  (.D(WX5830), .CP(CLK), .Q(WX5831) ) ;
AND2    gate1808  (.A(WX5332), .B(RESET), .Z(WX5832) ) ;
DFF     gate1809  (.D(WX5832), .CP(CLK), .Q(WX5833) ) ;
AND2    gate1810  (.A(WX5346), .B(RESET), .Z(WX5834) ) ;
DFF     gate1811  (.D(WX5834), .CP(CLK), .Q(WX5835) ) ;
AND2    gate1812  (.A(WX5360), .B(RESET), .Z(WX5836) ) ;
DFF     gate1813  (.D(WX5836), .CP(CLK), .Q(WX5837) ) ;
AND2    gate1814  (.A(WX5374), .B(RESET), .Z(WX5838) ) ;
DFF     gate1815  (.D(WX5838), .CP(CLK), .Q(WX5839) ) ;
AND2    gate1816  (.A(WX5388), .B(RESET), .Z(WX5840) ) ;
DFF     gate1817  (.D(WX5840), .CP(CLK), .Q(WX5841) ) ;
AND2    gate1818  (.A(WX5402), .B(RESET), .Z(WX5842) ) ;
DFF     gate1819  (.D(WX5842), .CP(CLK), .Q(WX5843) ) ;
AND2    gate1820  (.A(WX5416), .B(RESET), .Z(WX5844) ) ;
DFF     gate1821  (.D(WX5844), .CP(CLK), .Q(WX5845) ) ;
AND2    gate1822  (.A(WX5430), .B(RESET), .Z(WX5846) ) ;
DFF     gate1823  (.D(WX5846), .CP(CLK), .Q(WX5847) ) ;
AND2    gate1824  (.A(WX5444), .B(RESET), .Z(WX5848) ) ;
DFF     gate1825  (.D(WX5848), .CP(CLK), .Q(WX5849) ) ;
AND2    gate1826  (.A(WX5458), .B(RESET), .Z(WX5850) ) ;
DFF     gate1827  (.D(WX5850), .CP(CLK), .Q(WX5851) ) ;
AND2    gate1828  (.A(WX5472), .B(RESET), .Z(WX5852) ) ;
DFF     gate1829  (.D(WX5852), .CP(CLK), .Q(WX5853) ) ;
AND2    gate1830  (.A(WX5486), .B(RESET), .Z(WX5854) ) ;
DFF     gate1831  (.D(WX5854), .CP(CLK), .Q(WX5855) ) ;
AND2    gate1832  (.A(WX5500), .B(RESET), .Z(WX5856) ) ;
DFF     gate1833  (.D(WX5856), .CP(CLK), .Q(WX5857) ) ;
AND2    gate1834  (.A(WX5514), .B(RESET), .Z(WX5858) ) ;
DFF     gate1835  (.D(WX5858), .CP(CLK), .Q(WX5859) ) ;
AND2    gate1836  (.A(WX5528), .B(RESET), .Z(WX5860) ) ;
DFF     gate1837  (.D(WX5860), .CP(CLK), .Q(WX5861) ) ;
AND2    gate1838  (.A(WX5542), .B(RESET), .Z(WX5862) ) ;
DFF     gate1839  (.D(WX5862), .CP(CLK), .Q(WX5863) ) ;
AND2    gate1840  (.A(WX5556), .B(RESET), .Z(WX5864) ) ;
DFF     gate1841  (.D(WX5864), .CP(CLK), .Q(WX5865) ) ;
AND2    gate1842  (.A(WX5570), .B(RESET), .Z(WX5866) ) ;
DFF     gate1843  (.D(WX5866), .CP(CLK), .Q(WX5867) ) ;
AND2    gate1844  (.A(WX5584), .B(RESET), .Z(WX5868) ) ;
DFF     gate1845  (.D(WX5868), .CP(CLK), .Q(WX5869) ) ;
AND2    gate1846  (.A(WX5598), .B(RESET), .Z(WX5870) ) ;
DFF     gate1847  (.D(WX5870), .CP(CLK), .Q(WX5871) ) ;
AND2    gate1848  (.A(WX5612), .B(RESET), .Z(WX5872) ) ;
DFF     gate1849  (.D(WX5872), .CP(CLK), .Q(WX5873) ) ;
AND2    gate1850  (.A(WX5626), .B(RESET), .Z(WX5874) ) ;
DFF     gate1851  (.D(WX5874), .CP(CLK), .Q(WX5875) ) ;
AND2    gate1852  (.A(WX5640), .B(RESET), .Z(WX5876) ) ;
DFF     gate1853  (.D(WX5876), .CP(CLK), .Q(WX5877) ) ;
AND2    gate1854  (.A(WX5654), .B(RESET), .Z(WX5878) ) ;
DFF     gate1855  (.D(WX5878), .CP(CLK), .Q(WX5879) ) ;
AND2    gate1856  (.A(WX5817), .B(RESET), .Z(WX5880) ) ;
DFF     gate1857  (.D(WX5880), .CP(CLK), .Q(WX5881) ) ;
AND2    gate1858  (.A(WX5819), .B(RESET), .Z(WX5882) ) ;
DFF     gate1859  (.D(WX5882), .CP(CLK), .Q(WX5883) ) ;
AND2    gate1860  (.A(WX5821), .B(RESET), .Z(WX5884) ) ;
DFF     gate1861  (.D(WX5884), .CP(CLK), .Q(WX5885) ) ;
AND2    gate1862  (.A(WX5823), .B(RESET), .Z(WX5886) ) ;
DFF     gate1863  (.D(WX5886), .CP(CLK), .Q(WX5887) ) ;
AND2    gate1864  (.A(WX5825), .B(RESET), .Z(WX5888) ) ;
DFF     gate1865  (.D(WX5888), .CP(CLK), .Q(WX5889) ) ;
AND2    gate1866  (.A(WX5827), .B(RESET), .Z(WX5890) ) ;
DFF     gate1867  (.D(WX5890), .CP(CLK), .Q(WX5891) ) ;
AND2    gate1868  (.A(WX5829), .B(RESET), .Z(WX5892) ) ;
DFF     gate1869  (.D(WX5892), .CP(CLK), .Q(WX5893) ) ;
AND2    gate1870  (.A(WX5831), .B(RESET), .Z(WX5894) ) ;
DFF     gate1871  (.D(WX5894), .CP(CLK), .Q(WX5895) ) ;
AND2    gate1872  (.A(WX5833), .B(RESET), .Z(WX5896) ) ;
DFF     gate1873  (.D(WX5896), .CP(CLK), .Q(WX5897) ) ;
AND2    gate1874  (.A(WX5835), .B(RESET), .Z(WX5898) ) ;
DFF     gate1875  (.D(WX5898), .CP(CLK), .Q(WX5899) ) ;
AND2    gate1876  (.A(WX5837), .B(RESET), .Z(WX5900) ) ;
DFF     gate1877  (.D(WX5900), .CP(CLK), .Q(WX5901) ) ;
AND2    gate1878  (.A(WX5839), .B(RESET), .Z(WX5902) ) ;
DFF     gate1879  (.D(WX5902), .CP(CLK), .Q(WX5903) ) ;
AND2    gate1880  (.A(WX5841), .B(RESET), .Z(WX5904) ) ;
DFF     gate1881  (.D(WX5904), .CP(CLK), .Q(WX5905) ) ;
AND2    gate1882  (.A(WX5843), .B(RESET), .Z(WX5906) ) ;
DFF     gate1883  (.D(WX5906), .CP(CLK), .Q(WX5907) ) ;
AND2    gate1884  (.A(WX5845), .B(RESET), .Z(WX5908) ) ;
DFF     gate1885  (.D(WX5908), .CP(CLK), .Q(WX5909) ) ;
AND2    gate1886  (.A(WX5847), .B(RESET), .Z(WX5910) ) ;
DFF     gate1887  (.D(WX5910), .CP(CLK), .Q(WX5911) ) ;
AND2    gate1888  (.A(WX5849), .B(RESET), .Z(WX5912) ) ;
DFF     gate1889  (.D(WX5912), .CP(CLK), .Q(WX5913) ) ;
AND2    gate1890  (.A(WX5851), .B(RESET), .Z(WX5914) ) ;
DFF     gate1891  (.D(WX5914), .CP(CLK), .Q(WX5915) ) ;
AND2    gate1892  (.A(WX5853), .B(RESET), .Z(WX5916) ) ;
DFF     gate1893  (.D(WX5916), .CP(CLK), .Q(WX5917) ) ;
AND2    gate1894  (.A(WX5855), .B(RESET), .Z(WX5918) ) ;
DFF     gate1895  (.D(WX5918), .CP(CLK), .Q(WX5919) ) ;
AND2    gate1896  (.A(WX5857), .B(RESET), .Z(WX5920) ) ;
DFF     gate1897  (.D(WX5920), .CP(CLK), .Q(WX5921) ) ;
AND2    gate1898  (.A(WX5859), .B(RESET), .Z(WX5922) ) ;
DFF     gate1899  (.D(WX5922), .CP(CLK), .Q(WX5923) ) ;
AND2    gate1900  (.A(WX5861), .B(RESET), .Z(WX5924) ) ;
DFF     gate1901  (.D(WX5924), .CP(CLK), .Q(WX5925) ) ;
AND2    gate1902  (.A(WX5863), .B(RESET), .Z(WX5926) ) ;
DFF     gate1903  (.D(WX5926), .CP(CLK), .Q(WX5927) ) ;
AND2    gate1904  (.A(WX5865), .B(RESET), .Z(WX5928) ) ;
DFF     gate1905  (.D(WX5928), .CP(CLK), .Q(WX5929) ) ;
AND2    gate1906  (.A(WX5867), .B(RESET), .Z(WX5930) ) ;
DFF     gate1907  (.D(WX5930), .CP(CLK), .Q(WX5931) ) ;
AND2    gate1908  (.A(WX5869), .B(RESET), .Z(WX5932) ) ;
DFF     gate1909  (.D(WX5932), .CP(CLK), .Q(WX5933) ) ;
AND2    gate1910  (.A(WX5871), .B(RESET), .Z(WX5934) ) ;
DFF     gate1911  (.D(WX5934), .CP(CLK), .Q(WX5935) ) ;
AND2    gate1912  (.A(WX5873), .B(RESET), .Z(WX5936) ) ;
DFF     gate1913  (.D(WX5936), .CP(CLK), .Q(WX5937) ) ;
AND2    gate1914  (.A(WX5875), .B(RESET), .Z(WX5938) ) ;
DFF     gate1915  (.D(WX5938), .CP(CLK), .Q(WX5939) ) ;
AND2    gate1916  (.A(WX5877), .B(RESET), .Z(WX5940) ) ;
DFF     gate1917  (.D(WX5940), .CP(CLK), .Q(WX5941) ) ;
AND2    gate1918  (.A(WX5879), .B(RESET), .Z(WX5942) ) ;
DFF     gate1919  (.D(WX5942), .CP(CLK), .Q(WX5943) ) ;
AND2    gate1920  (.A(WX5881), .B(RESET), .Z(WX5944) ) ;
DFF     gate1921  (.D(WX5944), .CP(CLK), .Q(WX5945) ) ;
AND2    gate1922  (.A(WX5883), .B(RESET), .Z(WX5946) ) ;
DFF     gate1923  (.D(WX5946), .CP(CLK), .Q(WX5947) ) ;
AND2    gate1924  (.A(WX5885), .B(RESET), .Z(WX5948) ) ;
DFF     gate1925  (.D(WX5948), .CP(CLK), .Q(WX5949) ) ;
AND2    gate1926  (.A(WX5887), .B(RESET), .Z(WX5950) ) ;
DFF     gate1927  (.D(WX5950), .CP(CLK), .Q(WX5951) ) ;
AND2    gate1928  (.A(WX5889), .B(RESET), .Z(WX5952) ) ;
DFF     gate1929  (.D(WX5952), .CP(CLK), .Q(WX5953) ) ;
AND2    gate1930  (.A(WX5891), .B(RESET), .Z(WX5954) ) ;
DFF     gate1931  (.D(WX5954), .CP(CLK), .Q(WX5955) ) ;
AND2    gate1932  (.A(WX5893), .B(RESET), .Z(WX5956) ) ;
DFF     gate1933  (.D(WX5956), .CP(CLK), .Q(WX5957) ) ;
AND2    gate1934  (.A(WX5895), .B(RESET), .Z(WX5958) ) ;
DFF     gate1935  (.D(WX5958), .CP(CLK), .Q(WX5959) ) ;
AND2    gate1936  (.A(WX5897), .B(RESET), .Z(WX5960) ) ;
DFF     gate1937  (.D(WX5960), .CP(CLK), .Q(WX5961) ) ;
AND2    gate1938  (.A(WX5899), .B(RESET), .Z(WX5962) ) ;
DFF     gate1939  (.D(WX5962), .CP(CLK), .Q(WX5963) ) ;
AND2    gate1940  (.A(WX5901), .B(RESET), .Z(WX5964) ) ;
DFF     gate1941  (.D(WX5964), .CP(CLK), .Q(WX5965) ) ;
AND2    gate1942  (.A(WX5903), .B(RESET), .Z(WX5966) ) ;
DFF     gate1943  (.D(WX5966), .CP(CLK), .Q(WX5967) ) ;
AND2    gate1944  (.A(WX5905), .B(RESET), .Z(WX5968) ) ;
DFF     gate1945  (.D(WX5968), .CP(CLK), .Q(WX5969) ) ;
AND2    gate1946  (.A(WX5907), .B(RESET), .Z(WX5970) ) ;
DFF     gate1947  (.D(WX5970), .CP(CLK), .Q(WX5971) ) ;
AND2    gate1948  (.A(WX5909), .B(RESET), .Z(WX5972) ) ;
DFF     gate1949  (.D(WX5972), .CP(CLK), .Q(WX5973) ) ;
AND2    gate1950  (.A(WX5911), .B(RESET), .Z(WX5974) ) ;
DFF     gate1951  (.D(WX5974), .CP(CLK), .Q(WX5975) ) ;
AND2    gate1952  (.A(WX5913), .B(RESET), .Z(WX5976) ) ;
DFF     gate1953  (.D(WX5976), .CP(CLK), .Q(WX5977) ) ;
AND2    gate1954  (.A(WX5915), .B(RESET), .Z(WX5978) ) ;
DFF     gate1955  (.D(WX5978), .CP(CLK), .Q(WX5979) ) ;
AND2    gate1956  (.A(WX5917), .B(RESET), .Z(WX5980) ) ;
DFF     gate1957  (.D(WX5980), .CP(CLK), .Q(WX5981) ) ;
AND2    gate1958  (.A(WX5919), .B(RESET), .Z(WX5982) ) ;
DFF     gate1959  (.D(WX5982), .CP(CLK), .Q(WX5983) ) ;
AND2    gate1960  (.A(WX5921), .B(RESET), .Z(WX5984) ) ;
DFF     gate1961  (.D(WX5984), .CP(CLK), .Q(WX5985) ) ;
AND2    gate1962  (.A(WX5923), .B(RESET), .Z(WX5986) ) ;
DFF     gate1963  (.D(WX5986), .CP(CLK), .Q(WX5987) ) ;
AND2    gate1964  (.A(WX5925), .B(RESET), .Z(WX5988) ) ;
DFF     gate1965  (.D(WX5988), .CP(CLK), .Q(WX5989) ) ;
AND2    gate1966  (.A(WX5927), .B(RESET), .Z(WX5990) ) ;
DFF     gate1967  (.D(WX5990), .CP(CLK), .Q(WX5991) ) ;
AND2    gate1968  (.A(WX5929), .B(RESET), .Z(WX5992) ) ;
DFF     gate1969  (.D(WX5992), .CP(CLK), .Q(WX5993) ) ;
AND2    gate1970  (.A(WX5931), .B(RESET), .Z(WX5994) ) ;
DFF     gate1971  (.D(WX5994), .CP(CLK), .Q(WX5995) ) ;
AND2    gate1972  (.A(WX5933), .B(RESET), .Z(WX5996) ) ;
DFF     gate1973  (.D(WX5996), .CP(CLK), .Q(WX5997) ) ;
AND2    gate1974  (.A(WX5935), .B(RESET), .Z(WX5998) ) ;
DFF     gate1975  (.D(WX5998), .CP(CLK), .Q(WX5999) ) ;
AND2    gate1976  (.A(WX5937), .B(RESET), .Z(WX6000) ) ;
DFF     gate1977  (.D(WX6000), .CP(CLK), .Q(WX6001) ) ;
AND2    gate1978  (.A(WX5939), .B(RESET), .Z(WX6002) ) ;
DFF     gate1979  (.D(WX6002), .CP(CLK), .Q(WX6003) ) ;
AND2    gate1980  (.A(WX5941), .B(RESET), .Z(WX6004) ) ;
DFF     gate1981  (.D(WX6004), .CP(CLK), .Q(WX6005) ) ;
AND2    gate1982  (.A(WX5943), .B(RESET), .Z(WX6006) ) ;
DFF     gate1983  (.D(WX6006), .CP(CLK), .Q(WX6007) ) ;
AND2    gate1984  (.A(WX5945), .B(RESET), .Z(WX6008) ) ;
DFF     gate1985  (.D(WX6008), .CP(CLK), .Q(WX6009) ) ;
AND2    gate1986  (.A(WX5947), .B(RESET), .Z(WX6010) ) ;
DFF     gate1987  (.D(WX6010), .CP(CLK), .Q(WX6011) ) ;
AND2    gate1988  (.A(WX5949), .B(RESET), .Z(WX6012) ) ;
DFF     gate1989  (.D(WX6012), .CP(CLK), .Q(WX6013) ) ;
AND2    gate1990  (.A(WX5951), .B(RESET), .Z(WX6014) ) ;
DFF     gate1991  (.D(WX6014), .CP(CLK), .Q(WX6015) ) ;
AND2    gate1992  (.A(WX5953), .B(RESET), .Z(WX6016) ) ;
DFF     gate1993  (.D(WX6016), .CP(CLK), .Q(WX6017) ) ;
AND2    gate1994  (.A(WX5955), .B(RESET), .Z(WX6018) ) ;
DFF     gate1995  (.D(WX6018), .CP(CLK), .Q(WX6019) ) ;
AND2    gate1996  (.A(WX5957), .B(RESET), .Z(WX6020) ) ;
DFF     gate1997  (.D(WX6020), .CP(CLK), .Q(WX6021) ) ;
AND2    gate1998  (.A(WX5959), .B(RESET), .Z(WX6022) ) ;
DFF     gate1999  (.D(WX6022), .CP(CLK), .Q(WX6023) ) ;
AND2    gate2000  (.A(WX5961), .B(RESET), .Z(WX6024) ) ;
DFF     gate2001  (.D(WX6024), .CP(CLK), .Q(WX6025) ) ;
AND2    gate2002  (.A(WX5963), .B(RESET), .Z(WX6026) ) ;
DFF     gate2003  (.D(WX6026), .CP(CLK), .Q(WX6027) ) ;
AND2    gate2004  (.A(WX5965), .B(RESET), .Z(WX6028) ) ;
DFF     gate2005  (.D(WX6028), .CP(CLK), .Q(WX6029) ) ;
AND2    gate2006  (.A(WX5967), .B(RESET), .Z(WX6030) ) ;
DFF     gate2007  (.D(WX6030), .CP(CLK), .Q(WX6031) ) ;
AND2    gate2008  (.A(WX5969), .B(RESET), .Z(WX6032) ) ;
DFF     gate2009  (.D(WX6032), .CP(CLK), .Q(WX6033) ) ;
AND2    gate2010  (.A(WX5971), .B(RESET), .Z(WX6034) ) ;
DFF     gate2011  (.D(WX6034), .CP(CLK), .Q(WX6035) ) ;
AND2    gate2012  (.A(WX5973), .B(RESET), .Z(WX6036) ) ;
DFF     gate2013  (.D(WX6036), .CP(CLK), .Q(WX6037) ) ;
AND2    gate2014  (.A(WX5975), .B(RESET), .Z(WX6038) ) ;
DFF     gate2015  (.D(WX6038), .CP(CLK), .Q(WX6039) ) ;
AND2    gate2016  (.A(WX5977), .B(RESET), .Z(WX6040) ) ;
DFF     gate2017  (.D(WX6040), .CP(CLK), .Q(WX6041) ) ;
AND2    gate2018  (.A(WX5979), .B(RESET), .Z(WX6042) ) ;
DFF     gate2019  (.D(WX6042), .CP(CLK), .Q(WX6043) ) ;
AND2    gate2020  (.A(WX5981), .B(RESET), .Z(WX6044) ) ;
DFF     gate2021  (.D(WX6044), .CP(CLK), .Q(WX6045) ) ;
AND2    gate2022  (.A(WX5983), .B(RESET), .Z(WX6046) ) ;
DFF     gate2023  (.D(WX6046), .CP(CLK), .Q(WX6047) ) ;
AND2    gate2024  (.A(WX5985), .B(RESET), .Z(WX6048) ) ;
DFF     gate2025  (.D(WX6048), .CP(CLK), .Q(WX6049) ) ;
AND2    gate2026  (.A(WX5987), .B(RESET), .Z(WX6050) ) ;
DFF     gate2027  (.D(WX6050), .CP(CLK), .Q(WX6051) ) ;
AND2    gate2028  (.A(WX5989), .B(RESET), .Z(WX6052) ) ;
DFF     gate2029  (.D(WX6052), .CP(CLK), .Q(WX6053) ) ;
AND2    gate2030  (.A(WX5991), .B(RESET), .Z(WX6054) ) ;
DFF     gate2031  (.D(WX6054), .CP(CLK), .Q(WX6055) ) ;
AND2    gate2032  (.A(WX5993), .B(RESET), .Z(WX6056) ) ;
DFF     gate2033  (.D(WX6056), .CP(CLK), .Q(WX6057) ) ;
AND2    gate2034  (.A(WX5995), .B(RESET), .Z(WX6058) ) ;
DFF     gate2035  (.D(WX6058), .CP(CLK), .Q(WX6059) ) ;
AND2    gate2036  (.A(WX5997), .B(RESET), .Z(WX6060) ) ;
DFF     gate2037  (.D(WX6060), .CP(CLK), .Q(WX6061) ) ;
AND2    gate2038  (.A(WX5999), .B(RESET), .Z(WX6062) ) ;
DFF     gate2039  (.D(WX6062), .CP(CLK), .Q(WX6063) ) ;
AND2    gate2040  (.A(WX6001), .B(RESET), .Z(WX6064) ) ;
DFF     gate2041  (.D(WX6064), .CP(CLK), .Q(WX6065) ) ;
AND2    gate2042  (.A(WX6003), .B(RESET), .Z(WX6066) ) ;
DFF     gate2043  (.D(WX6066), .CP(CLK), .Q(WX6067) ) ;
AND2    gate2044  (.A(WX6005), .B(RESET), .Z(WX6068) ) ;
DFF     gate2045  (.D(WX6068), .CP(CLK), .Q(WX6069) ) ;
AND2    gate2046  (.A(WX6007), .B(RESET), .Z(WX6070) ) ;
DFF     gate2047  (.D(WX6070), .CP(CLK), .Q(WX6071) ) ;
AND2    gate2048  (.A(WX6406), .B(WX6435), .Z(WX6436) ) ;
AND2    gate2049  (.A(WX6434), .B(WX6435), .Z(WX6438) ) ;
AND2    gate2050  (.A(WX6433), .B(WX6435), .Z(WX6440) ) ;
AND2    gate2051  (.A(WX6432), .B(WX6435), .Z(WX6442) ) ;
AND2    gate2052  (.A(WX6405), .B(WX6435), .Z(WX6444) ) ;
AND2    gate2053  (.A(WX6431), .B(WX6435), .Z(WX6446) ) ;
AND2    gate2054  (.A(WX6430), .B(WX6435), .Z(WX6448) ) ;
AND2    gate2055  (.A(WX6429), .B(WX6435), .Z(WX6450) ) ;
AND2    gate2056  (.A(WX6428), .B(WX6435), .Z(WX6452) ) ;
AND2    gate2057  (.A(WX6427), .B(WX6435), .Z(WX6454) ) ;
AND2    gate2058  (.A(WX6426), .B(WX6435), .Z(WX6456) ) ;
AND2    gate2059  (.A(WX6404), .B(WX6435), .Z(WX6458) ) ;
AND2    gate2060  (.A(WX6425), .B(WX6435), .Z(WX6460) ) ;
AND2    gate2061  (.A(WX6424), .B(WX6435), .Z(WX6462) ) ;
AND2    gate2062  (.A(WX6423), .B(WX6435), .Z(WX6464) ) ;
AND2    gate2063  (.A(WX6422), .B(WX6435), .Z(WX6466) ) ;
AND2    gate2064  (.A(WX6403), .B(WX6435), .Z(WX6468) ) ;
AND2    gate2065  (.A(WX6421), .B(WX6435), .Z(WX6470) ) ;
AND2    gate2066  (.A(WX6420), .B(WX6435), .Z(WX6472) ) ;
AND2    gate2067  (.A(WX6419), .B(WX6435), .Z(WX6474) ) ;
AND2    gate2068  (.A(WX6418), .B(WX6435), .Z(WX6476) ) ;
AND2    gate2069  (.A(WX6417), .B(WX6435), .Z(WX6478) ) ;
AND2    gate2070  (.A(WX6416), .B(WX6435), .Z(WX6480) ) ;
AND2    gate2071  (.A(WX6415), .B(WX6435), .Z(WX6482) ) ;
AND2    gate2072  (.A(WX6414), .B(WX6435), .Z(WX6484) ) ;
AND2    gate2073  (.A(WX6413), .B(WX6435), .Z(WX6486) ) ;
AND2    gate2074  (.A(WX6412), .B(WX6435), .Z(WX6488) ) ;
AND2    gate2075  (.A(WX6411), .B(WX6435), .Z(WX6490) ) ;
AND2    gate2076  (.A(WX6410), .B(WX6435), .Z(WX6492) ) ;
AND2    gate2077  (.A(WX6409), .B(WX6435), .Z(WX6494) ) ;
AND2    gate2078  (.A(WX6408), .B(WX6435), .Z(WX6496) ) ;
AND2    gate2079  (.A(WX6407), .B(WX6435), .Z(WX6498) ) ;
AND2    gate2080  (.A(WX6952), .B(RESET), .Z(WX6949) ) ;
DFF     gate2081  (.D(WX6949), .CP(CLK), .Q(WX6950) ) ;
AND2    gate2082  (.A(WX6954), .B(RESET), .Z(WX6951) ) ;
DFF     gate2083  (.D(WX6951), .CP(CLK), .Q(WX6952) ) ;
AND2    gate2084  (.A(WX6956), .B(RESET), .Z(WX6953) ) ;
DFF     gate2085  (.D(WX6953), .CP(CLK), .Q(WX6954) ) ;
AND2    gate2086  (.A(WX6958), .B(RESET), .Z(WX6955) ) ;
DFF     gate2087  (.D(WX6955), .CP(CLK), .Q(WX6956) ) ;
AND2    gate2088  (.A(WX6960), .B(RESET), .Z(WX6957) ) ;
DFF     gate2089  (.D(WX6957), .CP(CLK), .Q(WX6958) ) ;
AND2    gate2090  (.A(WX6962), .B(RESET), .Z(WX6959) ) ;
DFF     gate2091  (.D(WX6959), .CP(CLK), .Q(WX6960) ) ;
AND2    gate2092  (.A(WX6964), .B(RESET), .Z(WX6961) ) ;
DFF     gate2093  (.D(WX6961), .CP(CLK), .Q(WX6962) ) ;
AND2    gate2094  (.A(WX6966), .B(RESET), .Z(WX6963) ) ;
DFF     gate2095  (.D(WX6963), .CP(CLK), .Q(WX6964) ) ;
AND2    gate2096  (.A(WX6968), .B(RESET), .Z(WX6965) ) ;
DFF     gate2097  (.D(WX6965), .CP(CLK), .Q(WX6966) ) ;
AND2    gate2098  (.A(WX6970), .B(RESET), .Z(WX6967) ) ;
DFF     gate2099  (.D(WX6967), .CP(CLK), .Q(WX6968) ) ;
AND2    gate2100  (.A(WX6972), .B(RESET), .Z(WX6969) ) ;
DFF     gate2101  (.D(WX6969), .CP(CLK), .Q(WX6970) ) ;
AND2    gate2102  (.A(WX6974), .B(RESET), .Z(WX6971) ) ;
DFF     gate2103  (.D(WX6971), .CP(CLK), .Q(WX6972) ) ;
AND2    gate2104  (.A(WX6976), .B(RESET), .Z(WX6973) ) ;
DFF     gate2105  (.D(WX6973), .CP(CLK), .Q(WX6974) ) ;
AND2    gate2106  (.A(WX6978), .B(RESET), .Z(WX6975) ) ;
DFF     gate2107  (.D(WX6975), .CP(CLK), .Q(WX6976) ) ;
AND2    gate2108  (.A(WX6980), .B(RESET), .Z(WX6977) ) ;
DFF     gate2109  (.D(WX6977), .CP(CLK), .Q(WX6978) ) ;
AND2    gate2110  (.A(WX6982), .B(RESET), .Z(WX6979) ) ;
DFF     gate2111  (.D(WX6979), .CP(CLK), .Q(WX6980) ) ;
AND2    gate2112  (.A(WX6984), .B(RESET), .Z(WX6981) ) ;
DFF     gate2113  (.D(WX6981), .CP(CLK), .Q(WX6982) ) ;
AND2    gate2114  (.A(WX6986), .B(RESET), .Z(WX6983) ) ;
DFF     gate2115  (.D(WX6983), .CP(CLK), .Q(WX6984) ) ;
AND2    gate2116  (.A(WX6988), .B(RESET), .Z(WX6985) ) ;
DFF     gate2117  (.D(WX6985), .CP(CLK), .Q(WX6986) ) ;
AND2    gate2118  (.A(WX6990), .B(RESET), .Z(WX6987) ) ;
DFF     gate2119  (.D(WX6987), .CP(CLK), .Q(WX6988) ) ;
AND2    gate2120  (.A(WX6992), .B(RESET), .Z(WX6989) ) ;
DFF     gate2121  (.D(WX6989), .CP(CLK), .Q(WX6990) ) ;
AND2    gate2122  (.A(WX6994), .B(RESET), .Z(WX6991) ) ;
DFF     gate2123  (.D(WX6991), .CP(CLK), .Q(WX6992) ) ;
AND2    gate2124  (.A(WX6996), .B(RESET), .Z(WX6993) ) ;
DFF     gate2125  (.D(WX6993), .CP(CLK), .Q(WX6994) ) ;
AND2    gate2126  (.A(WX6998), .B(RESET), .Z(WX6995) ) ;
DFF     gate2127  (.D(WX6995), .CP(CLK), .Q(WX6996) ) ;
AND2    gate2128  (.A(WX7000), .B(RESET), .Z(WX6997) ) ;
DFF     gate2129  (.D(WX6997), .CP(CLK), .Q(WX6998) ) ;
AND2    gate2130  (.A(WX7002), .B(RESET), .Z(WX6999) ) ;
DFF     gate2131  (.D(WX6999), .CP(CLK), .Q(WX7000) ) ;
AND2    gate2132  (.A(WX7004), .B(RESET), .Z(WX7001) ) ;
DFF     gate2133  (.D(WX7001), .CP(CLK), .Q(WX7002) ) ;
AND2    gate2134  (.A(WX7006), .B(RESET), .Z(WX7003) ) ;
DFF     gate2135  (.D(WX7003), .CP(CLK), .Q(WX7004) ) ;
AND2    gate2136  (.A(WX7008), .B(RESET), .Z(WX7005) ) ;
DFF     gate2137  (.D(WX7005), .CP(CLK), .Q(WX7006) ) ;
AND2    gate2138  (.A(WX7010), .B(RESET), .Z(WX7007) ) ;
DFF     gate2139  (.D(WX7007), .CP(CLK), .Q(WX7008) ) ;
AND2    gate2140  (.A(WX7012), .B(RESET), .Z(WX7009) ) ;
DFF     gate2141  (.D(WX7009), .CP(CLK), .Q(WX7010) ) ;
AND2    gate2142  (.A(WX6948), .B(RESET), .Z(WX7011) ) ;
DFF     gate2143  (.D(WX7011), .CP(CLK), .Q(WX7012) ) ;
AND2    gate2144  (.A(WX6513), .B(RESET), .Z(WX7109) ) ;
DFF     gate2145  (.D(WX7109), .CP(CLK), .Q(WX7110) ) ;
AND2    gate2146  (.A(WX6527), .B(RESET), .Z(WX7111) ) ;
DFF     gate2147  (.D(WX7111), .CP(CLK), .Q(WX7112) ) ;
AND2    gate2148  (.A(WX6541), .B(RESET), .Z(WX7113) ) ;
DFF     gate2149  (.D(WX7113), .CP(CLK), .Q(WX7114) ) ;
AND2    gate2150  (.A(WX6555), .B(RESET), .Z(WX7115) ) ;
DFF     gate2151  (.D(WX7115), .CP(CLK), .Q(WX7116) ) ;
AND2    gate2152  (.A(WX6569), .B(RESET), .Z(WX7117) ) ;
DFF     gate2153  (.D(WX7117), .CP(CLK), .Q(WX7118) ) ;
AND2    gate2154  (.A(WX6583), .B(RESET), .Z(WX7119) ) ;
DFF     gate2155  (.D(WX7119), .CP(CLK), .Q(WX7120) ) ;
AND2    gate2156  (.A(WX6597), .B(RESET), .Z(WX7121) ) ;
DFF     gate2157  (.D(WX7121), .CP(CLK), .Q(WX7122) ) ;
AND2    gate2158  (.A(WX6611), .B(RESET), .Z(WX7123) ) ;
DFF     gate2159  (.D(WX7123), .CP(CLK), .Q(WX7124) ) ;
AND2    gate2160  (.A(WX6625), .B(RESET), .Z(WX7125) ) ;
DFF     gate2161  (.D(WX7125), .CP(CLK), .Q(WX7126) ) ;
AND2    gate2162  (.A(WX6639), .B(RESET), .Z(WX7127) ) ;
DFF     gate2163  (.D(WX7127), .CP(CLK), .Q(WX7128) ) ;
AND2    gate2164  (.A(WX6653), .B(RESET), .Z(WX7129) ) ;
DFF     gate2165  (.D(WX7129), .CP(CLK), .Q(WX7130) ) ;
AND2    gate2166  (.A(WX6667), .B(RESET), .Z(WX7131) ) ;
DFF     gate2167  (.D(WX7131), .CP(CLK), .Q(WX7132) ) ;
AND2    gate2168  (.A(WX6681), .B(RESET), .Z(WX7133) ) ;
DFF     gate2169  (.D(WX7133), .CP(CLK), .Q(WX7134) ) ;
AND2    gate2170  (.A(WX6695), .B(RESET), .Z(WX7135) ) ;
DFF     gate2171  (.D(WX7135), .CP(CLK), .Q(WX7136) ) ;
AND2    gate2172  (.A(WX6709), .B(RESET), .Z(WX7137) ) ;
DFF     gate2173  (.D(WX7137), .CP(CLK), .Q(WX7138) ) ;
AND2    gate2174  (.A(WX6723), .B(RESET), .Z(WX7139) ) ;
DFF     gate2175  (.D(WX7139), .CP(CLK), .Q(WX7140) ) ;
AND2    gate2176  (.A(WX6737), .B(RESET), .Z(WX7141) ) ;
DFF     gate2177  (.D(WX7141), .CP(CLK), .Q(WX7142) ) ;
AND2    gate2178  (.A(WX6751), .B(RESET), .Z(WX7143) ) ;
DFF     gate2179  (.D(WX7143), .CP(CLK), .Q(WX7144) ) ;
AND2    gate2180  (.A(WX6765), .B(RESET), .Z(WX7145) ) ;
DFF     gate2181  (.D(WX7145), .CP(CLK), .Q(WX7146) ) ;
AND2    gate2182  (.A(WX6779), .B(RESET), .Z(WX7147) ) ;
DFF     gate2183  (.D(WX7147), .CP(CLK), .Q(WX7148) ) ;
AND2    gate2184  (.A(WX6793), .B(RESET), .Z(WX7149) ) ;
DFF     gate2185  (.D(WX7149), .CP(CLK), .Q(WX7150) ) ;
AND2    gate2186  (.A(WX6807), .B(RESET), .Z(WX7151) ) ;
DFF     gate2187  (.D(WX7151), .CP(CLK), .Q(WX7152) ) ;
AND2    gate2188  (.A(WX6821), .B(RESET), .Z(WX7153) ) ;
DFF     gate2189  (.D(WX7153), .CP(CLK), .Q(WX7154) ) ;
AND2    gate2190  (.A(WX6835), .B(RESET), .Z(WX7155) ) ;
DFF     gate2191  (.D(WX7155), .CP(CLK), .Q(WX7156) ) ;
AND2    gate2192  (.A(WX6849), .B(RESET), .Z(WX7157) ) ;
DFF     gate2193  (.D(WX7157), .CP(CLK), .Q(WX7158) ) ;
AND2    gate2194  (.A(WX6863), .B(RESET), .Z(WX7159) ) ;
DFF     gate2195  (.D(WX7159), .CP(CLK), .Q(WX7160) ) ;
AND2    gate2196  (.A(WX6877), .B(RESET), .Z(WX7161) ) ;
DFF     gate2197  (.D(WX7161), .CP(CLK), .Q(WX7162) ) ;
AND2    gate2198  (.A(WX6891), .B(RESET), .Z(WX7163) ) ;
DFF     gate2199  (.D(WX7163), .CP(CLK), .Q(WX7164) ) ;
AND2    gate2200  (.A(WX6905), .B(RESET), .Z(WX7165) ) ;
DFF     gate2201  (.D(WX7165), .CP(CLK), .Q(WX7166) ) ;
AND2    gate2202  (.A(WX6919), .B(RESET), .Z(WX7167) ) ;
DFF     gate2203  (.D(WX7167), .CP(CLK), .Q(WX7168) ) ;
AND2    gate2204  (.A(WX6933), .B(RESET), .Z(WX7169) ) ;
DFF     gate2205  (.D(WX7169), .CP(CLK), .Q(WX7170) ) ;
AND2    gate2206  (.A(WX6947), .B(RESET), .Z(WX7171) ) ;
DFF     gate2207  (.D(WX7171), .CP(CLK), .Q(WX7172) ) ;
AND2    gate2208  (.A(WX7110), .B(RESET), .Z(WX7173) ) ;
DFF     gate2209  (.D(WX7173), .CP(CLK), .Q(WX7174) ) ;
AND2    gate2210  (.A(WX7112), .B(RESET), .Z(WX7175) ) ;
DFF     gate2211  (.D(WX7175), .CP(CLK), .Q(WX7176) ) ;
AND2    gate2212  (.A(WX7114), .B(RESET), .Z(WX7177) ) ;
DFF     gate2213  (.D(WX7177), .CP(CLK), .Q(WX7178) ) ;
AND2    gate2214  (.A(WX7116), .B(RESET), .Z(WX7179) ) ;
DFF     gate2215  (.D(WX7179), .CP(CLK), .Q(WX7180) ) ;
AND2    gate2216  (.A(WX7118), .B(RESET), .Z(WX7181) ) ;
DFF     gate2217  (.D(WX7181), .CP(CLK), .Q(WX7182) ) ;
AND2    gate2218  (.A(WX7120), .B(RESET), .Z(WX7183) ) ;
DFF     gate2219  (.D(WX7183), .CP(CLK), .Q(WX7184) ) ;
AND2    gate2220  (.A(WX7122), .B(RESET), .Z(WX7185) ) ;
DFF     gate2221  (.D(WX7185), .CP(CLK), .Q(WX7186) ) ;
AND2    gate2222  (.A(WX7124), .B(RESET), .Z(WX7187) ) ;
DFF     gate2223  (.D(WX7187), .CP(CLK), .Q(WX7188) ) ;
AND2    gate2224  (.A(WX7126), .B(RESET), .Z(WX7189) ) ;
DFF     gate2225  (.D(WX7189), .CP(CLK), .Q(WX7190) ) ;
AND2    gate2226  (.A(WX7128), .B(RESET), .Z(WX7191) ) ;
DFF     gate2227  (.D(WX7191), .CP(CLK), .Q(WX7192) ) ;
AND2    gate2228  (.A(WX7130), .B(RESET), .Z(WX7193) ) ;
DFF     gate2229  (.D(WX7193), .CP(CLK), .Q(WX7194) ) ;
AND2    gate2230  (.A(WX7132), .B(RESET), .Z(WX7195) ) ;
DFF     gate2231  (.D(WX7195), .CP(CLK), .Q(WX7196) ) ;
AND2    gate2232  (.A(WX7134), .B(RESET), .Z(WX7197) ) ;
DFF     gate2233  (.D(WX7197), .CP(CLK), .Q(WX7198) ) ;
AND2    gate2234  (.A(WX7136), .B(RESET), .Z(WX7199) ) ;
DFF     gate2235  (.D(WX7199), .CP(CLK), .Q(WX7200) ) ;
AND2    gate2236  (.A(WX7138), .B(RESET), .Z(WX7201) ) ;
DFF     gate2237  (.D(WX7201), .CP(CLK), .Q(WX7202) ) ;
AND2    gate2238  (.A(WX7140), .B(RESET), .Z(WX7203) ) ;
DFF     gate2239  (.D(WX7203), .CP(CLK), .Q(WX7204) ) ;
AND2    gate2240  (.A(WX7142), .B(RESET), .Z(WX7205) ) ;
DFF     gate2241  (.D(WX7205), .CP(CLK), .Q(WX7206) ) ;
AND2    gate2242  (.A(WX7144), .B(RESET), .Z(WX7207) ) ;
DFF     gate2243  (.D(WX7207), .CP(CLK), .Q(WX7208) ) ;
AND2    gate2244  (.A(WX7146), .B(RESET), .Z(WX7209) ) ;
DFF     gate2245  (.D(WX7209), .CP(CLK), .Q(WX7210) ) ;
AND2    gate2246  (.A(WX7148), .B(RESET), .Z(WX7211) ) ;
DFF     gate2247  (.D(WX7211), .CP(CLK), .Q(WX7212) ) ;
AND2    gate2248  (.A(WX7150), .B(RESET), .Z(WX7213) ) ;
DFF     gate2249  (.D(WX7213), .CP(CLK), .Q(WX7214) ) ;
AND2    gate2250  (.A(WX7152), .B(RESET), .Z(WX7215) ) ;
DFF     gate2251  (.D(WX7215), .CP(CLK), .Q(WX7216) ) ;
AND2    gate2252  (.A(WX7154), .B(RESET), .Z(WX7217) ) ;
DFF     gate2253  (.D(WX7217), .CP(CLK), .Q(WX7218) ) ;
AND2    gate2254  (.A(WX7156), .B(RESET), .Z(WX7219) ) ;
DFF     gate2255  (.D(WX7219), .CP(CLK), .Q(WX7220) ) ;
AND2    gate2256  (.A(WX7158), .B(RESET), .Z(WX7221) ) ;
DFF     gate2257  (.D(WX7221), .CP(CLK), .Q(WX7222) ) ;
AND2    gate2258  (.A(WX7160), .B(RESET), .Z(WX7223) ) ;
DFF     gate2259  (.D(WX7223), .CP(CLK), .Q(WX7224) ) ;
AND2    gate2260  (.A(WX7162), .B(RESET), .Z(WX7225) ) ;
DFF     gate2261  (.D(WX7225), .CP(CLK), .Q(WX7226) ) ;
AND2    gate2262  (.A(WX7164), .B(RESET), .Z(WX7227) ) ;
DFF     gate2263  (.D(WX7227), .CP(CLK), .Q(WX7228) ) ;
AND2    gate2264  (.A(WX7166), .B(RESET), .Z(WX7229) ) ;
DFF     gate2265  (.D(WX7229), .CP(CLK), .Q(WX7230) ) ;
AND2    gate2266  (.A(WX7168), .B(RESET), .Z(WX7231) ) ;
DFF     gate2267  (.D(WX7231), .CP(CLK), .Q(WX7232) ) ;
AND2    gate2268  (.A(WX7170), .B(RESET), .Z(WX7233) ) ;
DFF     gate2269  (.D(WX7233), .CP(CLK), .Q(WX7234) ) ;
AND2    gate2270  (.A(WX7172), .B(RESET), .Z(WX7235) ) ;
DFF     gate2271  (.D(WX7235), .CP(CLK), .Q(WX7236) ) ;
AND2    gate2272  (.A(WX7174), .B(RESET), .Z(WX7237) ) ;
DFF     gate2273  (.D(WX7237), .CP(CLK), .Q(WX7238) ) ;
AND2    gate2274  (.A(WX7176), .B(RESET), .Z(WX7239) ) ;
DFF     gate2275  (.D(WX7239), .CP(CLK), .Q(WX7240) ) ;
AND2    gate2276  (.A(WX7178), .B(RESET), .Z(WX7241) ) ;
DFF     gate2277  (.D(WX7241), .CP(CLK), .Q(WX7242) ) ;
AND2    gate2278  (.A(WX7180), .B(RESET), .Z(WX7243) ) ;
DFF     gate2279  (.D(WX7243), .CP(CLK), .Q(WX7244) ) ;
AND2    gate2280  (.A(WX7182), .B(RESET), .Z(WX7245) ) ;
DFF     gate2281  (.D(WX7245), .CP(CLK), .Q(WX7246) ) ;
AND2    gate2282  (.A(WX7184), .B(RESET), .Z(WX7247) ) ;
DFF     gate2283  (.D(WX7247), .CP(CLK), .Q(WX7248) ) ;
AND2    gate2284  (.A(WX7186), .B(RESET), .Z(WX7249) ) ;
DFF     gate2285  (.D(WX7249), .CP(CLK), .Q(WX7250) ) ;
AND2    gate2286  (.A(WX7188), .B(RESET), .Z(WX7251) ) ;
DFF     gate2287  (.D(WX7251), .CP(CLK), .Q(WX7252) ) ;
AND2    gate2288  (.A(WX7190), .B(RESET), .Z(WX7253) ) ;
DFF     gate2289  (.D(WX7253), .CP(CLK), .Q(WX7254) ) ;
AND2    gate2290  (.A(WX7192), .B(RESET), .Z(WX7255) ) ;
DFF     gate2291  (.D(WX7255), .CP(CLK), .Q(WX7256) ) ;
AND2    gate2292  (.A(WX7194), .B(RESET), .Z(WX7257) ) ;
DFF     gate2293  (.D(WX7257), .CP(CLK), .Q(WX7258) ) ;
AND2    gate2294  (.A(WX7196), .B(RESET), .Z(WX7259) ) ;
DFF     gate2295  (.D(WX7259), .CP(CLK), .Q(WX7260) ) ;
AND2    gate2296  (.A(WX7198), .B(RESET), .Z(WX7261) ) ;
DFF     gate2297  (.D(WX7261), .CP(CLK), .Q(WX7262) ) ;
AND2    gate2298  (.A(WX7200), .B(RESET), .Z(WX7263) ) ;
DFF     gate2299  (.D(WX7263), .CP(CLK), .Q(WX7264) ) ;
AND2    gate2300  (.A(WX7202), .B(RESET), .Z(WX7265) ) ;
DFF     gate2301  (.D(WX7265), .CP(CLK), .Q(WX7266) ) ;
AND2    gate2302  (.A(WX7204), .B(RESET), .Z(WX7267) ) ;
DFF     gate2303  (.D(WX7267), .CP(CLK), .Q(WX7268) ) ;
AND2    gate2304  (.A(WX7206), .B(RESET), .Z(WX7269) ) ;
DFF     gate2305  (.D(WX7269), .CP(CLK), .Q(WX7270) ) ;
AND2    gate2306  (.A(WX7208), .B(RESET), .Z(WX7271) ) ;
DFF     gate2307  (.D(WX7271), .CP(CLK), .Q(WX7272) ) ;
AND2    gate2308  (.A(WX7210), .B(RESET), .Z(WX7273) ) ;
DFF     gate2309  (.D(WX7273), .CP(CLK), .Q(WX7274) ) ;
AND2    gate2310  (.A(WX7212), .B(RESET), .Z(WX7275) ) ;
DFF     gate2311  (.D(WX7275), .CP(CLK), .Q(WX7276) ) ;
AND2    gate2312  (.A(WX7214), .B(RESET), .Z(WX7277) ) ;
DFF     gate2313  (.D(WX7277), .CP(CLK), .Q(WX7278) ) ;
AND2    gate2314  (.A(WX7216), .B(RESET), .Z(WX7279) ) ;
DFF     gate2315  (.D(WX7279), .CP(CLK), .Q(WX7280) ) ;
AND2    gate2316  (.A(WX7218), .B(RESET), .Z(WX7281) ) ;
DFF     gate2317  (.D(WX7281), .CP(CLK), .Q(WX7282) ) ;
AND2    gate2318  (.A(WX7220), .B(RESET), .Z(WX7283) ) ;
DFF     gate2319  (.D(WX7283), .CP(CLK), .Q(WX7284) ) ;
AND2    gate2320  (.A(WX7222), .B(RESET), .Z(WX7285) ) ;
DFF     gate2321  (.D(WX7285), .CP(CLK), .Q(WX7286) ) ;
AND2    gate2322  (.A(WX7224), .B(RESET), .Z(WX7287) ) ;
DFF     gate2323  (.D(WX7287), .CP(CLK), .Q(WX7288) ) ;
AND2    gate2324  (.A(WX7226), .B(RESET), .Z(WX7289) ) ;
DFF     gate2325  (.D(WX7289), .CP(CLK), .Q(WX7290) ) ;
AND2    gate2326  (.A(WX7228), .B(RESET), .Z(WX7291) ) ;
DFF     gate2327  (.D(WX7291), .CP(CLK), .Q(WX7292) ) ;
AND2    gate2328  (.A(WX7230), .B(RESET), .Z(WX7293) ) ;
DFF     gate2329  (.D(WX7293), .CP(CLK), .Q(WX7294) ) ;
AND2    gate2330  (.A(WX7232), .B(RESET), .Z(WX7295) ) ;
DFF     gate2331  (.D(WX7295), .CP(CLK), .Q(WX7296) ) ;
AND2    gate2332  (.A(WX7234), .B(RESET), .Z(WX7297) ) ;
DFF     gate2333  (.D(WX7297), .CP(CLK), .Q(WX7298) ) ;
AND2    gate2334  (.A(WX7236), .B(RESET), .Z(WX7299) ) ;
DFF     gate2335  (.D(WX7299), .CP(CLK), .Q(WX7300) ) ;
AND2    gate2336  (.A(WX7238), .B(RESET), .Z(WX7301) ) ;
DFF     gate2337  (.D(WX7301), .CP(CLK), .Q(WX7302) ) ;
AND2    gate2338  (.A(WX7240), .B(RESET), .Z(WX7303) ) ;
DFF     gate2339  (.D(WX7303), .CP(CLK), .Q(WX7304) ) ;
AND2    gate2340  (.A(WX7242), .B(RESET), .Z(WX7305) ) ;
DFF     gate2341  (.D(WX7305), .CP(CLK), .Q(WX7306) ) ;
AND2    gate2342  (.A(WX7244), .B(RESET), .Z(WX7307) ) ;
DFF     gate2343  (.D(WX7307), .CP(CLK), .Q(WX7308) ) ;
AND2    gate2344  (.A(WX7246), .B(RESET), .Z(WX7309) ) ;
DFF     gate2345  (.D(WX7309), .CP(CLK), .Q(WX7310) ) ;
AND2    gate2346  (.A(WX7248), .B(RESET), .Z(WX7311) ) ;
DFF     gate2347  (.D(WX7311), .CP(CLK), .Q(WX7312) ) ;
AND2    gate2348  (.A(WX7250), .B(RESET), .Z(WX7313) ) ;
DFF     gate2349  (.D(WX7313), .CP(CLK), .Q(WX7314) ) ;
AND2    gate2350  (.A(WX7252), .B(RESET), .Z(WX7315) ) ;
DFF     gate2351  (.D(WX7315), .CP(CLK), .Q(WX7316) ) ;
AND2    gate2352  (.A(WX7254), .B(RESET), .Z(WX7317) ) ;
DFF     gate2353  (.D(WX7317), .CP(CLK), .Q(WX7318) ) ;
AND2    gate2354  (.A(WX7256), .B(RESET), .Z(WX7319) ) ;
DFF     gate2355  (.D(WX7319), .CP(CLK), .Q(WX7320) ) ;
AND2    gate2356  (.A(WX7258), .B(RESET), .Z(WX7321) ) ;
DFF     gate2357  (.D(WX7321), .CP(CLK), .Q(WX7322) ) ;
AND2    gate2358  (.A(WX7260), .B(RESET), .Z(WX7323) ) ;
DFF     gate2359  (.D(WX7323), .CP(CLK), .Q(WX7324) ) ;
AND2    gate2360  (.A(WX7262), .B(RESET), .Z(WX7325) ) ;
DFF     gate2361  (.D(WX7325), .CP(CLK), .Q(WX7326) ) ;
AND2    gate2362  (.A(WX7264), .B(RESET), .Z(WX7327) ) ;
DFF     gate2363  (.D(WX7327), .CP(CLK), .Q(WX7328) ) ;
AND2    gate2364  (.A(WX7266), .B(RESET), .Z(WX7329) ) ;
DFF     gate2365  (.D(WX7329), .CP(CLK), .Q(WX7330) ) ;
AND2    gate2366  (.A(WX7268), .B(RESET), .Z(WX7331) ) ;
DFF     gate2367  (.D(WX7331), .CP(CLK), .Q(WX7332) ) ;
AND2    gate2368  (.A(WX7270), .B(RESET), .Z(WX7333) ) ;
DFF     gate2369  (.D(WX7333), .CP(CLK), .Q(WX7334) ) ;
AND2    gate2370  (.A(WX7272), .B(RESET), .Z(WX7335) ) ;
DFF     gate2371  (.D(WX7335), .CP(CLK), .Q(WX7336) ) ;
AND2    gate2372  (.A(WX7274), .B(RESET), .Z(WX7337) ) ;
DFF     gate2373  (.D(WX7337), .CP(CLK), .Q(WX7338) ) ;
AND2    gate2374  (.A(WX7276), .B(RESET), .Z(WX7339) ) ;
DFF     gate2375  (.D(WX7339), .CP(CLK), .Q(WX7340) ) ;
AND2    gate2376  (.A(WX7278), .B(RESET), .Z(WX7341) ) ;
DFF     gate2377  (.D(WX7341), .CP(CLK), .Q(WX7342) ) ;
AND2    gate2378  (.A(WX7280), .B(RESET), .Z(WX7343) ) ;
DFF     gate2379  (.D(WX7343), .CP(CLK), .Q(WX7344) ) ;
AND2    gate2380  (.A(WX7282), .B(RESET), .Z(WX7345) ) ;
DFF     gate2381  (.D(WX7345), .CP(CLK), .Q(WX7346) ) ;
AND2    gate2382  (.A(WX7284), .B(RESET), .Z(WX7347) ) ;
DFF     gate2383  (.D(WX7347), .CP(CLK), .Q(WX7348) ) ;
AND2    gate2384  (.A(WX7286), .B(RESET), .Z(WX7349) ) ;
DFF     gate2385  (.D(WX7349), .CP(CLK), .Q(WX7350) ) ;
AND2    gate2386  (.A(WX7288), .B(RESET), .Z(WX7351) ) ;
DFF     gate2387  (.D(WX7351), .CP(CLK), .Q(WX7352) ) ;
AND2    gate2388  (.A(WX7290), .B(RESET), .Z(WX7353) ) ;
DFF     gate2389  (.D(WX7353), .CP(CLK), .Q(WX7354) ) ;
AND2    gate2390  (.A(WX7292), .B(RESET), .Z(WX7355) ) ;
DFF     gate2391  (.D(WX7355), .CP(CLK), .Q(WX7356) ) ;
AND2    gate2392  (.A(WX7294), .B(RESET), .Z(WX7357) ) ;
DFF     gate2393  (.D(WX7357), .CP(CLK), .Q(WX7358) ) ;
AND2    gate2394  (.A(WX7296), .B(RESET), .Z(WX7359) ) ;
DFF     gate2395  (.D(WX7359), .CP(CLK), .Q(WX7360) ) ;
AND2    gate2396  (.A(WX7298), .B(RESET), .Z(WX7361) ) ;
DFF     gate2397  (.D(WX7361), .CP(CLK), .Q(WX7362) ) ;
AND2    gate2398  (.A(WX7300), .B(RESET), .Z(WX7363) ) ;
DFF     gate2399  (.D(WX7363), .CP(CLK), .Q(WX7364) ) ;
AND2    gate2400  (.A(WX7699), .B(WX7728), .Z(WX7729) ) ;
AND2    gate2401  (.A(WX7727), .B(WX7728), .Z(WX7731) ) ;
AND2    gate2402  (.A(WX7726), .B(WX7728), .Z(WX7733) ) ;
AND2    gate2403  (.A(WX7725), .B(WX7728), .Z(WX7735) ) ;
AND2    gate2404  (.A(WX7698), .B(WX7728), .Z(WX7737) ) ;
AND2    gate2405  (.A(WX7724), .B(WX7728), .Z(WX7739) ) ;
AND2    gate2406  (.A(WX7723), .B(WX7728), .Z(WX7741) ) ;
AND2    gate2407  (.A(WX7722), .B(WX7728), .Z(WX7743) ) ;
AND2    gate2408  (.A(WX7721), .B(WX7728), .Z(WX7745) ) ;
AND2    gate2409  (.A(WX7720), .B(WX7728), .Z(WX7747) ) ;
AND2    gate2410  (.A(WX7719), .B(WX7728), .Z(WX7749) ) ;
AND2    gate2411  (.A(WX7697), .B(WX7728), .Z(WX7751) ) ;
AND2    gate2412  (.A(WX7718), .B(WX7728), .Z(WX7753) ) ;
AND2    gate2413  (.A(WX7717), .B(WX7728), .Z(WX7755) ) ;
AND2    gate2414  (.A(WX7716), .B(WX7728), .Z(WX7757) ) ;
AND2    gate2415  (.A(WX7715), .B(WX7728), .Z(WX7759) ) ;
AND2    gate2416  (.A(WX7696), .B(WX7728), .Z(WX7761) ) ;
AND2    gate2417  (.A(WX7714), .B(WX7728), .Z(WX7763) ) ;
AND2    gate2418  (.A(WX7713), .B(WX7728), .Z(WX7765) ) ;
AND2    gate2419  (.A(WX7712), .B(WX7728), .Z(WX7767) ) ;
AND2    gate2420  (.A(WX7711), .B(WX7728), .Z(WX7769) ) ;
AND2    gate2421  (.A(WX7710), .B(WX7728), .Z(WX7771) ) ;
AND2    gate2422  (.A(WX7709), .B(WX7728), .Z(WX7773) ) ;
AND2    gate2423  (.A(WX7708), .B(WX7728), .Z(WX7775) ) ;
AND2    gate2424  (.A(WX7707), .B(WX7728), .Z(WX7777) ) ;
AND2    gate2425  (.A(WX7706), .B(WX7728), .Z(WX7779) ) ;
AND2    gate2426  (.A(WX7705), .B(WX7728), .Z(WX7781) ) ;
AND2    gate2427  (.A(WX7704), .B(WX7728), .Z(WX7783) ) ;
AND2    gate2428  (.A(WX7703), .B(WX7728), .Z(WX7785) ) ;
AND2    gate2429  (.A(WX7702), .B(WX7728), .Z(WX7787) ) ;
AND2    gate2430  (.A(WX7701), .B(WX7728), .Z(WX7789) ) ;
AND2    gate2431  (.A(WX7700), .B(WX7728), .Z(WX7791) ) ;
AND2    gate2432  (.A(WX8245), .B(RESET), .Z(WX8242) ) ;
DFF     gate2433  (.D(WX8242), .CP(CLK), .Q(WX8243) ) ;
AND2    gate2434  (.A(WX8247), .B(RESET), .Z(WX8244) ) ;
DFF     gate2435  (.D(WX8244), .CP(CLK), .Q(WX8245) ) ;
AND2    gate2436  (.A(WX8249), .B(RESET), .Z(WX8246) ) ;
DFF     gate2437  (.D(WX8246), .CP(CLK), .Q(WX8247) ) ;
AND2    gate2438  (.A(WX8251), .B(RESET), .Z(WX8248) ) ;
DFF     gate2439  (.D(WX8248), .CP(CLK), .Q(WX8249) ) ;
AND2    gate2440  (.A(WX8253), .B(RESET), .Z(WX8250) ) ;
DFF     gate2441  (.D(WX8250), .CP(CLK), .Q(WX8251) ) ;
AND2    gate2442  (.A(WX8255), .B(RESET), .Z(WX8252) ) ;
DFF     gate2443  (.D(WX8252), .CP(CLK), .Q(WX8253) ) ;
AND2    gate2444  (.A(WX8257), .B(RESET), .Z(WX8254) ) ;
DFF     gate2445  (.D(WX8254), .CP(CLK), .Q(WX8255) ) ;
AND2    gate2446  (.A(WX8259), .B(RESET), .Z(WX8256) ) ;
DFF     gate2447  (.D(WX8256), .CP(CLK), .Q(WX8257) ) ;
AND2    gate2448  (.A(WX8261), .B(RESET), .Z(WX8258) ) ;
DFF     gate2449  (.D(WX8258), .CP(CLK), .Q(WX8259) ) ;
AND2    gate2450  (.A(WX8263), .B(RESET), .Z(WX8260) ) ;
DFF     gate2451  (.D(WX8260), .CP(CLK), .Q(WX8261) ) ;
AND2    gate2452  (.A(WX8265), .B(RESET), .Z(WX8262) ) ;
DFF     gate2453  (.D(WX8262), .CP(CLK), .Q(WX8263) ) ;
AND2    gate2454  (.A(WX8267), .B(RESET), .Z(WX8264) ) ;
DFF     gate2455  (.D(WX8264), .CP(CLK), .Q(WX8265) ) ;
AND2    gate2456  (.A(WX8269), .B(RESET), .Z(WX8266) ) ;
DFF     gate2457  (.D(WX8266), .CP(CLK), .Q(WX8267) ) ;
AND2    gate2458  (.A(WX8271), .B(RESET), .Z(WX8268) ) ;
DFF     gate2459  (.D(WX8268), .CP(CLK), .Q(WX8269) ) ;
AND2    gate2460  (.A(WX8273), .B(RESET), .Z(WX8270) ) ;
DFF     gate2461  (.D(WX8270), .CP(CLK), .Q(WX8271) ) ;
AND2    gate2462  (.A(WX8275), .B(RESET), .Z(WX8272) ) ;
DFF     gate2463  (.D(WX8272), .CP(CLK), .Q(WX8273) ) ;
AND2    gate2464  (.A(WX8277), .B(RESET), .Z(WX8274) ) ;
DFF     gate2465  (.D(WX8274), .CP(CLK), .Q(WX8275) ) ;
AND2    gate2466  (.A(WX8279), .B(RESET), .Z(WX8276) ) ;
DFF     gate2467  (.D(WX8276), .CP(CLK), .Q(WX8277) ) ;
AND2    gate2468  (.A(WX8281), .B(RESET), .Z(WX8278) ) ;
DFF     gate2469  (.D(WX8278), .CP(CLK), .Q(WX8279) ) ;
AND2    gate2470  (.A(WX8283), .B(RESET), .Z(WX8280) ) ;
DFF     gate2471  (.D(WX8280), .CP(CLK), .Q(WX8281) ) ;
AND2    gate2472  (.A(WX8285), .B(RESET), .Z(WX8282) ) ;
DFF     gate2473  (.D(WX8282), .CP(CLK), .Q(WX8283) ) ;
AND2    gate2474  (.A(WX8287), .B(RESET), .Z(WX8284) ) ;
DFF     gate2475  (.D(WX8284), .CP(CLK), .Q(WX8285) ) ;
AND2    gate2476  (.A(WX8289), .B(RESET), .Z(WX8286) ) ;
DFF     gate2477  (.D(WX8286), .CP(CLK), .Q(WX8287) ) ;
AND2    gate2478  (.A(WX8291), .B(RESET), .Z(WX8288) ) ;
DFF     gate2479  (.D(WX8288), .CP(CLK), .Q(WX8289) ) ;
AND2    gate2480  (.A(WX8293), .B(RESET), .Z(WX8290) ) ;
DFF     gate2481  (.D(WX8290), .CP(CLK), .Q(WX8291) ) ;
AND2    gate2482  (.A(WX8295), .B(RESET), .Z(WX8292) ) ;
DFF     gate2483  (.D(WX8292), .CP(CLK), .Q(WX8293) ) ;
AND2    gate2484  (.A(WX8297), .B(RESET), .Z(WX8294) ) ;
DFF     gate2485  (.D(WX8294), .CP(CLK), .Q(WX8295) ) ;
AND2    gate2486  (.A(WX8299), .B(RESET), .Z(WX8296) ) ;
DFF     gate2487  (.D(WX8296), .CP(CLK), .Q(WX8297) ) ;
AND2    gate2488  (.A(WX8301), .B(RESET), .Z(WX8298) ) ;
DFF     gate2489  (.D(WX8298), .CP(CLK), .Q(WX8299) ) ;
AND2    gate2490  (.A(WX8303), .B(RESET), .Z(WX8300) ) ;
DFF     gate2491  (.D(WX8300), .CP(CLK), .Q(WX8301) ) ;
AND2    gate2492  (.A(WX8305), .B(RESET), .Z(WX8302) ) ;
DFF     gate2493  (.D(WX8302), .CP(CLK), .Q(WX8303) ) ;
AND2    gate2494  (.A(WX8241), .B(RESET), .Z(WX8304) ) ;
DFF     gate2495  (.D(WX8304), .CP(CLK), .Q(WX8305) ) ;
AND2    gate2496  (.A(WX7806), .B(RESET), .Z(WX8402) ) ;
DFF     gate2497  (.D(WX8402), .CP(CLK), .Q(WX8403) ) ;
AND2    gate2498  (.A(WX7820), .B(RESET), .Z(WX8404) ) ;
DFF     gate2499  (.D(WX8404), .CP(CLK), .Q(WX8405) ) ;
AND2    gate2500  (.A(WX7834), .B(RESET), .Z(WX8406) ) ;
DFF     gate2501  (.D(WX8406), .CP(CLK), .Q(WX8407) ) ;
AND2    gate2502  (.A(WX7848), .B(RESET), .Z(WX8408) ) ;
DFF     gate2503  (.D(WX8408), .CP(CLK), .Q(WX8409) ) ;
AND2    gate2504  (.A(WX7862), .B(RESET), .Z(WX8410) ) ;
DFF     gate2505  (.D(WX8410), .CP(CLK), .Q(WX8411) ) ;
AND2    gate2506  (.A(WX7876), .B(RESET), .Z(WX8412) ) ;
DFF     gate2507  (.D(WX8412), .CP(CLK), .Q(WX8413) ) ;
AND2    gate2508  (.A(WX7890), .B(RESET), .Z(WX8414) ) ;
DFF     gate2509  (.D(WX8414), .CP(CLK), .Q(WX8415) ) ;
AND2    gate2510  (.A(WX7904), .B(RESET), .Z(WX8416) ) ;
DFF     gate2511  (.D(WX8416), .CP(CLK), .Q(WX8417) ) ;
AND2    gate2512  (.A(WX7918), .B(RESET), .Z(WX8418) ) ;
DFF     gate2513  (.D(WX8418), .CP(CLK), .Q(WX8419) ) ;
AND2    gate2514  (.A(WX7932), .B(RESET), .Z(WX8420) ) ;
DFF     gate2515  (.D(WX8420), .CP(CLK), .Q(WX8421) ) ;
AND2    gate2516  (.A(WX7946), .B(RESET), .Z(WX8422) ) ;
DFF     gate2517  (.D(WX8422), .CP(CLK), .Q(WX8423) ) ;
AND2    gate2518  (.A(WX7960), .B(RESET), .Z(WX8424) ) ;
DFF     gate2519  (.D(WX8424), .CP(CLK), .Q(WX8425) ) ;
AND2    gate2520  (.A(WX7974), .B(RESET), .Z(WX8426) ) ;
DFF     gate2521  (.D(WX8426), .CP(CLK), .Q(WX8427) ) ;
AND2    gate2522  (.A(WX7988), .B(RESET), .Z(WX8428) ) ;
DFF     gate2523  (.D(WX8428), .CP(CLK), .Q(WX8429) ) ;
AND2    gate2524  (.A(WX8002), .B(RESET), .Z(WX8430) ) ;
DFF     gate2525  (.D(WX8430), .CP(CLK), .Q(WX8431) ) ;
AND2    gate2526  (.A(WX8016), .B(RESET), .Z(WX8432) ) ;
DFF     gate2527  (.D(WX8432), .CP(CLK), .Q(WX8433) ) ;
AND2    gate2528  (.A(WX8030), .B(RESET), .Z(WX8434) ) ;
DFF     gate2529  (.D(WX8434), .CP(CLK), .Q(WX8435) ) ;
AND2    gate2530  (.A(WX8044), .B(RESET), .Z(WX8436) ) ;
DFF     gate2531  (.D(WX8436), .CP(CLK), .Q(WX8437) ) ;
AND2    gate2532  (.A(WX8058), .B(RESET), .Z(WX8438) ) ;
DFF     gate2533  (.D(WX8438), .CP(CLK), .Q(WX8439) ) ;
AND2    gate2534  (.A(WX8072), .B(RESET), .Z(WX8440) ) ;
DFF     gate2535  (.D(WX8440), .CP(CLK), .Q(WX8441) ) ;
AND2    gate2536  (.A(WX8086), .B(RESET), .Z(WX8442) ) ;
DFF     gate2537  (.D(WX8442), .CP(CLK), .Q(WX8443) ) ;
AND2    gate2538  (.A(WX8100), .B(RESET), .Z(WX8444) ) ;
DFF     gate2539  (.D(WX8444), .CP(CLK), .Q(WX8445) ) ;
AND2    gate2540  (.A(WX8114), .B(RESET), .Z(WX8446) ) ;
DFF     gate2541  (.D(WX8446), .CP(CLK), .Q(WX8447) ) ;
AND2    gate2542  (.A(WX8128), .B(RESET), .Z(WX8448) ) ;
DFF     gate2543  (.D(WX8448), .CP(CLK), .Q(WX8449) ) ;
AND2    gate2544  (.A(WX8142), .B(RESET), .Z(WX8450) ) ;
DFF     gate2545  (.D(WX8450), .CP(CLK), .Q(WX8451) ) ;
AND2    gate2546  (.A(WX8156), .B(RESET), .Z(WX8452) ) ;
DFF     gate2547  (.D(WX8452), .CP(CLK), .Q(WX8453) ) ;
AND2    gate2548  (.A(WX8170), .B(RESET), .Z(WX8454) ) ;
DFF     gate2549  (.D(WX8454), .CP(CLK), .Q(WX8455) ) ;
AND2    gate2550  (.A(WX8184), .B(RESET), .Z(WX8456) ) ;
DFF     gate2551  (.D(WX8456), .CP(CLK), .Q(WX8457) ) ;
AND2    gate2552  (.A(WX8198), .B(RESET), .Z(WX8458) ) ;
DFF     gate2553  (.D(WX8458), .CP(CLK), .Q(WX8459) ) ;
AND2    gate2554  (.A(WX8212), .B(RESET), .Z(WX8460) ) ;
DFF     gate2555  (.D(WX8460), .CP(CLK), .Q(WX8461) ) ;
AND2    gate2556  (.A(WX8226), .B(RESET), .Z(WX8462) ) ;
DFF     gate2557  (.D(WX8462), .CP(CLK), .Q(WX8463) ) ;
AND2    gate2558  (.A(WX8240), .B(RESET), .Z(WX8464) ) ;
DFF     gate2559  (.D(WX8464), .CP(CLK), .Q(WX8465) ) ;
AND2    gate2560  (.A(WX8403), .B(RESET), .Z(WX8466) ) ;
DFF     gate2561  (.D(WX8466), .CP(CLK), .Q(WX8467) ) ;
AND2    gate2562  (.A(WX8405), .B(RESET), .Z(WX8468) ) ;
DFF     gate2563  (.D(WX8468), .CP(CLK), .Q(WX8469) ) ;
AND2    gate2564  (.A(WX8407), .B(RESET), .Z(WX8470) ) ;
DFF     gate2565  (.D(WX8470), .CP(CLK), .Q(WX8471) ) ;
AND2    gate2566  (.A(WX8409), .B(RESET), .Z(WX8472) ) ;
DFF     gate2567  (.D(WX8472), .CP(CLK), .Q(WX8473) ) ;
AND2    gate2568  (.A(WX8411), .B(RESET), .Z(WX8474) ) ;
DFF     gate2569  (.D(WX8474), .CP(CLK), .Q(WX8475) ) ;
AND2    gate2570  (.A(WX8413), .B(RESET), .Z(WX8476) ) ;
DFF     gate2571  (.D(WX8476), .CP(CLK), .Q(WX8477) ) ;
AND2    gate2572  (.A(WX8415), .B(RESET), .Z(WX8478) ) ;
DFF     gate2573  (.D(WX8478), .CP(CLK), .Q(WX8479) ) ;
AND2    gate2574  (.A(WX8417), .B(RESET), .Z(WX8480) ) ;
DFF     gate2575  (.D(WX8480), .CP(CLK), .Q(WX8481) ) ;
AND2    gate2576  (.A(WX8419), .B(RESET), .Z(WX8482) ) ;
DFF     gate2577  (.D(WX8482), .CP(CLK), .Q(WX8483) ) ;
AND2    gate2578  (.A(WX8421), .B(RESET), .Z(WX8484) ) ;
DFF     gate2579  (.D(WX8484), .CP(CLK), .Q(WX8485) ) ;
AND2    gate2580  (.A(WX8423), .B(RESET), .Z(WX8486) ) ;
DFF     gate2581  (.D(WX8486), .CP(CLK), .Q(WX8487) ) ;
AND2    gate2582  (.A(WX8425), .B(RESET), .Z(WX8488) ) ;
DFF     gate2583  (.D(WX8488), .CP(CLK), .Q(WX8489) ) ;
AND2    gate2584  (.A(WX8427), .B(RESET), .Z(WX8490) ) ;
DFF     gate2585  (.D(WX8490), .CP(CLK), .Q(WX8491) ) ;
AND2    gate2586  (.A(WX8429), .B(RESET), .Z(WX8492) ) ;
DFF     gate2587  (.D(WX8492), .CP(CLK), .Q(WX8493) ) ;
AND2    gate2588  (.A(WX8431), .B(RESET), .Z(WX8494) ) ;
DFF     gate2589  (.D(WX8494), .CP(CLK), .Q(WX8495) ) ;
AND2    gate2590  (.A(WX8433), .B(RESET), .Z(WX8496) ) ;
DFF     gate2591  (.D(WX8496), .CP(CLK), .Q(WX8497) ) ;
AND2    gate2592  (.A(WX8435), .B(RESET), .Z(WX8498) ) ;
DFF     gate2593  (.D(WX8498), .CP(CLK), .Q(WX8499) ) ;
AND2    gate2594  (.A(WX8437), .B(RESET), .Z(WX8500) ) ;
DFF     gate2595  (.D(WX8500), .CP(CLK), .Q(WX8501) ) ;
AND2    gate2596  (.A(WX8439), .B(RESET), .Z(WX8502) ) ;
DFF     gate2597  (.D(WX8502), .CP(CLK), .Q(WX8503) ) ;
AND2    gate2598  (.A(WX8441), .B(RESET), .Z(WX8504) ) ;
DFF     gate2599  (.D(WX8504), .CP(CLK), .Q(WX8505) ) ;
AND2    gate2600  (.A(WX8443), .B(RESET), .Z(WX8506) ) ;
DFF     gate2601  (.D(WX8506), .CP(CLK), .Q(WX8507) ) ;
AND2    gate2602  (.A(WX8445), .B(RESET), .Z(WX8508) ) ;
DFF     gate2603  (.D(WX8508), .CP(CLK), .Q(WX8509) ) ;
AND2    gate2604  (.A(WX8447), .B(RESET), .Z(WX8510) ) ;
DFF     gate2605  (.D(WX8510), .CP(CLK), .Q(WX8511) ) ;
AND2    gate2606  (.A(WX8449), .B(RESET), .Z(WX8512) ) ;
DFF     gate2607  (.D(WX8512), .CP(CLK), .Q(WX8513) ) ;
AND2    gate2608  (.A(WX8451), .B(RESET), .Z(WX8514) ) ;
DFF     gate2609  (.D(WX8514), .CP(CLK), .Q(WX8515) ) ;
AND2    gate2610  (.A(WX8453), .B(RESET), .Z(WX8516) ) ;
DFF     gate2611  (.D(WX8516), .CP(CLK), .Q(WX8517) ) ;
AND2    gate2612  (.A(WX8455), .B(RESET), .Z(WX8518) ) ;
DFF     gate2613  (.D(WX8518), .CP(CLK), .Q(WX8519) ) ;
AND2    gate2614  (.A(WX8457), .B(RESET), .Z(WX8520) ) ;
DFF     gate2615  (.D(WX8520), .CP(CLK), .Q(WX8521) ) ;
AND2    gate2616  (.A(WX8459), .B(RESET), .Z(WX8522) ) ;
DFF     gate2617  (.D(WX8522), .CP(CLK), .Q(WX8523) ) ;
AND2    gate2618  (.A(WX8461), .B(RESET), .Z(WX8524) ) ;
DFF     gate2619  (.D(WX8524), .CP(CLK), .Q(WX8525) ) ;
AND2    gate2620  (.A(WX8463), .B(RESET), .Z(WX8526) ) ;
DFF     gate2621  (.D(WX8526), .CP(CLK), .Q(WX8527) ) ;
AND2    gate2622  (.A(WX8465), .B(RESET), .Z(WX8528) ) ;
DFF     gate2623  (.D(WX8528), .CP(CLK), .Q(WX8529) ) ;
AND2    gate2624  (.A(WX8467), .B(RESET), .Z(WX8530) ) ;
DFF     gate2625  (.D(WX8530), .CP(CLK), .Q(WX8531) ) ;
AND2    gate2626  (.A(WX8469), .B(RESET), .Z(WX8532) ) ;
DFF     gate2627  (.D(WX8532), .CP(CLK), .Q(WX8533) ) ;
AND2    gate2628  (.A(WX8471), .B(RESET), .Z(WX8534) ) ;
DFF     gate2629  (.D(WX8534), .CP(CLK), .Q(WX8535) ) ;
AND2    gate2630  (.A(WX8473), .B(RESET), .Z(WX8536) ) ;
DFF     gate2631  (.D(WX8536), .CP(CLK), .Q(WX8537) ) ;
AND2    gate2632  (.A(WX8475), .B(RESET), .Z(WX8538) ) ;
DFF     gate2633  (.D(WX8538), .CP(CLK), .Q(WX8539) ) ;
AND2    gate2634  (.A(WX8477), .B(RESET), .Z(WX8540) ) ;
DFF     gate2635  (.D(WX8540), .CP(CLK), .Q(WX8541) ) ;
AND2    gate2636  (.A(WX8479), .B(RESET), .Z(WX8542) ) ;
DFF     gate2637  (.D(WX8542), .CP(CLK), .Q(WX8543) ) ;
AND2    gate2638  (.A(WX8481), .B(RESET), .Z(WX8544) ) ;
DFF     gate2639  (.D(WX8544), .CP(CLK), .Q(WX8545) ) ;
AND2    gate2640  (.A(WX8483), .B(RESET), .Z(WX8546) ) ;
DFF     gate2641  (.D(WX8546), .CP(CLK), .Q(WX8547) ) ;
AND2    gate2642  (.A(WX8485), .B(RESET), .Z(WX8548) ) ;
DFF     gate2643  (.D(WX8548), .CP(CLK), .Q(WX8549) ) ;
AND2    gate2644  (.A(WX8487), .B(RESET), .Z(WX8550) ) ;
DFF     gate2645  (.D(WX8550), .CP(CLK), .Q(WX8551) ) ;
AND2    gate2646  (.A(WX8489), .B(RESET), .Z(WX8552) ) ;
DFF     gate2647  (.D(WX8552), .CP(CLK), .Q(WX8553) ) ;
AND2    gate2648  (.A(WX8491), .B(RESET), .Z(WX8554) ) ;
DFF     gate2649  (.D(WX8554), .CP(CLK), .Q(WX8555) ) ;
AND2    gate2650  (.A(WX8493), .B(RESET), .Z(WX8556) ) ;
DFF     gate2651  (.D(WX8556), .CP(CLK), .Q(WX8557) ) ;
AND2    gate2652  (.A(WX8495), .B(RESET), .Z(WX8558) ) ;
DFF     gate2653  (.D(WX8558), .CP(CLK), .Q(WX8559) ) ;
AND2    gate2654  (.A(WX8497), .B(RESET), .Z(WX8560) ) ;
DFF     gate2655  (.D(WX8560), .CP(CLK), .Q(WX8561) ) ;
AND2    gate2656  (.A(WX8499), .B(RESET), .Z(WX8562) ) ;
DFF     gate2657  (.D(WX8562), .CP(CLK), .Q(WX8563) ) ;
AND2    gate2658  (.A(WX8501), .B(RESET), .Z(WX8564) ) ;
DFF     gate2659  (.D(WX8564), .CP(CLK), .Q(WX8565) ) ;
AND2    gate2660  (.A(WX8503), .B(RESET), .Z(WX8566) ) ;
DFF     gate2661  (.D(WX8566), .CP(CLK), .Q(WX8567) ) ;
AND2    gate2662  (.A(WX8505), .B(RESET), .Z(WX8568) ) ;
DFF     gate2663  (.D(WX8568), .CP(CLK), .Q(WX8569) ) ;
AND2    gate2664  (.A(WX8507), .B(RESET), .Z(WX8570) ) ;
DFF     gate2665  (.D(WX8570), .CP(CLK), .Q(WX8571) ) ;
AND2    gate2666  (.A(WX8509), .B(RESET), .Z(WX8572) ) ;
DFF     gate2667  (.D(WX8572), .CP(CLK), .Q(WX8573) ) ;
AND2    gate2668  (.A(WX8511), .B(RESET), .Z(WX8574) ) ;
DFF     gate2669  (.D(WX8574), .CP(CLK), .Q(WX8575) ) ;
AND2    gate2670  (.A(WX8513), .B(RESET), .Z(WX8576) ) ;
DFF     gate2671  (.D(WX8576), .CP(CLK), .Q(WX8577) ) ;
AND2    gate2672  (.A(WX8515), .B(RESET), .Z(WX8578) ) ;
DFF     gate2673  (.D(WX8578), .CP(CLK), .Q(WX8579) ) ;
AND2    gate2674  (.A(WX8517), .B(RESET), .Z(WX8580) ) ;
DFF     gate2675  (.D(WX8580), .CP(CLK), .Q(WX8581) ) ;
AND2    gate2676  (.A(WX8519), .B(RESET), .Z(WX8582) ) ;
DFF     gate2677  (.D(WX8582), .CP(CLK), .Q(WX8583) ) ;
AND2    gate2678  (.A(WX8521), .B(RESET), .Z(WX8584) ) ;
DFF     gate2679  (.D(WX8584), .CP(CLK), .Q(WX8585) ) ;
AND2    gate2680  (.A(WX8523), .B(RESET), .Z(WX8586) ) ;
DFF     gate2681  (.D(WX8586), .CP(CLK), .Q(WX8587) ) ;
AND2    gate2682  (.A(WX8525), .B(RESET), .Z(WX8588) ) ;
DFF     gate2683  (.D(WX8588), .CP(CLK), .Q(WX8589) ) ;
AND2    gate2684  (.A(WX8527), .B(RESET), .Z(WX8590) ) ;
DFF     gate2685  (.D(WX8590), .CP(CLK), .Q(WX8591) ) ;
AND2    gate2686  (.A(WX8529), .B(RESET), .Z(WX8592) ) ;
DFF     gate2687  (.D(WX8592), .CP(CLK), .Q(WX8593) ) ;
AND2    gate2688  (.A(WX8531), .B(RESET), .Z(WX8594) ) ;
DFF     gate2689  (.D(WX8594), .CP(CLK), .Q(WX8595) ) ;
AND2    gate2690  (.A(WX8533), .B(RESET), .Z(WX8596) ) ;
DFF     gate2691  (.D(WX8596), .CP(CLK), .Q(WX8597) ) ;
AND2    gate2692  (.A(WX8535), .B(RESET), .Z(WX8598) ) ;
DFF     gate2693  (.D(WX8598), .CP(CLK), .Q(WX8599) ) ;
AND2    gate2694  (.A(WX8537), .B(RESET), .Z(WX8600) ) ;
DFF     gate2695  (.D(WX8600), .CP(CLK), .Q(WX8601) ) ;
AND2    gate2696  (.A(WX8539), .B(RESET), .Z(WX8602) ) ;
DFF     gate2697  (.D(WX8602), .CP(CLK), .Q(WX8603) ) ;
AND2    gate2698  (.A(WX8541), .B(RESET), .Z(WX8604) ) ;
DFF     gate2699  (.D(WX8604), .CP(CLK), .Q(WX8605) ) ;
AND2    gate2700  (.A(WX8543), .B(RESET), .Z(WX8606) ) ;
DFF     gate2701  (.D(WX8606), .CP(CLK), .Q(WX8607) ) ;
AND2    gate2702  (.A(WX8545), .B(RESET), .Z(WX8608) ) ;
DFF     gate2703  (.D(WX8608), .CP(CLK), .Q(WX8609) ) ;
AND2    gate2704  (.A(WX8547), .B(RESET), .Z(WX8610) ) ;
DFF     gate2705  (.D(WX8610), .CP(CLK), .Q(WX8611) ) ;
AND2    gate2706  (.A(WX8549), .B(RESET), .Z(WX8612) ) ;
DFF     gate2707  (.D(WX8612), .CP(CLK), .Q(WX8613) ) ;
AND2    gate2708  (.A(WX8551), .B(RESET), .Z(WX8614) ) ;
DFF     gate2709  (.D(WX8614), .CP(CLK), .Q(WX8615) ) ;
AND2    gate2710  (.A(WX8553), .B(RESET), .Z(WX8616) ) ;
DFF     gate2711  (.D(WX8616), .CP(CLK), .Q(WX8617) ) ;
AND2    gate2712  (.A(WX8555), .B(RESET), .Z(WX8618) ) ;
DFF     gate2713  (.D(WX8618), .CP(CLK), .Q(WX8619) ) ;
AND2    gate2714  (.A(WX8557), .B(RESET), .Z(WX8620) ) ;
DFF     gate2715  (.D(WX8620), .CP(CLK), .Q(WX8621) ) ;
AND2    gate2716  (.A(WX8559), .B(RESET), .Z(WX8622) ) ;
DFF     gate2717  (.D(WX8622), .CP(CLK), .Q(WX8623) ) ;
AND2    gate2718  (.A(WX8561), .B(RESET), .Z(WX8624) ) ;
DFF     gate2719  (.D(WX8624), .CP(CLK), .Q(WX8625) ) ;
AND2    gate2720  (.A(WX8563), .B(RESET), .Z(WX8626) ) ;
DFF     gate2721  (.D(WX8626), .CP(CLK), .Q(WX8627) ) ;
AND2    gate2722  (.A(WX8565), .B(RESET), .Z(WX8628) ) ;
DFF     gate2723  (.D(WX8628), .CP(CLK), .Q(WX8629) ) ;
AND2    gate2724  (.A(WX8567), .B(RESET), .Z(WX8630) ) ;
DFF     gate2725  (.D(WX8630), .CP(CLK), .Q(WX8631) ) ;
AND2    gate2726  (.A(WX8569), .B(RESET), .Z(WX8632) ) ;
DFF     gate2727  (.D(WX8632), .CP(CLK), .Q(WX8633) ) ;
AND2    gate2728  (.A(WX8571), .B(RESET), .Z(WX8634) ) ;
DFF     gate2729  (.D(WX8634), .CP(CLK), .Q(WX8635) ) ;
AND2    gate2730  (.A(WX8573), .B(RESET), .Z(WX8636) ) ;
DFF     gate2731  (.D(WX8636), .CP(CLK), .Q(WX8637) ) ;
AND2    gate2732  (.A(WX8575), .B(RESET), .Z(WX8638) ) ;
DFF     gate2733  (.D(WX8638), .CP(CLK), .Q(WX8639) ) ;
AND2    gate2734  (.A(WX8577), .B(RESET), .Z(WX8640) ) ;
DFF     gate2735  (.D(WX8640), .CP(CLK), .Q(WX8641) ) ;
AND2    gate2736  (.A(WX8579), .B(RESET), .Z(WX8642) ) ;
DFF     gate2737  (.D(WX8642), .CP(CLK), .Q(WX8643) ) ;
AND2    gate2738  (.A(WX8581), .B(RESET), .Z(WX8644) ) ;
DFF     gate2739  (.D(WX8644), .CP(CLK), .Q(WX8645) ) ;
AND2    gate2740  (.A(WX8583), .B(RESET), .Z(WX8646) ) ;
DFF     gate2741  (.D(WX8646), .CP(CLK), .Q(WX8647) ) ;
AND2    gate2742  (.A(WX8585), .B(RESET), .Z(WX8648) ) ;
DFF     gate2743  (.D(WX8648), .CP(CLK), .Q(WX8649) ) ;
AND2    gate2744  (.A(WX8587), .B(RESET), .Z(WX8650) ) ;
DFF     gate2745  (.D(WX8650), .CP(CLK), .Q(WX8651) ) ;
AND2    gate2746  (.A(WX8589), .B(RESET), .Z(WX8652) ) ;
DFF     gate2747  (.D(WX8652), .CP(CLK), .Q(WX8653) ) ;
AND2    gate2748  (.A(WX8591), .B(RESET), .Z(WX8654) ) ;
DFF     gate2749  (.D(WX8654), .CP(CLK), .Q(WX8655) ) ;
AND2    gate2750  (.A(WX8593), .B(RESET), .Z(WX8656) ) ;
DFF     gate2751  (.D(WX8656), .CP(CLK), .Q(WX8657) ) ;
AND2    gate2752  (.A(WX8992), .B(WX9021), .Z(WX9022) ) ;
AND2    gate2753  (.A(WX9020), .B(WX9021), .Z(WX9024) ) ;
AND2    gate2754  (.A(WX9019), .B(WX9021), .Z(WX9026) ) ;
AND2    gate2755  (.A(WX9018), .B(WX9021), .Z(WX9028) ) ;
AND2    gate2756  (.A(WX8991), .B(WX9021), .Z(WX9030) ) ;
AND2    gate2757  (.A(WX9017), .B(WX9021), .Z(WX9032) ) ;
AND2    gate2758  (.A(WX9016), .B(WX9021), .Z(WX9034) ) ;
AND2    gate2759  (.A(WX9015), .B(WX9021), .Z(WX9036) ) ;
AND2    gate2760  (.A(WX9014), .B(WX9021), .Z(WX9038) ) ;
AND2    gate2761  (.A(WX9013), .B(WX9021), .Z(WX9040) ) ;
AND2    gate2762  (.A(WX9012), .B(WX9021), .Z(WX9042) ) ;
AND2    gate2763  (.A(WX8990), .B(WX9021), .Z(WX9044) ) ;
AND2    gate2764  (.A(WX9011), .B(WX9021), .Z(WX9046) ) ;
AND2    gate2765  (.A(WX9010), .B(WX9021), .Z(WX9048) ) ;
AND2    gate2766  (.A(WX9009), .B(WX9021), .Z(WX9050) ) ;
AND2    gate2767  (.A(WX9008), .B(WX9021), .Z(WX9052) ) ;
AND2    gate2768  (.A(WX8989), .B(WX9021), .Z(WX9054) ) ;
AND2    gate2769  (.A(WX9007), .B(WX9021), .Z(WX9056) ) ;
AND2    gate2770  (.A(WX9006), .B(WX9021), .Z(WX9058) ) ;
AND2    gate2771  (.A(WX9005), .B(WX9021), .Z(WX9060) ) ;
AND2    gate2772  (.A(WX9004), .B(WX9021), .Z(WX9062) ) ;
AND2    gate2773  (.A(WX9003), .B(WX9021), .Z(WX9064) ) ;
AND2    gate2774  (.A(WX9002), .B(WX9021), .Z(WX9066) ) ;
AND2    gate2775  (.A(WX9001), .B(WX9021), .Z(WX9068) ) ;
AND2    gate2776  (.A(WX9000), .B(WX9021), .Z(WX9070) ) ;
AND2    gate2777  (.A(WX8999), .B(WX9021), .Z(WX9072) ) ;
AND2    gate2778  (.A(WX8998), .B(WX9021), .Z(WX9074) ) ;
AND2    gate2779  (.A(WX8997), .B(WX9021), .Z(WX9076) ) ;
AND2    gate2780  (.A(WX8996), .B(WX9021), .Z(WX9078) ) ;
AND2    gate2781  (.A(WX8995), .B(WX9021), .Z(WX9080) ) ;
AND2    gate2782  (.A(WX8994), .B(WX9021), .Z(WX9082) ) ;
AND2    gate2783  (.A(WX8993), .B(WX9021), .Z(WX9084) ) ;
AND2    gate2784  (.A(WX9538), .B(RESET), .Z(WX9535) ) ;
DFF     gate2785  (.D(WX9535), .CP(CLK), .Q(WX9536) ) ;
AND2    gate2786  (.A(WX9540), .B(RESET), .Z(WX9537) ) ;
DFF     gate2787  (.D(WX9537), .CP(CLK), .Q(WX9538) ) ;
AND2    gate2788  (.A(WX9542), .B(RESET), .Z(WX9539) ) ;
DFF     gate2789  (.D(WX9539), .CP(CLK), .Q(WX9540) ) ;
AND2    gate2790  (.A(WX9544), .B(RESET), .Z(WX9541) ) ;
DFF     gate2791  (.D(WX9541), .CP(CLK), .Q(WX9542) ) ;
AND2    gate2792  (.A(WX9546), .B(RESET), .Z(WX9543) ) ;
DFF     gate2793  (.D(WX9543), .CP(CLK), .Q(WX9544) ) ;
AND2    gate2794  (.A(WX9548), .B(RESET), .Z(WX9545) ) ;
DFF     gate2795  (.D(WX9545), .CP(CLK), .Q(WX9546) ) ;
AND2    gate2796  (.A(WX9550), .B(RESET), .Z(WX9547) ) ;
DFF     gate2797  (.D(WX9547), .CP(CLK), .Q(WX9548) ) ;
AND2    gate2798  (.A(WX9552), .B(RESET), .Z(WX9549) ) ;
DFF     gate2799  (.D(WX9549), .CP(CLK), .Q(WX9550) ) ;
AND2    gate2800  (.A(WX9554), .B(RESET), .Z(WX9551) ) ;
DFF     gate2801  (.D(WX9551), .CP(CLK), .Q(WX9552) ) ;
AND2    gate2802  (.A(WX9556), .B(RESET), .Z(WX9553) ) ;
DFF     gate2803  (.D(WX9553), .CP(CLK), .Q(WX9554) ) ;
AND2    gate2804  (.A(WX9558), .B(RESET), .Z(WX9555) ) ;
DFF     gate2805  (.D(WX9555), .CP(CLK), .Q(WX9556) ) ;
AND2    gate2806  (.A(WX9560), .B(RESET), .Z(WX9557) ) ;
DFF     gate2807  (.D(WX9557), .CP(CLK), .Q(WX9558) ) ;
AND2    gate2808  (.A(WX9562), .B(RESET), .Z(WX9559) ) ;
DFF     gate2809  (.D(WX9559), .CP(CLK), .Q(WX9560) ) ;
AND2    gate2810  (.A(WX9564), .B(RESET), .Z(WX9561) ) ;
DFF     gate2811  (.D(WX9561), .CP(CLK), .Q(WX9562) ) ;
AND2    gate2812  (.A(WX9566), .B(RESET), .Z(WX9563) ) ;
DFF     gate2813  (.D(WX9563), .CP(CLK), .Q(WX9564) ) ;
AND2    gate2814  (.A(WX9568), .B(RESET), .Z(WX9565) ) ;
DFF     gate2815  (.D(WX9565), .CP(CLK), .Q(WX9566) ) ;
AND2    gate2816  (.A(WX9570), .B(RESET), .Z(WX9567) ) ;
DFF     gate2817  (.D(WX9567), .CP(CLK), .Q(WX9568) ) ;
AND2    gate2818  (.A(WX9572), .B(RESET), .Z(WX9569) ) ;
DFF     gate2819  (.D(WX9569), .CP(CLK), .Q(WX9570) ) ;
AND2    gate2820  (.A(WX9574), .B(RESET), .Z(WX9571) ) ;
DFF     gate2821  (.D(WX9571), .CP(CLK), .Q(WX9572) ) ;
AND2    gate2822  (.A(WX9576), .B(RESET), .Z(WX9573) ) ;
DFF     gate2823  (.D(WX9573), .CP(CLK), .Q(WX9574) ) ;
AND2    gate2824  (.A(WX9578), .B(RESET), .Z(WX9575) ) ;
DFF     gate2825  (.D(WX9575), .CP(CLK), .Q(WX9576) ) ;
AND2    gate2826  (.A(WX9580), .B(RESET), .Z(WX9577) ) ;
DFF     gate2827  (.D(WX9577), .CP(CLK), .Q(WX9578) ) ;
AND2    gate2828  (.A(WX9582), .B(RESET), .Z(WX9579) ) ;
DFF     gate2829  (.D(WX9579), .CP(CLK), .Q(WX9580) ) ;
AND2    gate2830  (.A(WX9584), .B(RESET), .Z(WX9581) ) ;
DFF     gate2831  (.D(WX9581), .CP(CLK), .Q(WX9582) ) ;
AND2    gate2832  (.A(WX9586), .B(RESET), .Z(WX9583) ) ;
DFF     gate2833  (.D(WX9583), .CP(CLK), .Q(WX9584) ) ;
AND2    gate2834  (.A(WX9588), .B(RESET), .Z(WX9585) ) ;
DFF     gate2835  (.D(WX9585), .CP(CLK), .Q(WX9586) ) ;
AND2    gate2836  (.A(WX9590), .B(RESET), .Z(WX9587) ) ;
DFF     gate2837  (.D(WX9587), .CP(CLK), .Q(WX9588) ) ;
AND2    gate2838  (.A(WX9592), .B(RESET), .Z(WX9589) ) ;
DFF     gate2839  (.D(WX9589), .CP(CLK), .Q(WX9590) ) ;
AND2    gate2840  (.A(WX9594), .B(RESET), .Z(WX9591) ) ;
DFF     gate2841  (.D(WX9591), .CP(CLK), .Q(WX9592) ) ;
AND2    gate2842  (.A(WX9596), .B(RESET), .Z(WX9593) ) ;
DFF     gate2843  (.D(WX9593), .CP(CLK), .Q(WX9594) ) ;
AND2    gate2844  (.A(WX9598), .B(RESET), .Z(WX9595) ) ;
DFF     gate2845  (.D(WX9595), .CP(CLK), .Q(WX9596) ) ;
AND2    gate2846  (.A(WX9534), .B(RESET), .Z(WX9597) ) ;
DFF     gate2847  (.D(WX9597), .CP(CLK), .Q(WX9598) ) ;
AND2    gate2848  (.A(WX9099), .B(RESET), .Z(WX9695) ) ;
DFF     gate2849  (.D(WX9695), .CP(CLK), .Q(WX9696) ) ;
AND2    gate2850  (.A(WX9113), .B(RESET), .Z(WX9697) ) ;
DFF     gate2851  (.D(WX9697), .CP(CLK), .Q(WX9698) ) ;
AND2    gate2852  (.A(WX9127), .B(RESET), .Z(WX9699) ) ;
DFF     gate2853  (.D(WX9699), .CP(CLK), .Q(WX9700) ) ;
AND2    gate2854  (.A(WX9141), .B(RESET), .Z(WX9701) ) ;
DFF     gate2855  (.D(WX9701), .CP(CLK), .Q(WX9702) ) ;
AND2    gate2856  (.A(WX9155), .B(RESET), .Z(WX9703) ) ;
DFF     gate2857  (.D(WX9703), .CP(CLK), .Q(WX9704) ) ;
AND2    gate2858  (.A(WX9169), .B(RESET), .Z(WX9705) ) ;
DFF     gate2859  (.D(WX9705), .CP(CLK), .Q(WX9706) ) ;
AND2    gate2860  (.A(WX9183), .B(RESET), .Z(WX9707) ) ;
DFF     gate2861  (.D(WX9707), .CP(CLK), .Q(WX9708) ) ;
AND2    gate2862  (.A(WX9197), .B(RESET), .Z(WX9709) ) ;
DFF     gate2863  (.D(WX9709), .CP(CLK), .Q(WX9710) ) ;
AND2    gate2864  (.A(WX9211), .B(RESET), .Z(WX9711) ) ;
DFF     gate2865  (.D(WX9711), .CP(CLK), .Q(WX9712) ) ;
AND2    gate2866  (.A(WX9225), .B(RESET), .Z(WX9713) ) ;
DFF     gate2867  (.D(WX9713), .CP(CLK), .Q(WX9714) ) ;
AND2    gate2868  (.A(WX9239), .B(RESET), .Z(WX9715) ) ;
DFF     gate2869  (.D(WX9715), .CP(CLK), .Q(WX9716) ) ;
AND2    gate2870  (.A(WX9253), .B(RESET), .Z(WX9717) ) ;
DFF     gate2871  (.D(WX9717), .CP(CLK), .Q(WX9718) ) ;
AND2    gate2872  (.A(WX9267), .B(RESET), .Z(WX9719) ) ;
DFF     gate2873  (.D(WX9719), .CP(CLK), .Q(WX9720) ) ;
AND2    gate2874  (.A(WX9281), .B(RESET), .Z(WX9721) ) ;
DFF     gate2875  (.D(WX9721), .CP(CLK), .Q(WX9722) ) ;
AND2    gate2876  (.A(WX9295), .B(RESET), .Z(WX9723) ) ;
DFF     gate2877  (.D(WX9723), .CP(CLK), .Q(WX9724) ) ;
AND2    gate2878  (.A(WX9309), .B(RESET), .Z(WX9725) ) ;
DFF     gate2879  (.D(WX9725), .CP(CLK), .Q(WX9726) ) ;
AND2    gate2880  (.A(WX9323), .B(RESET), .Z(WX9727) ) ;
DFF     gate2881  (.D(WX9727), .CP(CLK), .Q(WX9728) ) ;
AND2    gate2882  (.A(WX9337), .B(RESET), .Z(WX9729) ) ;
DFF     gate2883  (.D(WX9729), .CP(CLK), .Q(WX9730) ) ;
AND2    gate2884  (.A(WX9351), .B(RESET), .Z(WX9731) ) ;
DFF     gate2885  (.D(WX9731), .CP(CLK), .Q(WX9732) ) ;
AND2    gate2886  (.A(WX9365), .B(RESET), .Z(WX9733) ) ;
DFF     gate2887  (.D(WX9733), .CP(CLK), .Q(WX9734) ) ;
AND2    gate2888  (.A(WX9379), .B(RESET), .Z(WX9735) ) ;
DFF     gate2889  (.D(WX9735), .CP(CLK), .Q(WX9736) ) ;
AND2    gate2890  (.A(WX9393), .B(RESET), .Z(WX9737) ) ;
DFF     gate2891  (.D(WX9737), .CP(CLK), .Q(WX9738) ) ;
AND2    gate2892  (.A(WX9407), .B(RESET), .Z(WX9739) ) ;
DFF     gate2893  (.D(WX9739), .CP(CLK), .Q(WX9740) ) ;
AND2    gate2894  (.A(WX9421), .B(RESET), .Z(WX9741) ) ;
DFF     gate2895  (.D(WX9741), .CP(CLK), .Q(WX9742) ) ;
AND2    gate2896  (.A(WX9435), .B(RESET), .Z(WX9743) ) ;
DFF     gate2897  (.D(WX9743), .CP(CLK), .Q(WX9744) ) ;
AND2    gate2898  (.A(WX9449), .B(RESET), .Z(WX9745) ) ;
DFF     gate2899  (.D(WX9745), .CP(CLK), .Q(WX9746) ) ;
AND2    gate2900  (.A(WX9463), .B(RESET), .Z(WX9747) ) ;
DFF     gate2901  (.D(WX9747), .CP(CLK), .Q(WX9748) ) ;
AND2    gate2902  (.A(WX9477), .B(RESET), .Z(WX9749) ) ;
DFF     gate2903  (.D(WX9749), .CP(CLK), .Q(WX9750) ) ;
AND2    gate2904  (.A(WX9491), .B(RESET), .Z(WX9751) ) ;
DFF     gate2905  (.D(WX9751), .CP(CLK), .Q(WX9752) ) ;
AND2    gate2906  (.A(WX9505), .B(RESET), .Z(WX9753) ) ;
DFF     gate2907  (.D(WX9753), .CP(CLK), .Q(WX9754) ) ;
AND2    gate2908  (.A(WX9519), .B(RESET), .Z(WX9755) ) ;
DFF     gate2909  (.D(WX9755), .CP(CLK), .Q(WX9756) ) ;
AND2    gate2910  (.A(WX9533), .B(RESET), .Z(WX9757) ) ;
DFF     gate2911  (.D(WX9757), .CP(CLK), .Q(WX9758) ) ;
AND2    gate2912  (.A(WX9696), .B(RESET), .Z(WX9759) ) ;
DFF     gate2913  (.D(WX9759), .CP(CLK), .Q(WX9760) ) ;
AND2    gate2914  (.A(WX9698), .B(RESET), .Z(WX9761) ) ;
DFF     gate2915  (.D(WX9761), .CP(CLK), .Q(WX9762) ) ;
AND2    gate2916  (.A(WX9700), .B(RESET), .Z(WX9763) ) ;
DFF     gate2917  (.D(WX9763), .CP(CLK), .Q(WX9764) ) ;
AND2    gate2918  (.A(WX9702), .B(RESET), .Z(WX9765) ) ;
DFF     gate2919  (.D(WX9765), .CP(CLK), .Q(WX9766) ) ;
AND2    gate2920  (.A(WX9704), .B(RESET), .Z(WX9767) ) ;
DFF     gate2921  (.D(WX9767), .CP(CLK), .Q(WX9768) ) ;
AND2    gate2922  (.A(WX9706), .B(RESET), .Z(WX9769) ) ;
DFF     gate2923  (.D(WX9769), .CP(CLK), .Q(WX9770) ) ;
AND2    gate2924  (.A(WX9708), .B(RESET), .Z(WX9771) ) ;
DFF     gate2925  (.D(WX9771), .CP(CLK), .Q(WX9772) ) ;
AND2    gate2926  (.A(WX9710), .B(RESET), .Z(WX9773) ) ;
DFF     gate2927  (.D(WX9773), .CP(CLK), .Q(WX9774) ) ;
AND2    gate2928  (.A(WX9712), .B(RESET), .Z(WX9775) ) ;
DFF     gate2929  (.D(WX9775), .CP(CLK), .Q(WX9776) ) ;
AND2    gate2930  (.A(WX9714), .B(RESET), .Z(WX9777) ) ;
DFF     gate2931  (.D(WX9777), .CP(CLK), .Q(WX9778) ) ;
AND2    gate2932  (.A(WX9716), .B(RESET), .Z(WX9779) ) ;
DFF     gate2933  (.D(WX9779), .CP(CLK), .Q(WX9780) ) ;
AND2    gate2934  (.A(WX9718), .B(RESET), .Z(WX9781) ) ;
DFF     gate2935  (.D(WX9781), .CP(CLK), .Q(WX9782) ) ;
AND2    gate2936  (.A(WX9720), .B(RESET), .Z(WX9783) ) ;
DFF     gate2937  (.D(WX9783), .CP(CLK), .Q(WX9784) ) ;
AND2    gate2938  (.A(WX9722), .B(RESET), .Z(WX9785) ) ;
DFF     gate2939  (.D(WX9785), .CP(CLK), .Q(WX9786) ) ;
AND2    gate2940  (.A(WX9724), .B(RESET), .Z(WX9787) ) ;
DFF     gate2941  (.D(WX9787), .CP(CLK), .Q(WX9788) ) ;
AND2    gate2942  (.A(WX9726), .B(RESET), .Z(WX9789) ) ;
DFF     gate2943  (.D(WX9789), .CP(CLK), .Q(WX9790) ) ;
AND2    gate2944  (.A(WX9728), .B(RESET), .Z(WX9791) ) ;
DFF     gate2945  (.D(WX9791), .CP(CLK), .Q(WX9792) ) ;
AND2    gate2946  (.A(WX9730), .B(RESET), .Z(WX9793) ) ;
DFF     gate2947  (.D(WX9793), .CP(CLK), .Q(WX9794) ) ;
AND2    gate2948  (.A(WX9732), .B(RESET), .Z(WX9795) ) ;
DFF     gate2949  (.D(WX9795), .CP(CLK), .Q(WX9796) ) ;
AND2    gate2950  (.A(WX9734), .B(RESET), .Z(WX9797) ) ;
DFF     gate2951  (.D(WX9797), .CP(CLK), .Q(WX9798) ) ;
AND2    gate2952  (.A(WX9736), .B(RESET), .Z(WX9799) ) ;
DFF     gate2953  (.D(WX9799), .CP(CLK), .Q(WX9800) ) ;
AND2    gate2954  (.A(WX9738), .B(RESET), .Z(WX9801) ) ;
DFF     gate2955  (.D(WX9801), .CP(CLK), .Q(WX9802) ) ;
AND2    gate2956  (.A(WX9740), .B(RESET), .Z(WX9803) ) ;
DFF     gate2957  (.D(WX9803), .CP(CLK), .Q(WX9804) ) ;
AND2    gate2958  (.A(WX9742), .B(RESET), .Z(WX9805) ) ;
DFF     gate2959  (.D(WX9805), .CP(CLK), .Q(WX9806) ) ;
AND2    gate2960  (.A(WX9744), .B(RESET), .Z(WX9807) ) ;
DFF     gate2961  (.D(WX9807), .CP(CLK), .Q(WX9808) ) ;
AND2    gate2962  (.A(WX9746), .B(RESET), .Z(WX9809) ) ;
DFF     gate2963  (.D(WX9809), .CP(CLK), .Q(WX9810) ) ;
AND2    gate2964  (.A(WX9748), .B(RESET), .Z(WX9811) ) ;
DFF     gate2965  (.D(WX9811), .CP(CLK), .Q(WX9812) ) ;
AND2    gate2966  (.A(WX9750), .B(RESET), .Z(WX9813) ) ;
DFF     gate2967  (.D(WX9813), .CP(CLK), .Q(WX9814) ) ;
AND2    gate2968  (.A(WX9752), .B(RESET), .Z(WX9815) ) ;
DFF     gate2969  (.D(WX9815), .CP(CLK), .Q(WX9816) ) ;
AND2    gate2970  (.A(WX9754), .B(RESET), .Z(WX9817) ) ;
DFF     gate2971  (.D(WX9817), .CP(CLK), .Q(WX9818) ) ;
AND2    gate2972  (.A(WX9756), .B(RESET), .Z(WX9819) ) ;
DFF     gate2973  (.D(WX9819), .CP(CLK), .Q(WX9820) ) ;
AND2    gate2974  (.A(WX9758), .B(RESET), .Z(WX9821) ) ;
DFF     gate2975  (.D(WX9821), .CP(CLK), .Q(WX9822) ) ;
AND2    gate2976  (.A(WX9760), .B(RESET), .Z(WX9823) ) ;
DFF     gate2977  (.D(WX9823), .CP(CLK), .Q(WX9824) ) ;
AND2    gate2978  (.A(WX9762), .B(RESET), .Z(WX9825) ) ;
DFF     gate2979  (.D(WX9825), .CP(CLK), .Q(WX9826) ) ;
AND2    gate2980  (.A(WX9764), .B(RESET), .Z(WX9827) ) ;
DFF     gate2981  (.D(WX9827), .CP(CLK), .Q(WX9828) ) ;
AND2    gate2982  (.A(WX9766), .B(RESET), .Z(WX9829) ) ;
DFF     gate2983  (.D(WX9829), .CP(CLK), .Q(WX9830) ) ;
AND2    gate2984  (.A(WX9768), .B(RESET), .Z(WX9831) ) ;
DFF     gate2985  (.D(WX9831), .CP(CLK), .Q(WX9832) ) ;
AND2    gate2986  (.A(WX9770), .B(RESET), .Z(WX9833) ) ;
DFF     gate2987  (.D(WX9833), .CP(CLK), .Q(WX9834) ) ;
AND2    gate2988  (.A(WX9772), .B(RESET), .Z(WX9835) ) ;
DFF     gate2989  (.D(WX9835), .CP(CLK), .Q(WX9836) ) ;
AND2    gate2990  (.A(WX9774), .B(RESET), .Z(WX9837) ) ;
DFF     gate2991  (.D(WX9837), .CP(CLK), .Q(WX9838) ) ;
AND2    gate2992  (.A(WX9776), .B(RESET), .Z(WX9839) ) ;
DFF     gate2993  (.D(WX9839), .CP(CLK), .Q(WX9840) ) ;
AND2    gate2994  (.A(WX9778), .B(RESET), .Z(WX9841) ) ;
DFF     gate2995  (.D(WX9841), .CP(CLK), .Q(WX9842) ) ;
AND2    gate2996  (.A(WX9780), .B(RESET), .Z(WX9843) ) ;
DFF     gate2997  (.D(WX9843), .CP(CLK), .Q(WX9844) ) ;
AND2    gate2998  (.A(WX9782), .B(RESET), .Z(WX9845) ) ;
DFF     gate2999  (.D(WX9845), .CP(CLK), .Q(WX9846) ) ;
AND2    gate3000  (.A(WX9784), .B(RESET), .Z(WX9847) ) ;
DFF     gate3001  (.D(WX9847), .CP(CLK), .Q(WX9848) ) ;
AND2    gate3002  (.A(WX9786), .B(RESET), .Z(WX9849) ) ;
DFF     gate3003  (.D(WX9849), .CP(CLK), .Q(WX9850) ) ;
AND2    gate3004  (.A(WX9788), .B(RESET), .Z(WX9851) ) ;
DFF     gate3005  (.D(WX9851), .CP(CLK), .Q(WX9852) ) ;
AND2    gate3006  (.A(WX9790), .B(RESET), .Z(WX9853) ) ;
DFF     gate3007  (.D(WX9853), .CP(CLK), .Q(WX9854) ) ;
AND2    gate3008  (.A(WX9792), .B(RESET), .Z(WX9855) ) ;
DFF     gate3009  (.D(WX9855), .CP(CLK), .Q(WX9856) ) ;
AND2    gate3010  (.A(WX9794), .B(RESET), .Z(WX9857) ) ;
DFF     gate3011  (.D(WX9857), .CP(CLK), .Q(WX9858) ) ;
AND2    gate3012  (.A(WX9796), .B(RESET), .Z(WX9859) ) ;
DFF     gate3013  (.D(WX9859), .CP(CLK), .Q(WX9860) ) ;
AND2    gate3014  (.A(WX9798), .B(RESET), .Z(WX9861) ) ;
DFF     gate3015  (.D(WX9861), .CP(CLK), .Q(WX9862) ) ;
AND2    gate3016  (.A(WX9800), .B(RESET), .Z(WX9863) ) ;
DFF     gate3017  (.D(WX9863), .CP(CLK), .Q(WX9864) ) ;
AND2    gate3018  (.A(WX9802), .B(RESET), .Z(WX9865) ) ;
DFF     gate3019  (.D(WX9865), .CP(CLK), .Q(WX9866) ) ;
AND2    gate3020  (.A(WX9804), .B(RESET), .Z(WX9867) ) ;
DFF     gate3021  (.D(WX9867), .CP(CLK), .Q(WX9868) ) ;
AND2    gate3022  (.A(WX9806), .B(RESET), .Z(WX9869) ) ;
DFF     gate3023  (.D(WX9869), .CP(CLK), .Q(WX9870) ) ;
AND2    gate3024  (.A(WX9808), .B(RESET), .Z(WX9871) ) ;
DFF     gate3025  (.D(WX9871), .CP(CLK), .Q(WX9872) ) ;
AND2    gate3026  (.A(WX9810), .B(RESET), .Z(WX9873) ) ;
DFF     gate3027  (.D(WX9873), .CP(CLK), .Q(WX9874) ) ;
AND2    gate3028  (.A(WX9812), .B(RESET), .Z(WX9875) ) ;
DFF     gate3029  (.D(WX9875), .CP(CLK), .Q(WX9876) ) ;
AND2    gate3030  (.A(WX9814), .B(RESET), .Z(WX9877) ) ;
DFF     gate3031  (.D(WX9877), .CP(CLK), .Q(WX9878) ) ;
AND2    gate3032  (.A(WX9816), .B(RESET), .Z(WX9879) ) ;
DFF     gate3033  (.D(WX9879), .CP(CLK), .Q(WX9880) ) ;
AND2    gate3034  (.A(WX9818), .B(RESET), .Z(WX9881) ) ;
DFF     gate3035  (.D(WX9881), .CP(CLK), .Q(WX9882) ) ;
AND2    gate3036  (.A(WX9820), .B(RESET), .Z(WX9883) ) ;
DFF     gate3037  (.D(WX9883), .CP(CLK), .Q(WX9884) ) ;
AND2    gate3038  (.A(WX9822), .B(RESET), .Z(WX9885) ) ;
DFF     gate3039  (.D(WX9885), .CP(CLK), .Q(WX9886) ) ;
AND2    gate3040  (.A(WX9824), .B(RESET), .Z(WX9887) ) ;
DFF     gate3041  (.D(WX9887), .CP(CLK), .Q(WX9888) ) ;
AND2    gate3042  (.A(WX9826), .B(RESET), .Z(WX9889) ) ;
DFF     gate3043  (.D(WX9889), .CP(CLK), .Q(WX9890) ) ;
AND2    gate3044  (.A(WX9828), .B(RESET), .Z(WX9891) ) ;
DFF     gate3045  (.D(WX9891), .CP(CLK), .Q(WX9892) ) ;
AND2    gate3046  (.A(WX9830), .B(RESET), .Z(WX9893) ) ;
DFF     gate3047  (.D(WX9893), .CP(CLK), .Q(WX9894) ) ;
AND2    gate3048  (.A(WX9832), .B(RESET), .Z(WX9895) ) ;
DFF     gate3049  (.D(WX9895), .CP(CLK), .Q(WX9896) ) ;
AND2    gate3050  (.A(WX9834), .B(RESET), .Z(WX9897) ) ;
DFF     gate3051  (.D(WX9897), .CP(CLK), .Q(WX9898) ) ;
AND2    gate3052  (.A(WX9836), .B(RESET), .Z(WX9899) ) ;
DFF     gate3053  (.D(WX9899), .CP(CLK), .Q(WX9900) ) ;
AND2    gate3054  (.A(WX9838), .B(RESET), .Z(WX9901) ) ;
DFF     gate3055  (.D(WX9901), .CP(CLK), .Q(WX9902) ) ;
AND2    gate3056  (.A(WX9840), .B(RESET), .Z(WX9903) ) ;
DFF     gate3057  (.D(WX9903), .CP(CLK), .Q(WX9904) ) ;
AND2    gate3058  (.A(WX9842), .B(RESET), .Z(WX9905) ) ;
DFF     gate3059  (.D(WX9905), .CP(CLK), .Q(WX9906) ) ;
AND2    gate3060  (.A(WX9844), .B(RESET), .Z(WX9907) ) ;
DFF     gate3061  (.D(WX9907), .CP(CLK), .Q(WX9908) ) ;
AND2    gate3062  (.A(WX9846), .B(RESET), .Z(WX9909) ) ;
DFF     gate3063  (.D(WX9909), .CP(CLK), .Q(WX9910) ) ;
AND2    gate3064  (.A(WX9848), .B(RESET), .Z(WX9911) ) ;
DFF     gate3065  (.D(WX9911), .CP(CLK), .Q(WX9912) ) ;
AND2    gate3066  (.A(WX9850), .B(RESET), .Z(WX9913) ) ;
DFF     gate3067  (.D(WX9913), .CP(CLK), .Q(WX9914) ) ;
AND2    gate3068  (.A(WX9852), .B(RESET), .Z(WX9915) ) ;
DFF     gate3069  (.D(WX9915), .CP(CLK), .Q(WX9916) ) ;
AND2    gate3070  (.A(WX9854), .B(RESET), .Z(WX9917) ) ;
DFF     gate3071  (.D(WX9917), .CP(CLK), .Q(WX9918) ) ;
AND2    gate3072  (.A(WX9856), .B(RESET), .Z(WX9919) ) ;
DFF     gate3073  (.D(WX9919), .CP(CLK), .Q(WX9920) ) ;
AND2    gate3074  (.A(WX9858), .B(RESET), .Z(WX9921) ) ;
DFF     gate3075  (.D(WX9921), .CP(CLK), .Q(WX9922) ) ;
AND2    gate3076  (.A(WX9860), .B(RESET), .Z(WX9923) ) ;
DFF     gate3077  (.D(WX9923), .CP(CLK), .Q(WX9924) ) ;
AND2    gate3078  (.A(WX9862), .B(RESET), .Z(WX9925) ) ;
DFF     gate3079  (.D(WX9925), .CP(CLK), .Q(WX9926) ) ;
AND2    gate3080  (.A(WX9864), .B(RESET), .Z(WX9927) ) ;
DFF     gate3081  (.D(WX9927), .CP(CLK), .Q(WX9928) ) ;
AND2    gate3082  (.A(WX9866), .B(RESET), .Z(WX9929) ) ;
DFF     gate3083  (.D(WX9929), .CP(CLK), .Q(WX9930) ) ;
AND2    gate3084  (.A(WX9868), .B(RESET), .Z(WX9931) ) ;
DFF     gate3085  (.D(WX9931), .CP(CLK), .Q(WX9932) ) ;
AND2    gate3086  (.A(WX9870), .B(RESET), .Z(WX9933) ) ;
DFF     gate3087  (.D(WX9933), .CP(CLK), .Q(WX9934) ) ;
AND2    gate3088  (.A(WX9872), .B(RESET), .Z(WX9935) ) ;
DFF     gate3089  (.D(WX9935), .CP(CLK), .Q(WX9936) ) ;
AND2    gate3090  (.A(WX9874), .B(RESET), .Z(WX9937) ) ;
DFF     gate3091  (.D(WX9937), .CP(CLK), .Q(WX9938) ) ;
AND2    gate3092  (.A(WX9876), .B(RESET), .Z(WX9939) ) ;
DFF     gate3093  (.D(WX9939), .CP(CLK), .Q(WX9940) ) ;
AND2    gate3094  (.A(WX9878), .B(RESET), .Z(WX9941) ) ;
DFF     gate3095  (.D(WX9941), .CP(CLK), .Q(WX9942) ) ;
AND2    gate3096  (.A(WX9880), .B(RESET), .Z(WX9943) ) ;
DFF     gate3097  (.D(WX9943), .CP(CLK), .Q(WX9944) ) ;
AND2    gate3098  (.A(WX9882), .B(RESET), .Z(WX9945) ) ;
DFF     gate3099  (.D(WX9945), .CP(CLK), .Q(WX9946) ) ;
AND2    gate3100  (.A(WX9884), .B(RESET), .Z(WX9947) ) ;
DFF     gate3101  (.D(WX9947), .CP(CLK), .Q(WX9948) ) ;
AND2    gate3102  (.A(WX9886), .B(RESET), .Z(WX9949) ) ;
DFF     gate3103  (.D(WX9949), .CP(CLK), .Q(WX9950) ) ;
AND2    gate3104  (.A(WX10285), .B(WX10314), .Z(WX10315) ) ;
AND2    gate3105  (.A(WX10313), .B(WX10314), .Z(WX10317) ) ;
AND2    gate3106  (.A(WX10312), .B(WX10314), .Z(WX10319) ) ;
AND2    gate3107  (.A(WX10311), .B(WX10314), .Z(WX10321) ) ;
AND2    gate3108  (.A(WX10284), .B(WX10314), .Z(WX10323) ) ;
AND2    gate3109  (.A(WX10310), .B(WX10314), .Z(WX10325) ) ;
AND2    gate3110  (.A(WX10309), .B(WX10314), .Z(WX10327) ) ;
AND2    gate3111  (.A(WX10308), .B(WX10314), .Z(WX10329) ) ;
AND2    gate3112  (.A(WX10307), .B(WX10314), .Z(WX10331) ) ;
AND2    gate3113  (.A(WX10306), .B(WX10314), .Z(WX10333) ) ;
AND2    gate3114  (.A(WX10305), .B(WX10314), .Z(WX10335) ) ;
AND2    gate3115  (.A(WX10283), .B(WX10314), .Z(WX10337) ) ;
AND2    gate3116  (.A(WX10304), .B(WX10314), .Z(WX10339) ) ;
AND2    gate3117  (.A(WX10303), .B(WX10314), .Z(WX10341) ) ;
AND2    gate3118  (.A(WX10302), .B(WX10314), .Z(WX10343) ) ;
AND2    gate3119  (.A(WX10301), .B(WX10314), .Z(WX10345) ) ;
AND2    gate3120  (.A(WX10282), .B(WX10314), .Z(WX10347) ) ;
AND2    gate3121  (.A(WX10300), .B(WX10314), .Z(WX10349) ) ;
AND2    gate3122  (.A(WX10299), .B(WX10314), .Z(WX10351) ) ;
AND2    gate3123  (.A(WX10298), .B(WX10314), .Z(WX10353) ) ;
AND2    gate3124  (.A(WX10297), .B(WX10314), .Z(WX10355) ) ;
AND2    gate3125  (.A(WX10296), .B(WX10314), .Z(WX10357) ) ;
AND2    gate3126  (.A(WX10295), .B(WX10314), .Z(WX10359) ) ;
AND2    gate3127  (.A(WX10294), .B(WX10314), .Z(WX10361) ) ;
AND2    gate3128  (.A(WX10293), .B(WX10314), .Z(WX10363) ) ;
AND2    gate3129  (.A(WX10292), .B(WX10314), .Z(WX10365) ) ;
AND2    gate3130  (.A(WX10291), .B(WX10314), .Z(WX10367) ) ;
AND2    gate3131  (.A(WX10290), .B(WX10314), .Z(WX10369) ) ;
AND2    gate3132  (.A(WX10289), .B(WX10314), .Z(WX10371) ) ;
AND2    gate3133  (.A(WX10288), .B(WX10314), .Z(WX10373) ) ;
AND2    gate3134  (.A(WX10287), .B(WX10314), .Z(WX10375) ) ;
AND2    gate3135  (.A(WX10286), .B(WX10314), .Z(WX10377) ) ;
AND2    gate3136  (.A(WX10831), .B(RESET), .Z(WX10828) ) ;
DFF     gate3137  (.D(WX10828), .CP(CLK), .Q(WX10829) ) ;
AND2    gate3138  (.A(WX10833), .B(RESET), .Z(WX10830) ) ;
DFF     gate3139  (.D(WX10830), .CP(CLK), .Q(WX10831) ) ;
AND2    gate3140  (.A(WX10835), .B(RESET), .Z(WX10832) ) ;
DFF     gate3141  (.D(WX10832), .CP(CLK), .Q(WX10833) ) ;
AND2    gate3142  (.A(WX10837), .B(RESET), .Z(WX10834) ) ;
DFF     gate3143  (.D(WX10834), .CP(CLK), .Q(WX10835) ) ;
AND2    gate3144  (.A(WX10839), .B(RESET), .Z(WX10836) ) ;
DFF     gate3145  (.D(WX10836), .CP(CLK), .Q(WX10837) ) ;
AND2    gate3146  (.A(WX10841), .B(RESET), .Z(WX10838) ) ;
DFF     gate3147  (.D(WX10838), .CP(CLK), .Q(WX10839) ) ;
AND2    gate3148  (.A(WX10843), .B(RESET), .Z(WX10840) ) ;
DFF     gate3149  (.D(WX10840), .CP(CLK), .Q(WX10841) ) ;
AND2    gate3150  (.A(WX10845), .B(RESET), .Z(WX10842) ) ;
DFF     gate3151  (.D(WX10842), .CP(CLK), .Q(WX10843) ) ;
AND2    gate3152  (.A(WX10847), .B(RESET), .Z(WX10844) ) ;
DFF     gate3153  (.D(WX10844), .CP(CLK), .Q(WX10845) ) ;
AND2    gate3154  (.A(WX10849), .B(RESET), .Z(WX10846) ) ;
DFF     gate3155  (.D(WX10846), .CP(CLK), .Q(WX10847) ) ;
AND2    gate3156  (.A(WX10851), .B(RESET), .Z(WX10848) ) ;
DFF     gate3157  (.D(WX10848), .CP(CLK), .Q(WX10849) ) ;
AND2    gate3158  (.A(WX10853), .B(RESET), .Z(WX10850) ) ;
DFF     gate3159  (.D(WX10850), .CP(CLK), .Q(WX10851) ) ;
AND2    gate3160  (.A(WX10855), .B(RESET), .Z(WX10852) ) ;
DFF     gate3161  (.D(WX10852), .CP(CLK), .Q(WX10853) ) ;
AND2    gate3162  (.A(WX10857), .B(RESET), .Z(WX10854) ) ;
DFF     gate3163  (.D(WX10854), .CP(CLK), .Q(WX10855) ) ;
AND2    gate3164  (.A(WX10859), .B(RESET), .Z(WX10856) ) ;
DFF     gate3165  (.D(WX10856), .CP(CLK), .Q(WX10857) ) ;
AND2    gate3166  (.A(WX10861), .B(RESET), .Z(WX10858) ) ;
DFF     gate3167  (.D(WX10858), .CP(CLK), .Q(WX10859) ) ;
AND2    gate3168  (.A(WX10863), .B(RESET), .Z(WX10860) ) ;
DFF     gate3169  (.D(WX10860), .CP(CLK), .Q(WX10861) ) ;
AND2    gate3170  (.A(WX10865), .B(RESET), .Z(WX10862) ) ;
DFF     gate3171  (.D(WX10862), .CP(CLK), .Q(WX10863) ) ;
AND2    gate3172  (.A(WX10867), .B(RESET), .Z(WX10864) ) ;
DFF     gate3173  (.D(WX10864), .CP(CLK), .Q(WX10865) ) ;
AND2    gate3174  (.A(WX10869), .B(RESET), .Z(WX10866) ) ;
DFF     gate3175  (.D(WX10866), .CP(CLK), .Q(WX10867) ) ;
AND2    gate3176  (.A(WX10871), .B(RESET), .Z(WX10868) ) ;
DFF     gate3177  (.D(WX10868), .CP(CLK), .Q(WX10869) ) ;
AND2    gate3178  (.A(WX10873), .B(RESET), .Z(WX10870) ) ;
DFF     gate3179  (.D(WX10870), .CP(CLK), .Q(WX10871) ) ;
AND2    gate3180  (.A(WX10875), .B(RESET), .Z(WX10872) ) ;
DFF     gate3181  (.D(WX10872), .CP(CLK), .Q(WX10873) ) ;
AND2    gate3182  (.A(WX10877), .B(RESET), .Z(WX10874) ) ;
DFF     gate3183  (.D(WX10874), .CP(CLK), .Q(WX10875) ) ;
AND2    gate3184  (.A(WX10879), .B(RESET), .Z(WX10876) ) ;
DFF     gate3185  (.D(WX10876), .CP(CLK), .Q(WX10877) ) ;
AND2    gate3186  (.A(WX10881), .B(RESET), .Z(WX10878) ) ;
DFF     gate3187  (.D(WX10878), .CP(CLK), .Q(WX10879) ) ;
AND2    gate3188  (.A(WX10883), .B(RESET), .Z(WX10880) ) ;
DFF     gate3189  (.D(WX10880), .CP(CLK), .Q(WX10881) ) ;
AND2    gate3190  (.A(WX10885), .B(RESET), .Z(WX10882) ) ;
DFF     gate3191  (.D(WX10882), .CP(CLK), .Q(WX10883) ) ;
AND2    gate3192  (.A(WX10887), .B(RESET), .Z(WX10884) ) ;
DFF     gate3193  (.D(WX10884), .CP(CLK), .Q(WX10885) ) ;
AND2    gate3194  (.A(WX10889), .B(RESET), .Z(WX10886) ) ;
DFF     gate3195  (.D(WX10886), .CP(CLK), .Q(WX10887) ) ;
AND2    gate3196  (.A(WX10891), .B(RESET), .Z(WX10888) ) ;
DFF     gate3197  (.D(WX10888), .CP(CLK), .Q(WX10889) ) ;
AND2    gate3198  (.A(WX10827), .B(RESET), .Z(WX10890) ) ;
DFF     gate3199  (.D(WX10890), .CP(CLK), .Q(WX10891) ) ;
AND2    gate3200  (.A(WX10392), .B(RESET), .Z(WX10988) ) ;
DFF     gate3201  (.D(WX10988), .CP(CLK), .Q(WX10989) ) ;
AND2    gate3202  (.A(WX10406), .B(RESET), .Z(WX10990) ) ;
DFF     gate3203  (.D(WX10990), .CP(CLK), .Q(WX10991) ) ;
AND2    gate3204  (.A(WX10420), .B(RESET), .Z(WX10992) ) ;
DFF     gate3205  (.D(WX10992), .CP(CLK), .Q(WX10993) ) ;
AND2    gate3206  (.A(WX10434), .B(RESET), .Z(WX10994) ) ;
DFF     gate3207  (.D(WX10994), .CP(CLK), .Q(WX10995) ) ;
AND2    gate3208  (.A(WX10448), .B(RESET), .Z(WX10996) ) ;
DFF     gate3209  (.D(WX10996), .CP(CLK), .Q(WX10997) ) ;
AND2    gate3210  (.A(WX10462), .B(RESET), .Z(WX10998) ) ;
DFF     gate3211  (.D(WX10998), .CP(CLK), .Q(WX10999) ) ;
AND2    gate3212  (.A(WX10476), .B(RESET), .Z(WX11000) ) ;
DFF     gate3213  (.D(WX11000), .CP(CLK), .Q(WX11001) ) ;
AND2    gate3214  (.A(WX10490), .B(RESET), .Z(WX11002) ) ;
DFF     gate3215  (.D(WX11002), .CP(CLK), .Q(WX11003) ) ;
AND2    gate3216  (.A(WX10504), .B(RESET), .Z(WX11004) ) ;
DFF     gate3217  (.D(WX11004), .CP(CLK), .Q(WX11005) ) ;
AND2    gate3218  (.A(WX10518), .B(RESET), .Z(WX11006) ) ;
DFF     gate3219  (.D(WX11006), .CP(CLK), .Q(WX11007) ) ;
AND2    gate3220  (.A(WX10532), .B(RESET), .Z(WX11008) ) ;
DFF     gate3221  (.D(WX11008), .CP(CLK), .Q(WX11009) ) ;
AND2    gate3222  (.A(WX10546), .B(RESET), .Z(WX11010) ) ;
DFF     gate3223  (.D(WX11010), .CP(CLK), .Q(WX11011) ) ;
AND2    gate3224  (.A(WX10560), .B(RESET), .Z(WX11012) ) ;
DFF     gate3225  (.D(WX11012), .CP(CLK), .Q(WX11013) ) ;
AND2    gate3226  (.A(WX10574), .B(RESET), .Z(WX11014) ) ;
DFF     gate3227  (.D(WX11014), .CP(CLK), .Q(WX11015) ) ;
AND2    gate3228  (.A(WX10588), .B(RESET), .Z(WX11016) ) ;
DFF     gate3229  (.D(WX11016), .CP(CLK), .Q(WX11017) ) ;
AND2    gate3230  (.A(WX10602), .B(RESET), .Z(WX11018) ) ;
DFF     gate3231  (.D(WX11018), .CP(CLK), .Q(WX11019) ) ;
AND2    gate3232  (.A(WX10616), .B(RESET), .Z(WX11020) ) ;
DFF     gate3233  (.D(WX11020), .CP(CLK), .Q(WX11021) ) ;
AND2    gate3234  (.A(WX10630), .B(RESET), .Z(WX11022) ) ;
DFF     gate3235  (.D(WX11022), .CP(CLK), .Q(WX11023) ) ;
AND2    gate3236  (.A(WX10644), .B(RESET), .Z(WX11024) ) ;
DFF     gate3237  (.D(WX11024), .CP(CLK), .Q(WX11025) ) ;
AND2    gate3238  (.A(WX10658), .B(RESET), .Z(WX11026) ) ;
DFF     gate3239  (.D(WX11026), .CP(CLK), .Q(WX11027) ) ;
AND2    gate3240  (.A(WX10672), .B(RESET), .Z(WX11028) ) ;
DFF     gate3241  (.D(WX11028), .CP(CLK), .Q(WX11029) ) ;
AND2    gate3242  (.A(WX10686), .B(RESET), .Z(WX11030) ) ;
DFF     gate3243  (.D(WX11030), .CP(CLK), .Q(WX11031) ) ;
AND2    gate3244  (.A(WX10700), .B(RESET), .Z(WX11032) ) ;
DFF     gate3245  (.D(WX11032), .CP(CLK), .Q(WX11033) ) ;
AND2    gate3246  (.A(WX10714), .B(RESET), .Z(WX11034) ) ;
DFF     gate3247  (.D(WX11034), .CP(CLK), .Q(WX11035) ) ;
AND2    gate3248  (.A(WX10728), .B(RESET), .Z(WX11036) ) ;
DFF     gate3249  (.D(WX11036), .CP(CLK), .Q(WX11037) ) ;
AND2    gate3250  (.A(WX10742), .B(RESET), .Z(WX11038) ) ;
DFF     gate3251  (.D(WX11038), .CP(CLK), .Q(WX11039) ) ;
AND2    gate3252  (.A(WX10756), .B(RESET), .Z(WX11040) ) ;
DFF     gate3253  (.D(WX11040), .CP(CLK), .Q(WX11041) ) ;
AND2    gate3254  (.A(WX10770), .B(RESET), .Z(WX11042) ) ;
DFF     gate3255  (.D(WX11042), .CP(CLK), .Q(WX11043) ) ;
AND2    gate3256  (.A(WX10784), .B(RESET), .Z(WX11044) ) ;
DFF     gate3257  (.D(WX11044), .CP(CLK), .Q(WX11045) ) ;
AND2    gate3258  (.A(WX10798), .B(RESET), .Z(WX11046) ) ;
DFF     gate3259  (.D(WX11046), .CP(CLK), .Q(WX11047) ) ;
AND2    gate3260  (.A(WX10812), .B(RESET), .Z(WX11048) ) ;
DFF     gate3261  (.D(WX11048), .CP(CLK), .Q(WX11049) ) ;
AND2    gate3262  (.A(WX10826), .B(RESET), .Z(WX11050) ) ;
DFF     gate3263  (.D(WX11050), .CP(CLK), .Q(WX11051) ) ;
AND2    gate3264  (.A(WX10989), .B(RESET), .Z(WX11052) ) ;
DFF     gate3265  (.D(WX11052), .CP(CLK), .Q(WX11053) ) ;
AND2    gate3266  (.A(WX10991), .B(RESET), .Z(WX11054) ) ;
DFF     gate3267  (.D(WX11054), .CP(CLK), .Q(WX11055) ) ;
AND2    gate3268  (.A(WX10993), .B(RESET), .Z(WX11056) ) ;
DFF     gate3269  (.D(WX11056), .CP(CLK), .Q(WX11057) ) ;
AND2    gate3270  (.A(WX10995), .B(RESET), .Z(WX11058) ) ;
DFF     gate3271  (.D(WX11058), .CP(CLK), .Q(WX11059) ) ;
AND2    gate3272  (.A(WX10997), .B(RESET), .Z(WX11060) ) ;
DFF     gate3273  (.D(WX11060), .CP(CLK), .Q(WX11061) ) ;
AND2    gate3274  (.A(WX10999), .B(RESET), .Z(WX11062) ) ;
DFF     gate3275  (.D(WX11062), .CP(CLK), .Q(WX11063) ) ;
AND2    gate3276  (.A(WX11001), .B(RESET), .Z(WX11064) ) ;
DFF     gate3277  (.D(WX11064), .CP(CLK), .Q(WX11065) ) ;
AND2    gate3278  (.A(WX11003), .B(RESET), .Z(WX11066) ) ;
DFF     gate3279  (.D(WX11066), .CP(CLK), .Q(WX11067) ) ;
AND2    gate3280  (.A(WX11005), .B(RESET), .Z(WX11068) ) ;
DFF     gate3281  (.D(WX11068), .CP(CLK), .Q(WX11069) ) ;
AND2    gate3282  (.A(WX11007), .B(RESET), .Z(WX11070) ) ;
DFF     gate3283  (.D(WX11070), .CP(CLK), .Q(WX11071) ) ;
AND2    gate3284  (.A(WX11009), .B(RESET), .Z(WX11072) ) ;
DFF     gate3285  (.D(WX11072), .CP(CLK), .Q(WX11073) ) ;
AND2    gate3286  (.A(WX11011), .B(RESET), .Z(WX11074) ) ;
DFF     gate3287  (.D(WX11074), .CP(CLK), .Q(WX11075) ) ;
AND2    gate3288  (.A(WX11013), .B(RESET), .Z(WX11076) ) ;
DFF     gate3289  (.D(WX11076), .CP(CLK), .Q(WX11077) ) ;
AND2    gate3290  (.A(WX11015), .B(RESET), .Z(WX11078) ) ;
DFF     gate3291  (.D(WX11078), .CP(CLK), .Q(WX11079) ) ;
AND2    gate3292  (.A(WX11017), .B(RESET), .Z(WX11080) ) ;
DFF     gate3293  (.D(WX11080), .CP(CLK), .Q(WX11081) ) ;
AND2    gate3294  (.A(WX11019), .B(RESET), .Z(WX11082) ) ;
DFF     gate3295  (.D(WX11082), .CP(CLK), .Q(WX11083) ) ;
AND2    gate3296  (.A(WX11021), .B(RESET), .Z(WX11084) ) ;
DFF     gate3297  (.D(WX11084), .CP(CLK), .Q(WX11085) ) ;
AND2    gate3298  (.A(WX11023), .B(RESET), .Z(WX11086) ) ;
DFF     gate3299  (.D(WX11086), .CP(CLK), .Q(WX11087) ) ;
AND2    gate3300  (.A(WX11025), .B(RESET), .Z(WX11088) ) ;
DFF     gate3301  (.D(WX11088), .CP(CLK), .Q(WX11089) ) ;
AND2    gate3302  (.A(WX11027), .B(RESET), .Z(WX11090) ) ;
DFF     gate3303  (.D(WX11090), .CP(CLK), .Q(WX11091) ) ;
AND2    gate3304  (.A(WX11029), .B(RESET), .Z(WX11092) ) ;
DFF     gate3305  (.D(WX11092), .CP(CLK), .Q(WX11093) ) ;
AND2    gate3306  (.A(WX11031), .B(RESET), .Z(WX11094) ) ;
DFF     gate3307  (.D(WX11094), .CP(CLK), .Q(WX11095) ) ;
AND2    gate3308  (.A(WX11033), .B(RESET), .Z(WX11096) ) ;
DFF     gate3309  (.D(WX11096), .CP(CLK), .Q(WX11097) ) ;
AND2    gate3310  (.A(WX11035), .B(RESET), .Z(WX11098) ) ;
DFF     gate3311  (.D(WX11098), .CP(CLK), .Q(WX11099) ) ;
AND2    gate3312  (.A(WX11037), .B(RESET), .Z(WX11100) ) ;
DFF     gate3313  (.D(WX11100), .CP(CLK), .Q(WX11101) ) ;
AND2    gate3314  (.A(WX11039), .B(RESET), .Z(WX11102) ) ;
DFF     gate3315  (.D(WX11102), .CP(CLK), .Q(WX11103) ) ;
AND2    gate3316  (.A(WX11041), .B(RESET), .Z(WX11104) ) ;
DFF     gate3317  (.D(WX11104), .CP(CLK), .Q(WX11105) ) ;
AND2    gate3318  (.A(WX11043), .B(RESET), .Z(WX11106) ) ;
DFF     gate3319  (.D(WX11106), .CP(CLK), .Q(WX11107) ) ;
AND2    gate3320  (.A(WX11045), .B(RESET), .Z(WX11108) ) ;
DFF     gate3321  (.D(WX11108), .CP(CLK), .Q(WX11109) ) ;
AND2    gate3322  (.A(WX11047), .B(RESET), .Z(WX11110) ) ;
DFF     gate3323  (.D(WX11110), .CP(CLK), .Q(WX11111) ) ;
AND2    gate3324  (.A(WX11049), .B(RESET), .Z(WX11112) ) ;
DFF     gate3325  (.D(WX11112), .CP(CLK), .Q(WX11113) ) ;
AND2    gate3326  (.A(WX11051), .B(RESET), .Z(WX11114) ) ;
DFF     gate3327  (.D(WX11114), .CP(CLK), .Q(WX11115) ) ;
AND2    gate3328  (.A(WX11053), .B(RESET), .Z(WX11116) ) ;
DFF     gate3329  (.D(WX11116), .CP(CLK), .Q(WX11117) ) ;
AND2    gate3330  (.A(WX11055), .B(RESET), .Z(WX11118) ) ;
DFF     gate3331  (.D(WX11118), .CP(CLK), .Q(WX11119) ) ;
AND2    gate3332  (.A(WX11057), .B(RESET), .Z(WX11120) ) ;
DFF     gate3333  (.D(WX11120), .CP(CLK), .Q(WX11121) ) ;
AND2    gate3334  (.A(WX11059), .B(RESET), .Z(WX11122) ) ;
DFF     gate3335  (.D(WX11122), .CP(CLK), .Q(WX11123) ) ;
AND2    gate3336  (.A(WX11061), .B(RESET), .Z(WX11124) ) ;
DFF     gate3337  (.D(WX11124), .CP(CLK), .Q(WX11125) ) ;
AND2    gate3338  (.A(WX11063), .B(RESET), .Z(WX11126) ) ;
DFF     gate3339  (.D(WX11126), .CP(CLK), .Q(WX11127) ) ;
AND2    gate3340  (.A(WX11065), .B(RESET), .Z(WX11128) ) ;
DFF     gate3341  (.D(WX11128), .CP(CLK), .Q(WX11129) ) ;
AND2    gate3342  (.A(WX11067), .B(RESET), .Z(WX11130) ) ;
DFF     gate3343  (.D(WX11130), .CP(CLK), .Q(WX11131) ) ;
AND2    gate3344  (.A(WX11069), .B(RESET), .Z(WX11132) ) ;
DFF     gate3345  (.D(WX11132), .CP(CLK), .Q(WX11133) ) ;
AND2    gate3346  (.A(WX11071), .B(RESET), .Z(WX11134) ) ;
DFF     gate3347  (.D(WX11134), .CP(CLK), .Q(WX11135) ) ;
AND2    gate3348  (.A(WX11073), .B(RESET), .Z(WX11136) ) ;
DFF     gate3349  (.D(WX11136), .CP(CLK), .Q(WX11137) ) ;
AND2    gate3350  (.A(WX11075), .B(RESET), .Z(WX11138) ) ;
DFF     gate3351  (.D(WX11138), .CP(CLK), .Q(WX11139) ) ;
AND2    gate3352  (.A(WX11077), .B(RESET), .Z(WX11140) ) ;
DFF     gate3353  (.D(WX11140), .CP(CLK), .Q(WX11141) ) ;
AND2    gate3354  (.A(WX11079), .B(RESET), .Z(WX11142) ) ;
DFF     gate3355  (.D(WX11142), .CP(CLK), .Q(WX11143) ) ;
AND2    gate3356  (.A(WX11081), .B(RESET), .Z(WX11144) ) ;
DFF     gate3357  (.D(WX11144), .CP(CLK), .Q(WX11145) ) ;
AND2    gate3358  (.A(WX11083), .B(RESET), .Z(WX11146) ) ;
DFF     gate3359  (.D(WX11146), .CP(CLK), .Q(WX11147) ) ;
AND2    gate3360  (.A(WX11085), .B(RESET), .Z(WX11148) ) ;
DFF     gate3361  (.D(WX11148), .CP(CLK), .Q(WX11149) ) ;
AND2    gate3362  (.A(WX11087), .B(RESET), .Z(WX11150) ) ;
DFF     gate3363  (.D(WX11150), .CP(CLK), .Q(WX11151) ) ;
AND2    gate3364  (.A(WX11089), .B(RESET), .Z(WX11152) ) ;
DFF     gate3365  (.D(WX11152), .CP(CLK), .Q(WX11153) ) ;
AND2    gate3366  (.A(WX11091), .B(RESET), .Z(WX11154) ) ;
DFF     gate3367  (.D(WX11154), .CP(CLK), .Q(WX11155) ) ;
AND2    gate3368  (.A(WX11093), .B(RESET), .Z(WX11156) ) ;
DFF     gate3369  (.D(WX11156), .CP(CLK), .Q(WX11157) ) ;
AND2    gate3370  (.A(WX11095), .B(RESET), .Z(WX11158) ) ;
DFF     gate3371  (.D(WX11158), .CP(CLK), .Q(WX11159) ) ;
AND2    gate3372  (.A(WX11097), .B(RESET), .Z(WX11160) ) ;
DFF     gate3373  (.D(WX11160), .CP(CLK), .Q(WX11161) ) ;
AND2    gate3374  (.A(WX11099), .B(RESET), .Z(WX11162) ) ;
DFF     gate3375  (.D(WX11162), .CP(CLK), .Q(WX11163) ) ;
AND2    gate3376  (.A(WX11101), .B(RESET), .Z(WX11164) ) ;
DFF     gate3377  (.D(WX11164), .CP(CLK), .Q(WX11165) ) ;
AND2    gate3378  (.A(WX11103), .B(RESET), .Z(WX11166) ) ;
DFF     gate3379  (.D(WX11166), .CP(CLK), .Q(WX11167) ) ;
AND2    gate3380  (.A(WX11105), .B(RESET), .Z(WX11168) ) ;
DFF     gate3381  (.D(WX11168), .CP(CLK), .Q(WX11169) ) ;
AND2    gate3382  (.A(WX11107), .B(RESET), .Z(WX11170) ) ;
DFF     gate3383  (.D(WX11170), .CP(CLK), .Q(WX11171) ) ;
AND2    gate3384  (.A(WX11109), .B(RESET), .Z(WX11172) ) ;
DFF     gate3385  (.D(WX11172), .CP(CLK), .Q(WX11173) ) ;
AND2    gate3386  (.A(WX11111), .B(RESET), .Z(WX11174) ) ;
DFF     gate3387  (.D(WX11174), .CP(CLK), .Q(WX11175) ) ;
AND2    gate3388  (.A(WX11113), .B(RESET), .Z(WX11176) ) ;
DFF     gate3389  (.D(WX11176), .CP(CLK), .Q(WX11177) ) ;
AND2    gate3390  (.A(WX11115), .B(RESET), .Z(WX11178) ) ;
DFF     gate3391  (.D(WX11178), .CP(CLK), .Q(WX11179) ) ;
AND2    gate3392  (.A(WX11117), .B(RESET), .Z(WX11180) ) ;
DFF     gate3393  (.D(WX11180), .CP(CLK), .Q(WX11181) ) ;
AND2    gate3394  (.A(WX11119), .B(RESET), .Z(WX11182) ) ;
DFF     gate3395  (.D(WX11182), .CP(CLK), .Q(WX11183) ) ;
AND2    gate3396  (.A(WX11121), .B(RESET), .Z(WX11184) ) ;
DFF     gate3397  (.D(WX11184), .CP(CLK), .Q(WX11185) ) ;
AND2    gate3398  (.A(WX11123), .B(RESET), .Z(WX11186) ) ;
DFF     gate3399  (.D(WX11186), .CP(CLK), .Q(WX11187) ) ;
AND2    gate3400  (.A(WX11125), .B(RESET), .Z(WX11188) ) ;
DFF     gate3401  (.D(WX11188), .CP(CLK), .Q(WX11189) ) ;
AND2    gate3402  (.A(WX11127), .B(RESET), .Z(WX11190) ) ;
DFF     gate3403  (.D(WX11190), .CP(CLK), .Q(WX11191) ) ;
AND2    gate3404  (.A(WX11129), .B(RESET), .Z(WX11192) ) ;
DFF     gate3405  (.D(WX11192), .CP(CLK), .Q(WX11193) ) ;
AND2    gate3406  (.A(WX11131), .B(RESET), .Z(WX11194) ) ;
DFF     gate3407  (.D(WX11194), .CP(CLK), .Q(WX11195) ) ;
AND2    gate3408  (.A(WX11133), .B(RESET), .Z(WX11196) ) ;
DFF     gate3409  (.D(WX11196), .CP(CLK), .Q(WX11197) ) ;
AND2    gate3410  (.A(WX11135), .B(RESET), .Z(WX11198) ) ;
DFF     gate3411  (.D(WX11198), .CP(CLK), .Q(WX11199) ) ;
AND2    gate3412  (.A(WX11137), .B(RESET), .Z(WX11200) ) ;
DFF     gate3413  (.D(WX11200), .CP(CLK), .Q(WX11201) ) ;
AND2    gate3414  (.A(WX11139), .B(RESET), .Z(WX11202) ) ;
DFF     gate3415  (.D(WX11202), .CP(CLK), .Q(WX11203) ) ;
AND2    gate3416  (.A(WX11141), .B(RESET), .Z(WX11204) ) ;
DFF     gate3417  (.D(WX11204), .CP(CLK), .Q(WX11205) ) ;
AND2    gate3418  (.A(WX11143), .B(RESET), .Z(WX11206) ) ;
DFF     gate3419  (.D(WX11206), .CP(CLK), .Q(WX11207) ) ;
AND2    gate3420  (.A(WX11145), .B(RESET), .Z(WX11208) ) ;
DFF     gate3421  (.D(WX11208), .CP(CLK), .Q(WX11209) ) ;
AND2    gate3422  (.A(WX11147), .B(RESET), .Z(WX11210) ) ;
DFF     gate3423  (.D(WX11210), .CP(CLK), .Q(WX11211) ) ;
AND2    gate3424  (.A(WX11149), .B(RESET), .Z(WX11212) ) ;
DFF     gate3425  (.D(WX11212), .CP(CLK), .Q(WX11213) ) ;
AND2    gate3426  (.A(WX11151), .B(RESET), .Z(WX11214) ) ;
DFF     gate3427  (.D(WX11214), .CP(CLK), .Q(WX11215) ) ;
AND2    gate3428  (.A(WX11153), .B(RESET), .Z(WX11216) ) ;
DFF     gate3429  (.D(WX11216), .CP(CLK), .Q(WX11217) ) ;
AND2    gate3430  (.A(WX11155), .B(RESET), .Z(WX11218) ) ;
DFF     gate3431  (.D(WX11218), .CP(CLK), .Q(WX11219) ) ;
AND2    gate3432  (.A(WX11157), .B(RESET), .Z(WX11220) ) ;
DFF     gate3433  (.D(WX11220), .CP(CLK), .Q(WX11221) ) ;
AND2    gate3434  (.A(WX11159), .B(RESET), .Z(WX11222) ) ;
DFF     gate3435  (.D(WX11222), .CP(CLK), .Q(WX11223) ) ;
AND2    gate3436  (.A(WX11161), .B(RESET), .Z(WX11224) ) ;
DFF     gate3437  (.D(WX11224), .CP(CLK), .Q(WX11225) ) ;
AND2    gate3438  (.A(WX11163), .B(RESET), .Z(WX11226) ) ;
DFF     gate3439  (.D(WX11226), .CP(CLK), .Q(WX11227) ) ;
AND2    gate3440  (.A(WX11165), .B(RESET), .Z(WX11228) ) ;
DFF     gate3441  (.D(WX11228), .CP(CLK), .Q(WX11229) ) ;
AND2    gate3442  (.A(WX11167), .B(RESET), .Z(WX11230) ) ;
DFF     gate3443  (.D(WX11230), .CP(CLK), .Q(WX11231) ) ;
AND2    gate3444  (.A(WX11169), .B(RESET), .Z(WX11232) ) ;
DFF     gate3445  (.D(WX11232), .CP(CLK), .Q(WX11233) ) ;
AND2    gate3446  (.A(WX11171), .B(RESET), .Z(WX11234) ) ;
DFF     gate3447  (.D(WX11234), .CP(CLK), .Q(WX11235) ) ;
AND2    gate3448  (.A(WX11173), .B(RESET), .Z(WX11236) ) ;
DFF     gate3449  (.D(WX11236), .CP(CLK), .Q(WX11237) ) ;
AND2    gate3450  (.A(WX11175), .B(RESET), .Z(WX11238) ) ;
DFF     gate3451  (.D(WX11238), .CP(CLK), .Q(WX11239) ) ;
AND2    gate3452  (.A(WX11177), .B(RESET), .Z(WX11240) ) ;
DFF     gate3453  (.D(WX11240), .CP(CLK), .Q(WX11241) ) ;
AND2    gate3454  (.A(WX11179), .B(RESET), .Z(WX11242) ) ;
DFF     gate3455  (.D(WX11242), .CP(CLK), .Q(WX11243) ) ;
AND2    gate3456  (.A(WX11578), .B(WX11607), .Z(WX11608) ) ;
AND2    gate3457  (.A(WX11606), .B(WX11607), .Z(WX11610) ) ;
AND2    gate3458  (.A(WX11605), .B(WX11607), .Z(WX11612) ) ;
AND2    gate3459  (.A(WX11604), .B(WX11607), .Z(WX11614) ) ;
AND2    gate3460  (.A(WX11577), .B(WX11607), .Z(WX11616) ) ;
AND2    gate3461  (.A(WX11603), .B(WX11607), .Z(WX11618) ) ;
AND2    gate3462  (.A(WX11602), .B(WX11607), .Z(WX11620) ) ;
AND2    gate3463  (.A(WX11601), .B(WX11607), .Z(WX11622) ) ;
AND2    gate3464  (.A(WX11600), .B(WX11607), .Z(WX11624) ) ;
AND2    gate3465  (.A(WX11599), .B(WX11607), .Z(WX11626) ) ;
AND2    gate3466  (.A(WX11598), .B(WX11607), .Z(WX11628) ) ;
AND2    gate3467  (.A(WX11576), .B(WX11607), .Z(WX11630) ) ;
AND2    gate3468  (.A(WX11597), .B(WX11607), .Z(WX11632) ) ;
AND2    gate3469  (.A(WX11596), .B(WX11607), .Z(WX11634) ) ;
AND2    gate3470  (.A(WX11595), .B(WX11607), .Z(WX11636) ) ;
AND2    gate3471  (.A(WX11594), .B(WX11607), .Z(WX11638) ) ;
AND2    gate3472  (.A(WX11575), .B(WX11607), .Z(WX11640) ) ;
AND2    gate3473  (.A(WX11593), .B(WX11607), .Z(WX11642) ) ;
AND2    gate3474  (.A(WX11592), .B(WX11607), .Z(WX11644) ) ;
AND2    gate3475  (.A(WX11591), .B(WX11607), .Z(WX11646) ) ;
AND2    gate3476  (.A(WX11590), .B(WX11607), .Z(WX11648) ) ;
AND2    gate3477  (.A(WX11589), .B(WX11607), .Z(WX11650) ) ;
AND2    gate3478  (.A(WX11588), .B(WX11607), .Z(WX11652) ) ;
AND2    gate3479  (.A(WX11587), .B(WX11607), .Z(WX11654) ) ;
AND2    gate3480  (.A(WX11586), .B(WX11607), .Z(WX11656) ) ;
AND2    gate3481  (.A(WX11585), .B(WX11607), .Z(WX11658) ) ;
AND2    gate3482  (.A(WX11584), .B(WX11607), .Z(WX11660) ) ;
AND2    gate3483  (.A(WX11583), .B(WX11607), .Z(WX11662) ) ;
AND2    gate3484  (.A(WX11582), .B(WX11607), .Z(WX11664) ) ;
AND2    gate3485  (.A(WX11581), .B(WX11607), .Z(WX11666) ) ;
AND2    gate3486  (.A(WX11580), .B(WX11607), .Z(WX11668) ) ;
AND2    gate3487  (.A(WX11579), .B(WX11607), .Z(WX11670) ) ;
INV     gate3488  (.A(WX999), .Z(WX1003) ) ;
INV     gate3489  (.A(WX1003), .Z(WX37) ) ;
INV     gate3490  (.A(WX997), .Z(WX1004) ) ;
INV     gate3491  (.A(WX1004), .Z(WX41) ) ;
INV     gate3492  (.A(WX1004), .Z(WX45) ) ;
OR2     gate3493  (.A(WX36), .B(WX35), .Z(WX38) ) ;
INV     gate3494  (.A(WX38), .Z(WX47) ) ;
INV     gate3495  (.A(WX47), .Z(WX48) ) ;
INV     gate3496  (.A(WX1003), .Z(WX51) ) ;
INV     gate3497  (.A(WX1004), .Z(WX55) ) ;
INV     gate3498  (.A(WX1004), .Z(WX59) ) ;
OR2     gate3499  (.A(WX50), .B(WX49), .Z(WX52) ) ;
INV     gate3500  (.A(WX52), .Z(WX61) ) ;
INV     gate3501  (.A(WX61), .Z(WX62) ) ;
INV     gate3502  (.A(WX1003), .Z(WX65) ) ;
INV     gate3503  (.A(WX1004), .Z(WX69) ) ;
INV     gate3504  (.A(WX1004), .Z(WX73) ) ;
OR2     gate3505  (.A(WX64), .B(WX63), .Z(WX66) ) ;
INV     gate3506  (.A(WX66), .Z(WX75) ) ;
INV     gate3507  (.A(WX75), .Z(WX76) ) ;
INV     gate3508  (.A(WX1003), .Z(WX79) ) ;
INV     gate3509  (.A(WX1004), .Z(WX83) ) ;
INV     gate3510  (.A(WX1004), .Z(WX87) ) ;
OR2     gate3511  (.A(WX78), .B(WX77), .Z(WX80) ) ;
INV     gate3512  (.A(WX80), .Z(WX89) ) ;
INV     gate3513  (.A(WX89), .Z(WX90) ) ;
INV     gate3514  (.A(WX1003), .Z(WX93) ) ;
INV     gate3515  (.A(WX1004), .Z(WX97) ) ;
INV     gate3516  (.A(WX1004), .Z(WX101) ) ;
OR2     gate3517  (.A(WX92), .B(WX91), .Z(WX94) ) ;
INV     gate3518  (.A(WX94), .Z(WX103) ) ;
INV     gate3519  (.A(WX103), .Z(WX104) ) ;
INV     gate3520  (.A(WX1003), .Z(WX107) ) ;
INV     gate3521  (.A(WX1004), .Z(WX111) ) ;
INV     gate3522  (.A(WX1004), .Z(WX115) ) ;
OR2     gate3523  (.A(WX106), .B(WX105), .Z(WX108) ) ;
INV     gate3524  (.A(WX108), .Z(WX117) ) ;
INV     gate3525  (.A(WX117), .Z(WX118) ) ;
INV     gate3526  (.A(WX1003), .Z(WX121) ) ;
INV     gate3527  (.A(WX1004), .Z(WX125) ) ;
INV     gate3528  (.A(WX1004), .Z(WX129) ) ;
OR2     gate3529  (.A(WX120), .B(WX119), .Z(WX122) ) ;
INV     gate3530  (.A(WX122), .Z(WX131) ) ;
INV     gate3531  (.A(WX131), .Z(WX132) ) ;
INV     gate3532  (.A(WX1003), .Z(WX135) ) ;
INV     gate3533  (.A(WX1004), .Z(WX139) ) ;
INV     gate3534  (.A(WX1004), .Z(WX143) ) ;
OR2     gate3535  (.A(WX134), .B(WX133), .Z(WX136) ) ;
INV     gate3536  (.A(WX136), .Z(WX145) ) ;
INV     gate3537  (.A(WX145), .Z(WX146) ) ;
INV     gate3538  (.A(WX1003), .Z(WX149) ) ;
INV     gate3539  (.A(WX1004), .Z(WX153) ) ;
INV     gate3540  (.A(WX1004), .Z(WX157) ) ;
OR2     gate3541  (.A(WX148), .B(WX147), .Z(WX150) ) ;
INV     gate3542  (.A(WX150), .Z(WX159) ) ;
INV     gate3543  (.A(WX159), .Z(WX160) ) ;
INV     gate3544  (.A(WX1003), .Z(WX163) ) ;
INV     gate3545  (.A(WX1004), .Z(WX167) ) ;
INV     gate3546  (.A(WX1004), .Z(WX171) ) ;
OR2     gate3547  (.A(WX162), .B(WX161), .Z(WX164) ) ;
INV     gate3548  (.A(WX164), .Z(WX173) ) ;
INV     gate3549  (.A(WX173), .Z(WX174) ) ;
INV     gate3550  (.A(WX1003), .Z(WX177) ) ;
INV     gate3551  (.A(WX1004), .Z(WX181) ) ;
INV     gate3552  (.A(WX1004), .Z(WX185) ) ;
OR2     gate3553  (.A(WX176), .B(WX175), .Z(WX178) ) ;
INV     gate3554  (.A(WX178), .Z(WX187) ) ;
INV     gate3555  (.A(WX187), .Z(WX188) ) ;
INV     gate3556  (.A(WX1003), .Z(WX191) ) ;
INV     gate3557  (.A(WX1004), .Z(WX195) ) ;
INV     gate3558  (.A(WX1004), .Z(WX199) ) ;
OR2     gate3559  (.A(WX190), .B(WX189), .Z(WX192) ) ;
INV     gate3560  (.A(WX192), .Z(WX201) ) ;
INV     gate3561  (.A(WX201), .Z(WX202) ) ;
INV     gate3562  (.A(WX1003), .Z(WX205) ) ;
INV     gate3563  (.A(WX1004), .Z(WX209) ) ;
INV     gate3564  (.A(WX1004), .Z(WX213) ) ;
OR2     gate3565  (.A(WX204), .B(WX203), .Z(WX206) ) ;
INV     gate3566  (.A(WX206), .Z(WX215) ) ;
INV     gate3567  (.A(WX215), .Z(WX216) ) ;
INV     gate3568  (.A(WX1003), .Z(WX219) ) ;
INV     gate3569  (.A(WX1004), .Z(WX223) ) ;
INV     gate3570  (.A(WX1004), .Z(WX227) ) ;
OR2     gate3571  (.A(WX218), .B(WX217), .Z(WX220) ) ;
INV     gate3572  (.A(WX220), .Z(WX229) ) ;
INV     gate3573  (.A(WX229), .Z(WX230) ) ;
INV     gate3574  (.A(WX1003), .Z(WX233) ) ;
INV     gate3575  (.A(WX1004), .Z(WX237) ) ;
INV     gate3576  (.A(WX1004), .Z(WX241) ) ;
OR2     gate3577  (.A(WX232), .B(WX231), .Z(WX234) ) ;
INV     gate3578  (.A(WX234), .Z(WX243) ) ;
INV     gate3579  (.A(WX243), .Z(WX244) ) ;
INV     gate3580  (.A(WX1003), .Z(WX247) ) ;
INV     gate3581  (.A(WX1004), .Z(WX251) ) ;
INV     gate3582  (.A(WX1004), .Z(WX255) ) ;
OR2     gate3583  (.A(WX246), .B(WX245), .Z(WX248) ) ;
INV     gate3584  (.A(WX248), .Z(WX257) ) ;
INV     gate3585  (.A(WX257), .Z(WX258) ) ;
INV     gate3586  (.A(WX1003), .Z(WX261) ) ;
INV     gate3587  (.A(WX1004), .Z(WX265) ) ;
INV     gate3588  (.A(WX1004), .Z(WX269) ) ;
OR2     gate3589  (.A(WX260), .B(WX259), .Z(WX262) ) ;
INV     gate3590  (.A(WX262), .Z(WX271) ) ;
INV     gate3591  (.A(WX271), .Z(WX272) ) ;
INV     gate3592  (.A(WX1003), .Z(WX275) ) ;
INV     gate3593  (.A(WX1004), .Z(WX279) ) ;
INV     gate3594  (.A(WX1004), .Z(WX283) ) ;
OR2     gate3595  (.A(WX274), .B(WX273), .Z(WX276) ) ;
INV     gate3596  (.A(WX276), .Z(WX285) ) ;
INV     gate3597  (.A(WX285), .Z(WX286) ) ;
INV     gate3598  (.A(WX1003), .Z(WX289) ) ;
INV     gate3599  (.A(WX1004), .Z(WX293) ) ;
INV     gate3600  (.A(WX1004), .Z(WX297) ) ;
OR2     gate3601  (.A(WX288), .B(WX287), .Z(WX290) ) ;
INV     gate3602  (.A(WX290), .Z(WX299) ) ;
INV     gate3603  (.A(WX299), .Z(WX300) ) ;
INV     gate3604  (.A(WX1003), .Z(WX303) ) ;
INV     gate3605  (.A(WX1004), .Z(WX307) ) ;
INV     gate3606  (.A(WX1004), .Z(WX311) ) ;
OR2     gate3607  (.A(WX302), .B(WX301), .Z(WX304) ) ;
INV     gate3608  (.A(WX304), .Z(WX313) ) ;
INV     gate3609  (.A(WX313), .Z(WX314) ) ;
INV     gate3610  (.A(WX1003), .Z(WX317) ) ;
INV     gate3611  (.A(WX1004), .Z(WX321) ) ;
INV     gate3612  (.A(WX1004), .Z(WX325) ) ;
OR2     gate3613  (.A(WX316), .B(WX315), .Z(WX318) ) ;
INV     gate3614  (.A(WX318), .Z(WX327) ) ;
INV     gate3615  (.A(WX327), .Z(WX328) ) ;
INV     gate3616  (.A(WX1003), .Z(WX331) ) ;
INV     gate3617  (.A(WX1004), .Z(WX335) ) ;
INV     gate3618  (.A(WX1004), .Z(WX339) ) ;
OR2     gate3619  (.A(WX330), .B(WX329), .Z(WX332) ) ;
INV     gate3620  (.A(WX332), .Z(WX341) ) ;
INV     gate3621  (.A(WX341), .Z(WX342) ) ;
INV     gate3622  (.A(WX1003), .Z(WX345) ) ;
INV     gate3623  (.A(WX1004), .Z(WX349) ) ;
INV     gate3624  (.A(WX1004), .Z(WX353) ) ;
OR2     gate3625  (.A(WX344), .B(WX343), .Z(WX346) ) ;
INV     gate3626  (.A(WX346), .Z(WX355) ) ;
INV     gate3627  (.A(WX355), .Z(WX356) ) ;
INV     gate3628  (.A(WX1003), .Z(WX359) ) ;
INV     gate3629  (.A(WX1004), .Z(WX363) ) ;
INV     gate3630  (.A(WX1004), .Z(WX367) ) ;
OR2     gate3631  (.A(WX358), .B(WX357), .Z(WX360) ) ;
INV     gate3632  (.A(WX360), .Z(WX369) ) ;
INV     gate3633  (.A(WX369), .Z(WX370) ) ;
INV     gate3634  (.A(WX1003), .Z(WX373) ) ;
INV     gate3635  (.A(WX1004), .Z(WX377) ) ;
INV     gate3636  (.A(WX1004), .Z(WX381) ) ;
OR2     gate3637  (.A(WX372), .B(WX371), .Z(WX374) ) ;
INV     gate3638  (.A(WX374), .Z(WX383) ) ;
INV     gate3639  (.A(WX383), .Z(WX384) ) ;
INV     gate3640  (.A(WX1003), .Z(WX387) ) ;
INV     gate3641  (.A(WX1004), .Z(WX391) ) ;
INV     gate3642  (.A(WX1004), .Z(WX395) ) ;
OR2     gate3643  (.A(WX386), .B(WX385), .Z(WX388) ) ;
INV     gate3644  (.A(WX388), .Z(WX397) ) ;
INV     gate3645  (.A(WX397), .Z(WX398) ) ;
INV     gate3646  (.A(WX1003), .Z(WX401) ) ;
INV     gate3647  (.A(WX1004), .Z(WX405) ) ;
INV     gate3648  (.A(WX1004), .Z(WX409) ) ;
OR2     gate3649  (.A(WX400), .B(WX399), .Z(WX402) ) ;
INV     gate3650  (.A(WX402), .Z(WX411) ) ;
INV     gate3651  (.A(WX411), .Z(WX412) ) ;
INV     gate3652  (.A(WX1003), .Z(WX415) ) ;
INV     gate3653  (.A(WX1004), .Z(WX419) ) ;
INV     gate3654  (.A(WX1004), .Z(WX423) ) ;
OR2     gate3655  (.A(WX414), .B(WX413), .Z(WX416) ) ;
INV     gate3656  (.A(WX416), .Z(WX425) ) ;
INV     gate3657  (.A(WX425), .Z(WX426) ) ;
INV     gate3658  (.A(WX1003), .Z(WX429) ) ;
INV     gate3659  (.A(WX1004), .Z(WX433) ) ;
INV     gate3660  (.A(WX1004), .Z(WX437) ) ;
OR2     gate3661  (.A(WX428), .B(WX427), .Z(WX430) ) ;
INV     gate3662  (.A(WX430), .Z(WX439) ) ;
INV     gate3663  (.A(WX439), .Z(WX440) ) ;
INV     gate3664  (.A(WX1003), .Z(WX443) ) ;
INV     gate3665  (.A(WX1004), .Z(WX447) ) ;
INV     gate3666  (.A(WX1004), .Z(WX451) ) ;
OR2     gate3667  (.A(WX442), .B(WX441), .Z(WX444) ) ;
INV     gate3668  (.A(WX444), .Z(WX453) ) ;
INV     gate3669  (.A(WX453), .Z(WX454) ) ;
INV     gate3670  (.A(WX1003), .Z(WX457) ) ;
INV     gate3671  (.A(WX1004), .Z(WX461) ) ;
INV     gate3672  (.A(WX1004), .Z(WX465) ) ;
OR2     gate3673  (.A(WX456), .B(WX455), .Z(WX458) ) ;
INV     gate3674  (.A(WX458), .Z(WX467) ) ;
INV     gate3675  (.A(WX467), .Z(WX468) ) ;
INV     gate3676  (.A(WX1003), .Z(WX471) ) ;
INV     gate3677  (.A(WX1004), .Z(WX475) ) ;
INV     gate3678  (.A(WX1004), .Z(WX479) ) ;
OR2     gate3679  (.A(WX470), .B(WX469), .Z(WX472) ) ;
INV     gate3680  (.A(WX472), .Z(WX481) ) ;
INV     gate3681  (.A(WX481), .Z(WX482) ) ;
INV     gate3682  (.A(WX485), .Z(WX483) ) ;
INV     gate3683  (.A(WX964), .Z(WX965) ) ;
INV     gate3684  (.A(WX965), .Z(WX548) ) ;
INV     gate3685  (.A(WX966), .Z(WX967) ) ;
INV     gate3686  (.A(WX967), .Z(WX549) ) ;
INV     gate3687  (.A(WX968), .Z(WX969) ) ;
INV     gate3688  (.A(WX969), .Z(WX550) ) ;
INV     gate3689  (.A(WX970), .Z(WX971) ) ;
INV     gate3690  (.A(WX971), .Z(WX551) ) ;
INV     gate3691  (.A(WX972), .Z(WX973) ) ;
INV     gate3692  (.A(WX973), .Z(WX552) ) ;
INV     gate3693  (.A(WX974), .Z(WX975) ) ;
INV     gate3694  (.A(WX975), .Z(WX553) ) ;
INV     gate3695  (.A(WX976), .Z(WX977) ) ;
INV     gate3696  (.A(WX977), .Z(WX554) ) ;
INV     gate3697  (.A(WX978), .Z(WX979) ) ;
INV     gate3698  (.A(WX979), .Z(WX555) ) ;
INV     gate3699  (.A(WX980), .Z(WX981) ) ;
INV     gate3700  (.A(WX981), .Z(WX556) ) ;
INV     gate3701  (.A(WX982), .Z(WX983) ) ;
INV     gate3702  (.A(WX983), .Z(WX557) ) ;
INV     gate3703  (.A(WX984), .Z(WX985) ) ;
INV     gate3704  (.A(WX985), .Z(WX558) ) ;
INV     gate3705  (.A(WX986), .Z(WX987) ) ;
INV     gate3706  (.A(WX987), .Z(WX559) ) ;
INV     gate3707  (.A(WX988), .Z(WX989) ) ;
INV     gate3708  (.A(WX989), .Z(WX560) ) ;
INV     gate3709  (.A(WX990), .Z(WX991) ) ;
INV     gate3710  (.A(WX991), .Z(WX561) ) ;
INV     gate3711  (.A(WX992), .Z(WX993) ) ;
INV     gate3712  (.A(WX993), .Z(WX562) ) ;
INV     gate3713  (.A(WX994), .Z(WX995) ) ;
INV     gate3714  (.A(WX995), .Z(WX563) ) ;
INV     gate3715  (.A(WX932), .Z(WX933) ) ;
INV     gate3716  (.A(WX933), .Z(WX564) ) ;
INV     gate3717  (.A(WX934), .Z(WX935) ) ;
INV     gate3718  (.A(WX935), .Z(WX565) ) ;
INV     gate3719  (.A(WX936), .Z(WX937) ) ;
INV     gate3720  (.A(WX937), .Z(WX566) ) ;
INV     gate3721  (.A(WX938), .Z(WX939) ) ;
INV     gate3722  (.A(WX939), .Z(WX567) ) ;
INV     gate3723  (.A(WX940), .Z(WX941) ) ;
INV     gate3724  (.A(WX941), .Z(WX568) ) ;
INV     gate3725  (.A(WX942), .Z(WX943) ) ;
INV     gate3726  (.A(WX943), .Z(WX569) ) ;
INV     gate3727  (.A(WX944), .Z(WX945) ) ;
INV     gate3728  (.A(WX945), .Z(WX570) ) ;
INV     gate3729  (.A(WX946), .Z(WX947) ) ;
INV     gate3730  (.A(WX947), .Z(WX571) ) ;
INV     gate3731  (.A(WX948), .Z(WX949) ) ;
INV     gate3732  (.A(WX949), .Z(WX572) ) ;
INV     gate3733  (.A(WX950), .Z(WX951) ) ;
INV     gate3734  (.A(WX951), .Z(WX573) ) ;
INV     gate3735  (.A(WX952), .Z(WX953) ) ;
INV     gate3736  (.A(WX953), .Z(WX574) ) ;
INV     gate3737  (.A(WX954), .Z(WX955) ) ;
INV     gate3738  (.A(WX955), .Z(WX575) ) ;
INV     gate3739  (.A(WX956), .Z(WX957) ) ;
INV     gate3740  (.A(WX957), .Z(WX576) ) ;
INV     gate3741  (.A(WX958), .Z(WX959) ) ;
INV     gate3742  (.A(WX959), .Z(WX577) ) ;
INV     gate3743  (.A(WX960), .Z(WX961) ) ;
INV     gate3744  (.A(WX961), .Z(WX578) ) ;
INV     gate3745  (.A(WX962), .Z(WX963) ) ;
INV     gate3746  (.A(WX963), .Z(WX579) ) ;
INV     gate3747  (.A(WX548), .Z(WX580) ) ;
INV     gate3748  (.A(WX549), .Z(WX581) ) ;
INV     gate3749  (.A(WX550), .Z(WX582) ) ;
INV     gate3750  (.A(WX551), .Z(WX583) ) ;
INV     gate3751  (.A(WX552), .Z(WX584) ) ;
INV     gate3752  (.A(WX553), .Z(WX585) ) ;
INV     gate3753  (.A(WX554), .Z(WX586) ) ;
INV     gate3754  (.A(WX555), .Z(WX587) ) ;
INV     gate3755  (.A(WX556), .Z(WX588) ) ;
INV     gate3756  (.A(WX557), .Z(WX589) ) ;
INV     gate3757  (.A(WX558), .Z(WX590) ) ;
INV     gate3758  (.A(WX559), .Z(WX591) ) ;
INV     gate3759  (.A(WX560), .Z(WX592) ) ;
INV     gate3760  (.A(WX561), .Z(WX593) ) ;
INV     gate3761  (.A(WX562), .Z(WX594) ) ;
INV     gate3762  (.A(WX563), .Z(WX595) ) ;
INV     gate3763  (.A(WX564), .Z(WX596) ) ;
INV     gate3764  (.A(WX565), .Z(WX597) ) ;
INV     gate3765  (.A(WX566), .Z(WX598) ) ;
INV     gate3766  (.A(WX567), .Z(WX599) ) ;
INV     gate3767  (.A(WX568), .Z(WX600) ) ;
INV     gate3768  (.A(WX569), .Z(WX601) ) ;
INV     gate3769  (.A(WX570), .Z(WX602) ) ;
INV     gate3770  (.A(WX571), .Z(WX603) ) ;
INV     gate3771  (.A(WX572), .Z(WX604) ) ;
INV     gate3772  (.A(WX573), .Z(WX605) ) ;
INV     gate3773  (.A(WX574), .Z(WX606) ) ;
INV     gate3774  (.A(WX575), .Z(WX607) ) ;
INV     gate3775  (.A(WX576), .Z(WX608) ) ;
INV     gate3776  (.A(WX577), .Z(WX609) ) ;
INV     gate3777  (.A(WX578), .Z(WX610) ) ;
INV     gate3778  (.A(WX579), .Z(WX611) ) ;
INV     gate3779  (.A(WX837), .Z(WX612) ) ;
INV     gate3780  (.A(WX839), .Z(WX613) ) ;
INV     gate3781  (.A(WX841), .Z(WX614) ) ;
INV     gate3782  (.A(WX843), .Z(WX615) ) ;
INV     gate3783  (.A(WX845), .Z(WX616) ) ;
INV     gate3784  (.A(WX847), .Z(WX617) ) ;
INV     gate3785  (.A(WX849), .Z(WX618) ) ;
INV     gate3786  (.A(WX851), .Z(WX619) ) ;
INV     gate3787  (.A(WX853), .Z(WX620) ) ;
INV     gate3788  (.A(WX855), .Z(WX621) ) ;
INV     gate3789  (.A(WX857), .Z(WX622) ) ;
INV     gate3790  (.A(WX859), .Z(WX623) ) ;
INV     gate3791  (.A(WX861), .Z(WX624) ) ;
INV     gate3792  (.A(WX863), .Z(WX625) ) ;
INV     gate3793  (.A(WX865), .Z(WX626) ) ;
INV     gate3794  (.A(WX867), .Z(WX627) ) ;
INV     gate3795  (.A(WX869), .Z(WX628) ) ;
INV     gate3796  (.A(WX871), .Z(WX629) ) ;
INV     gate3797  (.A(WX873), .Z(WX630) ) ;
INV     gate3798  (.A(WX875), .Z(WX631) ) ;
INV     gate3799  (.A(WX877), .Z(WX632) ) ;
INV     gate3800  (.A(WX879), .Z(WX633) ) ;
INV     gate3801  (.A(WX881), .Z(WX634) ) ;
INV     gate3802  (.A(WX883), .Z(WX635) ) ;
INV     gate3803  (.A(WX885), .Z(WX636) ) ;
INV     gate3804  (.A(WX887), .Z(WX637) ) ;
INV     gate3805  (.A(WX889), .Z(WX638) ) ;
INV     gate3806  (.A(WX891), .Z(WX639) ) ;
INV     gate3807  (.A(WX893), .Z(WX640) ) ;
INV     gate3808  (.A(WX895), .Z(WX641) ) ;
INV     gate3809  (.A(WX897), .Z(WX642) ) ;
INV     gate3810  (.A(WX899), .Z(WX643) ) ;
NAND2   gate3811  (.A(II2507), .B(II2508), .Z(WX916) ) ;
INV     gate3812  (.A(WX916), .Z(WX932) ) ;
NAND2   gate3813  (.A(II2538), .B(II2539), .Z(WX917) ) ;
INV     gate3814  (.A(WX917), .Z(WX934) ) ;
NAND2   gate3815  (.A(II2569), .B(II2570), .Z(WX918) ) ;
INV     gate3816  (.A(WX918), .Z(WX936) ) ;
NAND2   gate3817  (.A(II2600), .B(II2601), .Z(WX919) ) ;
INV     gate3818  (.A(WX919), .Z(WX938) ) ;
NAND2   gate3819  (.A(II2631), .B(II2632), .Z(WX920) ) ;
INV     gate3820  (.A(WX920), .Z(WX940) ) ;
NAND2   gate3821  (.A(II2662), .B(II2663), .Z(WX921) ) ;
INV     gate3822  (.A(WX921), .Z(WX942) ) ;
NAND2   gate3823  (.A(II2693), .B(II2694), .Z(WX922) ) ;
INV     gate3824  (.A(WX922), .Z(WX944) ) ;
NAND2   gate3825  (.A(II2724), .B(II2725), .Z(WX923) ) ;
INV     gate3826  (.A(WX923), .Z(WX946) ) ;
NAND2   gate3827  (.A(II2755), .B(II2756), .Z(WX924) ) ;
INV     gate3828  (.A(WX924), .Z(WX948) ) ;
NAND2   gate3829  (.A(II2786), .B(II2787), .Z(WX925) ) ;
INV     gate3830  (.A(WX925), .Z(WX950) ) ;
NAND2   gate3831  (.A(II2817), .B(II2818), .Z(WX926) ) ;
INV     gate3832  (.A(WX926), .Z(WX952) ) ;
NAND2   gate3833  (.A(II2848), .B(II2849), .Z(WX927) ) ;
INV     gate3834  (.A(WX927), .Z(WX954) ) ;
NAND2   gate3835  (.A(II2879), .B(II2880), .Z(WX928) ) ;
INV     gate3836  (.A(WX928), .Z(WX956) ) ;
NAND2   gate3837  (.A(II2910), .B(II2911), .Z(WX929) ) ;
INV     gate3838  (.A(WX929), .Z(WX958) ) ;
NAND2   gate3839  (.A(II2941), .B(II2942), .Z(WX930) ) ;
INV     gate3840  (.A(WX930), .Z(WX960) ) ;
NAND2   gate3841  (.A(II2972), .B(II2973), .Z(WX931) ) ;
INV     gate3842  (.A(WX931), .Z(WX962) ) ;
NAND2   gate3843  (.A(II2011), .B(II2012), .Z(WX900) ) ;
INV     gate3844  (.A(WX900), .Z(WX964) ) ;
NAND2   gate3845  (.A(II2042), .B(II2043), .Z(WX901) ) ;
INV     gate3846  (.A(WX901), .Z(WX966) ) ;
NAND2   gate3847  (.A(II2073), .B(II2074), .Z(WX902) ) ;
INV     gate3848  (.A(WX902), .Z(WX968) ) ;
NAND2   gate3849  (.A(II2104), .B(II2105), .Z(WX903) ) ;
INV     gate3850  (.A(WX903), .Z(WX970) ) ;
NAND2   gate3851  (.A(II2135), .B(II2136), .Z(WX904) ) ;
INV     gate3852  (.A(WX904), .Z(WX972) ) ;
NAND2   gate3853  (.A(II2166), .B(II2167), .Z(WX905) ) ;
INV     gate3854  (.A(WX905), .Z(WX974) ) ;
NAND2   gate3855  (.A(II2197), .B(II2198), .Z(WX906) ) ;
INV     gate3856  (.A(WX906), .Z(WX976) ) ;
NAND2   gate3857  (.A(II2228), .B(II2229), .Z(WX907) ) ;
INV     gate3858  (.A(WX907), .Z(WX978) ) ;
NAND2   gate3859  (.A(II2259), .B(II2260), .Z(WX908) ) ;
INV     gate3860  (.A(WX908), .Z(WX980) ) ;
NAND2   gate3861  (.A(II2290), .B(II2291), .Z(WX909) ) ;
INV     gate3862  (.A(WX909), .Z(WX982) ) ;
NAND2   gate3863  (.A(II2321), .B(II2322), .Z(WX910) ) ;
INV     gate3864  (.A(WX910), .Z(WX984) ) ;
NAND2   gate3865  (.A(II2352), .B(II2353), .Z(WX911) ) ;
INV     gate3866  (.A(WX911), .Z(WX986) ) ;
NAND2   gate3867  (.A(II2383), .B(II2384), .Z(WX912) ) ;
INV     gate3868  (.A(WX912), .Z(WX988) ) ;
NAND2   gate3869  (.A(II2414), .B(II2415), .Z(WX913) ) ;
INV     gate3870  (.A(WX913), .Z(WX990) ) ;
NAND2   gate3871  (.A(II2445), .B(II2446), .Z(WX914) ) ;
INV     gate3872  (.A(WX914), .Z(WX992) ) ;
NAND2   gate3873  (.A(II2476), .B(II2477), .Z(WX915) ) ;
INV     gate3874  (.A(WX915), .Z(WX994) ) ;
INV     gate3875  (.A(TM0), .Z(WX996) ) ;
INV     gate3876  (.A(TM0), .Z(WX997) ) ;
INV     gate3877  (.A(TM0), .Z(WX998) ) ;
INV     gate3878  (.A(TM1), .Z(WX999) ) ;
INV     gate3879  (.A(TM1), .Z(WX1000) ) ;
INV     gate3880  (.A(WX1000), .Z(WX1001) ) ;
INV     gate3881  (.A(WX998), .Z(WX1002) ) ;
INV     gate3882  (.A(WX996), .Z(WX1005) ) ;
INV     gate3883  (.A(WX1005), .Z(WX1009) ) ;
OR2     gate3884  (.A(WX1008), .B(WX1007), .Z(WX1010) ) ;
INV     gate3885  (.A(WX1010), .Z(WX1011) ) ;
INV     gate3886  (.A(WX1005), .Z(WX1016) ) ;
OR2     gate3887  (.A(WX1015), .B(WX1014), .Z(WX1017) ) ;
INV     gate3888  (.A(WX1017), .Z(WX1018) ) ;
INV     gate3889  (.A(WX1005), .Z(WX1023) ) ;
OR2     gate3890  (.A(WX1022), .B(WX1021), .Z(WX1024) ) ;
INV     gate3891  (.A(WX1024), .Z(WX1025) ) ;
INV     gate3892  (.A(WX1005), .Z(WX1030) ) ;
OR2     gate3893  (.A(WX1029), .B(WX1028), .Z(WX1031) ) ;
INV     gate3894  (.A(WX1031), .Z(WX1032) ) ;
INV     gate3895  (.A(WX1005), .Z(WX1037) ) ;
OR2     gate3896  (.A(WX1036), .B(WX1035), .Z(WX1038) ) ;
INV     gate3897  (.A(WX1038), .Z(WX1039) ) ;
INV     gate3898  (.A(WX1005), .Z(WX1044) ) ;
OR2     gate3899  (.A(WX1043), .B(WX1042), .Z(WX1045) ) ;
INV     gate3900  (.A(WX1045), .Z(WX1046) ) ;
INV     gate3901  (.A(WX1005), .Z(WX1051) ) ;
OR2     gate3902  (.A(WX1050), .B(WX1049), .Z(WX1052) ) ;
INV     gate3903  (.A(WX1052), .Z(WX1053) ) ;
INV     gate3904  (.A(WX1005), .Z(WX1058) ) ;
OR2     gate3905  (.A(WX1057), .B(WX1056), .Z(WX1059) ) ;
INV     gate3906  (.A(WX1059), .Z(WX1060) ) ;
INV     gate3907  (.A(WX1005), .Z(WX1065) ) ;
OR2     gate3908  (.A(WX1064), .B(WX1063), .Z(WX1066) ) ;
INV     gate3909  (.A(WX1066), .Z(WX1067) ) ;
INV     gate3910  (.A(WX1005), .Z(WX1072) ) ;
OR2     gate3911  (.A(WX1071), .B(WX1070), .Z(WX1073) ) ;
INV     gate3912  (.A(WX1073), .Z(WX1074) ) ;
INV     gate3913  (.A(WX1005), .Z(WX1079) ) ;
OR2     gate3914  (.A(WX1078), .B(WX1077), .Z(WX1080) ) ;
INV     gate3915  (.A(WX1080), .Z(WX1081) ) ;
INV     gate3916  (.A(WX1005), .Z(WX1086) ) ;
OR2     gate3917  (.A(WX1085), .B(WX1084), .Z(WX1087) ) ;
INV     gate3918  (.A(WX1087), .Z(WX1088) ) ;
INV     gate3919  (.A(WX1005), .Z(WX1093) ) ;
OR2     gate3920  (.A(WX1092), .B(WX1091), .Z(WX1094) ) ;
INV     gate3921  (.A(WX1094), .Z(WX1095) ) ;
INV     gate3922  (.A(WX1005), .Z(WX1100) ) ;
OR2     gate3923  (.A(WX1099), .B(WX1098), .Z(WX1101) ) ;
INV     gate3924  (.A(WX1101), .Z(WX1102) ) ;
INV     gate3925  (.A(WX1005), .Z(WX1107) ) ;
OR2     gate3926  (.A(WX1106), .B(WX1105), .Z(WX1108) ) ;
INV     gate3927  (.A(WX1108), .Z(WX1109) ) ;
INV     gate3928  (.A(WX1005), .Z(WX1114) ) ;
OR2     gate3929  (.A(WX1113), .B(WX1112), .Z(WX1115) ) ;
INV     gate3930  (.A(WX1115), .Z(WX1116) ) ;
INV     gate3931  (.A(WX1005), .Z(WX1121) ) ;
OR2     gate3932  (.A(WX1120), .B(WX1119), .Z(WX1122) ) ;
INV     gate3933  (.A(WX1122), .Z(WX1123) ) ;
INV     gate3934  (.A(WX1005), .Z(WX1128) ) ;
OR2     gate3935  (.A(WX1127), .B(WX1126), .Z(WX1129) ) ;
INV     gate3936  (.A(WX1129), .Z(WX1130) ) ;
INV     gate3937  (.A(WX1005), .Z(WX1135) ) ;
OR2     gate3938  (.A(WX1134), .B(WX1133), .Z(WX1136) ) ;
INV     gate3939  (.A(WX1136), .Z(WX1137) ) ;
INV     gate3940  (.A(WX1005), .Z(WX1142) ) ;
OR2     gate3941  (.A(WX1141), .B(WX1140), .Z(WX1143) ) ;
INV     gate3942  (.A(WX1143), .Z(WX1144) ) ;
INV     gate3943  (.A(WX1005), .Z(WX1149) ) ;
OR2     gate3944  (.A(WX1148), .B(WX1147), .Z(WX1150) ) ;
INV     gate3945  (.A(WX1150), .Z(WX1151) ) ;
INV     gate3946  (.A(WX1005), .Z(WX1156) ) ;
OR2     gate3947  (.A(WX1155), .B(WX1154), .Z(WX1157) ) ;
INV     gate3948  (.A(WX1157), .Z(WX1158) ) ;
INV     gate3949  (.A(WX1005), .Z(WX1163) ) ;
OR2     gate3950  (.A(WX1162), .B(WX1161), .Z(WX1164) ) ;
INV     gate3951  (.A(WX1164), .Z(WX1165) ) ;
INV     gate3952  (.A(WX1005), .Z(WX1170) ) ;
OR2     gate3953  (.A(WX1169), .B(WX1168), .Z(WX1171) ) ;
INV     gate3954  (.A(WX1171), .Z(WX1172) ) ;
INV     gate3955  (.A(WX1005), .Z(WX1177) ) ;
OR2     gate3956  (.A(WX1176), .B(WX1175), .Z(WX1178) ) ;
INV     gate3957  (.A(WX1178), .Z(WX1179) ) ;
INV     gate3958  (.A(WX1005), .Z(WX1184) ) ;
OR2     gate3959  (.A(WX1183), .B(WX1182), .Z(WX1185) ) ;
INV     gate3960  (.A(WX1185), .Z(WX1186) ) ;
INV     gate3961  (.A(WX1005), .Z(WX1191) ) ;
OR2     gate3962  (.A(WX1190), .B(WX1189), .Z(WX1192) ) ;
INV     gate3963  (.A(WX1192), .Z(WX1193) ) ;
INV     gate3964  (.A(WX1005), .Z(WX1198) ) ;
OR2     gate3965  (.A(WX1197), .B(WX1196), .Z(WX1199) ) ;
INV     gate3966  (.A(WX1199), .Z(WX1200) ) ;
INV     gate3967  (.A(WX1005), .Z(WX1205) ) ;
OR2     gate3968  (.A(WX1204), .B(WX1203), .Z(WX1206) ) ;
INV     gate3969  (.A(WX1206), .Z(WX1207) ) ;
INV     gate3970  (.A(WX1005), .Z(WX1212) ) ;
OR2     gate3971  (.A(WX1211), .B(WX1210), .Z(WX1213) ) ;
INV     gate3972  (.A(WX1213), .Z(WX1214) ) ;
INV     gate3973  (.A(WX1005), .Z(WX1219) ) ;
OR2     gate3974  (.A(WX1218), .B(WX1217), .Z(WX1220) ) ;
INV     gate3975  (.A(WX1220), .Z(WX1221) ) ;
INV     gate3976  (.A(WX1005), .Z(WX1226) ) ;
OR2     gate3977  (.A(WX1225), .B(WX1224), .Z(WX1227) ) ;
INV     gate3978  (.A(WX1227), .Z(WX1228) ) ;
INV     gate3979  (.A(RESET), .Z(WX1230) ) ;
INV     gate3980  (.A(WX1230), .Z(WX1263) ) ;
INV     gate3981  (.A(WX2292), .Z(WX2296) ) ;
INV     gate3982  (.A(WX2296), .Z(WX1330) ) ;
INV     gate3983  (.A(WX2290), .Z(WX2297) ) ;
INV     gate3984  (.A(WX2297), .Z(WX1334) ) ;
INV     gate3985  (.A(WX2297), .Z(WX1338) ) ;
OR2     gate3986  (.A(WX1329), .B(WX1328), .Z(WX1331) ) ;
INV     gate3987  (.A(WX1331), .Z(WX1340) ) ;
INV     gate3988  (.A(WX1340), .Z(WX1341) ) ;
INV     gate3989  (.A(WX2296), .Z(WX1344) ) ;
INV     gate3990  (.A(WX2297), .Z(WX1348) ) ;
INV     gate3991  (.A(WX2297), .Z(WX1352) ) ;
OR2     gate3992  (.A(WX1343), .B(WX1342), .Z(WX1345) ) ;
INV     gate3993  (.A(WX1345), .Z(WX1354) ) ;
INV     gate3994  (.A(WX1354), .Z(WX1355) ) ;
INV     gate3995  (.A(WX2296), .Z(WX1358) ) ;
INV     gate3996  (.A(WX2297), .Z(WX1362) ) ;
INV     gate3997  (.A(WX2297), .Z(WX1366) ) ;
OR2     gate3998  (.A(WX1357), .B(WX1356), .Z(WX1359) ) ;
INV     gate3999  (.A(WX1359), .Z(WX1368) ) ;
INV     gate4000  (.A(WX1368), .Z(WX1369) ) ;
INV     gate4001  (.A(WX2296), .Z(WX1372) ) ;
INV     gate4002  (.A(WX2297), .Z(WX1376) ) ;
INV     gate4003  (.A(WX2297), .Z(WX1380) ) ;
OR2     gate4004  (.A(WX1371), .B(WX1370), .Z(WX1373) ) ;
INV     gate4005  (.A(WX1373), .Z(WX1382) ) ;
INV     gate4006  (.A(WX1382), .Z(WX1383) ) ;
INV     gate4007  (.A(WX2296), .Z(WX1386) ) ;
INV     gate4008  (.A(WX2297), .Z(WX1390) ) ;
INV     gate4009  (.A(WX2297), .Z(WX1394) ) ;
OR2     gate4010  (.A(WX1385), .B(WX1384), .Z(WX1387) ) ;
INV     gate4011  (.A(WX1387), .Z(WX1396) ) ;
INV     gate4012  (.A(WX1396), .Z(WX1397) ) ;
INV     gate4013  (.A(WX2296), .Z(WX1400) ) ;
INV     gate4014  (.A(WX2297), .Z(WX1404) ) ;
INV     gate4015  (.A(WX2297), .Z(WX1408) ) ;
OR2     gate4016  (.A(WX1399), .B(WX1398), .Z(WX1401) ) ;
INV     gate4017  (.A(WX1401), .Z(WX1410) ) ;
INV     gate4018  (.A(WX1410), .Z(WX1411) ) ;
INV     gate4019  (.A(WX2296), .Z(WX1414) ) ;
INV     gate4020  (.A(WX2297), .Z(WX1418) ) ;
INV     gate4021  (.A(WX2297), .Z(WX1422) ) ;
OR2     gate4022  (.A(WX1413), .B(WX1412), .Z(WX1415) ) ;
INV     gate4023  (.A(WX1415), .Z(WX1424) ) ;
INV     gate4024  (.A(WX1424), .Z(WX1425) ) ;
INV     gate4025  (.A(WX2296), .Z(WX1428) ) ;
INV     gate4026  (.A(WX2297), .Z(WX1432) ) ;
INV     gate4027  (.A(WX2297), .Z(WX1436) ) ;
OR2     gate4028  (.A(WX1427), .B(WX1426), .Z(WX1429) ) ;
INV     gate4029  (.A(WX1429), .Z(WX1438) ) ;
INV     gate4030  (.A(WX1438), .Z(WX1439) ) ;
INV     gate4031  (.A(WX2296), .Z(WX1442) ) ;
INV     gate4032  (.A(WX2297), .Z(WX1446) ) ;
INV     gate4033  (.A(WX2297), .Z(WX1450) ) ;
OR2     gate4034  (.A(WX1441), .B(WX1440), .Z(WX1443) ) ;
INV     gate4035  (.A(WX1443), .Z(WX1452) ) ;
INV     gate4036  (.A(WX1452), .Z(WX1453) ) ;
INV     gate4037  (.A(WX2296), .Z(WX1456) ) ;
INV     gate4038  (.A(WX2297), .Z(WX1460) ) ;
INV     gate4039  (.A(WX2297), .Z(WX1464) ) ;
OR2     gate4040  (.A(WX1455), .B(WX1454), .Z(WX1457) ) ;
INV     gate4041  (.A(WX1457), .Z(WX1466) ) ;
INV     gate4042  (.A(WX1466), .Z(WX1467) ) ;
INV     gate4043  (.A(WX2296), .Z(WX1470) ) ;
INV     gate4044  (.A(WX2297), .Z(WX1474) ) ;
INV     gate4045  (.A(WX2297), .Z(WX1478) ) ;
OR2     gate4046  (.A(WX1469), .B(WX1468), .Z(WX1471) ) ;
INV     gate4047  (.A(WX1471), .Z(WX1480) ) ;
INV     gate4048  (.A(WX1480), .Z(WX1481) ) ;
INV     gate4049  (.A(WX2296), .Z(WX1484) ) ;
INV     gate4050  (.A(WX2297), .Z(WX1488) ) ;
INV     gate4051  (.A(WX2297), .Z(WX1492) ) ;
OR2     gate4052  (.A(WX1483), .B(WX1482), .Z(WX1485) ) ;
INV     gate4053  (.A(WX1485), .Z(WX1494) ) ;
INV     gate4054  (.A(WX1494), .Z(WX1495) ) ;
INV     gate4055  (.A(WX2296), .Z(WX1498) ) ;
INV     gate4056  (.A(WX2297), .Z(WX1502) ) ;
INV     gate4057  (.A(WX2297), .Z(WX1506) ) ;
OR2     gate4058  (.A(WX1497), .B(WX1496), .Z(WX1499) ) ;
INV     gate4059  (.A(WX1499), .Z(WX1508) ) ;
INV     gate4060  (.A(WX1508), .Z(WX1509) ) ;
INV     gate4061  (.A(WX2296), .Z(WX1512) ) ;
INV     gate4062  (.A(WX2297), .Z(WX1516) ) ;
INV     gate4063  (.A(WX2297), .Z(WX1520) ) ;
OR2     gate4064  (.A(WX1511), .B(WX1510), .Z(WX1513) ) ;
INV     gate4065  (.A(WX1513), .Z(WX1522) ) ;
INV     gate4066  (.A(WX1522), .Z(WX1523) ) ;
INV     gate4067  (.A(WX2296), .Z(WX1526) ) ;
INV     gate4068  (.A(WX2297), .Z(WX1530) ) ;
INV     gate4069  (.A(WX2297), .Z(WX1534) ) ;
OR2     gate4070  (.A(WX1525), .B(WX1524), .Z(WX1527) ) ;
INV     gate4071  (.A(WX1527), .Z(WX1536) ) ;
INV     gate4072  (.A(WX1536), .Z(WX1537) ) ;
INV     gate4073  (.A(WX2296), .Z(WX1540) ) ;
INV     gate4074  (.A(WX2297), .Z(WX1544) ) ;
INV     gate4075  (.A(WX2297), .Z(WX1548) ) ;
OR2     gate4076  (.A(WX1539), .B(WX1538), .Z(WX1541) ) ;
INV     gate4077  (.A(WX1541), .Z(WX1550) ) ;
INV     gate4078  (.A(WX1550), .Z(WX1551) ) ;
INV     gate4079  (.A(WX2296), .Z(WX1554) ) ;
INV     gate4080  (.A(WX2297), .Z(WX1558) ) ;
INV     gate4081  (.A(WX2297), .Z(WX1562) ) ;
OR2     gate4082  (.A(WX1553), .B(WX1552), .Z(WX1555) ) ;
INV     gate4083  (.A(WX1555), .Z(WX1564) ) ;
INV     gate4084  (.A(WX1564), .Z(WX1565) ) ;
INV     gate4085  (.A(WX2296), .Z(WX1568) ) ;
INV     gate4086  (.A(WX2297), .Z(WX1572) ) ;
INV     gate4087  (.A(WX2297), .Z(WX1576) ) ;
OR2     gate4088  (.A(WX1567), .B(WX1566), .Z(WX1569) ) ;
INV     gate4089  (.A(WX1569), .Z(WX1578) ) ;
INV     gate4090  (.A(WX1578), .Z(WX1579) ) ;
INV     gate4091  (.A(WX2296), .Z(WX1582) ) ;
INV     gate4092  (.A(WX2297), .Z(WX1586) ) ;
INV     gate4093  (.A(WX2297), .Z(WX1590) ) ;
OR2     gate4094  (.A(WX1581), .B(WX1580), .Z(WX1583) ) ;
INV     gate4095  (.A(WX1583), .Z(WX1592) ) ;
INV     gate4096  (.A(WX1592), .Z(WX1593) ) ;
INV     gate4097  (.A(WX2296), .Z(WX1596) ) ;
INV     gate4098  (.A(WX2297), .Z(WX1600) ) ;
INV     gate4099  (.A(WX2297), .Z(WX1604) ) ;
OR2     gate4100  (.A(WX1595), .B(WX1594), .Z(WX1597) ) ;
INV     gate4101  (.A(WX1597), .Z(WX1606) ) ;
INV     gate4102  (.A(WX1606), .Z(WX1607) ) ;
INV     gate4103  (.A(WX2296), .Z(WX1610) ) ;
INV     gate4104  (.A(WX2297), .Z(WX1614) ) ;
INV     gate4105  (.A(WX2297), .Z(WX1618) ) ;
OR2     gate4106  (.A(WX1609), .B(WX1608), .Z(WX1611) ) ;
INV     gate4107  (.A(WX1611), .Z(WX1620) ) ;
INV     gate4108  (.A(WX1620), .Z(WX1621) ) ;
INV     gate4109  (.A(WX2296), .Z(WX1624) ) ;
INV     gate4110  (.A(WX2297), .Z(WX1628) ) ;
INV     gate4111  (.A(WX2297), .Z(WX1632) ) ;
OR2     gate4112  (.A(WX1623), .B(WX1622), .Z(WX1625) ) ;
INV     gate4113  (.A(WX1625), .Z(WX1634) ) ;
INV     gate4114  (.A(WX1634), .Z(WX1635) ) ;
INV     gate4115  (.A(WX2296), .Z(WX1638) ) ;
INV     gate4116  (.A(WX2297), .Z(WX1642) ) ;
INV     gate4117  (.A(WX2297), .Z(WX1646) ) ;
OR2     gate4118  (.A(WX1637), .B(WX1636), .Z(WX1639) ) ;
INV     gate4119  (.A(WX1639), .Z(WX1648) ) ;
INV     gate4120  (.A(WX1648), .Z(WX1649) ) ;
INV     gate4121  (.A(WX2296), .Z(WX1652) ) ;
INV     gate4122  (.A(WX2297), .Z(WX1656) ) ;
INV     gate4123  (.A(WX2297), .Z(WX1660) ) ;
OR2     gate4124  (.A(WX1651), .B(WX1650), .Z(WX1653) ) ;
INV     gate4125  (.A(WX1653), .Z(WX1662) ) ;
INV     gate4126  (.A(WX1662), .Z(WX1663) ) ;
INV     gate4127  (.A(WX2296), .Z(WX1666) ) ;
INV     gate4128  (.A(WX2297), .Z(WX1670) ) ;
INV     gate4129  (.A(WX2297), .Z(WX1674) ) ;
OR2     gate4130  (.A(WX1665), .B(WX1664), .Z(WX1667) ) ;
INV     gate4131  (.A(WX1667), .Z(WX1676) ) ;
INV     gate4132  (.A(WX1676), .Z(WX1677) ) ;
INV     gate4133  (.A(WX2296), .Z(WX1680) ) ;
INV     gate4134  (.A(WX2297), .Z(WX1684) ) ;
INV     gate4135  (.A(WX2297), .Z(WX1688) ) ;
OR2     gate4136  (.A(WX1679), .B(WX1678), .Z(WX1681) ) ;
INV     gate4137  (.A(WX1681), .Z(WX1690) ) ;
INV     gate4138  (.A(WX1690), .Z(WX1691) ) ;
INV     gate4139  (.A(WX2296), .Z(WX1694) ) ;
INV     gate4140  (.A(WX2297), .Z(WX1698) ) ;
INV     gate4141  (.A(WX2297), .Z(WX1702) ) ;
OR2     gate4142  (.A(WX1693), .B(WX1692), .Z(WX1695) ) ;
INV     gate4143  (.A(WX1695), .Z(WX1704) ) ;
INV     gate4144  (.A(WX1704), .Z(WX1705) ) ;
INV     gate4145  (.A(WX2296), .Z(WX1708) ) ;
INV     gate4146  (.A(WX2297), .Z(WX1712) ) ;
INV     gate4147  (.A(WX2297), .Z(WX1716) ) ;
OR2     gate4148  (.A(WX1707), .B(WX1706), .Z(WX1709) ) ;
INV     gate4149  (.A(WX1709), .Z(WX1718) ) ;
INV     gate4150  (.A(WX1718), .Z(WX1719) ) ;
INV     gate4151  (.A(WX2296), .Z(WX1722) ) ;
INV     gate4152  (.A(WX2297), .Z(WX1726) ) ;
INV     gate4153  (.A(WX2297), .Z(WX1730) ) ;
OR2     gate4154  (.A(WX1721), .B(WX1720), .Z(WX1723) ) ;
INV     gate4155  (.A(WX1723), .Z(WX1732) ) ;
INV     gate4156  (.A(WX1732), .Z(WX1733) ) ;
INV     gate4157  (.A(WX2296), .Z(WX1736) ) ;
INV     gate4158  (.A(WX2297), .Z(WX1740) ) ;
INV     gate4159  (.A(WX2297), .Z(WX1744) ) ;
OR2     gate4160  (.A(WX1735), .B(WX1734), .Z(WX1737) ) ;
INV     gate4161  (.A(WX1737), .Z(WX1746) ) ;
INV     gate4162  (.A(WX1746), .Z(WX1747) ) ;
INV     gate4163  (.A(WX2296), .Z(WX1750) ) ;
INV     gate4164  (.A(WX2297), .Z(WX1754) ) ;
INV     gate4165  (.A(WX2297), .Z(WX1758) ) ;
OR2     gate4166  (.A(WX1749), .B(WX1748), .Z(WX1751) ) ;
INV     gate4167  (.A(WX1751), .Z(WX1760) ) ;
INV     gate4168  (.A(WX1760), .Z(WX1761) ) ;
INV     gate4169  (.A(WX2296), .Z(WX1764) ) ;
INV     gate4170  (.A(WX2297), .Z(WX1768) ) ;
INV     gate4171  (.A(WX2297), .Z(WX1772) ) ;
OR2     gate4172  (.A(WX1763), .B(WX1762), .Z(WX1765) ) ;
INV     gate4173  (.A(WX1765), .Z(WX1774) ) ;
INV     gate4174  (.A(WX1774), .Z(WX1775) ) ;
INV     gate4175  (.A(WX1778), .Z(WX1776) ) ;
INV     gate4176  (.A(WX2257), .Z(WX2258) ) ;
INV     gate4177  (.A(WX2258), .Z(WX1841) ) ;
INV     gate4178  (.A(WX2259), .Z(WX2260) ) ;
INV     gate4179  (.A(WX2260), .Z(WX1842) ) ;
INV     gate4180  (.A(WX2261), .Z(WX2262) ) ;
INV     gate4181  (.A(WX2262), .Z(WX1843) ) ;
INV     gate4182  (.A(WX2263), .Z(WX2264) ) ;
INV     gate4183  (.A(WX2264), .Z(WX1844) ) ;
INV     gate4184  (.A(WX2265), .Z(WX2266) ) ;
INV     gate4185  (.A(WX2266), .Z(WX1845) ) ;
INV     gate4186  (.A(WX2267), .Z(WX2268) ) ;
INV     gate4187  (.A(WX2268), .Z(WX1846) ) ;
INV     gate4188  (.A(WX2269), .Z(WX2270) ) ;
INV     gate4189  (.A(WX2270), .Z(WX1847) ) ;
INV     gate4190  (.A(WX2271), .Z(WX2272) ) ;
INV     gate4191  (.A(WX2272), .Z(WX1848) ) ;
INV     gate4192  (.A(WX2273), .Z(WX2274) ) ;
INV     gate4193  (.A(WX2274), .Z(WX1849) ) ;
INV     gate4194  (.A(WX2275), .Z(WX2276) ) ;
INV     gate4195  (.A(WX2276), .Z(WX1850) ) ;
INV     gate4196  (.A(WX2277), .Z(WX2278) ) ;
INV     gate4197  (.A(WX2278), .Z(WX1851) ) ;
INV     gate4198  (.A(WX2279), .Z(WX2280) ) ;
INV     gate4199  (.A(WX2280), .Z(WX1852) ) ;
INV     gate4200  (.A(WX2281), .Z(WX2282) ) ;
INV     gate4201  (.A(WX2282), .Z(WX1853) ) ;
INV     gate4202  (.A(WX2283), .Z(WX2284) ) ;
INV     gate4203  (.A(WX2284), .Z(WX1854) ) ;
INV     gate4204  (.A(WX2285), .Z(WX2286) ) ;
INV     gate4205  (.A(WX2286), .Z(WX1855) ) ;
INV     gate4206  (.A(WX2287), .Z(WX2288) ) ;
INV     gate4207  (.A(WX2288), .Z(WX1856) ) ;
INV     gate4208  (.A(WX2225), .Z(WX2226) ) ;
INV     gate4209  (.A(WX2226), .Z(WX1857) ) ;
INV     gate4210  (.A(WX2227), .Z(WX2228) ) ;
INV     gate4211  (.A(WX2228), .Z(WX1858) ) ;
INV     gate4212  (.A(WX2229), .Z(WX2230) ) ;
INV     gate4213  (.A(WX2230), .Z(WX1859) ) ;
INV     gate4214  (.A(WX2231), .Z(WX2232) ) ;
INV     gate4215  (.A(WX2232), .Z(WX1860) ) ;
INV     gate4216  (.A(WX2233), .Z(WX2234) ) ;
INV     gate4217  (.A(WX2234), .Z(WX1861) ) ;
INV     gate4218  (.A(WX2235), .Z(WX2236) ) ;
INV     gate4219  (.A(WX2236), .Z(WX1862) ) ;
INV     gate4220  (.A(WX2237), .Z(WX2238) ) ;
INV     gate4221  (.A(WX2238), .Z(WX1863) ) ;
INV     gate4222  (.A(WX2239), .Z(WX2240) ) ;
INV     gate4223  (.A(WX2240), .Z(WX1864) ) ;
INV     gate4224  (.A(WX2241), .Z(WX2242) ) ;
INV     gate4225  (.A(WX2242), .Z(WX1865) ) ;
INV     gate4226  (.A(WX2243), .Z(WX2244) ) ;
INV     gate4227  (.A(WX2244), .Z(WX1866) ) ;
INV     gate4228  (.A(WX2245), .Z(WX2246) ) ;
INV     gate4229  (.A(WX2246), .Z(WX1867) ) ;
INV     gate4230  (.A(WX2247), .Z(WX2248) ) ;
INV     gate4231  (.A(WX2248), .Z(WX1868) ) ;
INV     gate4232  (.A(WX2249), .Z(WX2250) ) ;
INV     gate4233  (.A(WX2250), .Z(WX1869) ) ;
INV     gate4234  (.A(WX2251), .Z(WX2252) ) ;
INV     gate4235  (.A(WX2252), .Z(WX1870) ) ;
INV     gate4236  (.A(WX2253), .Z(WX2254) ) ;
INV     gate4237  (.A(WX2254), .Z(WX1871) ) ;
INV     gate4238  (.A(WX2255), .Z(WX2256) ) ;
INV     gate4239  (.A(WX2256), .Z(WX1872) ) ;
INV     gate4240  (.A(WX1841), .Z(WX1873) ) ;
INV     gate4241  (.A(WX1842), .Z(WX1874) ) ;
INV     gate4242  (.A(WX1843), .Z(WX1875) ) ;
INV     gate4243  (.A(WX1844), .Z(WX1876) ) ;
INV     gate4244  (.A(WX1845), .Z(WX1877) ) ;
INV     gate4245  (.A(WX1846), .Z(WX1878) ) ;
INV     gate4246  (.A(WX1847), .Z(WX1879) ) ;
INV     gate4247  (.A(WX1848), .Z(WX1880) ) ;
INV     gate4248  (.A(WX1849), .Z(WX1881) ) ;
INV     gate4249  (.A(WX1850), .Z(WX1882) ) ;
INV     gate4250  (.A(WX1851), .Z(WX1883) ) ;
INV     gate4251  (.A(WX1852), .Z(WX1884) ) ;
INV     gate4252  (.A(WX1853), .Z(WX1885) ) ;
INV     gate4253  (.A(WX1854), .Z(WX1886) ) ;
INV     gate4254  (.A(WX1855), .Z(WX1887) ) ;
INV     gate4255  (.A(WX1856), .Z(WX1888) ) ;
INV     gate4256  (.A(WX1857), .Z(WX1889) ) ;
INV     gate4257  (.A(WX1858), .Z(WX1890) ) ;
INV     gate4258  (.A(WX1859), .Z(WX1891) ) ;
INV     gate4259  (.A(WX1860), .Z(WX1892) ) ;
INV     gate4260  (.A(WX1861), .Z(WX1893) ) ;
INV     gate4261  (.A(WX1862), .Z(WX1894) ) ;
INV     gate4262  (.A(WX1863), .Z(WX1895) ) ;
INV     gate4263  (.A(WX1864), .Z(WX1896) ) ;
INV     gate4264  (.A(WX1865), .Z(WX1897) ) ;
INV     gate4265  (.A(WX1866), .Z(WX1898) ) ;
INV     gate4266  (.A(WX1867), .Z(WX1899) ) ;
INV     gate4267  (.A(WX1868), .Z(WX1900) ) ;
INV     gate4268  (.A(WX1869), .Z(WX1901) ) ;
INV     gate4269  (.A(WX1870), .Z(WX1902) ) ;
INV     gate4270  (.A(WX1871), .Z(WX1903) ) ;
INV     gate4271  (.A(WX1872), .Z(WX1904) ) ;
INV     gate4272  (.A(WX2130), .Z(WX1905) ) ;
INV     gate4273  (.A(WX2132), .Z(WX1906) ) ;
INV     gate4274  (.A(WX2134), .Z(WX1907) ) ;
INV     gate4275  (.A(WX2136), .Z(WX1908) ) ;
INV     gate4276  (.A(WX2138), .Z(WX1909) ) ;
INV     gate4277  (.A(WX2140), .Z(WX1910) ) ;
INV     gate4278  (.A(WX2142), .Z(WX1911) ) ;
INV     gate4279  (.A(WX2144), .Z(WX1912) ) ;
INV     gate4280  (.A(WX2146), .Z(WX1913) ) ;
INV     gate4281  (.A(WX2148), .Z(WX1914) ) ;
INV     gate4282  (.A(WX2150), .Z(WX1915) ) ;
INV     gate4283  (.A(WX2152), .Z(WX1916) ) ;
INV     gate4284  (.A(WX2154), .Z(WX1917) ) ;
INV     gate4285  (.A(WX2156), .Z(WX1918) ) ;
INV     gate4286  (.A(WX2158), .Z(WX1919) ) ;
INV     gate4287  (.A(WX2160), .Z(WX1920) ) ;
INV     gate4288  (.A(WX2162), .Z(WX1921) ) ;
INV     gate4289  (.A(WX2164), .Z(WX1922) ) ;
INV     gate4290  (.A(WX2166), .Z(WX1923) ) ;
INV     gate4291  (.A(WX2168), .Z(WX1924) ) ;
INV     gate4292  (.A(WX2170), .Z(WX1925) ) ;
INV     gate4293  (.A(WX2172), .Z(WX1926) ) ;
INV     gate4294  (.A(WX2174), .Z(WX1927) ) ;
INV     gate4295  (.A(WX2176), .Z(WX1928) ) ;
INV     gate4296  (.A(WX2178), .Z(WX1929) ) ;
INV     gate4297  (.A(WX2180), .Z(WX1930) ) ;
INV     gate4298  (.A(WX2182), .Z(WX1931) ) ;
INV     gate4299  (.A(WX2184), .Z(WX1932) ) ;
INV     gate4300  (.A(WX2186), .Z(WX1933) ) ;
INV     gate4301  (.A(WX2188), .Z(WX1934) ) ;
INV     gate4302  (.A(WX2190), .Z(WX1935) ) ;
INV     gate4303  (.A(WX2192), .Z(WX1936) ) ;
NAND2   gate4304  (.A(II6512), .B(II6513), .Z(WX2209) ) ;
INV     gate4305  (.A(WX2209), .Z(WX2225) ) ;
NAND2   gate4306  (.A(II6543), .B(II6544), .Z(WX2210) ) ;
INV     gate4307  (.A(WX2210), .Z(WX2227) ) ;
NAND2   gate4308  (.A(II6574), .B(II6575), .Z(WX2211) ) ;
INV     gate4309  (.A(WX2211), .Z(WX2229) ) ;
NAND2   gate4310  (.A(II6605), .B(II6606), .Z(WX2212) ) ;
INV     gate4311  (.A(WX2212), .Z(WX2231) ) ;
NAND2   gate4312  (.A(II6636), .B(II6637), .Z(WX2213) ) ;
INV     gate4313  (.A(WX2213), .Z(WX2233) ) ;
NAND2   gate4314  (.A(II6667), .B(II6668), .Z(WX2214) ) ;
INV     gate4315  (.A(WX2214), .Z(WX2235) ) ;
NAND2   gate4316  (.A(II6698), .B(II6699), .Z(WX2215) ) ;
INV     gate4317  (.A(WX2215), .Z(WX2237) ) ;
NAND2   gate4318  (.A(II6729), .B(II6730), .Z(WX2216) ) ;
INV     gate4319  (.A(WX2216), .Z(WX2239) ) ;
NAND2   gate4320  (.A(II6760), .B(II6761), .Z(WX2217) ) ;
INV     gate4321  (.A(WX2217), .Z(WX2241) ) ;
NAND2   gate4322  (.A(II6791), .B(II6792), .Z(WX2218) ) ;
INV     gate4323  (.A(WX2218), .Z(WX2243) ) ;
NAND2   gate4324  (.A(II6822), .B(II6823), .Z(WX2219) ) ;
INV     gate4325  (.A(WX2219), .Z(WX2245) ) ;
NAND2   gate4326  (.A(II6853), .B(II6854), .Z(WX2220) ) ;
INV     gate4327  (.A(WX2220), .Z(WX2247) ) ;
NAND2   gate4328  (.A(II6884), .B(II6885), .Z(WX2221) ) ;
INV     gate4329  (.A(WX2221), .Z(WX2249) ) ;
NAND2   gate4330  (.A(II6915), .B(II6916), .Z(WX2222) ) ;
INV     gate4331  (.A(WX2222), .Z(WX2251) ) ;
NAND2   gate4332  (.A(II6946), .B(II6947), .Z(WX2223) ) ;
INV     gate4333  (.A(WX2223), .Z(WX2253) ) ;
NAND2   gate4334  (.A(II6977), .B(II6978), .Z(WX2224) ) ;
INV     gate4335  (.A(WX2224), .Z(WX2255) ) ;
NAND2   gate4336  (.A(II6016), .B(II6017), .Z(WX2193) ) ;
INV     gate4337  (.A(WX2193), .Z(WX2257) ) ;
NAND2   gate4338  (.A(II6047), .B(II6048), .Z(WX2194) ) ;
INV     gate4339  (.A(WX2194), .Z(WX2259) ) ;
NAND2   gate4340  (.A(II6078), .B(II6079), .Z(WX2195) ) ;
INV     gate4341  (.A(WX2195), .Z(WX2261) ) ;
NAND2   gate4342  (.A(II6109), .B(II6110), .Z(WX2196) ) ;
INV     gate4343  (.A(WX2196), .Z(WX2263) ) ;
NAND2   gate4344  (.A(II6140), .B(II6141), .Z(WX2197) ) ;
INV     gate4345  (.A(WX2197), .Z(WX2265) ) ;
NAND2   gate4346  (.A(II6171), .B(II6172), .Z(WX2198) ) ;
INV     gate4347  (.A(WX2198), .Z(WX2267) ) ;
NAND2   gate4348  (.A(II6202), .B(II6203), .Z(WX2199) ) ;
INV     gate4349  (.A(WX2199), .Z(WX2269) ) ;
NAND2   gate4350  (.A(II6233), .B(II6234), .Z(WX2200) ) ;
INV     gate4351  (.A(WX2200), .Z(WX2271) ) ;
NAND2   gate4352  (.A(II6264), .B(II6265), .Z(WX2201) ) ;
INV     gate4353  (.A(WX2201), .Z(WX2273) ) ;
NAND2   gate4354  (.A(II6295), .B(II6296), .Z(WX2202) ) ;
INV     gate4355  (.A(WX2202), .Z(WX2275) ) ;
NAND2   gate4356  (.A(II6326), .B(II6327), .Z(WX2203) ) ;
INV     gate4357  (.A(WX2203), .Z(WX2277) ) ;
NAND2   gate4358  (.A(II6357), .B(II6358), .Z(WX2204) ) ;
INV     gate4359  (.A(WX2204), .Z(WX2279) ) ;
NAND2   gate4360  (.A(II6388), .B(II6389), .Z(WX2205) ) ;
INV     gate4361  (.A(WX2205), .Z(WX2281) ) ;
NAND2   gate4362  (.A(II6419), .B(II6420), .Z(WX2206) ) ;
INV     gate4363  (.A(WX2206), .Z(WX2283) ) ;
NAND2   gate4364  (.A(II6450), .B(II6451), .Z(WX2207) ) ;
INV     gate4365  (.A(WX2207), .Z(WX2285) ) ;
NAND2   gate4366  (.A(II6481), .B(II6482), .Z(WX2208) ) ;
INV     gate4367  (.A(WX2208), .Z(WX2287) ) ;
INV     gate4368  (.A(TM0), .Z(WX2289) ) ;
INV     gate4369  (.A(TM0), .Z(WX2290) ) ;
INV     gate4370  (.A(TM0), .Z(WX2291) ) ;
INV     gate4371  (.A(TM1), .Z(WX2292) ) ;
INV     gate4372  (.A(TM1), .Z(WX2293) ) ;
INV     gate4373  (.A(WX2293), .Z(WX2294) ) ;
INV     gate4374  (.A(WX2291), .Z(WX2295) ) ;
INV     gate4375  (.A(WX2289), .Z(WX2298) ) ;
INV     gate4376  (.A(WX2298), .Z(WX2302) ) ;
OR2     gate4377  (.A(WX2301), .B(WX2300), .Z(WX2303) ) ;
INV     gate4378  (.A(WX2303), .Z(WX2304) ) ;
INV     gate4379  (.A(WX2304), .Z(WX2305) ) ;
INV     gate4380  (.A(WX2298), .Z(WX2309) ) ;
OR2     gate4381  (.A(WX2308), .B(WX2307), .Z(WX2310) ) ;
INV     gate4382  (.A(WX2310), .Z(WX2311) ) ;
INV     gate4383  (.A(WX2311), .Z(WX2312) ) ;
INV     gate4384  (.A(WX2298), .Z(WX2316) ) ;
OR2     gate4385  (.A(WX2315), .B(WX2314), .Z(WX2317) ) ;
INV     gate4386  (.A(WX2317), .Z(WX2318) ) ;
INV     gate4387  (.A(WX2318), .Z(WX2319) ) ;
INV     gate4388  (.A(WX2298), .Z(WX2323) ) ;
OR2     gate4389  (.A(WX2322), .B(WX2321), .Z(WX2324) ) ;
INV     gate4390  (.A(WX2324), .Z(WX2325) ) ;
INV     gate4391  (.A(WX2325), .Z(WX2326) ) ;
INV     gate4392  (.A(WX2298), .Z(WX2330) ) ;
OR2     gate4393  (.A(WX2329), .B(WX2328), .Z(WX2331) ) ;
INV     gate4394  (.A(WX2331), .Z(WX2332) ) ;
INV     gate4395  (.A(WX2332), .Z(WX2333) ) ;
INV     gate4396  (.A(WX2298), .Z(WX2337) ) ;
OR2     gate4397  (.A(WX2336), .B(WX2335), .Z(WX2338) ) ;
INV     gate4398  (.A(WX2338), .Z(WX2339) ) ;
INV     gate4399  (.A(WX2339), .Z(WX2340) ) ;
INV     gate4400  (.A(WX2298), .Z(WX2344) ) ;
OR2     gate4401  (.A(WX2343), .B(WX2342), .Z(WX2345) ) ;
INV     gate4402  (.A(WX2345), .Z(WX2346) ) ;
INV     gate4403  (.A(WX2346), .Z(WX2347) ) ;
INV     gate4404  (.A(WX2298), .Z(WX2351) ) ;
OR2     gate4405  (.A(WX2350), .B(WX2349), .Z(WX2352) ) ;
INV     gate4406  (.A(WX2352), .Z(WX2353) ) ;
INV     gate4407  (.A(WX2353), .Z(WX2354) ) ;
INV     gate4408  (.A(WX2298), .Z(WX2358) ) ;
OR2     gate4409  (.A(WX2357), .B(WX2356), .Z(WX2359) ) ;
INV     gate4410  (.A(WX2359), .Z(WX2360) ) ;
INV     gate4411  (.A(WX2360), .Z(WX2361) ) ;
INV     gate4412  (.A(WX2298), .Z(WX2365) ) ;
OR2     gate4413  (.A(WX2364), .B(WX2363), .Z(WX2366) ) ;
INV     gate4414  (.A(WX2366), .Z(WX2367) ) ;
INV     gate4415  (.A(WX2367), .Z(WX2368) ) ;
INV     gate4416  (.A(WX2298), .Z(WX2372) ) ;
OR2     gate4417  (.A(WX2371), .B(WX2370), .Z(WX2373) ) ;
INV     gate4418  (.A(WX2373), .Z(WX2374) ) ;
INV     gate4419  (.A(WX2374), .Z(WX2375) ) ;
INV     gate4420  (.A(WX2298), .Z(WX2379) ) ;
OR2     gate4421  (.A(WX2378), .B(WX2377), .Z(WX2380) ) ;
INV     gate4422  (.A(WX2380), .Z(WX2381) ) ;
INV     gate4423  (.A(WX2381), .Z(WX2382) ) ;
INV     gate4424  (.A(WX2298), .Z(WX2386) ) ;
OR2     gate4425  (.A(WX2385), .B(WX2384), .Z(WX2387) ) ;
INV     gate4426  (.A(WX2387), .Z(WX2388) ) ;
INV     gate4427  (.A(WX2388), .Z(WX2389) ) ;
INV     gate4428  (.A(WX2298), .Z(WX2393) ) ;
OR2     gate4429  (.A(WX2392), .B(WX2391), .Z(WX2394) ) ;
INV     gate4430  (.A(WX2394), .Z(WX2395) ) ;
INV     gate4431  (.A(WX2395), .Z(WX2396) ) ;
INV     gate4432  (.A(WX2298), .Z(WX2400) ) ;
OR2     gate4433  (.A(WX2399), .B(WX2398), .Z(WX2401) ) ;
INV     gate4434  (.A(WX2401), .Z(WX2402) ) ;
INV     gate4435  (.A(WX2402), .Z(WX2403) ) ;
INV     gate4436  (.A(WX2298), .Z(WX2407) ) ;
OR2     gate4437  (.A(WX2406), .B(WX2405), .Z(WX2408) ) ;
INV     gate4438  (.A(WX2408), .Z(WX2409) ) ;
INV     gate4439  (.A(WX2409), .Z(WX2410) ) ;
INV     gate4440  (.A(WX2298), .Z(WX2414) ) ;
OR2     gate4441  (.A(WX2413), .B(WX2412), .Z(WX2415) ) ;
INV     gate4442  (.A(WX2415), .Z(WX2416) ) ;
INV     gate4443  (.A(WX2416), .Z(WX2417) ) ;
INV     gate4444  (.A(WX2298), .Z(WX2421) ) ;
OR2     gate4445  (.A(WX2420), .B(WX2419), .Z(WX2422) ) ;
INV     gate4446  (.A(WX2422), .Z(WX2423) ) ;
INV     gate4447  (.A(WX2423), .Z(WX2424) ) ;
INV     gate4448  (.A(WX2298), .Z(WX2428) ) ;
OR2     gate4449  (.A(WX2427), .B(WX2426), .Z(WX2429) ) ;
INV     gate4450  (.A(WX2429), .Z(WX2430) ) ;
INV     gate4451  (.A(WX2430), .Z(WX2431) ) ;
INV     gate4452  (.A(WX2298), .Z(WX2435) ) ;
OR2     gate4453  (.A(WX2434), .B(WX2433), .Z(WX2436) ) ;
INV     gate4454  (.A(WX2436), .Z(WX2437) ) ;
INV     gate4455  (.A(WX2437), .Z(WX2438) ) ;
INV     gate4456  (.A(WX2298), .Z(WX2442) ) ;
OR2     gate4457  (.A(WX2441), .B(WX2440), .Z(WX2443) ) ;
INV     gate4458  (.A(WX2443), .Z(WX2444) ) ;
INV     gate4459  (.A(WX2444), .Z(WX2445) ) ;
INV     gate4460  (.A(WX2298), .Z(WX2449) ) ;
OR2     gate4461  (.A(WX2448), .B(WX2447), .Z(WX2450) ) ;
INV     gate4462  (.A(WX2450), .Z(WX2451) ) ;
INV     gate4463  (.A(WX2451), .Z(WX2452) ) ;
INV     gate4464  (.A(WX2298), .Z(WX2456) ) ;
OR2     gate4465  (.A(WX2455), .B(WX2454), .Z(WX2457) ) ;
INV     gate4466  (.A(WX2457), .Z(WX2458) ) ;
INV     gate4467  (.A(WX2458), .Z(WX2459) ) ;
INV     gate4468  (.A(WX2298), .Z(WX2463) ) ;
OR2     gate4469  (.A(WX2462), .B(WX2461), .Z(WX2464) ) ;
INV     gate4470  (.A(WX2464), .Z(WX2465) ) ;
INV     gate4471  (.A(WX2465), .Z(WX2466) ) ;
INV     gate4472  (.A(WX2298), .Z(WX2470) ) ;
OR2     gate4473  (.A(WX2469), .B(WX2468), .Z(WX2471) ) ;
INV     gate4474  (.A(WX2471), .Z(WX2472) ) ;
INV     gate4475  (.A(WX2472), .Z(WX2473) ) ;
INV     gate4476  (.A(WX2298), .Z(WX2477) ) ;
OR2     gate4477  (.A(WX2476), .B(WX2475), .Z(WX2478) ) ;
INV     gate4478  (.A(WX2478), .Z(WX2479) ) ;
INV     gate4479  (.A(WX2479), .Z(WX2480) ) ;
INV     gate4480  (.A(WX2298), .Z(WX2484) ) ;
OR2     gate4481  (.A(WX2483), .B(WX2482), .Z(WX2485) ) ;
INV     gate4482  (.A(WX2485), .Z(WX2486) ) ;
INV     gate4483  (.A(WX2486), .Z(WX2487) ) ;
INV     gate4484  (.A(WX2298), .Z(WX2491) ) ;
OR2     gate4485  (.A(WX2490), .B(WX2489), .Z(WX2492) ) ;
INV     gate4486  (.A(WX2492), .Z(WX2493) ) ;
INV     gate4487  (.A(WX2493), .Z(WX2494) ) ;
INV     gate4488  (.A(WX2298), .Z(WX2498) ) ;
OR2     gate4489  (.A(WX2497), .B(WX2496), .Z(WX2499) ) ;
INV     gate4490  (.A(WX2499), .Z(WX2500) ) ;
INV     gate4491  (.A(WX2500), .Z(WX2501) ) ;
INV     gate4492  (.A(WX2298), .Z(WX2505) ) ;
OR2     gate4493  (.A(WX2504), .B(WX2503), .Z(WX2506) ) ;
INV     gate4494  (.A(WX2506), .Z(WX2507) ) ;
INV     gate4495  (.A(WX2507), .Z(WX2508) ) ;
INV     gate4496  (.A(WX2298), .Z(WX2512) ) ;
OR2     gate4497  (.A(WX2511), .B(WX2510), .Z(WX2513) ) ;
INV     gate4498  (.A(WX2513), .Z(WX2514) ) ;
INV     gate4499  (.A(WX2514), .Z(WX2515) ) ;
INV     gate4500  (.A(WX2298), .Z(WX2519) ) ;
OR2     gate4501  (.A(WX2518), .B(WX2517), .Z(WX2520) ) ;
INV     gate4502  (.A(WX2520), .Z(WX2521) ) ;
INV     gate4503  (.A(WX2521), .Z(WX2522) ) ;
INV     gate4504  (.A(RESET), .Z(WX2523) ) ;
INV     gate4505  (.A(WX2523), .Z(WX2556) ) ;
INV     gate4506  (.A(WX3585), .Z(WX3589) ) ;
INV     gate4507  (.A(WX3589), .Z(WX2623) ) ;
INV     gate4508  (.A(WX3583), .Z(WX3590) ) ;
INV     gate4509  (.A(WX3590), .Z(WX2627) ) ;
INV     gate4510  (.A(WX3590), .Z(WX2631) ) ;
OR2     gate4511  (.A(WX2622), .B(WX2621), .Z(WX2624) ) ;
INV     gate4512  (.A(WX2624), .Z(WX2633) ) ;
INV     gate4513  (.A(WX2633), .Z(WX2634) ) ;
INV     gate4514  (.A(WX3589), .Z(WX2637) ) ;
INV     gate4515  (.A(WX3590), .Z(WX2641) ) ;
INV     gate4516  (.A(WX3590), .Z(WX2645) ) ;
OR2     gate4517  (.A(WX2636), .B(WX2635), .Z(WX2638) ) ;
INV     gate4518  (.A(WX2638), .Z(WX2647) ) ;
INV     gate4519  (.A(WX2647), .Z(WX2648) ) ;
INV     gate4520  (.A(WX3589), .Z(WX2651) ) ;
INV     gate4521  (.A(WX3590), .Z(WX2655) ) ;
INV     gate4522  (.A(WX3590), .Z(WX2659) ) ;
OR2     gate4523  (.A(WX2650), .B(WX2649), .Z(WX2652) ) ;
INV     gate4524  (.A(WX2652), .Z(WX2661) ) ;
INV     gate4525  (.A(WX2661), .Z(WX2662) ) ;
INV     gate4526  (.A(WX3589), .Z(WX2665) ) ;
INV     gate4527  (.A(WX3590), .Z(WX2669) ) ;
INV     gate4528  (.A(WX3590), .Z(WX2673) ) ;
OR2     gate4529  (.A(WX2664), .B(WX2663), .Z(WX2666) ) ;
INV     gate4530  (.A(WX2666), .Z(WX2675) ) ;
INV     gate4531  (.A(WX2675), .Z(WX2676) ) ;
INV     gate4532  (.A(WX3589), .Z(WX2679) ) ;
INV     gate4533  (.A(WX3590), .Z(WX2683) ) ;
INV     gate4534  (.A(WX3590), .Z(WX2687) ) ;
OR2     gate4535  (.A(WX2678), .B(WX2677), .Z(WX2680) ) ;
INV     gate4536  (.A(WX2680), .Z(WX2689) ) ;
INV     gate4537  (.A(WX2689), .Z(WX2690) ) ;
INV     gate4538  (.A(WX3589), .Z(WX2693) ) ;
INV     gate4539  (.A(WX3590), .Z(WX2697) ) ;
INV     gate4540  (.A(WX3590), .Z(WX2701) ) ;
OR2     gate4541  (.A(WX2692), .B(WX2691), .Z(WX2694) ) ;
INV     gate4542  (.A(WX2694), .Z(WX2703) ) ;
INV     gate4543  (.A(WX2703), .Z(WX2704) ) ;
INV     gate4544  (.A(WX3589), .Z(WX2707) ) ;
INV     gate4545  (.A(WX3590), .Z(WX2711) ) ;
INV     gate4546  (.A(WX3590), .Z(WX2715) ) ;
OR2     gate4547  (.A(WX2706), .B(WX2705), .Z(WX2708) ) ;
INV     gate4548  (.A(WX2708), .Z(WX2717) ) ;
INV     gate4549  (.A(WX2717), .Z(WX2718) ) ;
INV     gate4550  (.A(WX3589), .Z(WX2721) ) ;
INV     gate4551  (.A(WX3590), .Z(WX2725) ) ;
INV     gate4552  (.A(WX3590), .Z(WX2729) ) ;
OR2     gate4553  (.A(WX2720), .B(WX2719), .Z(WX2722) ) ;
INV     gate4554  (.A(WX2722), .Z(WX2731) ) ;
INV     gate4555  (.A(WX2731), .Z(WX2732) ) ;
INV     gate4556  (.A(WX3589), .Z(WX2735) ) ;
INV     gate4557  (.A(WX3590), .Z(WX2739) ) ;
INV     gate4558  (.A(WX3590), .Z(WX2743) ) ;
OR2     gate4559  (.A(WX2734), .B(WX2733), .Z(WX2736) ) ;
INV     gate4560  (.A(WX2736), .Z(WX2745) ) ;
INV     gate4561  (.A(WX2745), .Z(WX2746) ) ;
INV     gate4562  (.A(WX3589), .Z(WX2749) ) ;
INV     gate4563  (.A(WX3590), .Z(WX2753) ) ;
INV     gate4564  (.A(WX3590), .Z(WX2757) ) ;
OR2     gate4565  (.A(WX2748), .B(WX2747), .Z(WX2750) ) ;
INV     gate4566  (.A(WX2750), .Z(WX2759) ) ;
INV     gate4567  (.A(WX2759), .Z(WX2760) ) ;
INV     gate4568  (.A(WX3589), .Z(WX2763) ) ;
INV     gate4569  (.A(WX3590), .Z(WX2767) ) ;
INV     gate4570  (.A(WX3590), .Z(WX2771) ) ;
OR2     gate4571  (.A(WX2762), .B(WX2761), .Z(WX2764) ) ;
INV     gate4572  (.A(WX2764), .Z(WX2773) ) ;
INV     gate4573  (.A(WX2773), .Z(WX2774) ) ;
INV     gate4574  (.A(WX3589), .Z(WX2777) ) ;
INV     gate4575  (.A(WX3590), .Z(WX2781) ) ;
INV     gate4576  (.A(WX3590), .Z(WX2785) ) ;
OR2     gate4577  (.A(WX2776), .B(WX2775), .Z(WX2778) ) ;
INV     gate4578  (.A(WX2778), .Z(WX2787) ) ;
INV     gate4579  (.A(WX2787), .Z(WX2788) ) ;
INV     gate4580  (.A(WX3589), .Z(WX2791) ) ;
INV     gate4581  (.A(WX3590), .Z(WX2795) ) ;
INV     gate4582  (.A(WX3590), .Z(WX2799) ) ;
OR2     gate4583  (.A(WX2790), .B(WX2789), .Z(WX2792) ) ;
INV     gate4584  (.A(WX2792), .Z(WX2801) ) ;
INV     gate4585  (.A(WX2801), .Z(WX2802) ) ;
INV     gate4586  (.A(WX3589), .Z(WX2805) ) ;
INV     gate4587  (.A(WX3590), .Z(WX2809) ) ;
INV     gate4588  (.A(WX3590), .Z(WX2813) ) ;
OR2     gate4589  (.A(WX2804), .B(WX2803), .Z(WX2806) ) ;
INV     gate4590  (.A(WX2806), .Z(WX2815) ) ;
INV     gate4591  (.A(WX2815), .Z(WX2816) ) ;
INV     gate4592  (.A(WX3589), .Z(WX2819) ) ;
INV     gate4593  (.A(WX3590), .Z(WX2823) ) ;
INV     gate4594  (.A(WX3590), .Z(WX2827) ) ;
OR2     gate4595  (.A(WX2818), .B(WX2817), .Z(WX2820) ) ;
INV     gate4596  (.A(WX2820), .Z(WX2829) ) ;
INV     gate4597  (.A(WX2829), .Z(WX2830) ) ;
INV     gate4598  (.A(WX3589), .Z(WX2833) ) ;
INV     gate4599  (.A(WX3590), .Z(WX2837) ) ;
INV     gate4600  (.A(WX3590), .Z(WX2841) ) ;
OR2     gate4601  (.A(WX2832), .B(WX2831), .Z(WX2834) ) ;
INV     gate4602  (.A(WX2834), .Z(WX2843) ) ;
INV     gate4603  (.A(WX2843), .Z(WX2844) ) ;
INV     gate4604  (.A(WX3589), .Z(WX2847) ) ;
INV     gate4605  (.A(WX3590), .Z(WX2851) ) ;
INV     gate4606  (.A(WX3590), .Z(WX2855) ) ;
OR2     gate4607  (.A(WX2846), .B(WX2845), .Z(WX2848) ) ;
INV     gate4608  (.A(WX2848), .Z(WX2857) ) ;
INV     gate4609  (.A(WX2857), .Z(WX2858) ) ;
INV     gate4610  (.A(WX3589), .Z(WX2861) ) ;
INV     gate4611  (.A(WX3590), .Z(WX2865) ) ;
INV     gate4612  (.A(WX3590), .Z(WX2869) ) ;
OR2     gate4613  (.A(WX2860), .B(WX2859), .Z(WX2862) ) ;
INV     gate4614  (.A(WX2862), .Z(WX2871) ) ;
INV     gate4615  (.A(WX2871), .Z(WX2872) ) ;
INV     gate4616  (.A(WX3589), .Z(WX2875) ) ;
INV     gate4617  (.A(WX3590), .Z(WX2879) ) ;
INV     gate4618  (.A(WX3590), .Z(WX2883) ) ;
OR2     gate4619  (.A(WX2874), .B(WX2873), .Z(WX2876) ) ;
INV     gate4620  (.A(WX2876), .Z(WX2885) ) ;
INV     gate4621  (.A(WX2885), .Z(WX2886) ) ;
INV     gate4622  (.A(WX3589), .Z(WX2889) ) ;
INV     gate4623  (.A(WX3590), .Z(WX2893) ) ;
INV     gate4624  (.A(WX3590), .Z(WX2897) ) ;
OR2     gate4625  (.A(WX2888), .B(WX2887), .Z(WX2890) ) ;
INV     gate4626  (.A(WX2890), .Z(WX2899) ) ;
INV     gate4627  (.A(WX2899), .Z(WX2900) ) ;
INV     gate4628  (.A(WX3589), .Z(WX2903) ) ;
INV     gate4629  (.A(WX3590), .Z(WX2907) ) ;
INV     gate4630  (.A(WX3590), .Z(WX2911) ) ;
OR2     gate4631  (.A(WX2902), .B(WX2901), .Z(WX2904) ) ;
INV     gate4632  (.A(WX2904), .Z(WX2913) ) ;
INV     gate4633  (.A(WX2913), .Z(WX2914) ) ;
INV     gate4634  (.A(WX3589), .Z(WX2917) ) ;
INV     gate4635  (.A(WX3590), .Z(WX2921) ) ;
INV     gate4636  (.A(WX3590), .Z(WX2925) ) ;
OR2     gate4637  (.A(WX2916), .B(WX2915), .Z(WX2918) ) ;
INV     gate4638  (.A(WX2918), .Z(WX2927) ) ;
INV     gate4639  (.A(WX2927), .Z(WX2928) ) ;
INV     gate4640  (.A(WX3589), .Z(WX2931) ) ;
INV     gate4641  (.A(WX3590), .Z(WX2935) ) ;
INV     gate4642  (.A(WX3590), .Z(WX2939) ) ;
OR2     gate4643  (.A(WX2930), .B(WX2929), .Z(WX2932) ) ;
INV     gate4644  (.A(WX2932), .Z(WX2941) ) ;
INV     gate4645  (.A(WX2941), .Z(WX2942) ) ;
INV     gate4646  (.A(WX3589), .Z(WX2945) ) ;
INV     gate4647  (.A(WX3590), .Z(WX2949) ) ;
INV     gate4648  (.A(WX3590), .Z(WX2953) ) ;
OR2     gate4649  (.A(WX2944), .B(WX2943), .Z(WX2946) ) ;
INV     gate4650  (.A(WX2946), .Z(WX2955) ) ;
INV     gate4651  (.A(WX2955), .Z(WX2956) ) ;
INV     gate4652  (.A(WX3589), .Z(WX2959) ) ;
INV     gate4653  (.A(WX3590), .Z(WX2963) ) ;
INV     gate4654  (.A(WX3590), .Z(WX2967) ) ;
OR2     gate4655  (.A(WX2958), .B(WX2957), .Z(WX2960) ) ;
INV     gate4656  (.A(WX2960), .Z(WX2969) ) ;
INV     gate4657  (.A(WX2969), .Z(WX2970) ) ;
INV     gate4658  (.A(WX3589), .Z(WX2973) ) ;
INV     gate4659  (.A(WX3590), .Z(WX2977) ) ;
INV     gate4660  (.A(WX3590), .Z(WX2981) ) ;
OR2     gate4661  (.A(WX2972), .B(WX2971), .Z(WX2974) ) ;
INV     gate4662  (.A(WX2974), .Z(WX2983) ) ;
INV     gate4663  (.A(WX2983), .Z(WX2984) ) ;
INV     gate4664  (.A(WX3589), .Z(WX2987) ) ;
INV     gate4665  (.A(WX3590), .Z(WX2991) ) ;
INV     gate4666  (.A(WX3590), .Z(WX2995) ) ;
OR2     gate4667  (.A(WX2986), .B(WX2985), .Z(WX2988) ) ;
INV     gate4668  (.A(WX2988), .Z(WX2997) ) ;
INV     gate4669  (.A(WX2997), .Z(WX2998) ) ;
INV     gate4670  (.A(WX3589), .Z(WX3001) ) ;
INV     gate4671  (.A(WX3590), .Z(WX3005) ) ;
INV     gate4672  (.A(WX3590), .Z(WX3009) ) ;
OR2     gate4673  (.A(WX3000), .B(WX2999), .Z(WX3002) ) ;
INV     gate4674  (.A(WX3002), .Z(WX3011) ) ;
INV     gate4675  (.A(WX3011), .Z(WX3012) ) ;
INV     gate4676  (.A(WX3589), .Z(WX3015) ) ;
INV     gate4677  (.A(WX3590), .Z(WX3019) ) ;
INV     gate4678  (.A(WX3590), .Z(WX3023) ) ;
OR2     gate4679  (.A(WX3014), .B(WX3013), .Z(WX3016) ) ;
INV     gate4680  (.A(WX3016), .Z(WX3025) ) ;
INV     gate4681  (.A(WX3025), .Z(WX3026) ) ;
INV     gate4682  (.A(WX3589), .Z(WX3029) ) ;
INV     gate4683  (.A(WX3590), .Z(WX3033) ) ;
INV     gate4684  (.A(WX3590), .Z(WX3037) ) ;
OR2     gate4685  (.A(WX3028), .B(WX3027), .Z(WX3030) ) ;
INV     gate4686  (.A(WX3030), .Z(WX3039) ) ;
INV     gate4687  (.A(WX3039), .Z(WX3040) ) ;
INV     gate4688  (.A(WX3589), .Z(WX3043) ) ;
INV     gate4689  (.A(WX3590), .Z(WX3047) ) ;
INV     gate4690  (.A(WX3590), .Z(WX3051) ) ;
OR2     gate4691  (.A(WX3042), .B(WX3041), .Z(WX3044) ) ;
INV     gate4692  (.A(WX3044), .Z(WX3053) ) ;
INV     gate4693  (.A(WX3053), .Z(WX3054) ) ;
INV     gate4694  (.A(WX3589), .Z(WX3057) ) ;
INV     gate4695  (.A(WX3590), .Z(WX3061) ) ;
INV     gate4696  (.A(WX3590), .Z(WX3065) ) ;
OR2     gate4697  (.A(WX3056), .B(WX3055), .Z(WX3058) ) ;
INV     gate4698  (.A(WX3058), .Z(WX3067) ) ;
INV     gate4699  (.A(WX3067), .Z(WX3068) ) ;
INV     gate4700  (.A(WX3071), .Z(WX3069) ) ;
INV     gate4701  (.A(WX3550), .Z(WX3551) ) ;
INV     gate4702  (.A(WX3551), .Z(WX3134) ) ;
INV     gate4703  (.A(WX3552), .Z(WX3553) ) ;
INV     gate4704  (.A(WX3553), .Z(WX3135) ) ;
INV     gate4705  (.A(WX3554), .Z(WX3555) ) ;
INV     gate4706  (.A(WX3555), .Z(WX3136) ) ;
INV     gate4707  (.A(WX3556), .Z(WX3557) ) ;
INV     gate4708  (.A(WX3557), .Z(WX3137) ) ;
INV     gate4709  (.A(WX3558), .Z(WX3559) ) ;
INV     gate4710  (.A(WX3559), .Z(WX3138) ) ;
INV     gate4711  (.A(WX3560), .Z(WX3561) ) ;
INV     gate4712  (.A(WX3561), .Z(WX3139) ) ;
INV     gate4713  (.A(WX3562), .Z(WX3563) ) ;
INV     gate4714  (.A(WX3563), .Z(WX3140) ) ;
INV     gate4715  (.A(WX3564), .Z(WX3565) ) ;
INV     gate4716  (.A(WX3565), .Z(WX3141) ) ;
INV     gate4717  (.A(WX3566), .Z(WX3567) ) ;
INV     gate4718  (.A(WX3567), .Z(WX3142) ) ;
INV     gate4719  (.A(WX3568), .Z(WX3569) ) ;
INV     gate4720  (.A(WX3569), .Z(WX3143) ) ;
INV     gate4721  (.A(WX3570), .Z(WX3571) ) ;
INV     gate4722  (.A(WX3571), .Z(WX3144) ) ;
INV     gate4723  (.A(WX3572), .Z(WX3573) ) ;
INV     gate4724  (.A(WX3573), .Z(WX3145) ) ;
INV     gate4725  (.A(WX3574), .Z(WX3575) ) ;
INV     gate4726  (.A(WX3575), .Z(WX3146) ) ;
INV     gate4727  (.A(WX3576), .Z(WX3577) ) ;
INV     gate4728  (.A(WX3577), .Z(WX3147) ) ;
INV     gate4729  (.A(WX3578), .Z(WX3579) ) ;
INV     gate4730  (.A(WX3579), .Z(WX3148) ) ;
INV     gate4731  (.A(WX3580), .Z(WX3581) ) ;
INV     gate4732  (.A(WX3581), .Z(WX3149) ) ;
INV     gate4733  (.A(WX3518), .Z(WX3519) ) ;
INV     gate4734  (.A(WX3519), .Z(WX3150) ) ;
INV     gate4735  (.A(WX3520), .Z(WX3521) ) ;
INV     gate4736  (.A(WX3521), .Z(WX3151) ) ;
INV     gate4737  (.A(WX3522), .Z(WX3523) ) ;
INV     gate4738  (.A(WX3523), .Z(WX3152) ) ;
INV     gate4739  (.A(WX3524), .Z(WX3525) ) ;
INV     gate4740  (.A(WX3525), .Z(WX3153) ) ;
INV     gate4741  (.A(WX3526), .Z(WX3527) ) ;
INV     gate4742  (.A(WX3527), .Z(WX3154) ) ;
INV     gate4743  (.A(WX3528), .Z(WX3529) ) ;
INV     gate4744  (.A(WX3529), .Z(WX3155) ) ;
INV     gate4745  (.A(WX3530), .Z(WX3531) ) ;
INV     gate4746  (.A(WX3531), .Z(WX3156) ) ;
INV     gate4747  (.A(WX3532), .Z(WX3533) ) ;
INV     gate4748  (.A(WX3533), .Z(WX3157) ) ;
INV     gate4749  (.A(WX3534), .Z(WX3535) ) ;
INV     gate4750  (.A(WX3535), .Z(WX3158) ) ;
INV     gate4751  (.A(WX3536), .Z(WX3537) ) ;
INV     gate4752  (.A(WX3537), .Z(WX3159) ) ;
INV     gate4753  (.A(WX3538), .Z(WX3539) ) ;
INV     gate4754  (.A(WX3539), .Z(WX3160) ) ;
INV     gate4755  (.A(WX3540), .Z(WX3541) ) ;
INV     gate4756  (.A(WX3541), .Z(WX3161) ) ;
INV     gate4757  (.A(WX3542), .Z(WX3543) ) ;
INV     gate4758  (.A(WX3543), .Z(WX3162) ) ;
INV     gate4759  (.A(WX3544), .Z(WX3545) ) ;
INV     gate4760  (.A(WX3545), .Z(WX3163) ) ;
INV     gate4761  (.A(WX3546), .Z(WX3547) ) ;
INV     gate4762  (.A(WX3547), .Z(WX3164) ) ;
INV     gate4763  (.A(WX3548), .Z(WX3549) ) ;
INV     gate4764  (.A(WX3549), .Z(WX3165) ) ;
INV     gate4765  (.A(WX3134), .Z(WX3166) ) ;
INV     gate4766  (.A(WX3135), .Z(WX3167) ) ;
INV     gate4767  (.A(WX3136), .Z(WX3168) ) ;
INV     gate4768  (.A(WX3137), .Z(WX3169) ) ;
INV     gate4769  (.A(WX3138), .Z(WX3170) ) ;
INV     gate4770  (.A(WX3139), .Z(WX3171) ) ;
INV     gate4771  (.A(WX3140), .Z(WX3172) ) ;
INV     gate4772  (.A(WX3141), .Z(WX3173) ) ;
INV     gate4773  (.A(WX3142), .Z(WX3174) ) ;
INV     gate4774  (.A(WX3143), .Z(WX3175) ) ;
INV     gate4775  (.A(WX3144), .Z(WX3176) ) ;
INV     gate4776  (.A(WX3145), .Z(WX3177) ) ;
INV     gate4777  (.A(WX3146), .Z(WX3178) ) ;
INV     gate4778  (.A(WX3147), .Z(WX3179) ) ;
INV     gate4779  (.A(WX3148), .Z(WX3180) ) ;
INV     gate4780  (.A(WX3149), .Z(WX3181) ) ;
INV     gate4781  (.A(WX3150), .Z(WX3182) ) ;
INV     gate4782  (.A(WX3151), .Z(WX3183) ) ;
INV     gate4783  (.A(WX3152), .Z(WX3184) ) ;
INV     gate4784  (.A(WX3153), .Z(WX3185) ) ;
INV     gate4785  (.A(WX3154), .Z(WX3186) ) ;
INV     gate4786  (.A(WX3155), .Z(WX3187) ) ;
INV     gate4787  (.A(WX3156), .Z(WX3188) ) ;
INV     gate4788  (.A(WX3157), .Z(WX3189) ) ;
INV     gate4789  (.A(WX3158), .Z(WX3190) ) ;
INV     gate4790  (.A(WX3159), .Z(WX3191) ) ;
INV     gate4791  (.A(WX3160), .Z(WX3192) ) ;
INV     gate4792  (.A(WX3161), .Z(WX3193) ) ;
INV     gate4793  (.A(WX3162), .Z(WX3194) ) ;
INV     gate4794  (.A(WX3163), .Z(WX3195) ) ;
INV     gate4795  (.A(WX3164), .Z(WX3196) ) ;
INV     gate4796  (.A(WX3165), .Z(WX3197) ) ;
INV     gate4797  (.A(WX3423), .Z(WX3198) ) ;
INV     gate4798  (.A(WX3425), .Z(WX3199) ) ;
INV     gate4799  (.A(WX3427), .Z(WX3200) ) ;
INV     gate4800  (.A(WX3429), .Z(WX3201) ) ;
INV     gate4801  (.A(WX3431), .Z(WX3202) ) ;
INV     gate4802  (.A(WX3433), .Z(WX3203) ) ;
INV     gate4803  (.A(WX3435), .Z(WX3204) ) ;
INV     gate4804  (.A(WX3437), .Z(WX3205) ) ;
INV     gate4805  (.A(WX3439), .Z(WX3206) ) ;
INV     gate4806  (.A(WX3441), .Z(WX3207) ) ;
INV     gate4807  (.A(WX3443), .Z(WX3208) ) ;
INV     gate4808  (.A(WX3445), .Z(WX3209) ) ;
INV     gate4809  (.A(WX3447), .Z(WX3210) ) ;
INV     gate4810  (.A(WX3449), .Z(WX3211) ) ;
INV     gate4811  (.A(WX3451), .Z(WX3212) ) ;
INV     gate4812  (.A(WX3453), .Z(WX3213) ) ;
INV     gate4813  (.A(WX3455), .Z(WX3214) ) ;
INV     gate4814  (.A(WX3457), .Z(WX3215) ) ;
INV     gate4815  (.A(WX3459), .Z(WX3216) ) ;
INV     gate4816  (.A(WX3461), .Z(WX3217) ) ;
INV     gate4817  (.A(WX3463), .Z(WX3218) ) ;
INV     gate4818  (.A(WX3465), .Z(WX3219) ) ;
INV     gate4819  (.A(WX3467), .Z(WX3220) ) ;
INV     gate4820  (.A(WX3469), .Z(WX3221) ) ;
INV     gate4821  (.A(WX3471), .Z(WX3222) ) ;
INV     gate4822  (.A(WX3473), .Z(WX3223) ) ;
INV     gate4823  (.A(WX3475), .Z(WX3224) ) ;
INV     gate4824  (.A(WX3477), .Z(WX3225) ) ;
INV     gate4825  (.A(WX3479), .Z(WX3226) ) ;
INV     gate4826  (.A(WX3481), .Z(WX3227) ) ;
INV     gate4827  (.A(WX3483), .Z(WX3228) ) ;
INV     gate4828  (.A(WX3485), .Z(WX3229) ) ;
NAND2   gate4829  (.A(II10517), .B(II10518), .Z(WX3502) ) ;
INV     gate4830  (.A(WX3502), .Z(WX3518) ) ;
NAND2   gate4831  (.A(II10548), .B(II10549), .Z(WX3503) ) ;
INV     gate4832  (.A(WX3503), .Z(WX3520) ) ;
NAND2   gate4833  (.A(II10579), .B(II10580), .Z(WX3504) ) ;
INV     gate4834  (.A(WX3504), .Z(WX3522) ) ;
NAND2   gate4835  (.A(II10610), .B(II10611), .Z(WX3505) ) ;
INV     gate4836  (.A(WX3505), .Z(WX3524) ) ;
NAND2   gate4837  (.A(II10641), .B(II10642), .Z(WX3506) ) ;
INV     gate4838  (.A(WX3506), .Z(WX3526) ) ;
NAND2   gate4839  (.A(II10672), .B(II10673), .Z(WX3507) ) ;
INV     gate4840  (.A(WX3507), .Z(WX3528) ) ;
NAND2   gate4841  (.A(II10703), .B(II10704), .Z(WX3508) ) ;
INV     gate4842  (.A(WX3508), .Z(WX3530) ) ;
NAND2   gate4843  (.A(II10734), .B(II10735), .Z(WX3509) ) ;
INV     gate4844  (.A(WX3509), .Z(WX3532) ) ;
NAND2   gate4845  (.A(II10765), .B(II10766), .Z(WX3510) ) ;
INV     gate4846  (.A(WX3510), .Z(WX3534) ) ;
NAND2   gate4847  (.A(II10796), .B(II10797), .Z(WX3511) ) ;
INV     gate4848  (.A(WX3511), .Z(WX3536) ) ;
NAND2   gate4849  (.A(II10827), .B(II10828), .Z(WX3512) ) ;
INV     gate4850  (.A(WX3512), .Z(WX3538) ) ;
NAND2   gate4851  (.A(II10858), .B(II10859), .Z(WX3513) ) ;
INV     gate4852  (.A(WX3513), .Z(WX3540) ) ;
NAND2   gate4853  (.A(II10889), .B(II10890), .Z(WX3514) ) ;
INV     gate4854  (.A(WX3514), .Z(WX3542) ) ;
NAND2   gate4855  (.A(II10920), .B(II10921), .Z(WX3515) ) ;
INV     gate4856  (.A(WX3515), .Z(WX3544) ) ;
NAND2   gate4857  (.A(II10951), .B(II10952), .Z(WX3516) ) ;
INV     gate4858  (.A(WX3516), .Z(WX3546) ) ;
NAND2   gate4859  (.A(II10982), .B(II10983), .Z(WX3517) ) ;
INV     gate4860  (.A(WX3517), .Z(WX3548) ) ;
NAND2   gate4861  (.A(II10021), .B(II10022), .Z(WX3486) ) ;
INV     gate4862  (.A(WX3486), .Z(WX3550) ) ;
NAND2   gate4863  (.A(II10052), .B(II10053), .Z(WX3487) ) ;
INV     gate4864  (.A(WX3487), .Z(WX3552) ) ;
NAND2   gate4865  (.A(II10083), .B(II10084), .Z(WX3488) ) ;
INV     gate4866  (.A(WX3488), .Z(WX3554) ) ;
NAND2   gate4867  (.A(II10114), .B(II10115), .Z(WX3489) ) ;
INV     gate4868  (.A(WX3489), .Z(WX3556) ) ;
NAND2   gate4869  (.A(II10145), .B(II10146), .Z(WX3490) ) ;
INV     gate4870  (.A(WX3490), .Z(WX3558) ) ;
NAND2   gate4871  (.A(II10176), .B(II10177), .Z(WX3491) ) ;
INV     gate4872  (.A(WX3491), .Z(WX3560) ) ;
NAND2   gate4873  (.A(II10207), .B(II10208), .Z(WX3492) ) ;
INV     gate4874  (.A(WX3492), .Z(WX3562) ) ;
NAND2   gate4875  (.A(II10238), .B(II10239), .Z(WX3493) ) ;
INV     gate4876  (.A(WX3493), .Z(WX3564) ) ;
NAND2   gate4877  (.A(II10269), .B(II10270), .Z(WX3494) ) ;
INV     gate4878  (.A(WX3494), .Z(WX3566) ) ;
NAND2   gate4879  (.A(II10300), .B(II10301), .Z(WX3495) ) ;
INV     gate4880  (.A(WX3495), .Z(WX3568) ) ;
NAND2   gate4881  (.A(II10331), .B(II10332), .Z(WX3496) ) ;
INV     gate4882  (.A(WX3496), .Z(WX3570) ) ;
NAND2   gate4883  (.A(II10362), .B(II10363), .Z(WX3497) ) ;
INV     gate4884  (.A(WX3497), .Z(WX3572) ) ;
NAND2   gate4885  (.A(II10393), .B(II10394), .Z(WX3498) ) ;
INV     gate4886  (.A(WX3498), .Z(WX3574) ) ;
NAND2   gate4887  (.A(II10424), .B(II10425), .Z(WX3499) ) ;
INV     gate4888  (.A(WX3499), .Z(WX3576) ) ;
NAND2   gate4889  (.A(II10455), .B(II10456), .Z(WX3500) ) ;
INV     gate4890  (.A(WX3500), .Z(WX3578) ) ;
NAND2   gate4891  (.A(II10486), .B(II10487), .Z(WX3501) ) ;
INV     gate4892  (.A(WX3501), .Z(WX3580) ) ;
INV     gate4893  (.A(TM0), .Z(WX3582) ) ;
INV     gate4894  (.A(TM0), .Z(WX3583) ) ;
INV     gate4895  (.A(TM0), .Z(WX3584) ) ;
INV     gate4896  (.A(TM1), .Z(WX3585) ) ;
INV     gate4897  (.A(TM1), .Z(WX3586) ) ;
INV     gate4898  (.A(WX3586), .Z(WX3587) ) ;
INV     gate4899  (.A(WX3584), .Z(WX3588) ) ;
INV     gate4900  (.A(WX3582), .Z(WX3591) ) ;
INV     gate4901  (.A(WX3591), .Z(WX3595) ) ;
OR2     gate4902  (.A(WX3594), .B(WX3593), .Z(WX3596) ) ;
INV     gate4903  (.A(WX3596), .Z(WX3597) ) ;
INV     gate4904  (.A(WX3597), .Z(WX3598) ) ;
INV     gate4905  (.A(WX3591), .Z(WX3602) ) ;
OR2     gate4906  (.A(WX3601), .B(WX3600), .Z(WX3603) ) ;
INV     gate4907  (.A(WX3603), .Z(WX3604) ) ;
INV     gate4908  (.A(WX3604), .Z(WX3605) ) ;
INV     gate4909  (.A(WX3591), .Z(WX3609) ) ;
OR2     gate4910  (.A(WX3608), .B(WX3607), .Z(WX3610) ) ;
INV     gate4911  (.A(WX3610), .Z(WX3611) ) ;
INV     gate4912  (.A(WX3611), .Z(WX3612) ) ;
INV     gate4913  (.A(WX3591), .Z(WX3616) ) ;
OR2     gate4914  (.A(WX3615), .B(WX3614), .Z(WX3617) ) ;
INV     gate4915  (.A(WX3617), .Z(WX3618) ) ;
INV     gate4916  (.A(WX3618), .Z(WX3619) ) ;
INV     gate4917  (.A(WX3591), .Z(WX3623) ) ;
OR2     gate4918  (.A(WX3622), .B(WX3621), .Z(WX3624) ) ;
INV     gate4919  (.A(WX3624), .Z(WX3625) ) ;
INV     gate4920  (.A(WX3625), .Z(WX3626) ) ;
INV     gate4921  (.A(WX3591), .Z(WX3630) ) ;
OR2     gate4922  (.A(WX3629), .B(WX3628), .Z(WX3631) ) ;
INV     gate4923  (.A(WX3631), .Z(WX3632) ) ;
INV     gate4924  (.A(WX3632), .Z(WX3633) ) ;
INV     gate4925  (.A(WX3591), .Z(WX3637) ) ;
OR2     gate4926  (.A(WX3636), .B(WX3635), .Z(WX3638) ) ;
INV     gate4927  (.A(WX3638), .Z(WX3639) ) ;
INV     gate4928  (.A(WX3639), .Z(WX3640) ) ;
INV     gate4929  (.A(WX3591), .Z(WX3644) ) ;
OR2     gate4930  (.A(WX3643), .B(WX3642), .Z(WX3645) ) ;
INV     gate4931  (.A(WX3645), .Z(WX3646) ) ;
INV     gate4932  (.A(WX3646), .Z(WX3647) ) ;
INV     gate4933  (.A(WX3591), .Z(WX3651) ) ;
OR2     gate4934  (.A(WX3650), .B(WX3649), .Z(WX3652) ) ;
INV     gate4935  (.A(WX3652), .Z(WX3653) ) ;
INV     gate4936  (.A(WX3653), .Z(WX3654) ) ;
INV     gate4937  (.A(WX3591), .Z(WX3658) ) ;
OR2     gate4938  (.A(WX3657), .B(WX3656), .Z(WX3659) ) ;
INV     gate4939  (.A(WX3659), .Z(WX3660) ) ;
INV     gate4940  (.A(WX3660), .Z(WX3661) ) ;
INV     gate4941  (.A(WX3591), .Z(WX3665) ) ;
OR2     gate4942  (.A(WX3664), .B(WX3663), .Z(WX3666) ) ;
INV     gate4943  (.A(WX3666), .Z(WX3667) ) ;
INV     gate4944  (.A(WX3667), .Z(WX3668) ) ;
INV     gate4945  (.A(WX3591), .Z(WX3672) ) ;
OR2     gate4946  (.A(WX3671), .B(WX3670), .Z(WX3673) ) ;
INV     gate4947  (.A(WX3673), .Z(WX3674) ) ;
INV     gate4948  (.A(WX3674), .Z(WX3675) ) ;
INV     gate4949  (.A(WX3591), .Z(WX3679) ) ;
OR2     gate4950  (.A(WX3678), .B(WX3677), .Z(WX3680) ) ;
INV     gate4951  (.A(WX3680), .Z(WX3681) ) ;
INV     gate4952  (.A(WX3681), .Z(WX3682) ) ;
INV     gate4953  (.A(WX3591), .Z(WX3686) ) ;
OR2     gate4954  (.A(WX3685), .B(WX3684), .Z(WX3687) ) ;
INV     gate4955  (.A(WX3687), .Z(WX3688) ) ;
INV     gate4956  (.A(WX3688), .Z(WX3689) ) ;
INV     gate4957  (.A(WX3591), .Z(WX3693) ) ;
OR2     gate4958  (.A(WX3692), .B(WX3691), .Z(WX3694) ) ;
INV     gate4959  (.A(WX3694), .Z(WX3695) ) ;
INV     gate4960  (.A(WX3695), .Z(WX3696) ) ;
INV     gate4961  (.A(WX3591), .Z(WX3700) ) ;
OR2     gate4962  (.A(WX3699), .B(WX3698), .Z(WX3701) ) ;
INV     gate4963  (.A(WX3701), .Z(WX3702) ) ;
INV     gate4964  (.A(WX3702), .Z(WX3703) ) ;
INV     gate4965  (.A(WX3591), .Z(WX3707) ) ;
OR2     gate4966  (.A(WX3706), .B(WX3705), .Z(WX3708) ) ;
INV     gate4967  (.A(WX3708), .Z(WX3709) ) ;
INV     gate4968  (.A(WX3709), .Z(WX3710) ) ;
INV     gate4969  (.A(WX3591), .Z(WX3714) ) ;
OR2     gate4970  (.A(WX3713), .B(WX3712), .Z(WX3715) ) ;
INV     gate4971  (.A(WX3715), .Z(WX3716) ) ;
INV     gate4972  (.A(WX3716), .Z(WX3717) ) ;
INV     gate4973  (.A(WX3591), .Z(WX3721) ) ;
OR2     gate4974  (.A(WX3720), .B(WX3719), .Z(WX3722) ) ;
INV     gate4975  (.A(WX3722), .Z(WX3723) ) ;
INV     gate4976  (.A(WX3723), .Z(WX3724) ) ;
INV     gate4977  (.A(WX3591), .Z(WX3728) ) ;
OR2     gate4978  (.A(WX3727), .B(WX3726), .Z(WX3729) ) ;
INV     gate4979  (.A(WX3729), .Z(WX3730) ) ;
INV     gate4980  (.A(WX3730), .Z(WX3731) ) ;
INV     gate4981  (.A(WX3591), .Z(WX3735) ) ;
OR2     gate4982  (.A(WX3734), .B(WX3733), .Z(WX3736) ) ;
INV     gate4983  (.A(WX3736), .Z(WX3737) ) ;
INV     gate4984  (.A(WX3737), .Z(WX3738) ) ;
INV     gate4985  (.A(WX3591), .Z(WX3742) ) ;
OR2     gate4986  (.A(WX3741), .B(WX3740), .Z(WX3743) ) ;
INV     gate4987  (.A(WX3743), .Z(WX3744) ) ;
INV     gate4988  (.A(WX3744), .Z(WX3745) ) ;
INV     gate4989  (.A(WX3591), .Z(WX3749) ) ;
OR2     gate4990  (.A(WX3748), .B(WX3747), .Z(WX3750) ) ;
INV     gate4991  (.A(WX3750), .Z(WX3751) ) ;
INV     gate4992  (.A(WX3751), .Z(WX3752) ) ;
INV     gate4993  (.A(WX3591), .Z(WX3756) ) ;
OR2     gate4994  (.A(WX3755), .B(WX3754), .Z(WX3757) ) ;
INV     gate4995  (.A(WX3757), .Z(WX3758) ) ;
INV     gate4996  (.A(WX3758), .Z(WX3759) ) ;
INV     gate4997  (.A(WX3591), .Z(WX3763) ) ;
OR2     gate4998  (.A(WX3762), .B(WX3761), .Z(WX3764) ) ;
INV     gate4999  (.A(WX3764), .Z(WX3765) ) ;
INV     gate5000  (.A(WX3765), .Z(WX3766) ) ;
INV     gate5001  (.A(WX3591), .Z(WX3770) ) ;
OR2     gate5002  (.A(WX3769), .B(WX3768), .Z(WX3771) ) ;
INV     gate5003  (.A(WX3771), .Z(WX3772) ) ;
INV     gate5004  (.A(WX3772), .Z(WX3773) ) ;
INV     gate5005  (.A(WX3591), .Z(WX3777) ) ;
OR2     gate5006  (.A(WX3776), .B(WX3775), .Z(WX3778) ) ;
INV     gate5007  (.A(WX3778), .Z(WX3779) ) ;
INV     gate5008  (.A(WX3779), .Z(WX3780) ) ;
INV     gate5009  (.A(WX3591), .Z(WX3784) ) ;
OR2     gate5010  (.A(WX3783), .B(WX3782), .Z(WX3785) ) ;
INV     gate5011  (.A(WX3785), .Z(WX3786) ) ;
INV     gate5012  (.A(WX3786), .Z(WX3787) ) ;
INV     gate5013  (.A(WX3591), .Z(WX3791) ) ;
OR2     gate5014  (.A(WX3790), .B(WX3789), .Z(WX3792) ) ;
INV     gate5015  (.A(WX3792), .Z(WX3793) ) ;
INV     gate5016  (.A(WX3793), .Z(WX3794) ) ;
INV     gate5017  (.A(WX3591), .Z(WX3798) ) ;
OR2     gate5018  (.A(WX3797), .B(WX3796), .Z(WX3799) ) ;
INV     gate5019  (.A(WX3799), .Z(WX3800) ) ;
INV     gate5020  (.A(WX3800), .Z(WX3801) ) ;
INV     gate5021  (.A(WX3591), .Z(WX3805) ) ;
OR2     gate5022  (.A(WX3804), .B(WX3803), .Z(WX3806) ) ;
INV     gate5023  (.A(WX3806), .Z(WX3807) ) ;
INV     gate5024  (.A(WX3807), .Z(WX3808) ) ;
INV     gate5025  (.A(WX3591), .Z(WX3812) ) ;
OR2     gate5026  (.A(WX3811), .B(WX3810), .Z(WX3813) ) ;
INV     gate5027  (.A(WX3813), .Z(WX3814) ) ;
INV     gate5028  (.A(WX3814), .Z(WX3815) ) ;
INV     gate5029  (.A(RESET), .Z(WX3816) ) ;
INV     gate5030  (.A(WX3816), .Z(WX3849) ) ;
INV     gate5031  (.A(WX4878), .Z(WX4882) ) ;
INV     gate5032  (.A(WX4882), .Z(WX3916) ) ;
INV     gate5033  (.A(WX4876), .Z(WX4883) ) ;
INV     gate5034  (.A(WX4883), .Z(WX3920) ) ;
INV     gate5035  (.A(WX4883), .Z(WX3924) ) ;
OR2     gate5036  (.A(WX3915), .B(WX3914), .Z(WX3917) ) ;
INV     gate5037  (.A(WX3917), .Z(WX3926) ) ;
INV     gate5038  (.A(WX3926), .Z(WX3927) ) ;
INV     gate5039  (.A(WX4882), .Z(WX3930) ) ;
INV     gate5040  (.A(WX4883), .Z(WX3934) ) ;
INV     gate5041  (.A(WX4883), .Z(WX3938) ) ;
OR2     gate5042  (.A(WX3929), .B(WX3928), .Z(WX3931) ) ;
INV     gate5043  (.A(WX3931), .Z(WX3940) ) ;
INV     gate5044  (.A(WX3940), .Z(WX3941) ) ;
INV     gate5045  (.A(WX4882), .Z(WX3944) ) ;
INV     gate5046  (.A(WX4883), .Z(WX3948) ) ;
INV     gate5047  (.A(WX4883), .Z(WX3952) ) ;
OR2     gate5048  (.A(WX3943), .B(WX3942), .Z(WX3945) ) ;
INV     gate5049  (.A(WX3945), .Z(WX3954) ) ;
INV     gate5050  (.A(WX3954), .Z(WX3955) ) ;
INV     gate5051  (.A(WX4882), .Z(WX3958) ) ;
INV     gate5052  (.A(WX4883), .Z(WX3962) ) ;
INV     gate5053  (.A(WX4883), .Z(WX3966) ) ;
OR2     gate5054  (.A(WX3957), .B(WX3956), .Z(WX3959) ) ;
INV     gate5055  (.A(WX3959), .Z(WX3968) ) ;
INV     gate5056  (.A(WX3968), .Z(WX3969) ) ;
INV     gate5057  (.A(WX4882), .Z(WX3972) ) ;
INV     gate5058  (.A(WX4883), .Z(WX3976) ) ;
INV     gate5059  (.A(WX4883), .Z(WX3980) ) ;
OR2     gate5060  (.A(WX3971), .B(WX3970), .Z(WX3973) ) ;
INV     gate5061  (.A(WX3973), .Z(WX3982) ) ;
INV     gate5062  (.A(WX3982), .Z(WX3983) ) ;
INV     gate5063  (.A(WX4882), .Z(WX3986) ) ;
INV     gate5064  (.A(WX4883), .Z(WX3990) ) ;
INV     gate5065  (.A(WX4883), .Z(WX3994) ) ;
OR2     gate5066  (.A(WX3985), .B(WX3984), .Z(WX3987) ) ;
INV     gate5067  (.A(WX3987), .Z(WX3996) ) ;
INV     gate5068  (.A(WX3996), .Z(WX3997) ) ;
INV     gate5069  (.A(WX4882), .Z(WX4000) ) ;
INV     gate5070  (.A(WX4883), .Z(WX4004) ) ;
INV     gate5071  (.A(WX4883), .Z(WX4008) ) ;
OR2     gate5072  (.A(WX3999), .B(WX3998), .Z(WX4001) ) ;
INV     gate5073  (.A(WX4001), .Z(WX4010) ) ;
INV     gate5074  (.A(WX4010), .Z(WX4011) ) ;
INV     gate5075  (.A(WX4882), .Z(WX4014) ) ;
INV     gate5076  (.A(WX4883), .Z(WX4018) ) ;
INV     gate5077  (.A(WX4883), .Z(WX4022) ) ;
OR2     gate5078  (.A(WX4013), .B(WX4012), .Z(WX4015) ) ;
INV     gate5079  (.A(WX4015), .Z(WX4024) ) ;
INV     gate5080  (.A(WX4024), .Z(WX4025) ) ;
INV     gate5081  (.A(WX4882), .Z(WX4028) ) ;
INV     gate5082  (.A(WX4883), .Z(WX4032) ) ;
INV     gate5083  (.A(WX4883), .Z(WX4036) ) ;
OR2     gate5084  (.A(WX4027), .B(WX4026), .Z(WX4029) ) ;
INV     gate5085  (.A(WX4029), .Z(WX4038) ) ;
INV     gate5086  (.A(WX4038), .Z(WX4039) ) ;
INV     gate5087  (.A(WX4882), .Z(WX4042) ) ;
INV     gate5088  (.A(WX4883), .Z(WX4046) ) ;
INV     gate5089  (.A(WX4883), .Z(WX4050) ) ;
OR2     gate5090  (.A(WX4041), .B(WX4040), .Z(WX4043) ) ;
INV     gate5091  (.A(WX4043), .Z(WX4052) ) ;
INV     gate5092  (.A(WX4052), .Z(WX4053) ) ;
INV     gate5093  (.A(WX4882), .Z(WX4056) ) ;
INV     gate5094  (.A(WX4883), .Z(WX4060) ) ;
INV     gate5095  (.A(WX4883), .Z(WX4064) ) ;
OR2     gate5096  (.A(WX4055), .B(WX4054), .Z(WX4057) ) ;
INV     gate5097  (.A(WX4057), .Z(WX4066) ) ;
INV     gate5098  (.A(WX4066), .Z(WX4067) ) ;
INV     gate5099  (.A(WX4882), .Z(WX4070) ) ;
INV     gate5100  (.A(WX4883), .Z(WX4074) ) ;
INV     gate5101  (.A(WX4883), .Z(WX4078) ) ;
OR2     gate5102  (.A(WX4069), .B(WX4068), .Z(WX4071) ) ;
INV     gate5103  (.A(WX4071), .Z(WX4080) ) ;
INV     gate5104  (.A(WX4080), .Z(WX4081) ) ;
INV     gate5105  (.A(WX4882), .Z(WX4084) ) ;
INV     gate5106  (.A(WX4883), .Z(WX4088) ) ;
INV     gate5107  (.A(WX4883), .Z(WX4092) ) ;
OR2     gate5108  (.A(WX4083), .B(WX4082), .Z(WX4085) ) ;
INV     gate5109  (.A(WX4085), .Z(WX4094) ) ;
INV     gate5110  (.A(WX4094), .Z(WX4095) ) ;
INV     gate5111  (.A(WX4882), .Z(WX4098) ) ;
INV     gate5112  (.A(WX4883), .Z(WX4102) ) ;
INV     gate5113  (.A(WX4883), .Z(WX4106) ) ;
OR2     gate5114  (.A(WX4097), .B(WX4096), .Z(WX4099) ) ;
INV     gate5115  (.A(WX4099), .Z(WX4108) ) ;
INV     gate5116  (.A(WX4108), .Z(WX4109) ) ;
INV     gate5117  (.A(WX4882), .Z(WX4112) ) ;
INV     gate5118  (.A(WX4883), .Z(WX4116) ) ;
INV     gate5119  (.A(WX4883), .Z(WX4120) ) ;
OR2     gate5120  (.A(WX4111), .B(WX4110), .Z(WX4113) ) ;
INV     gate5121  (.A(WX4113), .Z(WX4122) ) ;
INV     gate5122  (.A(WX4122), .Z(WX4123) ) ;
INV     gate5123  (.A(WX4882), .Z(WX4126) ) ;
INV     gate5124  (.A(WX4883), .Z(WX4130) ) ;
INV     gate5125  (.A(WX4883), .Z(WX4134) ) ;
OR2     gate5126  (.A(WX4125), .B(WX4124), .Z(WX4127) ) ;
INV     gate5127  (.A(WX4127), .Z(WX4136) ) ;
INV     gate5128  (.A(WX4136), .Z(WX4137) ) ;
INV     gate5129  (.A(WX4882), .Z(WX4140) ) ;
INV     gate5130  (.A(WX4883), .Z(WX4144) ) ;
INV     gate5131  (.A(WX4883), .Z(WX4148) ) ;
OR2     gate5132  (.A(WX4139), .B(WX4138), .Z(WX4141) ) ;
INV     gate5133  (.A(WX4141), .Z(WX4150) ) ;
INV     gate5134  (.A(WX4150), .Z(WX4151) ) ;
INV     gate5135  (.A(WX4882), .Z(WX4154) ) ;
INV     gate5136  (.A(WX4883), .Z(WX4158) ) ;
INV     gate5137  (.A(WX4883), .Z(WX4162) ) ;
OR2     gate5138  (.A(WX4153), .B(WX4152), .Z(WX4155) ) ;
INV     gate5139  (.A(WX4155), .Z(WX4164) ) ;
INV     gate5140  (.A(WX4164), .Z(WX4165) ) ;
INV     gate5141  (.A(WX4882), .Z(WX4168) ) ;
INV     gate5142  (.A(WX4883), .Z(WX4172) ) ;
INV     gate5143  (.A(WX4883), .Z(WX4176) ) ;
OR2     gate5144  (.A(WX4167), .B(WX4166), .Z(WX4169) ) ;
INV     gate5145  (.A(WX4169), .Z(WX4178) ) ;
INV     gate5146  (.A(WX4178), .Z(WX4179) ) ;
INV     gate5147  (.A(WX4882), .Z(WX4182) ) ;
INV     gate5148  (.A(WX4883), .Z(WX4186) ) ;
INV     gate5149  (.A(WX4883), .Z(WX4190) ) ;
OR2     gate5150  (.A(WX4181), .B(WX4180), .Z(WX4183) ) ;
INV     gate5151  (.A(WX4183), .Z(WX4192) ) ;
INV     gate5152  (.A(WX4192), .Z(WX4193) ) ;
INV     gate5153  (.A(WX4882), .Z(WX4196) ) ;
INV     gate5154  (.A(WX4883), .Z(WX4200) ) ;
INV     gate5155  (.A(WX4883), .Z(WX4204) ) ;
OR2     gate5156  (.A(WX4195), .B(WX4194), .Z(WX4197) ) ;
INV     gate5157  (.A(WX4197), .Z(WX4206) ) ;
INV     gate5158  (.A(WX4206), .Z(WX4207) ) ;
INV     gate5159  (.A(WX4882), .Z(WX4210) ) ;
INV     gate5160  (.A(WX4883), .Z(WX4214) ) ;
INV     gate5161  (.A(WX4883), .Z(WX4218) ) ;
OR2     gate5162  (.A(WX4209), .B(WX4208), .Z(WX4211) ) ;
INV     gate5163  (.A(WX4211), .Z(WX4220) ) ;
INV     gate5164  (.A(WX4220), .Z(WX4221) ) ;
INV     gate5165  (.A(WX4882), .Z(WX4224) ) ;
INV     gate5166  (.A(WX4883), .Z(WX4228) ) ;
INV     gate5167  (.A(WX4883), .Z(WX4232) ) ;
OR2     gate5168  (.A(WX4223), .B(WX4222), .Z(WX4225) ) ;
INV     gate5169  (.A(WX4225), .Z(WX4234) ) ;
INV     gate5170  (.A(WX4234), .Z(WX4235) ) ;
INV     gate5171  (.A(WX4882), .Z(WX4238) ) ;
INV     gate5172  (.A(WX4883), .Z(WX4242) ) ;
INV     gate5173  (.A(WX4883), .Z(WX4246) ) ;
OR2     gate5174  (.A(WX4237), .B(WX4236), .Z(WX4239) ) ;
INV     gate5175  (.A(WX4239), .Z(WX4248) ) ;
INV     gate5176  (.A(WX4248), .Z(WX4249) ) ;
INV     gate5177  (.A(WX4882), .Z(WX4252) ) ;
INV     gate5178  (.A(WX4883), .Z(WX4256) ) ;
INV     gate5179  (.A(WX4883), .Z(WX4260) ) ;
OR2     gate5180  (.A(WX4251), .B(WX4250), .Z(WX4253) ) ;
INV     gate5181  (.A(WX4253), .Z(WX4262) ) ;
INV     gate5182  (.A(WX4262), .Z(WX4263) ) ;
INV     gate5183  (.A(WX4882), .Z(WX4266) ) ;
INV     gate5184  (.A(WX4883), .Z(WX4270) ) ;
INV     gate5185  (.A(WX4883), .Z(WX4274) ) ;
OR2     gate5186  (.A(WX4265), .B(WX4264), .Z(WX4267) ) ;
INV     gate5187  (.A(WX4267), .Z(WX4276) ) ;
INV     gate5188  (.A(WX4276), .Z(WX4277) ) ;
INV     gate5189  (.A(WX4882), .Z(WX4280) ) ;
INV     gate5190  (.A(WX4883), .Z(WX4284) ) ;
INV     gate5191  (.A(WX4883), .Z(WX4288) ) ;
OR2     gate5192  (.A(WX4279), .B(WX4278), .Z(WX4281) ) ;
INV     gate5193  (.A(WX4281), .Z(WX4290) ) ;
INV     gate5194  (.A(WX4290), .Z(WX4291) ) ;
INV     gate5195  (.A(WX4882), .Z(WX4294) ) ;
INV     gate5196  (.A(WX4883), .Z(WX4298) ) ;
INV     gate5197  (.A(WX4883), .Z(WX4302) ) ;
OR2     gate5198  (.A(WX4293), .B(WX4292), .Z(WX4295) ) ;
INV     gate5199  (.A(WX4295), .Z(WX4304) ) ;
INV     gate5200  (.A(WX4304), .Z(WX4305) ) ;
INV     gate5201  (.A(WX4882), .Z(WX4308) ) ;
INV     gate5202  (.A(WX4883), .Z(WX4312) ) ;
INV     gate5203  (.A(WX4883), .Z(WX4316) ) ;
OR2     gate5204  (.A(WX4307), .B(WX4306), .Z(WX4309) ) ;
INV     gate5205  (.A(WX4309), .Z(WX4318) ) ;
INV     gate5206  (.A(WX4318), .Z(WX4319) ) ;
INV     gate5207  (.A(WX4882), .Z(WX4322) ) ;
INV     gate5208  (.A(WX4883), .Z(WX4326) ) ;
INV     gate5209  (.A(WX4883), .Z(WX4330) ) ;
OR2     gate5210  (.A(WX4321), .B(WX4320), .Z(WX4323) ) ;
INV     gate5211  (.A(WX4323), .Z(WX4332) ) ;
INV     gate5212  (.A(WX4332), .Z(WX4333) ) ;
INV     gate5213  (.A(WX4882), .Z(WX4336) ) ;
INV     gate5214  (.A(WX4883), .Z(WX4340) ) ;
INV     gate5215  (.A(WX4883), .Z(WX4344) ) ;
OR2     gate5216  (.A(WX4335), .B(WX4334), .Z(WX4337) ) ;
INV     gate5217  (.A(WX4337), .Z(WX4346) ) ;
INV     gate5218  (.A(WX4346), .Z(WX4347) ) ;
INV     gate5219  (.A(WX4882), .Z(WX4350) ) ;
INV     gate5220  (.A(WX4883), .Z(WX4354) ) ;
INV     gate5221  (.A(WX4883), .Z(WX4358) ) ;
OR2     gate5222  (.A(WX4349), .B(WX4348), .Z(WX4351) ) ;
INV     gate5223  (.A(WX4351), .Z(WX4360) ) ;
INV     gate5224  (.A(WX4360), .Z(WX4361) ) ;
INV     gate5225  (.A(WX4364), .Z(WX4362) ) ;
INV     gate5226  (.A(WX4843), .Z(WX4844) ) ;
INV     gate5227  (.A(WX4844), .Z(WX4427) ) ;
INV     gate5228  (.A(WX4845), .Z(WX4846) ) ;
INV     gate5229  (.A(WX4846), .Z(WX4428) ) ;
INV     gate5230  (.A(WX4847), .Z(WX4848) ) ;
INV     gate5231  (.A(WX4848), .Z(WX4429) ) ;
INV     gate5232  (.A(WX4849), .Z(WX4850) ) ;
INV     gate5233  (.A(WX4850), .Z(WX4430) ) ;
INV     gate5234  (.A(WX4851), .Z(WX4852) ) ;
INV     gate5235  (.A(WX4852), .Z(WX4431) ) ;
INV     gate5236  (.A(WX4853), .Z(WX4854) ) ;
INV     gate5237  (.A(WX4854), .Z(WX4432) ) ;
INV     gate5238  (.A(WX4855), .Z(WX4856) ) ;
INV     gate5239  (.A(WX4856), .Z(WX4433) ) ;
INV     gate5240  (.A(WX4857), .Z(WX4858) ) ;
INV     gate5241  (.A(WX4858), .Z(WX4434) ) ;
INV     gate5242  (.A(WX4859), .Z(WX4860) ) ;
INV     gate5243  (.A(WX4860), .Z(WX4435) ) ;
INV     gate5244  (.A(WX4861), .Z(WX4862) ) ;
INV     gate5245  (.A(WX4862), .Z(WX4436) ) ;
INV     gate5246  (.A(WX4863), .Z(WX4864) ) ;
INV     gate5247  (.A(WX4864), .Z(WX4437) ) ;
INV     gate5248  (.A(WX4865), .Z(WX4866) ) ;
INV     gate5249  (.A(WX4866), .Z(WX4438) ) ;
INV     gate5250  (.A(WX4867), .Z(WX4868) ) ;
INV     gate5251  (.A(WX4868), .Z(WX4439) ) ;
INV     gate5252  (.A(WX4869), .Z(WX4870) ) ;
INV     gate5253  (.A(WX4870), .Z(WX4440) ) ;
INV     gate5254  (.A(WX4871), .Z(WX4872) ) ;
INV     gate5255  (.A(WX4872), .Z(WX4441) ) ;
INV     gate5256  (.A(WX4873), .Z(WX4874) ) ;
INV     gate5257  (.A(WX4874), .Z(WX4442) ) ;
INV     gate5258  (.A(WX4811), .Z(WX4812) ) ;
INV     gate5259  (.A(WX4812), .Z(WX4443) ) ;
INV     gate5260  (.A(WX4813), .Z(WX4814) ) ;
INV     gate5261  (.A(WX4814), .Z(WX4444) ) ;
INV     gate5262  (.A(WX4815), .Z(WX4816) ) ;
INV     gate5263  (.A(WX4816), .Z(WX4445) ) ;
INV     gate5264  (.A(WX4817), .Z(WX4818) ) ;
INV     gate5265  (.A(WX4818), .Z(WX4446) ) ;
INV     gate5266  (.A(WX4819), .Z(WX4820) ) ;
INV     gate5267  (.A(WX4820), .Z(WX4447) ) ;
INV     gate5268  (.A(WX4821), .Z(WX4822) ) ;
INV     gate5269  (.A(WX4822), .Z(WX4448) ) ;
INV     gate5270  (.A(WX4823), .Z(WX4824) ) ;
INV     gate5271  (.A(WX4824), .Z(WX4449) ) ;
INV     gate5272  (.A(WX4825), .Z(WX4826) ) ;
INV     gate5273  (.A(WX4826), .Z(WX4450) ) ;
INV     gate5274  (.A(WX4827), .Z(WX4828) ) ;
INV     gate5275  (.A(WX4828), .Z(WX4451) ) ;
INV     gate5276  (.A(WX4829), .Z(WX4830) ) ;
INV     gate5277  (.A(WX4830), .Z(WX4452) ) ;
INV     gate5278  (.A(WX4831), .Z(WX4832) ) ;
INV     gate5279  (.A(WX4832), .Z(WX4453) ) ;
INV     gate5280  (.A(WX4833), .Z(WX4834) ) ;
INV     gate5281  (.A(WX4834), .Z(WX4454) ) ;
INV     gate5282  (.A(WX4835), .Z(WX4836) ) ;
INV     gate5283  (.A(WX4836), .Z(WX4455) ) ;
INV     gate5284  (.A(WX4837), .Z(WX4838) ) ;
INV     gate5285  (.A(WX4838), .Z(WX4456) ) ;
INV     gate5286  (.A(WX4839), .Z(WX4840) ) ;
INV     gate5287  (.A(WX4840), .Z(WX4457) ) ;
INV     gate5288  (.A(WX4841), .Z(WX4842) ) ;
INV     gate5289  (.A(WX4842), .Z(WX4458) ) ;
INV     gate5290  (.A(WX4427), .Z(WX4459) ) ;
INV     gate5291  (.A(WX4428), .Z(WX4460) ) ;
INV     gate5292  (.A(WX4429), .Z(WX4461) ) ;
INV     gate5293  (.A(WX4430), .Z(WX4462) ) ;
INV     gate5294  (.A(WX4431), .Z(WX4463) ) ;
INV     gate5295  (.A(WX4432), .Z(WX4464) ) ;
INV     gate5296  (.A(WX4433), .Z(WX4465) ) ;
INV     gate5297  (.A(WX4434), .Z(WX4466) ) ;
INV     gate5298  (.A(WX4435), .Z(WX4467) ) ;
INV     gate5299  (.A(WX4436), .Z(WX4468) ) ;
INV     gate5300  (.A(WX4437), .Z(WX4469) ) ;
INV     gate5301  (.A(WX4438), .Z(WX4470) ) ;
INV     gate5302  (.A(WX4439), .Z(WX4471) ) ;
INV     gate5303  (.A(WX4440), .Z(WX4472) ) ;
INV     gate5304  (.A(WX4441), .Z(WX4473) ) ;
INV     gate5305  (.A(WX4442), .Z(WX4474) ) ;
INV     gate5306  (.A(WX4443), .Z(WX4475) ) ;
INV     gate5307  (.A(WX4444), .Z(WX4476) ) ;
INV     gate5308  (.A(WX4445), .Z(WX4477) ) ;
INV     gate5309  (.A(WX4446), .Z(WX4478) ) ;
INV     gate5310  (.A(WX4447), .Z(WX4479) ) ;
INV     gate5311  (.A(WX4448), .Z(WX4480) ) ;
INV     gate5312  (.A(WX4449), .Z(WX4481) ) ;
INV     gate5313  (.A(WX4450), .Z(WX4482) ) ;
INV     gate5314  (.A(WX4451), .Z(WX4483) ) ;
INV     gate5315  (.A(WX4452), .Z(WX4484) ) ;
INV     gate5316  (.A(WX4453), .Z(WX4485) ) ;
INV     gate5317  (.A(WX4454), .Z(WX4486) ) ;
INV     gate5318  (.A(WX4455), .Z(WX4487) ) ;
INV     gate5319  (.A(WX4456), .Z(WX4488) ) ;
INV     gate5320  (.A(WX4457), .Z(WX4489) ) ;
INV     gate5321  (.A(WX4458), .Z(WX4490) ) ;
INV     gate5322  (.A(WX4716), .Z(WX4491) ) ;
INV     gate5323  (.A(WX4718), .Z(WX4492) ) ;
INV     gate5324  (.A(WX4720), .Z(WX4493) ) ;
INV     gate5325  (.A(WX4722), .Z(WX4494) ) ;
INV     gate5326  (.A(WX4724), .Z(WX4495) ) ;
INV     gate5327  (.A(WX4726), .Z(WX4496) ) ;
INV     gate5328  (.A(WX4728), .Z(WX4497) ) ;
INV     gate5329  (.A(WX4730), .Z(WX4498) ) ;
INV     gate5330  (.A(WX4732), .Z(WX4499) ) ;
INV     gate5331  (.A(WX4734), .Z(WX4500) ) ;
INV     gate5332  (.A(WX4736), .Z(WX4501) ) ;
INV     gate5333  (.A(WX4738), .Z(WX4502) ) ;
INV     gate5334  (.A(WX4740), .Z(WX4503) ) ;
INV     gate5335  (.A(WX4742), .Z(WX4504) ) ;
INV     gate5336  (.A(WX4744), .Z(WX4505) ) ;
INV     gate5337  (.A(WX4746), .Z(WX4506) ) ;
INV     gate5338  (.A(WX4748), .Z(WX4507) ) ;
INV     gate5339  (.A(WX4750), .Z(WX4508) ) ;
INV     gate5340  (.A(WX4752), .Z(WX4509) ) ;
INV     gate5341  (.A(WX4754), .Z(WX4510) ) ;
INV     gate5342  (.A(WX4756), .Z(WX4511) ) ;
INV     gate5343  (.A(WX4758), .Z(WX4512) ) ;
INV     gate5344  (.A(WX4760), .Z(WX4513) ) ;
INV     gate5345  (.A(WX4762), .Z(WX4514) ) ;
INV     gate5346  (.A(WX4764), .Z(WX4515) ) ;
INV     gate5347  (.A(WX4766), .Z(WX4516) ) ;
INV     gate5348  (.A(WX4768), .Z(WX4517) ) ;
INV     gate5349  (.A(WX4770), .Z(WX4518) ) ;
INV     gate5350  (.A(WX4772), .Z(WX4519) ) ;
INV     gate5351  (.A(WX4774), .Z(WX4520) ) ;
INV     gate5352  (.A(WX4776), .Z(WX4521) ) ;
INV     gate5353  (.A(WX4778), .Z(WX4522) ) ;
NAND2   gate5354  (.A(II14522), .B(II14523), .Z(WX4795) ) ;
INV     gate5355  (.A(WX4795), .Z(WX4811) ) ;
NAND2   gate5356  (.A(II14553), .B(II14554), .Z(WX4796) ) ;
INV     gate5357  (.A(WX4796), .Z(WX4813) ) ;
NAND2   gate5358  (.A(II14584), .B(II14585), .Z(WX4797) ) ;
INV     gate5359  (.A(WX4797), .Z(WX4815) ) ;
NAND2   gate5360  (.A(II14615), .B(II14616), .Z(WX4798) ) ;
INV     gate5361  (.A(WX4798), .Z(WX4817) ) ;
NAND2   gate5362  (.A(II14646), .B(II14647), .Z(WX4799) ) ;
INV     gate5363  (.A(WX4799), .Z(WX4819) ) ;
NAND2   gate5364  (.A(II14677), .B(II14678), .Z(WX4800) ) ;
INV     gate5365  (.A(WX4800), .Z(WX4821) ) ;
NAND2   gate5366  (.A(II14708), .B(II14709), .Z(WX4801) ) ;
INV     gate5367  (.A(WX4801), .Z(WX4823) ) ;
NAND2   gate5368  (.A(II14739), .B(II14740), .Z(WX4802) ) ;
INV     gate5369  (.A(WX4802), .Z(WX4825) ) ;
NAND2   gate5370  (.A(II14770), .B(II14771), .Z(WX4803) ) ;
INV     gate5371  (.A(WX4803), .Z(WX4827) ) ;
NAND2   gate5372  (.A(II14801), .B(II14802), .Z(WX4804) ) ;
INV     gate5373  (.A(WX4804), .Z(WX4829) ) ;
NAND2   gate5374  (.A(II14832), .B(II14833), .Z(WX4805) ) ;
INV     gate5375  (.A(WX4805), .Z(WX4831) ) ;
NAND2   gate5376  (.A(II14863), .B(II14864), .Z(WX4806) ) ;
INV     gate5377  (.A(WX4806), .Z(WX4833) ) ;
NAND2   gate5378  (.A(II14894), .B(II14895), .Z(WX4807) ) ;
INV     gate5379  (.A(WX4807), .Z(WX4835) ) ;
NAND2   gate5380  (.A(II14925), .B(II14926), .Z(WX4808) ) ;
INV     gate5381  (.A(WX4808), .Z(WX4837) ) ;
NAND2   gate5382  (.A(II14956), .B(II14957), .Z(WX4809) ) ;
INV     gate5383  (.A(WX4809), .Z(WX4839) ) ;
NAND2   gate5384  (.A(II14987), .B(II14988), .Z(WX4810) ) ;
INV     gate5385  (.A(WX4810), .Z(WX4841) ) ;
NAND2   gate5386  (.A(II14026), .B(II14027), .Z(WX4779) ) ;
INV     gate5387  (.A(WX4779), .Z(WX4843) ) ;
NAND2   gate5388  (.A(II14057), .B(II14058), .Z(WX4780) ) ;
INV     gate5389  (.A(WX4780), .Z(WX4845) ) ;
NAND2   gate5390  (.A(II14088), .B(II14089), .Z(WX4781) ) ;
INV     gate5391  (.A(WX4781), .Z(WX4847) ) ;
NAND2   gate5392  (.A(II14119), .B(II14120), .Z(WX4782) ) ;
INV     gate5393  (.A(WX4782), .Z(WX4849) ) ;
NAND2   gate5394  (.A(II14150), .B(II14151), .Z(WX4783) ) ;
INV     gate5395  (.A(WX4783), .Z(WX4851) ) ;
NAND2   gate5396  (.A(II14181), .B(II14182), .Z(WX4784) ) ;
INV     gate5397  (.A(WX4784), .Z(WX4853) ) ;
NAND2   gate5398  (.A(II14212), .B(II14213), .Z(WX4785) ) ;
INV     gate5399  (.A(WX4785), .Z(WX4855) ) ;
NAND2   gate5400  (.A(II14243), .B(II14244), .Z(WX4786) ) ;
INV     gate5401  (.A(WX4786), .Z(WX4857) ) ;
NAND2   gate5402  (.A(II14274), .B(II14275), .Z(WX4787) ) ;
INV     gate5403  (.A(WX4787), .Z(WX4859) ) ;
NAND2   gate5404  (.A(II14305), .B(II14306), .Z(WX4788) ) ;
INV     gate5405  (.A(WX4788), .Z(WX4861) ) ;
NAND2   gate5406  (.A(II14336), .B(II14337), .Z(WX4789) ) ;
INV     gate5407  (.A(WX4789), .Z(WX4863) ) ;
NAND2   gate5408  (.A(II14367), .B(II14368), .Z(WX4790) ) ;
INV     gate5409  (.A(WX4790), .Z(WX4865) ) ;
NAND2   gate5410  (.A(II14398), .B(II14399), .Z(WX4791) ) ;
INV     gate5411  (.A(WX4791), .Z(WX4867) ) ;
NAND2   gate5412  (.A(II14429), .B(II14430), .Z(WX4792) ) ;
INV     gate5413  (.A(WX4792), .Z(WX4869) ) ;
NAND2   gate5414  (.A(II14460), .B(II14461), .Z(WX4793) ) ;
INV     gate5415  (.A(WX4793), .Z(WX4871) ) ;
NAND2   gate5416  (.A(II14491), .B(II14492), .Z(WX4794) ) ;
INV     gate5417  (.A(WX4794), .Z(WX4873) ) ;
INV     gate5418  (.A(TM0), .Z(WX4875) ) ;
INV     gate5419  (.A(TM0), .Z(WX4876) ) ;
INV     gate5420  (.A(TM0), .Z(WX4877) ) ;
INV     gate5421  (.A(TM1), .Z(WX4878) ) ;
INV     gate5422  (.A(TM1), .Z(WX4879) ) ;
INV     gate5423  (.A(WX4879), .Z(WX4880) ) ;
INV     gate5424  (.A(WX4877), .Z(WX4881) ) ;
INV     gate5425  (.A(WX4875), .Z(WX4884) ) ;
INV     gate5426  (.A(WX4884), .Z(WX4888) ) ;
OR2     gate5427  (.A(WX4887), .B(WX4886), .Z(WX4889) ) ;
INV     gate5428  (.A(WX4889), .Z(WX4890) ) ;
INV     gate5429  (.A(WX4890), .Z(WX4891) ) ;
INV     gate5430  (.A(WX4884), .Z(WX4895) ) ;
OR2     gate5431  (.A(WX4894), .B(WX4893), .Z(WX4896) ) ;
INV     gate5432  (.A(WX4896), .Z(WX4897) ) ;
INV     gate5433  (.A(WX4897), .Z(WX4898) ) ;
INV     gate5434  (.A(WX4884), .Z(WX4902) ) ;
OR2     gate5435  (.A(WX4901), .B(WX4900), .Z(WX4903) ) ;
INV     gate5436  (.A(WX4903), .Z(WX4904) ) ;
INV     gate5437  (.A(WX4904), .Z(WX4905) ) ;
INV     gate5438  (.A(WX4884), .Z(WX4909) ) ;
OR2     gate5439  (.A(WX4908), .B(WX4907), .Z(WX4910) ) ;
INV     gate5440  (.A(WX4910), .Z(WX4911) ) ;
INV     gate5441  (.A(WX4911), .Z(WX4912) ) ;
INV     gate5442  (.A(WX4884), .Z(WX4916) ) ;
OR2     gate5443  (.A(WX4915), .B(WX4914), .Z(WX4917) ) ;
INV     gate5444  (.A(WX4917), .Z(WX4918) ) ;
INV     gate5445  (.A(WX4918), .Z(WX4919) ) ;
INV     gate5446  (.A(WX4884), .Z(WX4923) ) ;
OR2     gate5447  (.A(WX4922), .B(WX4921), .Z(WX4924) ) ;
INV     gate5448  (.A(WX4924), .Z(WX4925) ) ;
INV     gate5449  (.A(WX4925), .Z(WX4926) ) ;
INV     gate5450  (.A(WX4884), .Z(WX4930) ) ;
OR2     gate5451  (.A(WX4929), .B(WX4928), .Z(WX4931) ) ;
INV     gate5452  (.A(WX4931), .Z(WX4932) ) ;
INV     gate5453  (.A(WX4932), .Z(WX4933) ) ;
INV     gate5454  (.A(WX4884), .Z(WX4937) ) ;
OR2     gate5455  (.A(WX4936), .B(WX4935), .Z(WX4938) ) ;
INV     gate5456  (.A(WX4938), .Z(WX4939) ) ;
INV     gate5457  (.A(WX4939), .Z(WX4940) ) ;
INV     gate5458  (.A(WX4884), .Z(WX4944) ) ;
OR2     gate5459  (.A(WX4943), .B(WX4942), .Z(WX4945) ) ;
INV     gate5460  (.A(WX4945), .Z(WX4946) ) ;
INV     gate5461  (.A(WX4946), .Z(WX4947) ) ;
INV     gate5462  (.A(WX4884), .Z(WX4951) ) ;
OR2     gate5463  (.A(WX4950), .B(WX4949), .Z(WX4952) ) ;
INV     gate5464  (.A(WX4952), .Z(WX4953) ) ;
INV     gate5465  (.A(WX4953), .Z(WX4954) ) ;
INV     gate5466  (.A(WX4884), .Z(WX4958) ) ;
OR2     gate5467  (.A(WX4957), .B(WX4956), .Z(WX4959) ) ;
INV     gate5468  (.A(WX4959), .Z(WX4960) ) ;
INV     gate5469  (.A(WX4960), .Z(WX4961) ) ;
INV     gate5470  (.A(WX4884), .Z(WX4965) ) ;
OR2     gate5471  (.A(WX4964), .B(WX4963), .Z(WX4966) ) ;
INV     gate5472  (.A(WX4966), .Z(WX4967) ) ;
INV     gate5473  (.A(WX4967), .Z(WX4968) ) ;
INV     gate5474  (.A(WX4884), .Z(WX4972) ) ;
OR2     gate5475  (.A(WX4971), .B(WX4970), .Z(WX4973) ) ;
INV     gate5476  (.A(WX4973), .Z(WX4974) ) ;
INV     gate5477  (.A(WX4974), .Z(WX4975) ) ;
INV     gate5478  (.A(WX4884), .Z(WX4979) ) ;
OR2     gate5479  (.A(WX4978), .B(WX4977), .Z(WX4980) ) ;
INV     gate5480  (.A(WX4980), .Z(WX4981) ) ;
INV     gate5481  (.A(WX4981), .Z(WX4982) ) ;
INV     gate5482  (.A(WX4884), .Z(WX4986) ) ;
OR2     gate5483  (.A(WX4985), .B(WX4984), .Z(WX4987) ) ;
INV     gate5484  (.A(WX4987), .Z(WX4988) ) ;
INV     gate5485  (.A(WX4988), .Z(WX4989) ) ;
INV     gate5486  (.A(WX4884), .Z(WX4993) ) ;
OR2     gate5487  (.A(WX4992), .B(WX4991), .Z(WX4994) ) ;
INV     gate5488  (.A(WX4994), .Z(WX4995) ) ;
INV     gate5489  (.A(WX4995), .Z(WX4996) ) ;
INV     gate5490  (.A(WX4884), .Z(WX5000) ) ;
OR2     gate5491  (.A(WX4999), .B(WX4998), .Z(WX5001) ) ;
INV     gate5492  (.A(WX5001), .Z(WX5002) ) ;
INV     gate5493  (.A(WX5002), .Z(WX5003) ) ;
INV     gate5494  (.A(WX4884), .Z(WX5007) ) ;
OR2     gate5495  (.A(WX5006), .B(WX5005), .Z(WX5008) ) ;
INV     gate5496  (.A(WX5008), .Z(WX5009) ) ;
INV     gate5497  (.A(WX5009), .Z(WX5010) ) ;
INV     gate5498  (.A(WX4884), .Z(WX5014) ) ;
OR2     gate5499  (.A(WX5013), .B(WX5012), .Z(WX5015) ) ;
INV     gate5500  (.A(WX5015), .Z(WX5016) ) ;
INV     gate5501  (.A(WX5016), .Z(WX5017) ) ;
INV     gate5502  (.A(WX4884), .Z(WX5021) ) ;
OR2     gate5503  (.A(WX5020), .B(WX5019), .Z(WX5022) ) ;
INV     gate5504  (.A(WX5022), .Z(WX5023) ) ;
INV     gate5505  (.A(WX5023), .Z(WX5024) ) ;
INV     gate5506  (.A(WX4884), .Z(WX5028) ) ;
OR2     gate5507  (.A(WX5027), .B(WX5026), .Z(WX5029) ) ;
INV     gate5508  (.A(WX5029), .Z(WX5030) ) ;
INV     gate5509  (.A(WX5030), .Z(WX5031) ) ;
INV     gate5510  (.A(WX4884), .Z(WX5035) ) ;
OR2     gate5511  (.A(WX5034), .B(WX5033), .Z(WX5036) ) ;
INV     gate5512  (.A(WX5036), .Z(WX5037) ) ;
INV     gate5513  (.A(WX5037), .Z(WX5038) ) ;
INV     gate5514  (.A(WX4884), .Z(WX5042) ) ;
OR2     gate5515  (.A(WX5041), .B(WX5040), .Z(WX5043) ) ;
INV     gate5516  (.A(WX5043), .Z(WX5044) ) ;
INV     gate5517  (.A(WX5044), .Z(WX5045) ) ;
INV     gate5518  (.A(WX4884), .Z(WX5049) ) ;
OR2     gate5519  (.A(WX5048), .B(WX5047), .Z(WX5050) ) ;
INV     gate5520  (.A(WX5050), .Z(WX5051) ) ;
INV     gate5521  (.A(WX5051), .Z(WX5052) ) ;
INV     gate5522  (.A(WX4884), .Z(WX5056) ) ;
OR2     gate5523  (.A(WX5055), .B(WX5054), .Z(WX5057) ) ;
INV     gate5524  (.A(WX5057), .Z(WX5058) ) ;
INV     gate5525  (.A(WX5058), .Z(WX5059) ) ;
INV     gate5526  (.A(WX4884), .Z(WX5063) ) ;
OR2     gate5527  (.A(WX5062), .B(WX5061), .Z(WX5064) ) ;
INV     gate5528  (.A(WX5064), .Z(WX5065) ) ;
INV     gate5529  (.A(WX5065), .Z(WX5066) ) ;
INV     gate5530  (.A(WX4884), .Z(WX5070) ) ;
OR2     gate5531  (.A(WX5069), .B(WX5068), .Z(WX5071) ) ;
INV     gate5532  (.A(WX5071), .Z(WX5072) ) ;
INV     gate5533  (.A(WX5072), .Z(WX5073) ) ;
INV     gate5534  (.A(WX4884), .Z(WX5077) ) ;
OR2     gate5535  (.A(WX5076), .B(WX5075), .Z(WX5078) ) ;
INV     gate5536  (.A(WX5078), .Z(WX5079) ) ;
INV     gate5537  (.A(WX5079), .Z(WX5080) ) ;
INV     gate5538  (.A(WX4884), .Z(WX5084) ) ;
OR2     gate5539  (.A(WX5083), .B(WX5082), .Z(WX5085) ) ;
INV     gate5540  (.A(WX5085), .Z(WX5086) ) ;
INV     gate5541  (.A(WX5086), .Z(WX5087) ) ;
INV     gate5542  (.A(WX4884), .Z(WX5091) ) ;
OR2     gate5543  (.A(WX5090), .B(WX5089), .Z(WX5092) ) ;
INV     gate5544  (.A(WX5092), .Z(WX5093) ) ;
INV     gate5545  (.A(WX5093), .Z(WX5094) ) ;
INV     gate5546  (.A(WX4884), .Z(WX5098) ) ;
OR2     gate5547  (.A(WX5097), .B(WX5096), .Z(WX5099) ) ;
INV     gate5548  (.A(WX5099), .Z(WX5100) ) ;
INV     gate5549  (.A(WX5100), .Z(WX5101) ) ;
INV     gate5550  (.A(WX4884), .Z(WX5105) ) ;
OR2     gate5551  (.A(WX5104), .B(WX5103), .Z(WX5106) ) ;
INV     gate5552  (.A(WX5106), .Z(WX5107) ) ;
INV     gate5553  (.A(WX5107), .Z(WX5108) ) ;
INV     gate5554  (.A(RESET), .Z(WX5109) ) ;
INV     gate5555  (.A(WX5109), .Z(WX5142) ) ;
INV     gate5556  (.A(WX6171), .Z(WX6175) ) ;
INV     gate5557  (.A(WX6175), .Z(WX5209) ) ;
INV     gate5558  (.A(WX6169), .Z(WX6176) ) ;
INV     gate5559  (.A(WX6176), .Z(WX5213) ) ;
INV     gate5560  (.A(WX6176), .Z(WX5217) ) ;
OR2     gate5561  (.A(WX5208), .B(WX5207), .Z(WX5210) ) ;
INV     gate5562  (.A(WX5210), .Z(WX5219) ) ;
INV     gate5563  (.A(WX5219), .Z(WX5220) ) ;
INV     gate5564  (.A(WX6175), .Z(WX5223) ) ;
INV     gate5565  (.A(WX6176), .Z(WX5227) ) ;
INV     gate5566  (.A(WX6176), .Z(WX5231) ) ;
OR2     gate5567  (.A(WX5222), .B(WX5221), .Z(WX5224) ) ;
INV     gate5568  (.A(WX5224), .Z(WX5233) ) ;
INV     gate5569  (.A(WX5233), .Z(WX5234) ) ;
INV     gate5570  (.A(WX6175), .Z(WX5237) ) ;
INV     gate5571  (.A(WX6176), .Z(WX5241) ) ;
INV     gate5572  (.A(WX6176), .Z(WX5245) ) ;
OR2     gate5573  (.A(WX5236), .B(WX5235), .Z(WX5238) ) ;
INV     gate5574  (.A(WX5238), .Z(WX5247) ) ;
INV     gate5575  (.A(WX5247), .Z(WX5248) ) ;
INV     gate5576  (.A(WX6175), .Z(WX5251) ) ;
INV     gate5577  (.A(WX6176), .Z(WX5255) ) ;
INV     gate5578  (.A(WX6176), .Z(WX5259) ) ;
OR2     gate5579  (.A(WX5250), .B(WX5249), .Z(WX5252) ) ;
INV     gate5580  (.A(WX5252), .Z(WX5261) ) ;
INV     gate5581  (.A(WX5261), .Z(WX5262) ) ;
INV     gate5582  (.A(WX6175), .Z(WX5265) ) ;
INV     gate5583  (.A(WX6176), .Z(WX5269) ) ;
INV     gate5584  (.A(WX6176), .Z(WX5273) ) ;
OR2     gate5585  (.A(WX5264), .B(WX5263), .Z(WX5266) ) ;
INV     gate5586  (.A(WX5266), .Z(WX5275) ) ;
INV     gate5587  (.A(WX5275), .Z(WX5276) ) ;
INV     gate5588  (.A(WX6175), .Z(WX5279) ) ;
INV     gate5589  (.A(WX6176), .Z(WX5283) ) ;
INV     gate5590  (.A(WX6176), .Z(WX5287) ) ;
OR2     gate5591  (.A(WX5278), .B(WX5277), .Z(WX5280) ) ;
INV     gate5592  (.A(WX5280), .Z(WX5289) ) ;
INV     gate5593  (.A(WX5289), .Z(WX5290) ) ;
INV     gate5594  (.A(WX6175), .Z(WX5293) ) ;
INV     gate5595  (.A(WX6176), .Z(WX5297) ) ;
INV     gate5596  (.A(WX6176), .Z(WX5301) ) ;
OR2     gate5597  (.A(WX5292), .B(WX5291), .Z(WX5294) ) ;
INV     gate5598  (.A(WX5294), .Z(WX5303) ) ;
INV     gate5599  (.A(WX5303), .Z(WX5304) ) ;
INV     gate5600  (.A(WX6175), .Z(WX5307) ) ;
INV     gate5601  (.A(WX6176), .Z(WX5311) ) ;
INV     gate5602  (.A(WX6176), .Z(WX5315) ) ;
OR2     gate5603  (.A(WX5306), .B(WX5305), .Z(WX5308) ) ;
INV     gate5604  (.A(WX5308), .Z(WX5317) ) ;
INV     gate5605  (.A(WX5317), .Z(WX5318) ) ;
INV     gate5606  (.A(WX6175), .Z(WX5321) ) ;
INV     gate5607  (.A(WX6176), .Z(WX5325) ) ;
INV     gate5608  (.A(WX6176), .Z(WX5329) ) ;
OR2     gate5609  (.A(WX5320), .B(WX5319), .Z(WX5322) ) ;
INV     gate5610  (.A(WX5322), .Z(WX5331) ) ;
INV     gate5611  (.A(WX5331), .Z(WX5332) ) ;
INV     gate5612  (.A(WX6175), .Z(WX5335) ) ;
INV     gate5613  (.A(WX6176), .Z(WX5339) ) ;
INV     gate5614  (.A(WX6176), .Z(WX5343) ) ;
OR2     gate5615  (.A(WX5334), .B(WX5333), .Z(WX5336) ) ;
INV     gate5616  (.A(WX5336), .Z(WX5345) ) ;
INV     gate5617  (.A(WX5345), .Z(WX5346) ) ;
INV     gate5618  (.A(WX6175), .Z(WX5349) ) ;
INV     gate5619  (.A(WX6176), .Z(WX5353) ) ;
INV     gate5620  (.A(WX6176), .Z(WX5357) ) ;
OR2     gate5621  (.A(WX5348), .B(WX5347), .Z(WX5350) ) ;
INV     gate5622  (.A(WX5350), .Z(WX5359) ) ;
INV     gate5623  (.A(WX5359), .Z(WX5360) ) ;
INV     gate5624  (.A(WX6175), .Z(WX5363) ) ;
INV     gate5625  (.A(WX6176), .Z(WX5367) ) ;
INV     gate5626  (.A(WX6176), .Z(WX5371) ) ;
OR2     gate5627  (.A(WX5362), .B(WX5361), .Z(WX5364) ) ;
INV     gate5628  (.A(WX5364), .Z(WX5373) ) ;
INV     gate5629  (.A(WX5373), .Z(WX5374) ) ;
INV     gate5630  (.A(WX6175), .Z(WX5377) ) ;
INV     gate5631  (.A(WX6176), .Z(WX5381) ) ;
INV     gate5632  (.A(WX6176), .Z(WX5385) ) ;
OR2     gate5633  (.A(WX5376), .B(WX5375), .Z(WX5378) ) ;
INV     gate5634  (.A(WX5378), .Z(WX5387) ) ;
INV     gate5635  (.A(WX5387), .Z(WX5388) ) ;
INV     gate5636  (.A(WX6175), .Z(WX5391) ) ;
INV     gate5637  (.A(WX6176), .Z(WX5395) ) ;
INV     gate5638  (.A(WX6176), .Z(WX5399) ) ;
OR2     gate5639  (.A(WX5390), .B(WX5389), .Z(WX5392) ) ;
INV     gate5640  (.A(WX5392), .Z(WX5401) ) ;
INV     gate5641  (.A(WX5401), .Z(WX5402) ) ;
INV     gate5642  (.A(WX6175), .Z(WX5405) ) ;
INV     gate5643  (.A(WX6176), .Z(WX5409) ) ;
INV     gate5644  (.A(WX6176), .Z(WX5413) ) ;
OR2     gate5645  (.A(WX5404), .B(WX5403), .Z(WX5406) ) ;
INV     gate5646  (.A(WX5406), .Z(WX5415) ) ;
INV     gate5647  (.A(WX5415), .Z(WX5416) ) ;
INV     gate5648  (.A(WX6175), .Z(WX5419) ) ;
INV     gate5649  (.A(WX6176), .Z(WX5423) ) ;
INV     gate5650  (.A(WX6176), .Z(WX5427) ) ;
OR2     gate5651  (.A(WX5418), .B(WX5417), .Z(WX5420) ) ;
INV     gate5652  (.A(WX5420), .Z(WX5429) ) ;
INV     gate5653  (.A(WX5429), .Z(WX5430) ) ;
INV     gate5654  (.A(WX6175), .Z(WX5433) ) ;
INV     gate5655  (.A(WX6176), .Z(WX5437) ) ;
INV     gate5656  (.A(WX6176), .Z(WX5441) ) ;
OR2     gate5657  (.A(WX5432), .B(WX5431), .Z(WX5434) ) ;
INV     gate5658  (.A(WX5434), .Z(WX5443) ) ;
INV     gate5659  (.A(WX5443), .Z(WX5444) ) ;
INV     gate5660  (.A(WX6175), .Z(WX5447) ) ;
INV     gate5661  (.A(WX6176), .Z(WX5451) ) ;
INV     gate5662  (.A(WX6176), .Z(WX5455) ) ;
OR2     gate5663  (.A(WX5446), .B(WX5445), .Z(WX5448) ) ;
INV     gate5664  (.A(WX5448), .Z(WX5457) ) ;
INV     gate5665  (.A(WX5457), .Z(WX5458) ) ;
INV     gate5666  (.A(WX6175), .Z(WX5461) ) ;
INV     gate5667  (.A(WX6176), .Z(WX5465) ) ;
INV     gate5668  (.A(WX6176), .Z(WX5469) ) ;
OR2     gate5669  (.A(WX5460), .B(WX5459), .Z(WX5462) ) ;
INV     gate5670  (.A(WX5462), .Z(WX5471) ) ;
INV     gate5671  (.A(WX5471), .Z(WX5472) ) ;
INV     gate5672  (.A(WX6175), .Z(WX5475) ) ;
INV     gate5673  (.A(WX6176), .Z(WX5479) ) ;
INV     gate5674  (.A(WX6176), .Z(WX5483) ) ;
OR2     gate5675  (.A(WX5474), .B(WX5473), .Z(WX5476) ) ;
INV     gate5676  (.A(WX5476), .Z(WX5485) ) ;
INV     gate5677  (.A(WX5485), .Z(WX5486) ) ;
INV     gate5678  (.A(WX6175), .Z(WX5489) ) ;
INV     gate5679  (.A(WX6176), .Z(WX5493) ) ;
INV     gate5680  (.A(WX6176), .Z(WX5497) ) ;
OR2     gate5681  (.A(WX5488), .B(WX5487), .Z(WX5490) ) ;
INV     gate5682  (.A(WX5490), .Z(WX5499) ) ;
INV     gate5683  (.A(WX5499), .Z(WX5500) ) ;
INV     gate5684  (.A(WX6175), .Z(WX5503) ) ;
INV     gate5685  (.A(WX6176), .Z(WX5507) ) ;
INV     gate5686  (.A(WX6176), .Z(WX5511) ) ;
OR2     gate5687  (.A(WX5502), .B(WX5501), .Z(WX5504) ) ;
INV     gate5688  (.A(WX5504), .Z(WX5513) ) ;
INV     gate5689  (.A(WX5513), .Z(WX5514) ) ;
INV     gate5690  (.A(WX6175), .Z(WX5517) ) ;
INV     gate5691  (.A(WX6176), .Z(WX5521) ) ;
INV     gate5692  (.A(WX6176), .Z(WX5525) ) ;
OR2     gate5693  (.A(WX5516), .B(WX5515), .Z(WX5518) ) ;
INV     gate5694  (.A(WX5518), .Z(WX5527) ) ;
INV     gate5695  (.A(WX5527), .Z(WX5528) ) ;
INV     gate5696  (.A(WX6175), .Z(WX5531) ) ;
INV     gate5697  (.A(WX6176), .Z(WX5535) ) ;
INV     gate5698  (.A(WX6176), .Z(WX5539) ) ;
OR2     gate5699  (.A(WX5530), .B(WX5529), .Z(WX5532) ) ;
INV     gate5700  (.A(WX5532), .Z(WX5541) ) ;
INV     gate5701  (.A(WX5541), .Z(WX5542) ) ;
INV     gate5702  (.A(WX6175), .Z(WX5545) ) ;
INV     gate5703  (.A(WX6176), .Z(WX5549) ) ;
INV     gate5704  (.A(WX6176), .Z(WX5553) ) ;
OR2     gate5705  (.A(WX5544), .B(WX5543), .Z(WX5546) ) ;
INV     gate5706  (.A(WX5546), .Z(WX5555) ) ;
INV     gate5707  (.A(WX5555), .Z(WX5556) ) ;
INV     gate5708  (.A(WX6175), .Z(WX5559) ) ;
INV     gate5709  (.A(WX6176), .Z(WX5563) ) ;
INV     gate5710  (.A(WX6176), .Z(WX5567) ) ;
OR2     gate5711  (.A(WX5558), .B(WX5557), .Z(WX5560) ) ;
INV     gate5712  (.A(WX5560), .Z(WX5569) ) ;
INV     gate5713  (.A(WX5569), .Z(WX5570) ) ;
INV     gate5714  (.A(WX6175), .Z(WX5573) ) ;
INV     gate5715  (.A(WX6176), .Z(WX5577) ) ;
INV     gate5716  (.A(WX6176), .Z(WX5581) ) ;
OR2     gate5717  (.A(WX5572), .B(WX5571), .Z(WX5574) ) ;
INV     gate5718  (.A(WX5574), .Z(WX5583) ) ;
INV     gate5719  (.A(WX5583), .Z(WX5584) ) ;
INV     gate5720  (.A(WX6175), .Z(WX5587) ) ;
INV     gate5721  (.A(WX6176), .Z(WX5591) ) ;
INV     gate5722  (.A(WX6176), .Z(WX5595) ) ;
OR2     gate5723  (.A(WX5586), .B(WX5585), .Z(WX5588) ) ;
INV     gate5724  (.A(WX5588), .Z(WX5597) ) ;
INV     gate5725  (.A(WX5597), .Z(WX5598) ) ;
INV     gate5726  (.A(WX6175), .Z(WX5601) ) ;
INV     gate5727  (.A(WX6176), .Z(WX5605) ) ;
INV     gate5728  (.A(WX6176), .Z(WX5609) ) ;
OR2     gate5729  (.A(WX5600), .B(WX5599), .Z(WX5602) ) ;
INV     gate5730  (.A(WX5602), .Z(WX5611) ) ;
INV     gate5731  (.A(WX5611), .Z(WX5612) ) ;
INV     gate5732  (.A(WX6175), .Z(WX5615) ) ;
INV     gate5733  (.A(WX6176), .Z(WX5619) ) ;
INV     gate5734  (.A(WX6176), .Z(WX5623) ) ;
OR2     gate5735  (.A(WX5614), .B(WX5613), .Z(WX5616) ) ;
INV     gate5736  (.A(WX5616), .Z(WX5625) ) ;
INV     gate5737  (.A(WX5625), .Z(WX5626) ) ;
INV     gate5738  (.A(WX6175), .Z(WX5629) ) ;
INV     gate5739  (.A(WX6176), .Z(WX5633) ) ;
INV     gate5740  (.A(WX6176), .Z(WX5637) ) ;
OR2     gate5741  (.A(WX5628), .B(WX5627), .Z(WX5630) ) ;
INV     gate5742  (.A(WX5630), .Z(WX5639) ) ;
INV     gate5743  (.A(WX5639), .Z(WX5640) ) ;
INV     gate5744  (.A(WX6175), .Z(WX5643) ) ;
INV     gate5745  (.A(WX6176), .Z(WX5647) ) ;
INV     gate5746  (.A(WX6176), .Z(WX5651) ) ;
OR2     gate5747  (.A(WX5642), .B(WX5641), .Z(WX5644) ) ;
INV     gate5748  (.A(WX5644), .Z(WX5653) ) ;
INV     gate5749  (.A(WX5653), .Z(WX5654) ) ;
INV     gate5750  (.A(WX5657), .Z(WX5655) ) ;
INV     gate5751  (.A(WX6136), .Z(WX6137) ) ;
INV     gate5752  (.A(WX6137), .Z(WX5720) ) ;
INV     gate5753  (.A(WX6138), .Z(WX6139) ) ;
INV     gate5754  (.A(WX6139), .Z(WX5721) ) ;
INV     gate5755  (.A(WX6140), .Z(WX6141) ) ;
INV     gate5756  (.A(WX6141), .Z(WX5722) ) ;
INV     gate5757  (.A(WX6142), .Z(WX6143) ) ;
INV     gate5758  (.A(WX6143), .Z(WX5723) ) ;
INV     gate5759  (.A(WX6144), .Z(WX6145) ) ;
INV     gate5760  (.A(WX6145), .Z(WX5724) ) ;
INV     gate5761  (.A(WX6146), .Z(WX6147) ) ;
INV     gate5762  (.A(WX6147), .Z(WX5725) ) ;
INV     gate5763  (.A(WX6148), .Z(WX6149) ) ;
INV     gate5764  (.A(WX6149), .Z(WX5726) ) ;
INV     gate5765  (.A(WX6150), .Z(WX6151) ) ;
INV     gate5766  (.A(WX6151), .Z(WX5727) ) ;
INV     gate5767  (.A(WX6152), .Z(WX6153) ) ;
INV     gate5768  (.A(WX6153), .Z(WX5728) ) ;
INV     gate5769  (.A(WX6154), .Z(WX6155) ) ;
INV     gate5770  (.A(WX6155), .Z(WX5729) ) ;
INV     gate5771  (.A(WX6156), .Z(WX6157) ) ;
INV     gate5772  (.A(WX6157), .Z(WX5730) ) ;
INV     gate5773  (.A(WX6158), .Z(WX6159) ) ;
INV     gate5774  (.A(WX6159), .Z(WX5731) ) ;
INV     gate5775  (.A(WX6160), .Z(WX6161) ) ;
INV     gate5776  (.A(WX6161), .Z(WX5732) ) ;
INV     gate5777  (.A(WX6162), .Z(WX6163) ) ;
INV     gate5778  (.A(WX6163), .Z(WX5733) ) ;
INV     gate5779  (.A(WX6164), .Z(WX6165) ) ;
INV     gate5780  (.A(WX6165), .Z(WX5734) ) ;
INV     gate5781  (.A(WX6166), .Z(WX6167) ) ;
INV     gate5782  (.A(WX6167), .Z(WX5735) ) ;
INV     gate5783  (.A(WX6104), .Z(WX6105) ) ;
INV     gate5784  (.A(WX6105), .Z(WX5736) ) ;
INV     gate5785  (.A(WX6106), .Z(WX6107) ) ;
INV     gate5786  (.A(WX6107), .Z(WX5737) ) ;
INV     gate5787  (.A(WX6108), .Z(WX6109) ) ;
INV     gate5788  (.A(WX6109), .Z(WX5738) ) ;
INV     gate5789  (.A(WX6110), .Z(WX6111) ) ;
INV     gate5790  (.A(WX6111), .Z(WX5739) ) ;
INV     gate5791  (.A(WX6112), .Z(WX6113) ) ;
INV     gate5792  (.A(WX6113), .Z(WX5740) ) ;
INV     gate5793  (.A(WX6114), .Z(WX6115) ) ;
INV     gate5794  (.A(WX6115), .Z(WX5741) ) ;
INV     gate5795  (.A(WX6116), .Z(WX6117) ) ;
INV     gate5796  (.A(WX6117), .Z(WX5742) ) ;
INV     gate5797  (.A(WX6118), .Z(WX6119) ) ;
INV     gate5798  (.A(WX6119), .Z(WX5743) ) ;
INV     gate5799  (.A(WX6120), .Z(WX6121) ) ;
INV     gate5800  (.A(WX6121), .Z(WX5744) ) ;
INV     gate5801  (.A(WX6122), .Z(WX6123) ) ;
INV     gate5802  (.A(WX6123), .Z(WX5745) ) ;
INV     gate5803  (.A(WX6124), .Z(WX6125) ) ;
INV     gate5804  (.A(WX6125), .Z(WX5746) ) ;
INV     gate5805  (.A(WX6126), .Z(WX6127) ) ;
INV     gate5806  (.A(WX6127), .Z(WX5747) ) ;
INV     gate5807  (.A(WX6128), .Z(WX6129) ) ;
INV     gate5808  (.A(WX6129), .Z(WX5748) ) ;
INV     gate5809  (.A(WX6130), .Z(WX6131) ) ;
INV     gate5810  (.A(WX6131), .Z(WX5749) ) ;
INV     gate5811  (.A(WX6132), .Z(WX6133) ) ;
INV     gate5812  (.A(WX6133), .Z(WX5750) ) ;
INV     gate5813  (.A(WX6134), .Z(WX6135) ) ;
INV     gate5814  (.A(WX6135), .Z(WX5751) ) ;
INV     gate5815  (.A(WX5720), .Z(WX5752) ) ;
INV     gate5816  (.A(WX5721), .Z(WX5753) ) ;
INV     gate5817  (.A(WX5722), .Z(WX5754) ) ;
INV     gate5818  (.A(WX5723), .Z(WX5755) ) ;
INV     gate5819  (.A(WX5724), .Z(WX5756) ) ;
INV     gate5820  (.A(WX5725), .Z(WX5757) ) ;
INV     gate5821  (.A(WX5726), .Z(WX5758) ) ;
INV     gate5822  (.A(WX5727), .Z(WX5759) ) ;
INV     gate5823  (.A(WX5728), .Z(WX5760) ) ;
INV     gate5824  (.A(WX5729), .Z(WX5761) ) ;
INV     gate5825  (.A(WX5730), .Z(WX5762) ) ;
INV     gate5826  (.A(WX5731), .Z(WX5763) ) ;
INV     gate5827  (.A(WX5732), .Z(WX5764) ) ;
INV     gate5828  (.A(WX5733), .Z(WX5765) ) ;
INV     gate5829  (.A(WX5734), .Z(WX5766) ) ;
INV     gate5830  (.A(WX5735), .Z(WX5767) ) ;
INV     gate5831  (.A(WX5736), .Z(WX5768) ) ;
INV     gate5832  (.A(WX5737), .Z(WX5769) ) ;
INV     gate5833  (.A(WX5738), .Z(WX5770) ) ;
INV     gate5834  (.A(WX5739), .Z(WX5771) ) ;
INV     gate5835  (.A(WX5740), .Z(WX5772) ) ;
INV     gate5836  (.A(WX5741), .Z(WX5773) ) ;
INV     gate5837  (.A(WX5742), .Z(WX5774) ) ;
INV     gate5838  (.A(WX5743), .Z(WX5775) ) ;
INV     gate5839  (.A(WX5744), .Z(WX5776) ) ;
INV     gate5840  (.A(WX5745), .Z(WX5777) ) ;
INV     gate5841  (.A(WX5746), .Z(WX5778) ) ;
INV     gate5842  (.A(WX5747), .Z(WX5779) ) ;
INV     gate5843  (.A(WX5748), .Z(WX5780) ) ;
INV     gate5844  (.A(WX5749), .Z(WX5781) ) ;
INV     gate5845  (.A(WX5750), .Z(WX5782) ) ;
INV     gate5846  (.A(WX5751), .Z(WX5783) ) ;
INV     gate5847  (.A(WX6009), .Z(WX5784) ) ;
INV     gate5848  (.A(WX6011), .Z(WX5785) ) ;
INV     gate5849  (.A(WX6013), .Z(WX5786) ) ;
INV     gate5850  (.A(WX6015), .Z(WX5787) ) ;
INV     gate5851  (.A(WX6017), .Z(WX5788) ) ;
INV     gate5852  (.A(WX6019), .Z(WX5789) ) ;
INV     gate5853  (.A(WX6021), .Z(WX5790) ) ;
INV     gate5854  (.A(WX6023), .Z(WX5791) ) ;
INV     gate5855  (.A(WX6025), .Z(WX5792) ) ;
INV     gate5856  (.A(WX6027), .Z(WX5793) ) ;
INV     gate5857  (.A(WX6029), .Z(WX5794) ) ;
INV     gate5858  (.A(WX6031), .Z(WX5795) ) ;
INV     gate5859  (.A(WX6033), .Z(WX5796) ) ;
INV     gate5860  (.A(WX6035), .Z(WX5797) ) ;
INV     gate5861  (.A(WX6037), .Z(WX5798) ) ;
INV     gate5862  (.A(WX6039), .Z(WX5799) ) ;
INV     gate5863  (.A(WX6041), .Z(WX5800) ) ;
INV     gate5864  (.A(WX6043), .Z(WX5801) ) ;
INV     gate5865  (.A(WX6045), .Z(WX5802) ) ;
INV     gate5866  (.A(WX6047), .Z(WX5803) ) ;
INV     gate5867  (.A(WX6049), .Z(WX5804) ) ;
INV     gate5868  (.A(WX6051), .Z(WX5805) ) ;
INV     gate5869  (.A(WX6053), .Z(WX5806) ) ;
INV     gate5870  (.A(WX6055), .Z(WX5807) ) ;
INV     gate5871  (.A(WX6057), .Z(WX5808) ) ;
INV     gate5872  (.A(WX6059), .Z(WX5809) ) ;
INV     gate5873  (.A(WX6061), .Z(WX5810) ) ;
INV     gate5874  (.A(WX6063), .Z(WX5811) ) ;
INV     gate5875  (.A(WX6065), .Z(WX5812) ) ;
INV     gate5876  (.A(WX6067), .Z(WX5813) ) ;
INV     gate5877  (.A(WX6069), .Z(WX5814) ) ;
INV     gate5878  (.A(WX6071), .Z(WX5815) ) ;
NAND2   gate5879  (.A(II18527), .B(II18528), .Z(WX6088) ) ;
INV     gate5880  (.A(WX6088), .Z(WX6104) ) ;
NAND2   gate5881  (.A(II18558), .B(II18559), .Z(WX6089) ) ;
INV     gate5882  (.A(WX6089), .Z(WX6106) ) ;
NAND2   gate5883  (.A(II18589), .B(II18590), .Z(WX6090) ) ;
INV     gate5884  (.A(WX6090), .Z(WX6108) ) ;
NAND2   gate5885  (.A(II18620), .B(II18621), .Z(WX6091) ) ;
INV     gate5886  (.A(WX6091), .Z(WX6110) ) ;
NAND2   gate5887  (.A(II18651), .B(II18652), .Z(WX6092) ) ;
INV     gate5888  (.A(WX6092), .Z(WX6112) ) ;
NAND2   gate5889  (.A(II18682), .B(II18683), .Z(WX6093) ) ;
INV     gate5890  (.A(WX6093), .Z(WX6114) ) ;
NAND2   gate5891  (.A(II18713), .B(II18714), .Z(WX6094) ) ;
INV     gate5892  (.A(WX6094), .Z(WX6116) ) ;
NAND2   gate5893  (.A(II18744), .B(II18745), .Z(WX6095) ) ;
INV     gate5894  (.A(WX6095), .Z(WX6118) ) ;
NAND2   gate5895  (.A(II18775), .B(II18776), .Z(WX6096) ) ;
INV     gate5896  (.A(WX6096), .Z(WX6120) ) ;
NAND2   gate5897  (.A(II18806), .B(II18807), .Z(WX6097) ) ;
INV     gate5898  (.A(WX6097), .Z(WX6122) ) ;
NAND2   gate5899  (.A(II18837), .B(II18838), .Z(WX6098) ) ;
INV     gate5900  (.A(WX6098), .Z(WX6124) ) ;
NAND2   gate5901  (.A(II18868), .B(II18869), .Z(WX6099) ) ;
INV     gate5902  (.A(WX6099), .Z(WX6126) ) ;
NAND2   gate5903  (.A(II18899), .B(II18900), .Z(WX6100) ) ;
INV     gate5904  (.A(WX6100), .Z(WX6128) ) ;
NAND2   gate5905  (.A(II18930), .B(II18931), .Z(WX6101) ) ;
INV     gate5906  (.A(WX6101), .Z(WX6130) ) ;
NAND2   gate5907  (.A(II18961), .B(II18962), .Z(WX6102) ) ;
INV     gate5908  (.A(WX6102), .Z(WX6132) ) ;
NAND2   gate5909  (.A(II18992), .B(II18993), .Z(WX6103) ) ;
INV     gate5910  (.A(WX6103), .Z(WX6134) ) ;
NAND2   gate5911  (.A(II18031), .B(II18032), .Z(WX6072) ) ;
INV     gate5912  (.A(WX6072), .Z(WX6136) ) ;
NAND2   gate5913  (.A(II18062), .B(II18063), .Z(WX6073) ) ;
INV     gate5914  (.A(WX6073), .Z(WX6138) ) ;
NAND2   gate5915  (.A(II18093), .B(II18094), .Z(WX6074) ) ;
INV     gate5916  (.A(WX6074), .Z(WX6140) ) ;
NAND2   gate5917  (.A(II18124), .B(II18125), .Z(WX6075) ) ;
INV     gate5918  (.A(WX6075), .Z(WX6142) ) ;
NAND2   gate5919  (.A(II18155), .B(II18156), .Z(WX6076) ) ;
INV     gate5920  (.A(WX6076), .Z(WX6144) ) ;
NAND2   gate5921  (.A(II18186), .B(II18187), .Z(WX6077) ) ;
INV     gate5922  (.A(WX6077), .Z(WX6146) ) ;
NAND2   gate5923  (.A(II18217), .B(II18218), .Z(WX6078) ) ;
INV     gate5924  (.A(WX6078), .Z(WX6148) ) ;
NAND2   gate5925  (.A(II18248), .B(II18249), .Z(WX6079) ) ;
INV     gate5926  (.A(WX6079), .Z(WX6150) ) ;
NAND2   gate5927  (.A(II18279), .B(II18280), .Z(WX6080) ) ;
INV     gate5928  (.A(WX6080), .Z(WX6152) ) ;
NAND2   gate5929  (.A(II18310), .B(II18311), .Z(WX6081) ) ;
INV     gate5930  (.A(WX6081), .Z(WX6154) ) ;
NAND2   gate5931  (.A(II18341), .B(II18342), .Z(WX6082) ) ;
INV     gate5932  (.A(WX6082), .Z(WX6156) ) ;
NAND2   gate5933  (.A(II18372), .B(II18373), .Z(WX6083) ) ;
INV     gate5934  (.A(WX6083), .Z(WX6158) ) ;
NAND2   gate5935  (.A(II18403), .B(II18404), .Z(WX6084) ) ;
INV     gate5936  (.A(WX6084), .Z(WX6160) ) ;
NAND2   gate5937  (.A(II18434), .B(II18435), .Z(WX6085) ) ;
INV     gate5938  (.A(WX6085), .Z(WX6162) ) ;
NAND2   gate5939  (.A(II18465), .B(II18466), .Z(WX6086) ) ;
INV     gate5940  (.A(WX6086), .Z(WX6164) ) ;
NAND2   gate5941  (.A(II18496), .B(II18497), .Z(WX6087) ) ;
INV     gate5942  (.A(WX6087), .Z(WX6166) ) ;
INV     gate5943  (.A(TM0), .Z(WX6168) ) ;
INV     gate5944  (.A(TM0), .Z(WX6169) ) ;
INV     gate5945  (.A(TM0), .Z(WX6170) ) ;
INV     gate5946  (.A(TM1), .Z(WX6171) ) ;
INV     gate5947  (.A(TM1), .Z(WX6172) ) ;
INV     gate5948  (.A(WX6172), .Z(WX6173) ) ;
INV     gate5949  (.A(WX6170), .Z(WX6174) ) ;
INV     gate5950  (.A(WX6168), .Z(WX6177) ) ;
INV     gate5951  (.A(WX6177), .Z(WX6181) ) ;
OR2     gate5952  (.A(WX6180), .B(WX6179), .Z(WX6182) ) ;
INV     gate5953  (.A(WX6182), .Z(WX6183) ) ;
INV     gate5954  (.A(WX6183), .Z(WX6184) ) ;
INV     gate5955  (.A(WX6177), .Z(WX6188) ) ;
OR2     gate5956  (.A(WX6187), .B(WX6186), .Z(WX6189) ) ;
INV     gate5957  (.A(WX6189), .Z(WX6190) ) ;
INV     gate5958  (.A(WX6190), .Z(WX6191) ) ;
INV     gate5959  (.A(WX6177), .Z(WX6195) ) ;
OR2     gate5960  (.A(WX6194), .B(WX6193), .Z(WX6196) ) ;
INV     gate5961  (.A(WX6196), .Z(WX6197) ) ;
INV     gate5962  (.A(WX6197), .Z(WX6198) ) ;
INV     gate5963  (.A(WX6177), .Z(WX6202) ) ;
OR2     gate5964  (.A(WX6201), .B(WX6200), .Z(WX6203) ) ;
INV     gate5965  (.A(WX6203), .Z(WX6204) ) ;
INV     gate5966  (.A(WX6204), .Z(WX6205) ) ;
INV     gate5967  (.A(WX6177), .Z(WX6209) ) ;
OR2     gate5968  (.A(WX6208), .B(WX6207), .Z(WX6210) ) ;
INV     gate5969  (.A(WX6210), .Z(WX6211) ) ;
INV     gate5970  (.A(WX6211), .Z(WX6212) ) ;
INV     gate5971  (.A(WX6177), .Z(WX6216) ) ;
OR2     gate5972  (.A(WX6215), .B(WX6214), .Z(WX6217) ) ;
INV     gate5973  (.A(WX6217), .Z(WX6218) ) ;
INV     gate5974  (.A(WX6218), .Z(WX6219) ) ;
INV     gate5975  (.A(WX6177), .Z(WX6223) ) ;
OR2     gate5976  (.A(WX6222), .B(WX6221), .Z(WX6224) ) ;
INV     gate5977  (.A(WX6224), .Z(WX6225) ) ;
INV     gate5978  (.A(WX6225), .Z(WX6226) ) ;
INV     gate5979  (.A(WX6177), .Z(WX6230) ) ;
OR2     gate5980  (.A(WX6229), .B(WX6228), .Z(WX6231) ) ;
INV     gate5981  (.A(WX6231), .Z(WX6232) ) ;
INV     gate5982  (.A(WX6232), .Z(WX6233) ) ;
INV     gate5983  (.A(WX6177), .Z(WX6237) ) ;
OR2     gate5984  (.A(WX6236), .B(WX6235), .Z(WX6238) ) ;
INV     gate5985  (.A(WX6238), .Z(WX6239) ) ;
INV     gate5986  (.A(WX6239), .Z(WX6240) ) ;
INV     gate5987  (.A(WX6177), .Z(WX6244) ) ;
OR2     gate5988  (.A(WX6243), .B(WX6242), .Z(WX6245) ) ;
INV     gate5989  (.A(WX6245), .Z(WX6246) ) ;
INV     gate5990  (.A(WX6246), .Z(WX6247) ) ;
INV     gate5991  (.A(WX6177), .Z(WX6251) ) ;
OR2     gate5992  (.A(WX6250), .B(WX6249), .Z(WX6252) ) ;
INV     gate5993  (.A(WX6252), .Z(WX6253) ) ;
INV     gate5994  (.A(WX6253), .Z(WX6254) ) ;
INV     gate5995  (.A(WX6177), .Z(WX6258) ) ;
OR2     gate5996  (.A(WX6257), .B(WX6256), .Z(WX6259) ) ;
INV     gate5997  (.A(WX6259), .Z(WX6260) ) ;
INV     gate5998  (.A(WX6260), .Z(WX6261) ) ;
INV     gate5999  (.A(WX6177), .Z(WX6265) ) ;
OR2     gate6000  (.A(WX6264), .B(WX6263), .Z(WX6266) ) ;
INV     gate6001  (.A(WX6266), .Z(WX6267) ) ;
INV     gate6002  (.A(WX6267), .Z(WX6268) ) ;
INV     gate6003  (.A(WX6177), .Z(WX6272) ) ;
OR2     gate6004  (.A(WX6271), .B(WX6270), .Z(WX6273) ) ;
INV     gate6005  (.A(WX6273), .Z(WX6274) ) ;
INV     gate6006  (.A(WX6274), .Z(WX6275) ) ;
INV     gate6007  (.A(WX6177), .Z(WX6279) ) ;
OR2     gate6008  (.A(WX6278), .B(WX6277), .Z(WX6280) ) ;
INV     gate6009  (.A(WX6280), .Z(WX6281) ) ;
INV     gate6010  (.A(WX6281), .Z(WX6282) ) ;
INV     gate6011  (.A(WX6177), .Z(WX6286) ) ;
OR2     gate6012  (.A(WX6285), .B(WX6284), .Z(WX6287) ) ;
INV     gate6013  (.A(WX6287), .Z(WX6288) ) ;
INV     gate6014  (.A(WX6288), .Z(WX6289) ) ;
INV     gate6015  (.A(WX6177), .Z(WX6293) ) ;
OR2     gate6016  (.A(WX6292), .B(WX6291), .Z(WX6294) ) ;
INV     gate6017  (.A(WX6294), .Z(WX6295) ) ;
INV     gate6018  (.A(WX6295), .Z(WX6296) ) ;
INV     gate6019  (.A(WX6177), .Z(WX6300) ) ;
OR2     gate6020  (.A(WX6299), .B(WX6298), .Z(WX6301) ) ;
INV     gate6021  (.A(WX6301), .Z(WX6302) ) ;
INV     gate6022  (.A(WX6302), .Z(WX6303) ) ;
INV     gate6023  (.A(WX6177), .Z(WX6307) ) ;
OR2     gate6024  (.A(WX6306), .B(WX6305), .Z(WX6308) ) ;
INV     gate6025  (.A(WX6308), .Z(WX6309) ) ;
INV     gate6026  (.A(WX6309), .Z(WX6310) ) ;
INV     gate6027  (.A(WX6177), .Z(WX6314) ) ;
OR2     gate6028  (.A(WX6313), .B(WX6312), .Z(WX6315) ) ;
INV     gate6029  (.A(WX6315), .Z(WX6316) ) ;
INV     gate6030  (.A(WX6316), .Z(WX6317) ) ;
INV     gate6031  (.A(WX6177), .Z(WX6321) ) ;
OR2     gate6032  (.A(WX6320), .B(WX6319), .Z(WX6322) ) ;
INV     gate6033  (.A(WX6322), .Z(WX6323) ) ;
INV     gate6034  (.A(WX6323), .Z(WX6324) ) ;
INV     gate6035  (.A(WX6177), .Z(WX6328) ) ;
OR2     gate6036  (.A(WX6327), .B(WX6326), .Z(WX6329) ) ;
INV     gate6037  (.A(WX6329), .Z(WX6330) ) ;
INV     gate6038  (.A(WX6330), .Z(WX6331) ) ;
INV     gate6039  (.A(WX6177), .Z(WX6335) ) ;
OR2     gate6040  (.A(WX6334), .B(WX6333), .Z(WX6336) ) ;
INV     gate6041  (.A(WX6336), .Z(WX6337) ) ;
INV     gate6042  (.A(WX6337), .Z(WX6338) ) ;
INV     gate6043  (.A(WX6177), .Z(WX6342) ) ;
OR2     gate6044  (.A(WX6341), .B(WX6340), .Z(WX6343) ) ;
INV     gate6045  (.A(WX6343), .Z(WX6344) ) ;
INV     gate6046  (.A(WX6344), .Z(WX6345) ) ;
INV     gate6047  (.A(WX6177), .Z(WX6349) ) ;
OR2     gate6048  (.A(WX6348), .B(WX6347), .Z(WX6350) ) ;
INV     gate6049  (.A(WX6350), .Z(WX6351) ) ;
INV     gate6050  (.A(WX6351), .Z(WX6352) ) ;
INV     gate6051  (.A(WX6177), .Z(WX6356) ) ;
OR2     gate6052  (.A(WX6355), .B(WX6354), .Z(WX6357) ) ;
INV     gate6053  (.A(WX6357), .Z(WX6358) ) ;
INV     gate6054  (.A(WX6358), .Z(WX6359) ) ;
INV     gate6055  (.A(WX6177), .Z(WX6363) ) ;
OR2     gate6056  (.A(WX6362), .B(WX6361), .Z(WX6364) ) ;
INV     gate6057  (.A(WX6364), .Z(WX6365) ) ;
INV     gate6058  (.A(WX6365), .Z(WX6366) ) ;
INV     gate6059  (.A(WX6177), .Z(WX6370) ) ;
OR2     gate6060  (.A(WX6369), .B(WX6368), .Z(WX6371) ) ;
INV     gate6061  (.A(WX6371), .Z(WX6372) ) ;
INV     gate6062  (.A(WX6372), .Z(WX6373) ) ;
INV     gate6063  (.A(WX6177), .Z(WX6377) ) ;
OR2     gate6064  (.A(WX6376), .B(WX6375), .Z(WX6378) ) ;
INV     gate6065  (.A(WX6378), .Z(WX6379) ) ;
INV     gate6066  (.A(WX6379), .Z(WX6380) ) ;
INV     gate6067  (.A(WX6177), .Z(WX6384) ) ;
OR2     gate6068  (.A(WX6383), .B(WX6382), .Z(WX6385) ) ;
INV     gate6069  (.A(WX6385), .Z(WX6386) ) ;
INV     gate6070  (.A(WX6386), .Z(WX6387) ) ;
INV     gate6071  (.A(WX6177), .Z(WX6391) ) ;
OR2     gate6072  (.A(WX6390), .B(WX6389), .Z(WX6392) ) ;
INV     gate6073  (.A(WX6392), .Z(WX6393) ) ;
INV     gate6074  (.A(WX6393), .Z(WX6394) ) ;
INV     gate6075  (.A(WX6177), .Z(WX6398) ) ;
OR2     gate6076  (.A(WX6397), .B(WX6396), .Z(WX6399) ) ;
INV     gate6077  (.A(WX6399), .Z(WX6400) ) ;
INV     gate6078  (.A(WX6400), .Z(WX6401) ) ;
INV     gate6079  (.A(RESET), .Z(WX6402) ) ;
INV     gate6080  (.A(WX6402), .Z(WX6435) ) ;
INV     gate6081  (.A(WX7464), .Z(WX7468) ) ;
INV     gate6082  (.A(WX7468), .Z(WX6502) ) ;
INV     gate6083  (.A(WX7462), .Z(WX7469) ) ;
INV     gate6084  (.A(WX7469), .Z(WX6506) ) ;
INV     gate6085  (.A(WX7469), .Z(WX6510) ) ;
OR2     gate6086  (.A(WX6501), .B(WX6500), .Z(WX6503) ) ;
INV     gate6087  (.A(WX6503), .Z(WX6512) ) ;
INV     gate6088  (.A(WX6512), .Z(WX6513) ) ;
INV     gate6089  (.A(WX7468), .Z(WX6516) ) ;
INV     gate6090  (.A(WX7469), .Z(WX6520) ) ;
INV     gate6091  (.A(WX7469), .Z(WX6524) ) ;
OR2     gate6092  (.A(WX6515), .B(WX6514), .Z(WX6517) ) ;
INV     gate6093  (.A(WX6517), .Z(WX6526) ) ;
INV     gate6094  (.A(WX6526), .Z(WX6527) ) ;
INV     gate6095  (.A(WX7468), .Z(WX6530) ) ;
INV     gate6096  (.A(WX7469), .Z(WX6534) ) ;
INV     gate6097  (.A(WX7469), .Z(WX6538) ) ;
OR2     gate6098  (.A(WX6529), .B(WX6528), .Z(WX6531) ) ;
INV     gate6099  (.A(WX6531), .Z(WX6540) ) ;
INV     gate6100  (.A(WX6540), .Z(WX6541) ) ;
INV     gate6101  (.A(WX7468), .Z(WX6544) ) ;
INV     gate6102  (.A(WX7469), .Z(WX6548) ) ;
INV     gate6103  (.A(WX7469), .Z(WX6552) ) ;
OR2     gate6104  (.A(WX6543), .B(WX6542), .Z(WX6545) ) ;
INV     gate6105  (.A(WX6545), .Z(WX6554) ) ;
INV     gate6106  (.A(WX6554), .Z(WX6555) ) ;
INV     gate6107  (.A(WX7468), .Z(WX6558) ) ;
INV     gate6108  (.A(WX7469), .Z(WX6562) ) ;
INV     gate6109  (.A(WX7469), .Z(WX6566) ) ;
OR2     gate6110  (.A(WX6557), .B(WX6556), .Z(WX6559) ) ;
INV     gate6111  (.A(WX6559), .Z(WX6568) ) ;
INV     gate6112  (.A(WX6568), .Z(WX6569) ) ;
INV     gate6113  (.A(WX7468), .Z(WX6572) ) ;
INV     gate6114  (.A(WX7469), .Z(WX6576) ) ;
INV     gate6115  (.A(WX7469), .Z(WX6580) ) ;
OR2     gate6116  (.A(WX6571), .B(WX6570), .Z(WX6573) ) ;
INV     gate6117  (.A(WX6573), .Z(WX6582) ) ;
INV     gate6118  (.A(WX6582), .Z(WX6583) ) ;
INV     gate6119  (.A(WX7468), .Z(WX6586) ) ;
INV     gate6120  (.A(WX7469), .Z(WX6590) ) ;
INV     gate6121  (.A(WX7469), .Z(WX6594) ) ;
OR2     gate6122  (.A(WX6585), .B(WX6584), .Z(WX6587) ) ;
INV     gate6123  (.A(WX6587), .Z(WX6596) ) ;
INV     gate6124  (.A(WX6596), .Z(WX6597) ) ;
INV     gate6125  (.A(WX7468), .Z(WX6600) ) ;
INV     gate6126  (.A(WX7469), .Z(WX6604) ) ;
INV     gate6127  (.A(WX7469), .Z(WX6608) ) ;
OR2     gate6128  (.A(WX6599), .B(WX6598), .Z(WX6601) ) ;
INV     gate6129  (.A(WX6601), .Z(WX6610) ) ;
INV     gate6130  (.A(WX6610), .Z(WX6611) ) ;
INV     gate6131  (.A(WX7468), .Z(WX6614) ) ;
INV     gate6132  (.A(WX7469), .Z(WX6618) ) ;
INV     gate6133  (.A(WX7469), .Z(WX6622) ) ;
OR2     gate6134  (.A(WX6613), .B(WX6612), .Z(WX6615) ) ;
INV     gate6135  (.A(WX6615), .Z(WX6624) ) ;
INV     gate6136  (.A(WX6624), .Z(WX6625) ) ;
INV     gate6137  (.A(WX7468), .Z(WX6628) ) ;
INV     gate6138  (.A(WX7469), .Z(WX6632) ) ;
INV     gate6139  (.A(WX7469), .Z(WX6636) ) ;
OR2     gate6140  (.A(WX6627), .B(WX6626), .Z(WX6629) ) ;
INV     gate6141  (.A(WX6629), .Z(WX6638) ) ;
INV     gate6142  (.A(WX6638), .Z(WX6639) ) ;
INV     gate6143  (.A(WX7468), .Z(WX6642) ) ;
INV     gate6144  (.A(WX7469), .Z(WX6646) ) ;
INV     gate6145  (.A(WX7469), .Z(WX6650) ) ;
OR2     gate6146  (.A(WX6641), .B(WX6640), .Z(WX6643) ) ;
INV     gate6147  (.A(WX6643), .Z(WX6652) ) ;
INV     gate6148  (.A(WX6652), .Z(WX6653) ) ;
INV     gate6149  (.A(WX7468), .Z(WX6656) ) ;
INV     gate6150  (.A(WX7469), .Z(WX6660) ) ;
INV     gate6151  (.A(WX7469), .Z(WX6664) ) ;
OR2     gate6152  (.A(WX6655), .B(WX6654), .Z(WX6657) ) ;
INV     gate6153  (.A(WX6657), .Z(WX6666) ) ;
INV     gate6154  (.A(WX6666), .Z(WX6667) ) ;
INV     gate6155  (.A(WX7468), .Z(WX6670) ) ;
INV     gate6156  (.A(WX7469), .Z(WX6674) ) ;
INV     gate6157  (.A(WX7469), .Z(WX6678) ) ;
OR2     gate6158  (.A(WX6669), .B(WX6668), .Z(WX6671) ) ;
INV     gate6159  (.A(WX6671), .Z(WX6680) ) ;
INV     gate6160  (.A(WX6680), .Z(WX6681) ) ;
INV     gate6161  (.A(WX7468), .Z(WX6684) ) ;
INV     gate6162  (.A(WX7469), .Z(WX6688) ) ;
INV     gate6163  (.A(WX7469), .Z(WX6692) ) ;
OR2     gate6164  (.A(WX6683), .B(WX6682), .Z(WX6685) ) ;
INV     gate6165  (.A(WX6685), .Z(WX6694) ) ;
INV     gate6166  (.A(WX6694), .Z(WX6695) ) ;
INV     gate6167  (.A(WX7468), .Z(WX6698) ) ;
INV     gate6168  (.A(WX7469), .Z(WX6702) ) ;
INV     gate6169  (.A(WX7469), .Z(WX6706) ) ;
OR2     gate6170  (.A(WX6697), .B(WX6696), .Z(WX6699) ) ;
INV     gate6171  (.A(WX6699), .Z(WX6708) ) ;
INV     gate6172  (.A(WX6708), .Z(WX6709) ) ;
INV     gate6173  (.A(WX7468), .Z(WX6712) ) ;
INV     gate6174  (.A(WX7469), .Z(WX6716) ) ;
INV     gate6175  (.A(WX7469), .Z(WX6720) ) ;
OR2     gate6176  (.A(WX6711), .B(WX6710), .Z(WX6713) ) ;
INV     gate6177  (.A(WX6713), .Z(WX6722) ) ;
INV     gate6178  (.A(WX6722), .Z(WX6723) ) ;
INV     gate6179  (.A(WX7468), .Z(WX6726) ) ;
INV     gate6180  (.A(WX7469), .Z(WX6730) ) ;
INV     gate6181  (.A(WX7469), .Z(WX6734) ) ;
OR2     gate6182  (.A(WX6725), .B(WX6724), .Z(WX6727) ) ;
INV     gate6183  (.A(WX6727), .Z(WX6736) ) ;
INV     gate6184  (.A(WX6736), .Z(WX6737) ) ;
INV     gate6185  (.A(WX7468), .Z(WX6740) ) ;
INV     gate6186  (.A(WX7469), .Z(WX6744) ) ;
INV     gate6187  (.A(WX7469), .Z(WX6748) ) ;
OR2     gate6188  (.A(WX6739), .B(WX6738), .Z(WX6741) ) ;
INV     gate6189  (.A(WX6741), .Z(WX6750) ) ;
INV     gate6190  (.A(WX6750), .Z(WX6751) ) ;
INV     gate6191  (.A(WX7468), .Z(WX6754) ) ;
INV     gate6192  (.A(WX7469), .Z(WX6758) ) ;
INV     gate6193  (.A(WX7469), .Z(WX6762) ) ;
OR2     gate6194  (.A(WX6753), .B(WX6752), .Z(WX6755) ) ;
INV     gate6195  (.A(WX6755), .Z(WX6764) ) ;
INV     gate6196  (.A(WX6764), .Z(WX6765) ) ;
INV     gate6197  (.A(WX7468), .Z(WX6768) ) ;
INV     gate6198  (.A(WX7469), .Z(WX6772) ) ;
INV     gate6199  (.A(WX7469), .Z(WX6776) ) ;
OR2     gate6200  (.A(WX6767), .B(WX6766), .Z(WX6769) ) ;
INV     gate6201  (.A(WX6769), .Z(WX6778) ) ;
INV     gate6202  (.A(WX6778), .Z(WX6779) ) ;
INV     gate6203  (.A(WX7468), .Z(WX6782) ) ;
INV     gate6204  (.A(WX7469), .Z(WX6786) ) ;
INV     gate6205  (.A(WX7469), .Z(WX6790) ) ;
OR2     gate6206  (.A(WX6781), .B(WX6780), .Z(WX6783) ) ;
INV     gate6207  (.A(WX6783), .Z(WX6792) ) ;
INV     gate6208  (.A(WX6792), .Z(WX6793) ) ;
INV     gate6209  (.A(WX7468), .Z(WX6796) ) ;
INV     gate6210  (.A(WX7469), .Z(WX6800) ) ;
INV     gate6211  (.A(WX7469), .Z(WX6804) ) ;
OR2     gate6212  (.A(WX6795), .B(WX6794), .Z(WX6797) ) ;
INV     gate6213  (.A(WX6797), .Z(WX6806) ) ;
INV     gate6214  (.A(WX6806), .Z(WX6807) ) ;
INV     gate6215  (.A(WX7468), .Z(WX6810) ) ;
INV     gate6216  (.A(WX7469), .Z(WX6814) ) ;
INV     gate6217  (.A(WX7469), .Z(WX6818) ) ;
OR2     gate6218  (.A(WX6809), .B(WX6808), .Z(WX6811) ) ;
INV     gate6219  (.A(WX6811), .Z(WX6820) ) ;
INV     gate6220  (.A(WX6820), .Z(WX6821) ) ;
INV     gate6221  (.A(WX7468), .Z(WX6824) ) ;
INV     gate6222  (.A(WX7469), .Z(WX6828) ) ;
INV     gate6223  (.A(WX7469), .Z(WX6832) ) ;
OR2     gate6224  (.A(WX6823), .B(WX6822), .Z(WX6825) ) ;
INV     gate6225  (.A(WX6825), .Z(WX6834) ) ;
INV     gate6226  (.A(WX6834), .Z(WX6835) ) ;
INV     gate6227  (.A(WX7468), .Z(WX6838) ) ;
INV     gate6228  (.A(WX7469), .Z(WX6842) ) ;
INV     gate6229  (.A(WX7469), .Z(WX6846) ) ;
OR2     gate6230  (.A(WX6837), .B(WX6836), .Z(WX6839) ) ;
INV     gate6231  (.A(WX6839), .Z(WX6848) ) ;
INV     gate6232  (.A(WX6848), .Z(WX6849) ) ;
INV     gate6233  (.A(WX7468), .Z(WX6852) ) ;
INV     gate6234  (.A(WX7469), .Z(WX6856) ) ;
INV     gate6235  (.A(WX7469), .Z(WX6860) ) ;
OR2     gate6236  (.A(WX6851), .B(WX6850), .Z(WX6853) ) ;
INV     gate6237  (.A(WX6853), .Z(WX6862) ) ;
INV     gate6238  (.A(WX6862), .Z(WX6863) ) ;
INV     gate6239  (.A(WX7468), .Z(WX6866) ) ;
INV     gate6240  (.A(WX7469), .Z(WX6870) ) ;
INV     gate6241  (.A(WX7469), .Z(WX6874) ) ;
OR2     gate6242  (.A(WX6865), .B(WX6864), .Z(WX6867) ) ;
INV     gate6243  (.A(WX6867), .Z(WX6876) ) ;
INV     gate6244  (.A(WX6876), .Z(WX6877) ) ;
INV     gate6245  (.A(WX7468), .Z(WX6880) ) ;
INV     gate6246  (.A(WX7469), .Z(WX6884) ) ;
INV     gate6247  (.A(WX7469), .Z(WX6888) ) ;
OR2     gate6248  (.A(WX6879), .B(WX6878), .Z(WX6881) ) ;
INV     gate6249  (.A(WX6881), .Z(WX6890) ) ;
INV     gate6250  (.A(WX6890), .Z(WX6891) ) ;
INV     gate6251  (.A(WX7468), .Z(WX6894) ) ;
INV     gate6252  (.A(WX7469), .Z(WX6898) ) ;
INV     gate6253  (.A(WX7469), .Z(WX6902) ) ;
OR2     gate6254  (.A(WX6893), .B(WX6892), .Z(WX6895) ) ;
INV     gate6255  (.A(WX6895), .Z(WX6904) ) ;
INV     gate6256  (.A(WX6904), .Z(WX6905) ) ;
INV     gate6257  (.A(WX7468), .Z(WX6908) ) ;
INV     gate6258  (.A(WX7469), .Z(WX6912) ) ;
INV     gate6259  (.A(WX7469), .Z(WX6916) ) ;
OR2     gate6260  (.A(WX6907), .B(WX6906), .Z(WX6909) ) ;
INV     gate6261  (.A(WX6909), .Z(WX6918) ) ;
INV     gate6262  (.A(WX6918), .Z(WX6919) ) ;
INV     gate6263  (.A(WX7468), .Z(WX6922) ) ;
INV     gate6264  (.A(WX7469), .Z(WX6926) ) ;
INV     gate6265  (.A(WX7469), .Z(WX6930) ) ;
OR2     gate6266  (.A(WX6921), .B(WX6920), .Z(WX6923) ) ;
INV     gate6267  (.A(WX6923), .Z(WX6932) ) ;
INV     gate6268  (.A(WX6932), .Z(WX6933) ) ;
INV     gate6269  (.A(WX7468), .Z(WX6936) ) ;
INV     gate6270  (.A(WX7469), .Z(WX6940) ) ;
INV     gate6271  (.A(WX7469), .Z(WX6944) ) ;
OR2     gate6272  (.A(WX6935), .B(WX6934), .Z(WX6937) ) ;
INV     gate6273  (.A(WX6937), .Z(WX6946) ) ;
INV     gate6274  (.A(WX6946), .Z(WX6947) ) ;
INV     gate6275  (.A(WX6950), .Z(WX6948) ) ;
INV     gate6276  (.A(WX7429), .Z(WX7430) ) ;
INV     gate6277  (.A(WX7430), .Z(WX7013) ) ;
INV     gate6278  (.A(WX7431), .Z(WX7432) ) ;
INV     gate6279  (.A(WX7432), .Z(WX7014) ) ;
INV     gate6280  (.A(WX7433), .Z(WX7434) ) ;
INV     gate6281  (.A(WX7434), .Z(WX7015) ) ;
INV     gate6282  (.A(WX7435), .Z(WX7436) ) ;
INV     gate6283  (.A(WX7436), .Z(WX7016) ) ;
INV     gate6284  (.A(WX7437), .Z(WX7438) ) ;
INV     gate6285  (.A(WX7438), .Z(WX7017) ) ;
INV     gate6286  (.A(WX7439), .Z(WX7440) ) ;
INV     gate6287  (.A(WX7440), .Z(WX7018) ) ;
INV     gate6288  (.A(WX7441), .Z(WX7442) ) ;
INV     gate6289  (.A(WX7442), .Z(WX7019) ) ;
INV     gate6290  (.A(WX7443), .Z(WX7444) ) ;
INV     gate6291  (.A(WX7444), .Z(WX7020) ) ;
INV     gate6292  (.A(WX7445), .Z(WX7446) ) ;
INV     gate6293  (.A(WX7446), .Z(WX7021) ) ;
INV     gate6294  (.A(WX7447), .Z(WX7448) ) ;
INV     gate6295  (.A(WX7448), .Z(WX7022) ) ;
INV     gate6296  (.A(WX7449), .Z(WX7450) ) ;
INV     gate6297  (.A(WX7450), .Z(WX7023) ) ;
INV     gate6298  (.A(WX7451), .Z(WX7452) ) ;
INV     gate6299  (.A(WX7452), .Z(WX7024) ) ;
INV     gate6300  (.A(WX7453), .Z(WX7454) ) ;
INV     gate6301  (.A(WX7454), .Z(WX7025) ) ;
INV     gate6302  (.A(WX7455), .Z(WX7456) ) ;
INV     gate6303  (.A(WX7456), .Z(WX7026) ) ;
INV     gate6304  (.A(WX7457), .Z(WX7458) ) ;
INV     gate6305  (.A(WX7458), .Z(WX7027) ) ;
INV     gate6306  (.A(WX7459), .Z(WX7460) ) ;
INV     gate6307  (.A(WX7460), .Z(WX7028) ) ;
INV     gate6308  (.A(WX7397), .Z(WX7398) ) ;
INV     gate6309  (.A(WX7398), .Z(WX7029) ) ;
INV     gate6310  (.A(WX7399), .Z(WX7400) ) ;
INV     gate6311  (.A(WX7400), .Z(WX7030) ) ;
INV     gate6312  (.A(WX7401), .Z(WX7402) ) ;
INV     gate6313  (.A(WX7402), .Z(WX7031) ) ;
INV     gate6314  (.A(WX7403), .Z(WX7404) ) ;
INV     gate6315  (.A(WX7404), .Z(WX7032) ) ;
INV     gate6316  (.A(WX7405), .Z(WX7406) ) ;
INV     gate6317  (.A(WX7406), .Z(WX7033) ) ;
INV     gate6318  (.A(WX7407), .Z(WX7408) ) ;
INV     gate6319  (.A(WX7408), .Z(WX7034) ) ;
INV     gate6320  (.A(WX7409), .Z(WX7410) ) ;
INV     gate6321  (.A(WX7410), .Z(WX7035) ) ;
INV     gate6322  (.A(WX7411), .Z(WX7412) ) ;
INV     gate6323  (.A(WX7412), .Z(WX7036) ) ;
INV     gate6324  (.A(WX7413), .Z(WX7414) ) ;
INV     gate6325  (.A(WX7414), .Z(WX7037) ) ;
INV     gate6326  (.A(WX7415), .Z(WX7416) ) ;
INV     gate6327  (.A(WX7416), .Z(WX7038) ) ;
INV     gate6328  (.A(WX7417), .Z(WX7418) ) ;
INV     gate6329  (.A(WX7418), .Z(WX7039) ) ;
INV     gate6330  (.A(WX7419), .Z(WX7420) ) ;
INV     gate6331  (.A(WX7420), .Z(WX7040) ) ;
INV     gate6332  (.A(WX7421), .Z(WX7422) ) ;
INV     gate6333  (.A(WX7422), .Z(WX7041) ) ;
INV     gate6334  (.A(WX7423), .Z(WX7424) ) ;
INV     gate6335  (.A(WX7424), .Z(WX7042) ) ;
INV     gate6336  (.A(WX7425), .Z(WX7426) ) ;
INV     gate6337  (.A(WX7426), .Z(WX7043) ) ;
INV     gate6338  (.A(WX7427), .Z(WX7428) ) ;
INV     gate6339  (.A(WX7428), .Z(WX7044) ) ;
INV     gate6340  (.A(WX7013), .Z(WX7045) ) ;
INV     gate6341  (.A(WX7014), .Z(WX7046) ) ;
INV     gate6342  (.A(WX7015), .Z(WX7047) ) ;
INV     gate6343  (.A(WX7016), .Z(WX7048) ) ;
INV     gate6344  (.A(WX7017), .Z(WX7049) ) ;
INV     gate6345  (.A(WX7018), .Z(WX7050) ) ;
INV     gate6346  (.A(WX7019), .Z(WX7051) ) ;
INV     gate6347  (.A(WX7020), .Z(WX7052) ) ;
INV     gate6348  (.A(WX7021), .Z(WX7053) ) ;
INV     gate6349  (.A(WX7022), .Z(WX7054) ) ;
INV     gate6350  (.A(WX7023), .Z(WX7055) ) ;
INV     gate6351  (.A(WX7024), .Z(WX7056) ) ;
INV     gate6352  (.A(WX7025), .Z(WX7057) ) ;
INV     gate6353  (.A(WX7026), .Z(WX7058) ) ;
INV     gate6354  (.A(WX7027), .Z(WX7059) ) ;
INV     gate6355  (.A(WX7028), .Z(WX7060) ) ;
INV     gate6356  (.A(WX7029), .Z(WX7061) ) ;
INV     gate6357  (.A(WX7030), .Z(WX7062) ) ;
INV     gate6358  (.A(WX7031), .Z(WX7063) ) ;
INV     gate6359  (.A(WX7032), .Z(WX7064) ) ;
INV     gate6360  (.A(WX7033), .Z(WX7065) ) ;
INV     gate6361  (.A(WX7034), .Z(WX7066) ) ;
INV     gate6362  (.A(WX7035), .Z(WX7067) ) ;
INV     gate6363  (.A(WX7036), .Z(WX7068) ) ;
INV     gate6364  (.A(WX7037), .Z(WX7069) ) ;
INV     gate6365  (.A(WX7038), .Z(WX7070) ) ;
INV     gate6366  (.A(WX7039), .Z(WX7071) ) ;
INV     gate6367  (.A(WX7040), .Z(WX7072) ) ;
INV     gate6368  (.A(WX7041), .Z(WX7073) ) ;
INV     gate6369  (.A(WX7042), .Z(WX7074) ) ;
INV     gate6370  (.A(WX7043), .Z(WX7075) ) ;
INV     gate6371  (.A(WX7044), .Z(WX7076) ) ;
INV     gate6372  (.A(WX7302), .Z(WX7077) ) ;
INV     gate6373  (.A(WX7304), .Z(WX7078) ) ;
INV     gate6374  (.A(WX7306), .Z(WX7079) ) ;
INV     gate6375  (.A(WX7308), .Z(WX7080) ) ;
INV     gate6376  (.A(WX7310), .Z(WX7081) ) ;
INV     gate6377  (.A(WX7312), .Z(WX7082) ) ;
INV     gate6378  (.A(WX7314), .Z(WX7083) ) ;
INV     gate6379  (.A(WX7316), .Z(WX7084) ) ;
INV     gate6380  (.A(WX7318), .Z(WX7085) ) ;
INV     gate6381  (.A(WX7320), .Z(WX7086) ) ;
INV     gate6382  (.A(WX7322), .Z(WX7087) ) ;
INV     gate6383  (.A(WX7324), .Z(WX7088) ) ;
INV     gate6384  (.A(WX7326), .Z(WX7089) ) ;
INV     gate6385  (.A(WX7328), .Z(WX7090) ) ;
INV     gate6386  (.A(WX7330), .Z(WX7091) ) ;
INV     gate6387  (.A(WX7332), .Z(WX7092) ) ;
INV     gate6388  (.A(WX7334), .Z(WX7093) ) ;
INV     gate6389  (.A(WX7336), .Z(WX7094) ) ;
INV     gate6390  (.A(WX7338), .Z(WX7095) ) ;
INV     gate6391  (.A(WX7340), .Z(WX7096) ) ;
INV     gate6392  (.A(WX7342), .Z(WX7097) ) ;
INV     gate6393  (.A(WX7344), .Z(WX7098) ) ;
INV     gate6394  (.A(WX7346), .Z(WX7099) ) ;
INV     gate6395  (.A(WX7348), .Z(WX7100) ) ;
INV     gate6396  (.A(WX7350), .Z(WX7101) ) ;
INV     gate6397  (.A(WX7352), .Z(WX7102) ) ;
INV     gate6398  (.A(WX7354), .Z(WX7103) ) ;
INV     gate6399  (.A(WX7356), .Z(WX7104) ) ;
INV     gate6400  (.A(WX7358), .Z(WX7105) ) ;
INV     gate6401  (.A(WX7360), .Z(WX7106) ) ;
INV     gate6402  (.A(WX7362), .Z(WX7107) ) ;
INV     gate6403  (.A(WX7364), .Z(WX7108) ) ;
NAND2   gate6404  (.A(II22532), .B(II22533), .Z(WX7381) ) ;
INV     gate6405  (.A(WX7381), .Z(WX7397) ) ;
NAND2   gate6406  (.A(II22563), .B(II22564), .Z(WX7382) ) ;
INV     gate6407  (.A(WX7382), .Z(WX7399) ) ;
NAND2   gate6408  (.A(II22594), .B(II22595), .Z(WX7383) ) ;
INV     gate6409  (.A(WX7383), .Z(WX7401) ) ;
NAND2   gate6410  (.A(II22625), .B(II22626), .Z(WX7384) ) ;
INV     gate6411  (.A(WX7384), .Z(WX7403) ) ;
NAND2   gate6412  (.A(II22656), .B(II22657), .Z(WX7385) ) ;
INV     gate6413  (.A(WX7385), .Z(WX7405) ) ;
NAND2   gate6414  (.A(II22687), .B(II22688), .Z(WX7386) ) ;
INV     gate6415  (.A(WX7386), .Z(WX7407) ) ;
NAND2   gate6416  (.A(II22718), .B(II22719), .Z(WX7387) ) ;
INV     gate6417  (.A(WX7387), .Z(WX7409) ) ;
NAND2   gate6418  (.A(II22749), .B(II22750), .Z(WX7388) ) ;
INV     gate6419  (.A(WX7388), .Z(WX7411) ) ;
NAND2   gate6420  (.A(II22780), .B(II22781), .Z(WX7389) ) ;
INV     gate6421  (.A(WX7389), .Z(WX7413) ) ;
NAND2   gate6422  (.A(II22811), .B(II22812), .Z(WX7390) ) ;
INV     gate6423  (.A(WX7390), .Z(WX7415) ) ;
NAND2   gate6424  (.A(II22842), .B(II22843), .Z(WX7391) ) ;
INV     gate6425  (.A(WX7391), .Z(WX7417) ) ;
NAND2   gate6426  (.A(II22873), .B(II22874), .Z(WX7392) ) ;
INV     gate6427  (.A(WX7392), .Z(WX7419) ) ;
NAND2   gate6428  (.A(II22904), .B(II22905), .Z(WX7393) ) ;
INV     gate6429  (.A(WX7393), .Z(WX7421) ) ;
NAND2   gate6430  (.A(II22935), .B(II22936), .Z(WX7394) ) ;
INV     gate6431  (.A(WX7394), .Z(WX7423) ) ;
NAND2   gate6432  (.A(II22966), .B(II22967), .Z(WX7395) ) ;
INV     gate6433  (.A(WX7395), .Z(WX7425) ) ;
NAND2   gate6434  (.A(II22997), .B(II22998), .Z(WX7396) ) ;
INV     gate6435  (.A(WX7396), .Z(WX7427) ) ;
NAND2   gate6436  (.A(II22036), .B(II22037), .Z(WX7365) ) ;
INV     gate6437  (.A(WX7365), .Z(WX7429) ) ;
NAND2   gate6438  (.A(II22067), .B(II22068), .Z(WX7366) ) ;
INV     gate6439  (.A(WX7366), .Z(WX7431) ) ;
NAND2   gate6440  (.A(II22098), .B(II22099), .Z(WX7367) ) ;
INV     gate6441  (.A(WX7367), .Z(WX7433) ) ;
NAND2   gate6442  (.A(II22129), .B(II22130), .Z(WX7368) ) ;
INV     gate6443  (.A(WX7368), .Z(WX7435) ) ;
NAND2   gate6444  (.A(II22160), .B(II22161), .Z(WX7369) ) ;
INV     gate6445  (.A(WX7369), .Z(WX7437) ) ;
NAND2   gate6446  (.A(II22191), .B(II22192), .Z(WX7370) ) ;
INV     gate6447  (.A(WX7370), .Z(WX7439) ) ;
NAND2   gate6448  (.A(II22222), .B(II22223), .Z(WX7371) ) ;
INV     gate6449  (.A(WX7371), .Z(WX7441) ) ;
NAND2   gate6450  (.A(II22253), .B(II22254), .Z(WX7372) ) ;
INV     gate6451  (.A(WX7372), .Z(WX7443) ) ;
NAND2   gate6452  (.A(II22284), .B(II22285), .Z(WX7373) ) ;
INV     gate6453  (.A(WX7373), .Z(WX7445) ) ;
NAND2   gate6454  (.A(II22315), .B(II22316), .Z(WX7374) ) ;
INV     gate6455  (.A(WX7374), .Z(WX7447) ) ;
NAND2   gate6456  (.A(II22346), .B(II22347), .Z(WX7375) ) ;
INV     gate6457  (.A(WX7375), .Z(WX7449) ) ;
NAND2   gate6458  (.A(II22377), .B(II22378), .Z(WX7376) ) ;
INV     gate6459  (.A(WX7376), .Z(WX7451) ) ;
NAND2   gate6460  (.A(II22408), .B(II22409), .Z(WX7377) ) ;
INV     gate6461  (.A(WX7377), .Z(WX7453) ) ;
NAND2   gate6462  (.A(II22439), .B(II22440), .Z(WX7378) ) ;
INV     gate6463  (.A(WX7378), .Z(WX7455) ) ;
NAND2   gate6464  (.A(II22470), .B(II22471), .Z(WX7379) ) ;
INV     gate6465  (.A(WX7379), .Z(WX7457) ) ;
NAND2   gate6466  (.A(II22501), .B(II22502), .Z(WX7380) ) ;
INV     gate6467  (.A(WX7380), .Z(WX7459) ) ;
INV     gate6468  (.A(TM0), .Z(WX7461) ) ;
INV     gate6469  (.A(TM0), .Z(WX7462) ) ;
INV     gate6470  (.A(TM0), .Z(WX7463) ) ;
INV     gate6471  (.A(TM1), .Z(WX7464) ) ;
INV     gate6472  (.A(TM1), .Z(WX7465) ) ;
INV     gate6473  (.A(WX7465), .Z(WX7466) ) ;
INV     gate6474  (.A(WX7463), .Z(WX7467) ) ;
INV     gate6475  (.A(WX7461), .Z(WX7470) ) ;
INV     gate6476  (.A(WX7470), .Z(WX7474) ) ;
OR2     gate6477  (.A(WX7473), .B(WX7472), .Z(WX7475) ) ;
INV     gate6478  (.A(WX7475), .Z(WX7476) ) ;
INV     gate6479  (.A(WX7476), .Z(WX7477) ) ;
INV     gate6480  (.A(WX7470), .Z(WX7481) ) ;
OR2     gate6481  (.A(WX7480), .B(WX7479), .Z(WX7482) ) ;
INV     gate6482  (.A(WX7482), .Z(WX7483) ) ;
INV     gate6483  (.A(WX7483), .Z(WX7484) ) ;
INV     gate6484  (.A(WX7470), .Z(WX7488) ) ;
OR2     gate6485  (.A(WX7487), .B(WX7486), .Z(WX7489) ) ;
INV     gate6486  (.A(WX7489), .Z(WX7490) ) ;
INV     gate6487  (.A(WX7490), .Z(WX7491) ) ;
INV     gate6488  (.A(WX7470), .Z(WX7495) ) ;
OR2     gate6489  (.A(WX7494), .B(WX7493), .Z(WX7496) ) ;
INV     gate6490  (.A(WX7496), .Z(WX7497) ) ;
INV     gate6491  (.A(WX7497), .Z(WX7498) ) ;
INV     gate6492  (.A(WX7470), .Z(WX7502) ) ;
OR2     gate6493  (.A(WX7501), .B(WX7500), .Z(WX7503) ) ;
INV     gate6494  (.A(WX7503), .Z(WX7504) ) ;
INV     gate6495  (.A(WX7504), .Z(WX7505) ) ;
INV     gate6496  (.A(WX7470), .Z(WX7509) ) ;
OR2     gate6497  (.A(WX7508), .B(WX7507), .Z(WX7510) ) ;
INV     gate6498  (.A(WX7510), .Z(WX7511) ) ;
INV     gate6499  (.A(WX7511), .Z(WX7512) ) ;
INV     gate6500  (.A(WX7470), .Z(WX7516) ) ;
OR2     gate6501  (.A(WX7515), .B(WX7514), .Z(WX7517) ) ;
INV     gate6502  (.A(WX7517), .Z(WX7518) ) ;
INV     gate6503  (.A(WX7518), .Z(WX7519) ) ;
INV     gate6504  (.A(WX7470), .Z(WX7523) ) ;
OR2     gate6505  (.A(WX7522), .B(WX7521), .Z(WX7524) ) ;
INV     gate6506  (.A(WX7524), .Z(WX7525) ) ;
INV     gate6507  (.A(WX7525), .Z(WX7526) ) ;
INV     gate6508  (.A(WX7470), .Z(WX7530) ) ;
OR2     gate6509  (.A(WX7529), .B(WX7528), .Z(WX7531) ) ;
INV     gate6510  (.A(WX7531), .Z(WX7532) ) ;
INV     gate6511  (.A(WX7532), .Z(WX7533) ) ;
INV     gate6512  (.A(WX7470), .Z(WX7537) ) ;
OR2     gate6513  (.A(WX7536), .B(WX7535), .Z(WX7538) ) ;
INV     gate6514  (.A(WX7538), .Z(WX7539) ) ;
INV     gate6515  (.A(WX7539), .Z(WX7540) ) ;
INV     gate6516  (.A(WX7470), .Z(WX7544) ) ;
OR2     gate6517  (.A(WX7543), .B(WX7542), .Z(WX7545) ) ;
INV     gate6518  (.A(WX7545), .Z(WX7546) ) ;
INV     gate6519  (.A(WX7546), .Z(WX7547) ) ;
INV     gate6520  (.A(WX7470), .Z(WX7551) ) ;
OR2     gate6521  (.A(WX7550), .B(WX7549), .Z(WX7552) ) ;
INV     gate6522  (.A(WX7552), .Z(WX7553) ) ;
INV     gate6523  (.A(WX7553), .Z(WX7554) ) ;
INV     gate6524  (.A(WX7470), .Z(WX7558) ) ;
OR2     gate6525  (.A(WX7557), .B(WX7556), .Z(WX7559) ) ;
INV     gate6526  (.A(WX7559), .Z(WX7560) ) ;
INV     gate6527  (.A(WX7560), .Z(WX7561) ) ;
INV     gate6528  (.A(WX7470), .Z(WX7565) ) ;
OR2     gate6529  (.A(WX7564), .B(WX7563), .Z(WX7566) ) ;
INV     gate6530  (.A(WX7566), .Z(WX7567) ) ;
INV     gate6531  (.A(WX7567), .Z(WX7568) ) ;
INV     gate6532  (.A(WX7470), .Z(WX7572) ) ;
OR2     gate6533  (.A(WX7571), .B(WX7570), .Z(WX7573) ) ;
INV     gate6534  (.A(WX7573), .Z(WX7574) ) ;
INV     gate6535  (.A(WX7574), .Z(WX7575) ) ;
INV     gate6536  (.A(WX7470), .Z(WX7579) ) ;
OR2     gate6537  (.A(WX7578), .B(WX7577), .Z(WX7580) ) ;
INV     gate6538  (.A(WX7580), .Z(WX7581) ) ;
INV     gate6539  (.A(WX7581), .Z(WX7582) ) ;
INV     gate6540  (.A(WX7470), .Z(WX7586) ) ;
OR2     gate6541  (.A(WX7585), .B(WX7584), .Z(WX7587) ) ;
INV     gate6542  (.A(WX7587), .Z(WX7588) ) ;
INV     gate6543  (.A(WX7588), .Z(WX7589) ) ;
INV     gate6544  (.A(WX7470), .Z(WX7593) ) ;
OR2     gate6545  (.A(WX7592), .B(WX7591), .Z(WX7594) ) ;
INV     gate6546  (.A(WX7594), .Z(WX7595) ) ;
INV     gate6547  (.A(WX7595), .Z(WX7596) ) ;
INV     gate6548  (.A(WX7470), .Z(WX7600) ) ;
OR2     gate6549  (.A(WX7599), .B(WX7598), .Z(WX7601) ) ;
INV     gate6550  (.A(WX7601), .Z(WX7602) ) ;
INV     gate6551  (.A(WX7602), .Z(WX7603) ) ;
INV     gate6552  (.A(WX7470), .Z(WX7607) ) ;
OR2     gate6553  (.A(WX7606), .B(WX7605), .Z(WX7608) ) ;
INV     gate6554  (.A(WX7608), .Z(WX7609) ) ;
INV     gate6555  (.A(WX7609), .Z(WX7610) ) ;
INV     gate6556  (.A(WX7470), .Z(WX7614) ) ;
OR2     gate6557  (.A(WX7613), .B(WX7612), .Z(WX7615) ) ;
INV     gate6558  (.A(WX7615), .Z(WX7616) ) ;
INV     gate6559  (.A(WX7616), .Z(WX7617) ) ;
INV     gate6560  (.A(WX7470), .Z(WX7621) ) ;
OR2     gate6561  (.A(WX7620), .B(WX7619), .Z(WX7622) ) ;
INV     gate6562  (.A(WX7622), .Z(WX7623) ) ;
INV     gate6563  (.A(WX7623), .Z(WX7624) ) ;
INV     gate6564  (.A(WX7470), .Z(WX7628) ) ;
OR2     gate6565  (.A(WX7627), .B(WX7626), .Z(WX7629) ) ;
INV     gate6566  (.A(WX7629), .Z(WX7630) ) ;
INV     gate6567  (.A(WX7630), .Z(WX7631) ) ;
INV     gate6568  (.A(WX7470), .Z(WX7635) ) ;
OR2     gate6569  (.A(WX7634), .B(WX7633), .Z(WX7636) ) ;
INV     gate6570  (.A(WX7636), .Z(WX7637) ) ;
INV     gate6571  (.A(WX7637), .Z(WX7638) ) ;
INV     gate6572  (.A(WX7470), .Z(WX7642) ) ;
OR2     gate6573  (.A(WX7641), .B(WX7640), .Z(WX7643) ) ;
INV     gate6574  (.A(WX7643), .Z(WX7644) ) ;
INV     gate6575  (.A(WX7644), .Z(WX7645) ) ;
INV     gate6576  (.A(WX7470), .Z(WX7649) ) ;
OR2     gate6577  (.A(WX7648), .B(WX7647), .Z(WX7650) ) ;
INV     gate6578  (.A(WX7650), .Z(WX7651) ) ;
INV     gate6579  (.A(WX7651), .Z(WX7652) ) ;
INV     gate6580  (.A(WX7470), .Z(WX7656) ) ;
OR2     gate6581  (.A(WX7655), .B(WX7654), .Z(WX7657) ) ;
INV     gate6582  (.A(WX7657), .Z(WX7658) ) ;
INV     gate6583  (.A(WX7658), .Z(WX7659) ) ;
INV     gate6584  (.A(WX7470), .Z(WX7663) ) ;
OR2     gate6585  (.A(WX7662), .B(WX7661), .Z(WX7664) ) ;
INV     gate6586  (.A(WX7664), .Z(WX7665) ) ;
INV     gate6587  (.A(WX7665), .Z(WX7666) ) ;
INV     gate6588  (.A(WX7470), .Z(WX7670) ) ;
OR2     gate6589  (.A(WX7669), .B(WX7668), .Z(WX7671) ) ;
INV     gate6590  (.A(WX7671), .Z(WX7672) ) ;
INV     gate6591  (.A(WX7672), .Z(WX7673) ) ;
INV     gate6592  (.A(WX7470), .Z(WX7677) ) ;
OR2     gate6593  (.A(WX7676), .B(WX7675), .Z(WX7678) ) ;
INV     gate6594  (.A(WX7678), .Z(WX7679) ) ;
INV     gate6595  (.A(WX7679), .Z(WX7680) ) ;
INV     gate6596  (.A(WX7470), .Z(WX7684) ) ;
OR2     gate6597  (.A(WX7683), .B(WX7682), .Z(WX7685) ) ;
INV     gate6598  (.A(WX7685), .Z(WX7686) ) ;
INV     gate6599  (.A(WX7686), .Z(WX7687) ) ;
INV     gate6600  (.A(WX7470), .Z(WX7691) ) ;
OR2     gate6601  (.A(WX7690), .B(WX7689), .Z(WX7692) ) ;
INV     gate6602  (.A(WX7692), .Z(WX7693) ) ;
INV     gate6603  (.A(WX7693), .Z(WX7694) ) ;
INV     gate6604  (.A(RESET), .Z(WX7695) ) ;
INV     gate6605  (.A(WX7695), .Z(WX7728) ) ;
INV     gate6606  (.A(WX8757), .Z(WX8761) ) ;
INV     gate6607  (.A(WX8761), .Z(WX7795) ) ;
INV     gate6608  (.A(WX8755), .Z(WX8762) ) ;
INV     gate6609  (.A(WX8762), .Z(WX7799) ) ;
INV     gate6610  (.A(WX8762), .Z(WX7803) ) ;
OR2     gate6611  (.A(WX7794), .B(WX7793), .Z(WX7796) ) ;
INV     gate6612  (.A(WX7796), .Z(WX7805) ) ;
INV     gate6613  (.A(WX7805), .Z(WX7806) ) ;
INV     gate6614  (.A(WX8761), .Z(WX7809) ) ;
INV     gate6615  (.A(WX8762), .Z(WX7813) ) ;
INV     gate6616  (.A(WX8762), .Z(WX7817) ) ;
OR2     gate6617  (.A(WX7808), .B(WX7807), .Z(WX7810) ) ;
INV     gate6618  (.A(WX7810), .Z(WX7819) ) ;
INV     gate6619  (.A(WX7819), .Z(WX7820) ) ;
INV     gate6620  (.A(WX8761), .Z(WX7823) ) ;
INV     gate6621  (.A(WX8762), .Z(WX7827) ) ;
INV     gate6622  (.A(WX8762), .Z(WX7831) ) ;
OR2     gate6623  (.A(WX7822), .B(WX7821), .Z(WX7824) ) ;
INV     gate6624  (.A(WX7824), .Z(WX7833) ) ;
INV     gate6625  (.A(WX7833), .Z(WX7834) ) ;
INV     gate6626  (.A(WX8761), .Z(WX7837) ) ;
INV     gate6627  (.A(WX8762), .Z(WX7841) ) ;
INV     gate6628  (.A(WX8762), .Z(WX7845) ) ;
OR2     gate6629  (.A(WX7836), .B(WX7835), .Z(WX7838) ) ;
INV     gate6630  (.A(WX7838), .Z(WX7847) ) ;
INV     gate6631  (.A(WX7847), .Z(WX7848) ) ;
INV     gate6632  (.A(WX8761), .Z(WX7851) ) ;
INV     gate6633  (.A(WX8762), .Z(WX7855) ) ;
INV     gate6634  (.A(WX8762), .Z(WX7859) ) ;
OR2     gate6635  (.A(WX7850), .B(WX7849), .Z(WX7852) ) ;
INV     gate6636  (.A(WX7852), .Z(WX7861) ) ;
INV     gate6637  (.A(WX7861), .Z(WX7862) ) ;
INV     gate6638  (.A(WX8761), .Z(WX7865) ) ;
INV     gate6639  (.A(WX8762), .Z(WX7869) ) ;
INV     gate6640  (.A(WX8762), .Z(WX7873) ) ;
OR2     gate6641  (.A(WX7864), .B(WX7863), .Z(WX7866) ) ;
INV     gate6642  (.A(WX7866), .Z(WX7875) ) ;
INV     gate6643  (.A(WX7875), .Z(WX7876) ) ;
INV     gate6644  (.A(WX8761), .Z(WX7879) ) ;
INV     gate6645  (.A(WX8762), .Z(WX7883) ) ;
INV     gate6646  (.A(WX8762), .Z(WX7887) ) ;
OR2     gate6647  (.A(WX7878), .B(WX7877), .Z(WX7880) ) ;
INV     gate6648  (.A(WX7880), .Z(WX7889) ) ;
INV     gate6649  (.A(WX7889), .Z(WX7890) ) ;
INV     gate6650  (.A(WX8761), .Z(WX7893) ) ;
INV     gate6651  (.A(WX8762), .Z(WX7897) ) ;
INV     gate6652  (.A(WX8762), .Z(WX7901) ) ;
OR2     gate6653  (.A(WX7892), .B(WX7891), .Z(WX7894) ) ;
INV     gate6654  (.A(WX7894), .Z(WX7903) ) ;
INV     gate6655  (.A(WX7903), .Z(WX7904) ) ;
INV     gate6656  (.A(WX8761), .Z(WX7907) ) ;
INV     gate6657  (.A(WX8762), .Z(WX7911) ) ;
INV     gate6658  (.A(WX8762), .Z(WX7915) ) ;
OR2     gate6659  (.A(WX7906), .B(WX7905), .Z(WX7908) ) ;
INV     gate6660  (.A(WX7908), .Z(WX7917) ) ;
INV     gate6661  (.A(WX7917), .Z(WX7918) ) ;
INV     gate6662  (.A(WX8761), .Z(WX7921) ) ;
INV     gate6663  (.A(WX8762), .Z(WX7925) ) ;
INV     gate6664  (.A(WX8762), .Z(WX7929) ) ;
OR2     gate6665  (.A(WX7920), .B(WX7919), .Z(WX7922) ) ;
INV     gate6666  (.A(WX7922), .Z(WX7931) ) ;
INV     gate6667  (.A(WX7931), .Z(WX7932) ) ;
INV     gate6668  (.A(WX8761), .Z(WX7935) ) ;
INV     gate6669  (.A(WX8762), .Z(WX7939) ) ;
INV     gate6670  (.A(WX8762), .Z(WX7943) ) ;
OR2     gate6671  (.A(WX7934), .B(WX7933), .Z(WX7936) ) ;
INV     gate6672  (.A(WX7936), .Z(WX7945) ) ;
INV     gate6673  (.A(WX7945), .Z(WX7946) ) ;
INV     gate6674  (.A(WX8761), .Z(WX7949) ) ;
INV     gate6675  (.A(WX8762), .Z(WX7953) ) ;
INV     gate6676  (.A(WX8762), .Z(WX7957) ) ;
OR2     gate6677  (.A(WX7948), .B(WX7947), .Z(WX7950) ) ;
INV     gate6678  (.A(WX7950), .Z(WX7959) ) ;
INV     gate6679  (.A(WX7959), .Z(WX7960) ) ;
INV     gate6680  (.A(WX8761), .Z(WX7963) ) ;
INV     gate6681  (.A(WX8762), .Z(WX7967) ) ;
INV     gate6682  (.A(WX8762), .Z(WX7971) ) ;
OR2     gate6683  (.A(WX7962), .B(WX7961), .Z(WX7964) ) ;
INV     gate6684  (.A(WX7964), .Z(WX7973) ) ;
INV     gate6685  (.A(WX7973), .Z(WX7974) ) ;
INV     gate6686  (.A(WX8761), .Z(WX7977) ) ;
INV     gate6687  (.A(WX8762), .Z(WX7981) ) ;
INV     gate6688  (.A(WX8762), .Z(WX7985) ) ;
OR2     gate6689  (.A(WX7976), .B(WX7975), .Z(WX7978) ) ;
INV     gate6690  (.A(WX7978), .Z(WX7987) ) ;
INV     gate6691  (.A(WX7987), .Z(WX7988) ) ;
INV     gate6692  (.A(WX8761), .Z(WX7991) ) ;
INV     gate6693  (.A(WX8762), .Z(WX7995) ) ;
INV     gate6694  (.A(WX8762), .Z(WX7999) ) ;
OR2     gate6695  (.A(WX7990), .B(WX7989), .Z(WX7992) ) ;
INV     gate6696  (.A(WX7992), .Z(WX8001) ) ;
INV     gate6697  (.A(WX8001), .Z(WX8002) ) ;
INV     gate6698  (.A(WX8761), .Z(WX8005) ) ;
INV     gate6699  (.A(WX8762), .Z(WX8009) ) ;
INV     gate6700  (.A(WX8762), .Z(WX8013) ) ;
OR2     gate6701  (.A(WX8004), .B(WX8003), .Z(WX8006) ) ;
INV     gate6702  (.A(WX8006), .Z(WX8015) ) ;
INV     gate6703  (.A(WX8015), .Z(WX8016) ) ;
INV     gate6704  (.A(WX8761), .Z(WX8019) ) ;
INV     gate6705  (.A(WX8762), .Z(WX8023) ) ;
INV     gate6706  (.A(WX8762), .Z(WX8027) ) ;
OR2     gate6707  (.A(WX8018), .B(WX8017), .Z(WX8020) ) ;
INV     gate6708  (.A(WX8020), .Z(WX8029) ) ;
INV     gate6709  (.A(WX8029), .Z(WX8030) ) ;
INV     gate6710  (.A(WX8761), .Z(WX8033) ) ;
INV     gate6711  (.A(WX8762), .Z(WX8037) ) ;
INV     gate6712  (.A(WX8762), .Z(WX8041) ) ;
OR2     gate6713  (.A(WX8032), .B(WX8031), .Z(WX8034) ) ;
INV     gate6714  (.A(WX8034), .Z(WX8043) ) ;
INV     gate6715  (.A(WX8043), .Z(WX8044) ) ;
INV     gate6716  (.A(WX8761), .Z(WX8047) ) ;
INV     gate6717  (.A(WX8762), .Z(WX8051) ) ;
INV     gate6718  (.A(WX8762), .Z(WX8055) ) ;
OR2     gate6719  (.A(WX8046), .B(WX8045), .Z(WX8048) ) ;
INV     gate6720  (.A(WX8048), .Z(WX8057) ) ;
INV     gate6721  (.A(WX8057), .Z(WX8058) ) ;
INV     gate6722  (.A(WX8761), .Z(WX8061) ) ;
INV     gate6723  (.A(WX8762), .Z(WX8065) ) ;
INV     gate6724  (.A(WX8762), .Z(WX8069) ) ;
OR2     gate6725  (.A(WX8060), .B(WX8059), .Z(WX8062) ) ;
INV     gate6726  (.A(WX8062), .Z(WX8071) ) ;
INV     gate6727  (.A(WX8071), .Z(WX8072) ) ;
INV     gate6728  (.A(WX8761), .Z(WX8075) ) ;
INV     gate6729  (.A(WX8762), .Z(WX8079) ) ;
INV     gate6730  (.A(WX8762), .Z(WX8083) ) ;
OR2     gate6731  (.A(WX8074), .B(WX8073), .Z(WX8076) ) ;
INV     gate6732  (.A(WX8076), .Z(WX8085) ) ;
INV     gate6733  (.A(WX8085), .Z(WX8086) ) ;
INV     gate6734  (.A(WX8761), .Z(WX8089) ) ;
INV     gate6735  (.A(WX8762), .Z(WX8093) ) ;
INV     gate6736  (.A(WX8762), .Z(WX8097) ) ;
OR2     gate6737  (.A(WX8088), .B(WX8087), .Z(WX8090) ) ;
INV     gate6738  (.A(WX8090), .Z(WX8099) ) ;
INV     gate6739  (.A(WX8099), .Z(WX8100) ) ;
INV     gate6740  (.A(WX8761), .Z(WX8103) ) ;
INV     gate6741  (.A(WX8762), .Z(WX8107) ) ;
INV     gate6742  (.A(WX8762), .Z(WX8111) ) ;
OR2     gate6743  (.A(WX8102), .B(WX8101), .Z(WX8104) ) ;
INV     gate6744  (.A(WX8104), .Z(WX8113) ) ;
INV     gate6745  (.A(WX8113), .Z(WX8114) ) ;
INV     gate6746  (.A(WX8761), .Z(WX8117) ) ;
INV     gate6747  (.A(WX8762), .Z(WX8121) ) ;
INV     gate6748  (.A(WX8762), .Z(WX8125) ) ;
OR2     gate6749  (.A(WX8116), .B(WX8115), .Z(WX8118) ) ;
INV     gate6750  (.A(WX8118), .Z(WX8127) ) ;
INV     gate6751  (.A(WX8127), .Z(WX8128) ) ;
INV     gate6752  (.A(WX8761), .Z(WX8131) ) ;
INV     gate6753  (.A(WX8762), .Z(WX8135) ) ;
INV     gate6754  (.A(WX8762), .Z(WX8139) ) ;
OR2     gate6755  (.A(WX8130), .B(WX8129), .Z(WX8132) ) ;
INV     gate6756  (.A(WX8132), .Z(WX8141) ) ;
INV     gate6757  (.A(WX8141), .Z(WX8142) ) ;
INV     gate6758  (.A(WX8761), .Z(WX8145) ) ;
INV     gate6759  (.A(WX8762), .Z(WX8149) ) ;
INV     gate6760  (.A(WX8762), .Z(WX8153) ) ;
OR2     gate6761  (.A(WX8144), .B(WX8143), .Z(WX8146) ) ;
INV     gate6762  (.A(WX8146), .Z(WX8155) ) ;
INV     gate6763  (.A(WX8155), .Z(WX8156) ) ;
INV     gate6764  (.A(WX8761), .Z(WX8159) ) ;
INV     gate6765  (.A(WX8762), .Z(WX8163) ) ;
INV     gate6766  (.A(WX8762), .Z(WX8167) ) ;
OR2     gate6767  (.A(WX8158), .B(WX8157), .Z(WX8160) ) ;
INV     gate6768  (.A(WX8160), .Z(WX8169) ) ;
INV     gate6769  (.A(WX8169), .Z(WX8170) ) ;
INV     gate6770  (.A(WX8761), .Z(WX8173) ) ;
INV     gate6771  (.A(WX8762), .Z(WX8177) ) ;
INV     gate6772  (.A(WX8762), .Z(WX8181) ) ;
OR2     gate6773  (.A(WX8172), .B(WX8171), .Z(WX8174) ) ;
INV     gate6774  (.A(WX8174), .Z(WX8183) ) ;
INV     gate6775  (.A(WX8183), .Z(WX8184) ) ;
INV     gate6776  (.A(WX8761), .Z(WX8187) ) ;
INV     gate6777  (.A(WX8762), .Z(WX8191) ) ;
INV     gate6778  (.A(WX8762), .Z(WX8195) ) ;
OR2     gate6779  (.A(WX8186), .B(WX8185), .Z(WX8188) ) ;
INV     gate6780  (.A(WX8188), .Z(WX8197) ) ;
INV     gate6781  (.A(WX8197), .Z(WX8198) ) ;
INV     gate6782  (.A(WX8761), .Z(WX8201) ) ;
INV     gate6783  (.A(WX8762), .Z(WX8205) ) ;
INV     gate6784  (.A(WX8762), .Z(WX8209) ) ;
OR2     gate6785  (.A(WX8200), .B(WX8199), .Z(WX8202) ) ;
INV     gate6786  (.A(WX8202), .Z(WX8211) ) ;
INV     gate6787  (.A(WX8211), .Z(WX8212) ) ;
INV     gate6788  (.A(WX8761), .Z(WX8215) ) ;
INV     gate6789  (.A(WX8762), .Z(WX8219) ) ;
INV     gate6790  (.A(WX8762), .Z(WX8223) ) ;
OR2     gate6791  (.A(WX8214), .B(WX8213), .Z(WX8216) ) ;
INV     gate6792  (.A(WX8216), .Z(WX8225) ) ;
INV     gate6793  (.A(WX8225), .Z(WX8226) ) ;
INV     gate6794  (.A(WX8761), .Z(WX8229) ) ;
INV     gate6795  (.A(WX8762), .Z(WX8233) ) ;
INV     gate6796  (.A(WX8762), .Z(WX8237) ) ;
OR2     gate6797  (.A(WX8228), .B(WX8227), .Z(WX8230) ) ;
INV     gate6798  (.A(WX8230), .Z(WX8239) ) ;
INV     gate6799  (.A(WX8239), .Z(WX8240) ) ;
INV     gate6800  (.A(WX8243), .Z(WX8241) ) ;
INV     gate6801  (.A(WX8722), .Z(WX8723) ) ;
INV     gate6802  (.A(WX8723), .Z(WX8306) ) ;
INV     gate6803  (.A(WX8724), .Z(WX8725) ) ;
INV     gate6804  (.A(WX8725), .Z(WX8307) ) ;
INV     gate6805  (.A(WX8726), .Z(WX8727) ) ;
INV     gate6806  (.A(WX8727), .Z(WX8308) ) ;
INV     gate6807  (.A(WX8728), .Z(WX8729) ) ;
INV     gate6808  (.A(WX8729), .Z(WX8309) ) ;
INV     gate6809  (.A(WX8730), .Z(WX8731) ) ;
INV     gate6810  (.A(WX8731), .Z(WX8310) ) ;
INV     gate6811  (.A(WX8732), .Z(WX8733) ) ;
INV     gate6812  (.A(WX8733), .Z(WX8311) ) ;
INV     gate6813  (.A(WX8734), .Z(WX8735) ) ;
INV     gate6814  (.A(WX8735), .Z(WX8312) ) ;
INV     gate6815  (.A(WX8736), .Z(WX8737) ) ;
INV     gate6816  (.A(WX8737), .Z(WX8313) ) ;
INV     gate6817  (.A(WX8738), .Z(WX8739) ) ;
INV     gate6818  (.A(WX8739), .Z(WX8314) ) ;
INV     gate6819  (.A(WX8740), .Z(WX8741) ) ;
INV     gate6820  (.A(WX8741), .Z(WX8315) ) ;
INV     gate6821  (.A(WX8742), .Z(WX8743) ) ;
INV     gate6822  (.A(WX8743), .Z(WX8316) ) ;
INV     gate6823  (.A(WX8744), .Z(WX8745) ) ;
INV     gate6824  (.A(WX8745), .Z(WX8317) ) ;
INV     gate6825  (.A(WX8746), .Z(WX8747) ) ;
INV     gate6826  (.A(WX8747), .Z(WX8318) ) ;
INV     gate6827  (.A(WX8748), .Z(WX8749) ) ;
INV     gate6828  (.A(WX8749), .Z(WX8319) ) ;
INV     gate6829  (.A(WX8750), .Z(WX8751) ) ;
INV     gate6830  (.A(WX8751), .Z(WX8320) ) ;
INV     gate6831  (.A(WX8752), .Z(WX8753) ) ;
INV     gate6832  (.A(WX8753), .Z(WX8321) ) ;
INV     gate6833  (.A(WX8690), .Z(WX8691) ) ;
INV     gate6834  (.A(WX8691), .Z(WX8322) ) ;
INV     gate6835  (.A(WX8692), .Z(WX8693) ) ;
INV     gate6836  (.A(WX8693), .Z(WX8323) ) ;
INV     gate6837  (.A(WX8694), .Z(WX8695) ) ;
INV     gate6838  (.A(WX8695), .Z(WX8324) ) ;
INV     gate6839  (.A(WX8696), .Z(WX8697) ) ;
INV     gate6840  (.A(WX8697), .Z(WX8325) ) ;
INV     gate6841  (.A(WX8698), .Z(WX8699) ) ;
INV     gate6842  (.A(WX8699), .Z(WX8326) ) ;
INV     gate6843  (.A(WX8700), .Z(WX8701) ) ;
INV     gate6844  (.A(WX8701), .Z(WX8327) ) ;
INV     gate6845  (.A(WX8702), .Z(WX8703) ) ;
INV     gate6846  (.A(WX8703), .Z(WX8328) ) ;
INV     gate6847  (.A(WX8704), .Z(WX8705) ) ;
INV     gate6848  (.A(WX8705), .Z(WX8329) ) ;
INV     gate6849  (.A(WX8706), .Z(WX8707) ) ;
INV     gate6850  (.A(WX8707), .Z(WX8330) ) ;
INV     gate6851  (.A(WX8708), .Z(WX8709) ) ;
INV     gate6852  (.A(WX8709), .Z(WX8331) ) ;
INV     gate6853  (.A(WX8710), .Z(WX8711) ) ;
INV     gate6854  (.A(WX8711), .Z(WX8332) ) ;
INV     gate6855  (.A(WX8712), .Z(WX8713) ) ;
INV     gate6856  (.A(WX8713), .Z(WX8333) ) ;
INV     gate6857  (.A(WX8714), .Z(WX8715) ) ;
INV     gate6858  (.A(WX8715), .Z(WX8334) ) ;
INV     gate6859  (.A(WX8716), .Z(WX8717) ) ;
INV     gate6860  (.A(WX8717), .Z(WX8335) ) ;
INV     gate6861  (.A(WX8718), .Z(WX8719) ) ;
INV     gate6862  (.A(WX8719), .Z(WX8336) ) ;
INV     gate6863  (.A(WX8720), .Z(WX8721) ) ;
INV     gate6864  (.A(WX8721), .Z(WX8337) ) ;
INV     gate6865  (.A(WX8306), .Z(WX8338) ) ;
INV     gate6866  (.A(WX8307), .Z(WX8339) ) ;
INV     gate6867  (.A(WX8308), .Z(WX8340) ) ;
INV     gate6868  (.A(WX8309), .Z(WX8341) ) ;
INV     gate6869  (.A(WX8310), .Z(WX8342) ) ;
INV     gate6870  (.A(WX8311), .Z(WX8343) ) ;
INV     gate6871  (.A(WX8312), .Z(WX8344) ) ;
INV     gate6872  (.A(WX8313), .Z(WX8345) ) ;
INV     gate6873  (.A(WX8314), .Z(WX8346) ) ;
INV     gate6874  (.A(WX8315), .Z(WX8347) ) ;
INV     gate6875  (.A(WX8316), .Z(WX8348) ) ;
INV     gate6876  (.A(WX8317), .Z(WX8349) ) ;
INV     gate6877  (.A(WX8318), .Z(WX8350) ) ;
INV     gate6878  (.A(WX8319), .Z(WX8351) ) ;
INV     gate6879  (.A(WX8320), .Z(WX8352) ) ;
INV     gate6880  (.A(WX8321), .Z(WX8353) ) ;
INV     gate6881  (.A(WX8322), .Z(WX8354) ) ;
INV     gate6882  (.A(WX8323), .Z(WX8355) ) ;
INV     gate6883  (.A(WX8324), .Z(WX8356) ) ;
INV     gate6884  (.A(WX8325), .Z(WX8357) ) ;
INV     gate6885  (.A(WX8326), .Z(WX8358) ) ;
INV     gate6886  (.A(WX8327), .Z(WX8359) ) ;
INV     gate6887  (.A(WX8328), .Z(WX8360) ) ;
INV     gate6888  (.A(WX8329), .Z(WX8361) ) ;
INV     gate6889  (.A(WX8330), .Z(WX8362) ) ;
INV     gate6890  (.A(WX8331), .Z(WX8363) ) ;
INV     gate6891  (.A(WX8332), .Z(WX8364) ) ;
INV     gate6892  (.A(WX8333), .Z(WX8365) ) ;
INV     gate6893  (.A(WX8334), .Z(WX8366) ) ;
INV     gate6894  (.A(WX8335), .Z(WX8367) ) ;
INV     gate6895  (.A(WX8336), .Z(WX8368) ) ;
INV     gate6896  (.A(WX8337), .Z(WX8369) ) ;
INV     gate6897  (.A(WX8595), .Z(WX8370) ) ;
INV     gate6898  (.A(WX8597), .Z(WX8371) ) ;
INV     gate6899  (.A(WX8599), .Z(WX8372) ) ;
INV     gate6900  (.A(WX8601), .Z(WX8373) ) ;
INV     gate6901  (.A(WX8603), .Z(WX8374) ) ;
INV     gate6902  (.A(WX8605), .Z(WX8375) ) ;
INV     gate6903  (.A(WX8607), .Z(WX8376) ) ;
INV     gate6904  (.A(WX8609), .Z(WX8377) ) ;
INV     gate6905  (.A(WX8611), .Z(WX8378) ) ;
INV     gate6906  (.A(WX8613), .Z(WX8379) ) ;
INV     gate6907  (.A(WX8615), .Z(WX8380) ) ;
INV     gate6908  (.A(WX8617), .Z(WX8381) ) ;
INV     gate6909  (.A(WX8619), .Z(WX8382) ) ;
INV     gate6910  (.A(WX8621), .Z(WX8383) ) ;
INV     gate6911  (.A(WX8623), .Z(WX8384) ) ;
INV     gate6912  (.A(WX8625), .Z(WX8385) ) ;
INV     gate6913  (.A(WX8627), .Z(WX8386) ) ;
INV     gate6914  (.A(WX8629), .Z(WX8387) ) ;
INV     gate6915  (.A(WX8631), .Z(WX8388) ) ;
INV     gate6916  (.A(WX8633), .Z(WX8389) ) ;
INV     gate6917  (.A(WX8635), .Z(WX8390) ) ;
INV     gate6918  (.A(WX8637), .Z(WX8391) ) ;
INV     gate6919  (.A(WX8639), .Z(WX8392) ) ;
INV     gate6920  (.A(WX8641), .Z(WX8393) ) ;
INV     gate6921  (.A(WX8643), .Z(WX8394) ) ;
INV     gate6922  (.A(WX8645), .Z(WX8395) ) ;
INV     gate6923  (.A(WX8647), .Z(WX8396) ) ;
INV     gate6924  (.A(WX8649), .Z(WX8397) ) ;
INV     gate6925  (.A(WX8651), .Z(WX8398) ) ;
INV     gate6926  (.A(WX8653), .Z(WX8399) ) ;
INV     gate6927  (.A(WX8655), .Z(WX8400) ) ;
INV     gate6928  (.A(WX8657), .Z(WX8401) ) ;
NAND2   gate6929  (.A(II26537), .B(II26538), .Z(WX8674) ) ;
INV     gate6930  (.A(WX8674), .Z(WX8690) ) ;
NAND2   gate6931  (.A(II26568), .B(II26569), .Z(WX8675) ) ;
INV     gate6932  (.A(WX8675), .Z(WX8692) ) ;
NAND2   gate6933  (.A(II26599), .B(II26600), .Z(WX8676) ) ;
INV     gate6934  (.A(WX8676), .Z(WX8694) ) ;
NAND2   gate6935  (.A(II26630), .B(II26631), .Z(WX8677) ) ;
INV     gate6936  (.A(WX8677), .Z(WX8696) ) ;
NAND2   gate6937  (.A(II26661), .B(II26662), .Z(WX8678) ) ;
INV     gate6938  (.A(WX8678), .Z(WX8698) ) ;
NAND2   gate6939  (.A(II26692), .B(II26693), .Z(WX8679) ) ;
INV     gate6940  (.A(WX8679), .Z(WX8700) ) ;
NAND2   gate6941  (.A(II26723), .B(II26724), .Z(WX8680) ) ;
INV     gate6942  (.A(WX8680), .Z(WX8702) ) ;
NAND2   gate6943  (.A(II26754), .B(II26755), .Z(WX8681) ) ;
INV     gate6944  (.A(WX8681), .Z(WX8704) ) ;
NAND2   gate6945  (.A(II26785), .B(II26786), .Z(WX8682) ) ;
INV     gate6946  (.A(WX8682), .Z(WX8706) ) ;
NAND2   gate6947  (.A(II26816), .B(II26817), .Z(WX8683) ) ;
INV     gate6948  (.A(WX8683), .Z(WX8708) ) ;
NAND2   gate6949  (.A(II26847), .B(II26848), .Z(WX8684) ) ;
INV     gate6950  (.A(WX8684), .Z(WX8710) ) ;
NAND2   gate6951  (.A(II26878), .B(II26879), .Z(WX8685) ) ;
INV     gate6952  (.A(WX8685), .Z(WX8712) ) ;
NAND2   gate6953  (.A(II26909), .B(II26910), .Z(WX8686) ) ;
INV     gate6954  (.A(WX8686), .Z(WX8714) ) ;
NAND2   gate6955  (.A(II26940), .B(II26941), .Z(WX8687) ) ;
INV     gate6956  (.A(WX8687), .Z(WX8716) ) ;
NAND2   gate6957  (.A(II26971), .B(II26972), .Z(WX8688) ) ;
INV     gate6958  (.A(WX8688), .Z(WX8718) ) ;
NAND2   gate6959  (.A(II27002), .B(II27003), .Z(WX8689) ) ;
INV     gate6960  (.A(WX8689), .Z(WX8720) ) ;
NAND2   gate6961  (.A(II26041), .B(II26042), .Z(WX8658) ) ;
INV     gate6962  (.A(WX8658), .Z(WX8722) ) ;
NAND2   gate6963  (.A(II26072), .B(II26073), .Z(WX8659) ) ;
INV     gate6964  (.A(WX8659), .Z(WX8724) ) ;
NAND2   gate6965  (.A(II26103), .B(II26104), .Z(WX8660) ) ;
INV     gate6966  (.A(WX8660), .Z(WX8726) ) ;
NAND2   gate6967  (.A(II26134), .B(II26135), .Z(WX8661) ) ;
INV     gate6968  (.A(WX8661), .Z(WX8728) ) ;
NAND2   gate6969  (.A(II26165), .B(II26166), .Z(WX8662) ) ;
INV     gate6970  (.A(WX8662), .Z(WX8730) ) ;
NAND2   gate6971  (.A(II26196), .B(II26197), .Z(WX8663) ) ;
INV     gate6972  (.A(WX8663), .Z(WX8732) ) ;
NAND2   gate6973  (.A(II26227), .B(II26228), .Z(WX8664) ) ;
INV     gate6974  (.A(WX8664), .Z(WX8734) ) ;
NAND2   gate6975  (.A(II26258), .B(II26259), .Z(WX8665) ) ;
INV     gate6976  (.A(WX8665), .Z(WX8736) ) ;
NAND2   gate6977  (.A(II26289), .B(II26290), .Z(WX8666) ) ;
INV     gate6978  (.A(WX8666), .Z(WX8738) ) ;
NAND2   gate6979  (.A(II26320), .B(II26321), .Z(WX8667) ) ;
INV     gate6980  (.A(WX8667), .Z(WX8740) ) ;
NAND2   gate6981  (.A(II26351), .B(II26352), .Z(WX8668) ) ;
INV     gate6982  (.A(WX8668), .Z(WX8742) ) ;
NAND2   gate6983  (.A(II26382), .B(II26383), .Z(WX8669) ) ;
INV     gate6984  (.A(WX8669), .Z(WX8744) ) ;
NAND2   gate6985  (.A(II26413), .B(II26414), .Z(WX8670) ) ;
INV     gate6986  (.A(WX8670), .Z(WX8746) ) ;
NAND2   gate6987  (.A(II26444), .B(II26445), .Z(WX8671) ) ;
INV     gate6988  (.A(WX8671), .Z(WX8748) ) ;
NAND2   gate6989  (.A(II26475), .B(II26476), .Z(WX8672) ) ;
INV     gate6990  (.A(WX8672), .Z(WX8750) ) ;
NAND2   gate6991  (.A(II26506), .B(II26507), .Z(WX8673) ) ;
INV     gate6992  (.A(WX8673), .Z(WX8752) ) ;
INV     gate6993  (.A(TM0), .Z(WX8754) ) ;
INV     gate6994  (.A(TM0), .Z(WX8755) ) ;
INV     gate6995  (.A(TM0), .Z(WX8756) ) ;
INV     gate6996  (.A(TM1), .Z(WX8757) ) ;
INV     gate6997  (.A(TM1), .Z(WX8758) ) ;
INV     gate6998  (.A(WX8758), .Z(WX8759) ) ;
INV     gate6999  (.A(WX8756), .Z(WX8760) ) ;
INV     gate7000  (.A(WX8754), .Z(WX8763) ) ;
INV     gate7001  (.A(WX8763), .Z(WX8767) ) ;
OR2     gate7002  (.A(WX8766), .B(WX8765), .Z(WX8768) ) ;
INV     gate7003  (.A(WX8768), .Z(WX8769) ) ;
INV     gate7004  (.A(WX8769), .Z(WX8770) ) ;
INV     gate7005  (.A(WX8763), .Z(WX8774) ) ;
OR2     gate7006  (.A(WX8773), .B(WX8772), .Z(WX8775) ) ;
INV     gate7007  (.A(WX8775), .Z(WX8776) ) ;
INV     gate7008  (.A(WX8776), .Z(WX8777) ) ;
INV     gate7009  (.A(WX8763), .Z(WX8781) ) ;
OR2     gate7010  (.A(WX8780), .B(WX8779), .Z(WX8782) ) ;
INV     gate7011  (.A(WX8782), .Z(WX8783) ) ;
INV     gate7012  (.A(WX8783), .Z(WX8784) ) ;
INV     gate7013  (.A(WX8763), .Z(WX8788) ) ;
OR2     gate7014  (.A(WX8787), .B(WX8786), .Z(WX8789) ) ;
INV     gate7015  (.A(WX8789), .Z(WX8790) ) ;
INV     gate7016  (.A(WX8790), .Z(WX8791) ) ;
INV     gate7017  (.A(WX8763), .Z(WX8795) ) ;
OR2     gate7018  (.A(WX8794), .B(WX8793), .Z(WX8796) ) ;
INV     gate7019  (.A(WX8796), .Z(WX8797) ) ;
INV     gate7020  (.A(WX8797), .Z(WX8798) ) ;
INV     gate7021  (.A(WX8763), .Z(WX8802) ) ;
OR2     gate7022  (.A(WX8801), .B(WX8800), .Z(WX8803) ) ;
INV     gate7023  (.A(WX8803), .Z(WX8804) ) ;
INV     gate7024  (.A(WX8804), .Z(WX8805) ) ;
INV     gate7025  (.A(WX8763), .Z(WX8809) ) ;
OR2     gate7026  (.A(WX8808), .B(WX8807), .Z(WX8810) ) ;
INV     gate7027  (.A(WX8810), .Z(WX8811) ) ;
INV     gate7028  (.A(WX8811), .Z(WX8812) ) ;
INV     gate7029  (.A(WX8763), .Z(WX8816) ) ;
OR2     gate7030  (.A(WX8815), .B(WX8814), .Z(WX8817) ) ;
INV     gate7031  (.A(WX8817), .Z(WX8818) ) ;
INV     gate7032  (.A(WX8818), .Z(WX8819) ) ;
INV     gate7033  (.A(WX8763), .Z(WX8823) ) ;
OR2     gate7034  (.A(WX8822), .B(WX8821), .Z(WX8824) ) ;
INV     gate7035  (.A(WX8824), .Z(WX8825) ) ;
INV     gate7036  (.A(WX8825), .Z(WX8826) ) ;
INV     gate7037  (.A(WX8763), .Z(WX8830) ) ;
OR2     gate7038  (.A(WX8829), .B(WX8828), .Z(WX8831) ) ;
INV     gate7039  (.A(WX8831), .Z(WX8832) ) ;
INV     gate7040  (.A(WX8832), .Z(WX8833) ) ;
INV     gate7041  (.A(WX8763), .Z(WX8837) ) ;
OR2     gate7042  (.A(WX8836), .B(WX8835), .Z(WX8838) ) ;
INV     gate7043  (.A(WX8838), .Z(WX8839) ) ;
INV     gate7044  (.A(WX8839), .Z(WX8840) ) ;
INV     gate7045  (.A(WX8763), .Z(WX8844) ) ;
OR2     gate7046  (.A(WX8843), .B(WX8842), .Z(WX8845) ) ;
INV     gate7047  (.A(WX8845), .Z(WX8846) ) ;
INV     gate7048  (.A(WX8846), .Z(WX8847) ) ;
INV     gate7049  (.A(WX8763), .Z(WX8851) ) ;
OR2     gate7050  (.A(WX8850), .B(WX8849), .Z(WX8852) ) ;
INV     gate7051  (.A(WX8852), .Z(WX8853) ) ;
INV     gate7052  (.A(WX8853), .Z(WX8854) ) ;
INV     gate7053  (.A(WX8763), .Z(WX8858) ) ;
OR2     gate7054  (.A(WX8857), .B(WX8856), .Z(WX8859) ) ;
INV     gate7055  (.A(WX8859), .Z(WX8860) ) ;
INV     gate7056  (.A(WX8860), .Z(WX8861) ) ;
INV     gate7057  (.A(WX8763), .Z(WX8865) ) ;
OR2     gate7058  (.A(WX8864), .B(WX8863), .Z(WX8866) ) ;
INV     gate7059  (.A(WX8866), .Z(WX8867) ) ;
INV     gate7060  (.A(WX8867), .Z(WX8868) ) ;
INV     gate7061  (.A(WX8763), .Z(WX8872) ) ;
OR2     gate7062  (.A(WX8871), .B(WX8870), .Z(WX8873) ) ;
INV     gate7063  (.A(WX8873), .Z(WX8874) ) ;
INV     gate7064  (.A(WX8874), .Z(WX8875) ) ;
INV     gate7065  (.A(WX8763), .Z(WX8879) ) ;
OR2     gate7066  (.A(WX8878), .B(WX8877), .Z(WX8880) ) ;
INV     gate7067  (.A(WX8880), .Z(WX8881) ) ;
INV     gate7068  (.A(WX8881), .Z(WX8882) ) ;
INV     gate7069  (.A(WX8763), .Z(WX8886) ) ;
OR2     gate7070  (.A(WX8885), .B(WX8884), .Z(WX8887) ) ;
INV     gate7071  (.A(WX8887), .Z(WX8888) ) ;
INV     gate7072  (.A(WX8888), .Z(WX8889) ) ;
INV     gate7073  (.A(WX8763), .Z(WX8893) ) ;
OR2     gate7074  (.A(WX8892), .B(WX8891), .Z(WX8894) ) ;
INV     gate7075  (.A(WX8894), .Z(WX8895) ) ;
INV     gate7076  (.A(WX8895), .Z(WX8896) ) ;
INV     gate7077  (.A(WX8763), .Z(WX8900) ) ;
OR2     gate7078  (.A(WX8899), .B(WX8898), .Z(WX8901) ) ;
INV     gate7079  (.A(WX8901), .Z(WX8902) ) ;
INV     gate7080  (.A(WX8902), .Z(WX8903) ) ;
INV     gate7081  (.A(WX8763), .Z(WX8907) ) ;
OR2     gate7082  (.A(WX8906), .B(WX8905), .Z(WX8908) ) ;
INV     gate7083  (.A(WX8908), .Z(WX8909) ) ;
INV     gate7084  (.A(WX8909), .Z(WX8910) ) ;
INV     gate7085  (.A(WX8763), .Z(WX8914) ) ;
OR2     gate7086  (.A(WX8913), .B(WX8912), .Z(WX8915) ) ;
INV     gate7087  (.A(WX8915), .Z(WX8916) ) ;
INV     gate7088  (.A(WX8916), .Z(WX8917) ) ;
INV     gate7089  (.A(WX8763), .Z(WX8921) ) ;
OR2     gate7090  (.A(WX8920), .B(WX8919), .Z(WX8922) ) ;
INV     gate7091  (.A(WX8922), .Z(WX8923) ) ;
INV     gate7092  (.A(WX8923), .Z(WX8924) ) ;
INV     gate7093  (.A(WX8763), .Z(WX8928) ) ;
OR2     gate7094  (.A(WX8927), .B(WX8926), .Z(WX8929) ) ;
INV     gate7095  (.A(WX8929), .Z(WX8930) ) ;
INV     gate7096  (.A(WX8930), .Z(WX8931) ) ;
INV     gate7097  (.A(WX8763), .Z(WX8935) ) ;
OR2     gate7098  (.A(WX8934), .B(WX8933), .Z(WX8936) ) ;
INV     gate7099  (.A(WX8936), .Z(WX8937) ) ;
INV     gate7100  (.A(WX8937), .Z(WX8938) ) ;
INV     gate7101  (.A(WX8763), .Z(WX8942) ) ;
OR2     gate7102  (.A(WX8941), .B(WX8940), .Z(WX8943) ) ;
INV     gate7103  (.A(WX8943), .Z(WX8944) ) ;
INV     gate7104  (.A(WX8944), .Z(WX8945) ) ;
INV     gate7105  (.A(WX8763), .Z(WX8949) ) ;
OR2     gate7106  (.A(WX8948), .B(WX8947), .Z(WX8950) ) ;
INV     gate7107  (.A(WX8950), .Z(WX8951) ) ;
INV     gate7108  (.A(WX8951), .Z(WX8952) ) ;
INV     gate7109  (.A(WX8763), .Z(WX8956) ) ;
OR2     gate7110  (.A(WX8955), .B(WX8954), .Z(WX8957) ) ;
INV     gate7111  (.A(WX8957), .Z(WX8958) ) ;
INV     gate7112  (.A(WX8958), .Z(WX8959) ) ;
INV     gate7113  (.A(WX8763), .Z(WX8963) ) ;
OR2     gate7114  (.A(WX8962), .B(WX8961), .Z(WX8964) ) ;
INV     gate7115  (.A(WX8964), .Z(WX8965) ) ;
INV     gate7116  (.A(WX8965), .Z(WX8966) ) ;
INV     gate7117  (.A(WX8763), .Z(WX8970) ) ;
OR2     gate7118  (.A(WX8969), .B(WX8968), .Z(WX8971) ) ;
INV     gate7119  (.A(WX8971), .Z(WX8972) ) ;
INV     gate7120  (.A(WX8972), .Z(WX8973) ) ;
INV     gate7121  (.A(WX8763), .Z(WX8977) ) ;
OR2     gate7122  (.A(WX8976), .B(WX8975), .Z(WX8978) ) ;
INV     gate7123  (.A(WX8978), .Z(WX8979) ) ;
INV     gate7124  (.A(WX8979), .Z(WX8980) ) ;
INV     gate7125  (.A(WX8763), .Z(WX8984) ) ;
OR2     gate7126  (.A(WX8983), .B(WX8982), .Z(WX8985) ) ;
INV     gate7127  (.A(WX8985), .Z(WX8986) ) ;
INV     gate7128  (.A(WX8986), .Z(WX8987) ) ;
INV     gate7129  (.A(RESET), .Z(WX8988) ) ;
INV     gate7130  (.A(WX8988), .Z(WX9021) ) ;
INV     gate7131  (.A(WX10050), .Z(WX10054) ) ;
INV     gate7132  (.A(WX10054), .Z(WX9088) ) ;
INV     gate7133  (.A(WX10048), .Z(WX10055) ) ;
INV     gate7134  (.A(WX10055), .Z(WX9092) ) ;
INV     gate7135  (.A(WX10055), .Z(WX9096) ) ;
OR2     gate7136  (.A(WX9087), .B(WX9086), .Z(WX9089) ) ;
INV     gate7137  (.A(WX9089), .Z(WX9098) ) ;
INV     gate7138  (.A(WX9098), .Z(WX9099) ) ;
INV     gate7139  (.A(WX10054), .Z(WX9102) ) ;
INV     gate7140  (.A(WX10055), .Z(WX9106) ) ;
INV     gate7141  (.A(WX10055), .Z(WX9110) ) ;
OR2     gate7142  (.A(WX9101), .B(WX9100), .Z(WX9103) ) ;
INV     gate7143  (.A(WX9103), .Z(WX9112) ) ;
INV     gate7144  (.A(WX9112), .Z(WX9113) ) ;
INV     gate7145  (.A(WX10054), .Z(WX9116) ) ;
INV     gate7146  (.A(WX10055), .Z(WX9120) ) ;
INV     gate7147  (.A(WX10055), .Z(WX9124) ) ;
OR2     gate7148  (.A(WX9115), .B(WX9114), .Z(WX9117) ) ;
INV     gate7149  (.A(WX9117), .Z(WX9126) ) ;
INV     gate7150  (.A(WX9126), .Z(WX9127) ) ;
INV     gate7151  (.A(WX10054), .Z(WX9130) ) ;
INV     gate7152  (.A(WX10055), .Z(WX9134) ) ;
INV     gate7153  (.A(WX10055), .Z(WX9138) ) ;
OR2     gate7154  (.A(WX9129), .B(WX9128), .Z(WX9131) ) ;
INV     gate7155  (.A(WX9131), .Z(WX9140) ) ;
INV     gate7156  (.A(WX9140), .Z(WX9141) ) ;
INV     gate7157  (.A(WX10054), .Z(WX9144) ) ;
INV     gate7158  (.A(WX10055), .Z(WX9148) ) ;
INV     gate7159  (.A(WX10055), .Z(WX9152) ) ;
OR2     gate7160  (.A(WX9143), .B(WX9142), .Z(WX9145) ) ;
INV     gate7161  (.A(WX9145), .Z(WX9154) ) ;
INV     gate7162  (.A(WX9154), .Z(WX9155) ) ;
INV     gate7163  (.A(WX10054), .Z(WX9158) ) ;
INV     gate7164  (.A(WX10055), .Z(WX9162) ) ;
INV     gate7165  (.A(WX10055), .Z(WX9166) ) ;
OR2     gate7166  (.A(WX9157), .B(WX9156), .Z(WX9159) ) ;
INV     gate7167  (.A(WX9159), .Z(WX9168) ) ;
INV     gate7168  (.A(WX9168), .Z(WX9169) ) ;
INV     gate7169  (.A(WX10054), .Z(WX9172) ) ;
INV     gate7170  (.A(WX10055), .Z(WX9176) ) ;
INV     gate7171  (.A(WX10055), .Z(WX9180) ) ;
OR2     gate7172  (.A(WX9171), .B(WX9170), .Z(WX9173) ) ;
INV     gate7173  (.A(WX9173), .Z(WX9182) ) ;
INV     gate7174  (.A(WX9182), .Z(WX9183) ) ;
INV     gate7175  (.A(WX10054), .Z(WX9186) ) ;
INV     gate7176  (.A(WX10055), .Z(WX9190) ) ;
INV     gate7177  (.A(WX10055), .Z(WX9194) ) ;
OR2     gate7178  (.A(WX9185), .B(WX9184), .Z(WX9187) ) ;
INV     gate7179  (.A(WX9187), .Z(WX9196) ) ;
INV     gate7180  (.A(WX9196), .Z(WX9197) ) ;
INV     gate7181  (.A(WX10054), .Z(WX9200) ) ;
INV     gate7182  (.A(WX10055), .Z(WX9204) ) ;
INV     gate7183  (.A(WX10055), .Z(WX9208) ) ;
OR2     gate7184  (.A(WX9199), .B(WX9198), .Z(WX9201) ) ;
INV     gate7185  (.A(WX9201), .Z(WX9210) ) ;
INV     gate7186  (.A(WX9210), .Z(WX9211) ) ;
INV     gate7187  (.A(WX10054), .Z(WX9214) ) ;
INV     gate7188  (.A(WX10055), .Z(WX9218) ) ;
INV     gate7189  (.A(WX10055), .Z(WX9222) ) ;
OR2     gate7190  (.A(WX9213), .B(WX9212), .Z(WX9215) ) ;
INV     gate7191  (.A(WX9215), .Z(WX9224) ) ;
INV     gate7192  (.A(WX9224), .Z(WX9225) ) ;
INV     gate7193  (.A(WX10054), .Z(WX9228) ) ;
INV     gate7194  (.A(WX10055), .Z(WX9232) ) ;
INV     gate7195  (.A(WX10055), .Z(WX9236) ) ;
OR2     gate7196  (.A(WX9227), .B(WX9226), .Z(WX9229) ) ;
INV     gate7197  (.A(WX9229), .Z(WX9238) ) ;
INV     gate7198  (.A(WX9238), .Z(WX9239) ) ;
INV     gate7199  (.A(WX10054), .Z(WX9242) ) ;
INV     gate7200  (.A(WX10055), .Z(WX9246) ) ;
INV     gate7201  (.A(WX10055), .Z(WX9250) ) ;
OR2     gate7202  (.A(WX9241), .B(WX9240), .Z(WX9243) ) ;
INV     gate7203  (.A(WX9243), .Z(WX9252) ) ;
INV     gate7204  (.A(WX9252), .Z(WX9253) ) ;
INV     gate7205  (.A(WX10054), .Z(WX9256) ) ;
INV     gate7206  (.A(WX10055), .Z(WX9260) ) ;
INV     gate7207  (.A(WX10055), .Z(WX9264) ) ;
OR2     gate7208  (.A(WX9255), .B(WX9254), .Z(WX9257) ) ;
INV     gate7209  (.A(WX9257), .Z(WX9266) ) ;
INV     gate7210  (.A(WX9266), .Z(WX9267) ) ;
INV     gate7211  (.A(WX10054), .Z(WX9270) ) ;
INV     gate7212  (.A(WX10055), .Z(WX9274) ) ;
INV     gate7213  (.A(WX10055), .Z(WX9278) ) ;
OR2     gate7214  (.A(WX9269), .B(WX9268), .Z(WX9271) ) ;
INV     gate7215  (.A(WX9271), .Z(WX9280) ) ;
INV     gate7216  (.A(WX9280), .Z(WX9281) ) ;
INV     gate7217  (.A(WX10054), .Z(WX9284) ) ;
INV     gate7218  (.A(WX10055), .Z(WX9288) ) ;
INV     gate7219  (.A(WX10055), .Z(WX9292) ) ;
OR2     gate7220  (.A(WX9283), .B(WX9282), .Z(WX9285) ) ;
INV     gate7221  (.A(WX9285), .Z(WX9294) ) ;
INV     gate7222  (.A(WX9294), .Z(WX9295) ) ;
INV     gate7223  (.A(WX10054), .Z(WX9298) ) ;
INV     gate7224  (.A(WX10055), .Z(WX9302) ) ;
INV     gate7225  (.A(WX10055), .Z(WX9306) ) ;
OR2     gate7226  (.A(WX9297), .B(WX9296), .Z(WX9299) ) ;
INV     gate7227  (.A(WX9299), .Z(WX9308) ) ;
INV     gate7228  (.A(WX9308), .Z(WX9309) ) ;
INV     gate7229  (.A(WX10054), .Z(WX9312) ) ;
INV     gate7230  (.A(WX10055), .Z(WX9316) ) ;
INV     gate7231  (.A(WX10055), .Z(WX9320) ) ;
OR2     gate7232  (.A(WX9311), .B(WX9310), .Z(WX9313) ) ;
INV     gate7233  (.A(WX9313), .Z(WX9322) ) ;
INV     gate7234  (.A(WX9322), .Z(WX9323) ) ;
INV     gate7235  (.A(WX10054), .Z(WX9326) ) ;
INV     gate7236  (.A(WX10055), .Z(WX9330) ) ;
INV     gate7237  (.A(WX10055), .Z(WX9334) ) ;
OR2     gate7238  (.A(WX9325), .B(WX9324), .Z(WX9327) ) ;
INV     gate7239  (.A(WX9327), .Z(WX9336) ) ;
INV     gate7240  (.A(WX9336), .Z(WX9337) ) ;
INV     gate7241  (.A(WX10054), .Z(WX9340) ) ;
INV     gate7242  (.A(WX10055), .Z(WX9344) ) ;
INV     gate7243  (.A(WX10055), .Z(WX9348) ) ;
OR2     gate7244  (.A(WX9339), .B(WX9338), .Z(WX9341) ) ;
INV     gate7245  (.A(WX9341), .Z(WX9350) ) ;
INV     gate7246  (.A(WX9350), .Z(WX9351) ) ;
INV     gate7247  (.A(WX10054), .Z(WX9354) ) ;
INV     gate7248  (.A(WX10055), .Z(WX9358) ) ;
INV     gate7249  (.A(WX10055), .Z(WX9362) ) ;
OR2     gate7250  (.A(WX9353), .B(WX9352), .Z(WX9355) ) ;
INV     gate7251  (.A(WX9355), .Z(WX9364) ) ;
INV     gate7252  (.A(WX9364), .Z(WX9365) ) ;
INV     gate7253  (.A(WX10054), .Z(WX9368) ) ;
INV     gate7254  (.A(WX10055), .Z(WX9372) ) ;
INV     gate7255  (.A(WX10055), .Z(WX9376) ) ;
OR2     gate7256  (.A(WX9367), .B(WX9366), .Z(WX9369) ) ;
INV     gate7257  (.A(WX9369), .Z(WX9378) ) ;
INV     gate7258  (.A(WX9378), .Z(WX9379) ) ;
INV     gate7259  (.A(WX10054), .Z(WX9382) ) ;
INV     gate7260  (.A(WX10055), .Z(WX9386) ) ;
INV     gate7261  (.A(WX10055), .Z(WX9390) ) ;
OR2     gate7262  (.A(WX9381), .B(WX9380), .Z(WX9383) ) ;
INV     gate7263  (.A(WX9383), .Z(WX9392) ) ;
INV     gate7264  (.A(WX9392), .Z(WX9393) ) ;
INV     gate7265  (.A(WX10054), .Z(WX9396) ) ;
INV     gate7266  (.A(WX10055), .Z(WX9400) ) ;
INV     gate7267  (.A(WX10055), .Z(WX9404) ) ;
OR2     gate7268  (.A(WX9395), .B(WX9394), .Z(WX9397) ) ;
INV     gate7269  (.A(WX9397), .Z(WX9406) ) ;
INV     gate7270  (.A(WX9406), .Z(WX9407) ) ;
INV     gate7271  (.A(WX10054), .Z(WX9410) ) ;
INV     gate7272  (.A(WX10055), .Z(WX9414) ) ;
INV     gate7273  (.A(WX10055), .Z(WX9418) ) ;
OR2     gate7274  (.A(WX9409), .B(WX9408), .Z(WX9411) ) ;
INV     gate7275  (.A(WX9411), .Z(WX9420) ) ;
INV     gate7276  (.A(WX9420), .Z(WX9421) ) ;
INV     gate7277  (.A(WX10054), .Z(WX9424) ) ;
INV     gate7278  (.A(WX10055), .Z(WX9428) ) ;
INV     gate7279  (.A(WX10055), .Z(WX9432) ) ;
OR2     gate7280  (.A(WX9423), .B(WX9422), .Z(WX9425) ) ;
INV     gate7281  (.A(WX9425), .Z(WX9434) ) ;
INV     gate7282  (.A(WX9434), .Z(WX9435) ) ;
INV     gate7283  (.A(WX10054), .Z(WX9438) ) ;
INV     gate7284  (.A(WX10055), .Z(WX9442) ) ;
INV     gate7285  (.A(WX10055), .Z(WX9446) ) ;
OR2     gate7286  (.A(WX9437), .B(WX9436), .Z(WX9439) ) ;
INV     gate7287  (.A(WX9439), .Z(WX9448) ) ;
INV     gate7288  (.A(WX9448), .Z(WX9449) ) ;
INV     gate7289  (.A(WX10054), .Z(WX9452) ) ;
INV     gate7290  (.A(WX10055), .Z(WX9456) ) ;
INV     gate7291  (.A(WX10055), .Z(WX9460) ) ;
OR2     gate7292  (.A(WX9451), .B(WX9450), .Z(WX9453) ) ;
INV     gate7293  (.A(WX9453), .Z(WX9462) ) ;
INV     gate7294  (.A(WX9462), .Z(WX9463) ) ;
INV     gate7295  (.A(WX10054), .Z(WX9466) ) ;
INV     gate7296  (.A(WX10055), .Z(WX9470) ) ;
INV     gate7297  (.A(WX10055), .Z(WX9474) ) ;
OR2     gate7298  (.A(WX9465), .B(WX9464), .Z(WX9467) ) ;
INV     gate7299  (.A(WX9467), .Z(WX9476) ) ;
INV     gate7300  (.A(WX9476), .Z(WX9477) ) ;
INV     gate7301  (.A(WX10054), .Z(WX9480) ) ;
INV     gate7302  (.A(WX10055), .Z(WX9484) ) ;
INV     gate7303  (.A(WX10055), .Z(WX9488) ) ;
OR2     gate7304  (.A(WX9479), .B(WX9478), .Z(WX9481) ) ;
INV     gate7305  (.A(WX9481), .Z(WX9490) ) ;
INV     gate7306  (.A(WX9490), .Z(WX9491) ) ;
INV     gate7307  (.A(WX10054), .Z(WX9494) ) ;
INV     gate7308  (.A(WX10055), .Z(WX9498) ) ;
INV     gate7309  (.A(WX10055), .Z(WX9502) ) ;
OR2     gate7310  (.A(WX9493), .B(WX9492), .Z(WX9495) ) ;
INV     gate7311  (.A(WX9495), .Z(WX9504) ) ;
INV     gate7312  (.A(WX9504), .Z(WX9505) ) ;
INV     gate7313  (.A(WX10054), .Z(WX9508) ) ;
INV     gate7314  (.A(WX10055), .Z(WX9512) ) ;
INV     gate7315  (.A(WX10055), .Z(WX9516) ) ;
OR2     gate7316  (.A(WX9507), .B(WX9506), .Z(WX9509) ) ;
INV     gate7317  (.A(WX9509), .Z(WX9518) ) ;
INV     gate7318  (.A(WX9518), .Z(WX9519) ) ;
INV     gate7319  (.A(WX10054), .Z(WX9522) ) ;
INV     gate7320  (.A(WX10055), .Z(WX9526) ) ;
INV     gate7321  (.A(WX10055), .Z(WX9530) ) ;
OR2     gate7322  (.A(WX9521), .B(WX9520), .Z(WX9523) ) ;
INV     gate7323  (.A(WX9523), .Z(WX9532) ) ;
INV     gate7324  (.A(WX9532), .Z(WX9533) ) ;
INV     gate7325  (.A(WX9536), .Z(WX9534) ) ;
INV     gate7326  (.A(WX10015), .Z(WX10016) ) ;
INV     gate7327  (.A(WX10016), .Z(WX9599) ) ;
INV     gate7328  (.A(WX10017), .Z(WX10018) ) ;
INV     gate7329  (.A(WX10018), .Z(WX9600) ) ;
INV     gate7330  (.A(WX10019), .Z(WX10020) ) ;
INV     gate7331  (.A(WX10020), .Z(WX9601) ) ;
INV     gate7332  (.A(WX10021), .Z(WX10022) ) ;
INV     gate7333  (.A(WX10022), .Z(WX9602) ) ;
INV     gate7334  (.A(WX10023), .Z(WX10024) ) ;
INV     gate7335  (.A(WX10024), .Z(WX9603) ) ;
INV     gate7336  (.A(WX10025), .Z(WX10026) ) ;
INV     gate7337  (.A(WX10026), .Z(WX9604) ) ;
INV     gate7338  (.A(WX10027), .Z(WX10028) ) ;
INV     gate7339  (.A(WX10028), .Z(WX9605) ) ;
INV     gate7340  (.A(WX10029), .Z(WX10030) ) ;
INV     gate7341  (.A(WX10030), .Z(WX9606) ) ;
INV     gate7342  (.A(WX10031), .Z(WX10032) ) ;
INV     gate7343  (.A(WX10032), .Z(WX9607) ) ;
INV     gate7344  (.A(WX10033), .Z(WX10034) ) ;
INV     gate7345  (.A(WX10034), .Z(WX9608) ) ;
INV     gate7346  (.A(WX10035), .Z(WX10036) ) ;
INV     gate7347  (.A(WX10036), .Z(WX9609) ) ;
INV     gate7348  (.A(WX10037), .Z(WX10038) ) ;
INV     gate7349  (.A(WX10038), .Z(WX9610) ) ;
INV     gate7350  (.A(WX10039), .Z(WX10040) ) ;
INV     gate7351  (.A(WX10040), .Z(WX9611) ) ;
INV     gate7352  (.A(WX10041), .Z(WX10042) ) ;
INV     gate7353  (.A(WX10042), .Z(WX9612) ) ;
INV     gate7354  (.A(WX10043), .Z(WX10044) ) ;
INV     gate7355  (.A(WX10044), .Z(WX9613) ) ;
INV     gate7356  (.A(WX10045), .Z(WX10046) ) ;
INV     gate7357  (.A(WX10046), .Z(WX9614) ) ;
INV     gate7358  (.A(WX9983), .Z(WX9984) ) ;
INV     gate7359  (.A(WX9984), .Z(WX9615) ) ;
INV     gate7360  (.A(WX9985), .Z(WX9986) ) ;
INV     gate7361  (.A(WX9986), .Z(WX9616) ) ;
INV     gate7362  (.A(WX9987), .Z(WX9988) ) ;
INV     gate7363  (.A(WX9988), .Z(WX9617) ) ;
INV     gate7364  (.A(WX9989), .Z(WX9990) ) ;
INV     gate7365  (.A(WX9990), .Z(WX9618) ) ;
INV     gate7366  (.A(WX9991), .Z(WX9992) ) ;
INV     gate7367  (.A(WX9992), .Z(WX9619) ) ;
INV     gate7368  (.A(WX9993), .Z(WX9994) ) ;
INV     gate7369  (.A(WX9994), .Z(WX9620) ) ;
INV     gate7370  (.A(WX9995), .Z(WX9996) ) ;
INV     gate7371  (.A(WX9996), .Z(WX9621) ) ;
INV     gate7372  (.A(WX9997), .Z(WX9998) ) ;
INV     gate7373  (.A(WX9998), .Z(WX9622) ) ;
INV     gate7374  (.A(WX9999), .Z(WX10000) ) ;
INV     gate7375  (.A(WX10000), .Z(WX9623) ) ;
INV     gate7376  (.A(WX10001), .Z(WX10002) ) ;
INV     gate7377  (.A(WX10002), .Z(WX9624) ) ;
INV     gate7378  (.A(WX10003), .Z(WX10004) ) ;
INV     gate7379  (.A(WX10004), .Z(WX9625) ) ;
INV     gate7380  (.A(WX10005), .Z(WX10006) ) ;
INV     gate7381  (.A(WX10006), .Z(WX9626) ) ;
INV     gate7382  (.A(WX10007), .Z(WX10008) ) ;
INV     gate7383  (.A(WX10008), .Z(WX9627) ) ;
INV     gate7384  (.A(WX10009), .Z(WX10010) ) ;
INV     gate7385  (.A(WX10010), .Z(WX9628) ) ;
INV     gate7386  (.A(WX10011), .Z(WX10012) ) ;
INV     gate7387  (.A(WX10012), .Z(WX9629) ) ;
INV     gate7388  (.A(WX10013), .Z(WX10014) ) ;
INV     gate7389  (.A(WX10014), .Z(WX9630) ) ;
INV     gate7390  (.A(WX9599), .Z(WX9631) ) ;
INV     gate7391  (.A(WX9600), .Z(WX9632) ) ;
INV     gate7392  (.A(WX9601), .Z(WX9633) ) ;
INV     gate7393  (.A(WX9602), .Z(WX9634) ) ;
INV     gate7394  (.A(WX9603), .Z(WX9635) ) ;
INV     gate7395  (.A(WX9604), .Z(WX9636) ) ;
INV     gate7396  (.A(WX9605), .Z(WX9637) ) ;
INV     gate7397  (.A(WX9606), .Z(WX9638) ) ;
INV     gate7398  (.A(WX9607), .Z(WX9639) ) ;
INV     gate7399  (.A(WX9608), .Z(WX9640) ) ;
INV     gate7400  (.A(WX9609), .Z(WX9641) ) ;
INV     gate7401  (.A(WX9610), .Z(WX9642) ) ;
INV     gate7402  (.A(WX9611), .Z(WX9643) ) ;
INV     gate7403  (.A(WX9612), .Z(WX9644) ) ;
INV     gate7404  (.A(WX9613), .Z(WX9645) ) ;
INV     gate7405  (.A(WX9614), .Z(WX9646) ) ;
INV     gate7406  (.A(WX9615), .Z(WX9647) ) ;
INV     gate7407  (.A(WX9616), .Z(WX9648) ) ;
INV     gate7408  (.A(WX9617), .Z(WX9649) ) ;
INV     gate7409  (.A(WX9618), .Z(WX9650) ) ;
INV     gate7410  (.A(WX9619), .Z(WX9651) ) ;
INV     gate7411  (.A(WX9620), .Z(WX9652) ) ;
INV     gate7412  (.A(WX9621), .Z(WX9653) ) ;
INV     gate7413  (.A(WX9622), .Z(WX9654) ) ;
INV     gate7414  (.A(WX9623), .Z(WX9655) ) ;
INV     gate7415  (.A(WX9624), .Z(WX9656) ) ;
INV     gate7416  (.A(WX9625), .Z(WX9657) ) ;
INV     gate7417  (.A(WX9626), .Z(WX9658) ) ;
INV     gate7418  (.A(WX9627), .Z(WX9659) ) ;
INV     gate7419  (.A(WX9628), .Z(WX9660) ) ;
INV     gate7420  (.A(WX9629), .Z(WX9661) ) ;
INV     gate7421  (.A(WX9630), .Z(WX9662) ) ;
INV     gate7422  (.A(WX9888), .Z(WX9663) ) ;
INV     gate7423  (.A(WX9890), .Z(WX9664) ) ;
INV     gate7424  (.A(WX9892), .Z(WX9665) ) ;
INV     gate7425  (.A(WX9894), .Z(WX9666) ) ;
INV     gate7426  (.A(WX9896), .Z(WX9667) ) ;
INV     gate7427  (.A(WX9898), .Z(WX9668) ) ;
INV     gate7428  (.A(WX9900), .Z(WX9669) ) ;
INV     gate7429  (.A(WX9902), .Z(WX9670) ) ;
INV     gate7430  (.A(WX9904), .Z(WX9671) ) ;
INV     gate7431  (.A(WX9906), .Z(WX9672) ) ;
INV     gate7432  (.A(WX9908), .Z(WX9673) ) ;
INV     gate7433  (.A(WX9910), .Z(WX9674) ) ;
INV     gate7434  (.A(WX9912), .Z(WX9675) ) ;
INV     gate7435  (.A(WX9914), .Z(WX9676) ) ;
INV     gate7436  (.A(WX9916), .Z(WX9677) ) ;
INV     gate7437  (.A(WX9918), .Z(WX9678) ) ;
INV     gate7438  (.A(WX9920), .Z(WX9679) ) ;
INV     gate7439  (.A(WX9922), .Z(WX9680) ) ;
INV     gate7440  (.A(WX9924), .Z(WX9681) ) ;
INV     gate7441  (.A(WX9926), .Z(WX9682) ) ;
INV     gate7442  (.A(WX9928), .Z(WX9683) ) ;
INV     gate7443  (.A(WX9930), .Z(WX9684) ) ;
INV     gate7444  (.A(WX9932), .Z(WX9685) ) ;
INV     gate7445  (.A(WX9934), .Z(WX9686) ) ;
INV     gate7446  (.A(WX9936), .Z(WX9687) ) ;
INV     gate7447  (.A(WX9938), .Z(WX9688) ) ;
INV     gate7448  (.A(WX9940), .Z(WX9689) ) ;
INV     gate7449  (.A(WX9942), .Z(WX9690) ) ;
INV     gate7450  (.A(WX9944), .Z(WX9691) ) ;
INV     gate7451  (.A(WX9946), .Z(WX9692) ) ;
INV     gate7452  (.A(WX9948), .Z(WX9693) ) ;
INV     gate7453  (.A(WX9950), .Z(WX9694) ) ;
NAND2   gate7454  (.A(II30542), .B(II30543), .Z(WX9967) ) ;
INV     gate7455  (.A(WX9967), .Z(WX9983) ) ;
NAND2   gate7456  (.A(II30573), .B(II30574), .Z(WX9968) ) ;
INV     gate7457  (.A(WX9968), .Z(WX9985) ) ;
NAND2   gate7458  (.A(II30604), .B(II30605), .Z(WX9969) ) ;
INV     gate7459  (.A(WX9969), .Z(WX9987) ) ;
NAND2   gate7460  (.A(II30635), .B(II30636), .Z(WX9970) ) ;
INV     gate7461  (.A(WX9970), .Z(WX9989) ) ;
NAND2   gate7462  (.A(II30666), .B(II30667), .Z(WX9971) ) ;
INV     gate7463  (.A(WX9971), .Z(WX9991) ) ;
NAND2   gate7464  (.A(II30697), .B(II30698), .Z(WX9972) ) ;
INV     gate7465  (.A(WX9972), .Z(WX9993) ) ;
NAND2   gate7466  (.A(II30728), .B(II30729), .Z(WX9973) ) ;
INV     gate7467  (.A(WX9973), .Z(WX9995) ) ;
NAND2   gate7468  (.A(II30759), .B(II30760), .Z(WX9974) ) ;
INV     gate7469  (.A(WX9974), .Z(WX9997) ) ;
NAND2   gate7470  (.A(II30790), .B(II30791), .Z(WX9975) ) ;
INV     gate7471  (.A(WX9975), .Z(WX9999) ) ;
NAND2   gate7472  (.A(II30821), .B(II30822), .Z(WX9976) ) ;
INV     gate7473  (.A(WX9976), .Z(WX10001) ) ;
NAND2   gate7474  (.A(II30852), .B(II30853), .Z(WX9977) ) ;
INV     gate7475  (.A(WX9977), .Z(WX10003) ) ;
NAND2   gate7476  (.A(II30883), .B(II30884), .Z(WX9978) ) ;
INV     gate7477  (.A(WX9978), .Z(WX10005) ) ;
NAND2   gate7478  (.A(II30914), .B(II30915), .Z(WX9979) ) ;
INV     gate7479  (.A(WX9979), .Z(WX10007) ) ;
NAND2   gate7480  (.A(II30945), .B(II30946), .Z(WX9980) ) ;
INV     gate7481  (.A(WX9980), .Z(WX10009) ) ;
NAND2   gate7482  (.A(II30976), .B(II30977), .Z(WX9981) ) ;
INV     gate7483  (.A(WX9981), .Z(WX10011) ) ;
NAND2   gate7484  (.A(II31007), .B(II31008), .Z(WX9982) ) ;
INV     gate7485  (.A(WX9982), .Z(WX10013) ) ;
NAND2   gate7486  (.A(II30046), .B(II30047), .Z(WX9951) ) ;
INV     gate7487  (.A(WX9951), .Z(WX10015) ) ;
NAND2   gate7488  (.A(II30077), .B(II30078), .Z(WX9952) ) ;
INV     gate7489  (.A(WX9952), .Z(WX10017) ) ;
NAND2   gate7490  (.A(II30108), .B(II30109), .Z(WX9953) ) ;
INV     gate7491  (.A(WX9953), .Z(WX10019) ) ;
NAND2   gate7492  (.A(II30139), .B(II30140), .Z(WX9954) ) ;
INV     gate7493  (.A(WX9954), .Z(WX10021) ) ;
NAND2   gate7494  (.A(II30170), .B(II30171), .Z(WX9955) ) ;
INV     gate7495  (.A(WX9955), .Z(WX10023) ) ;
NAND2   gate7496  (.A(II30201), .B(II30202), .Z(WX9956) ) ;
INV     gate7497  (.A(WX9956), .Z(WX10025) ) ;
NAND2   gate7498  (.A(II30232), .B(II30233), .Z(WX9957) ) ;
INV     gate7499  (.A(WX9957), .Z(WX10027) ) ;
NAND2   gate7500  (.A(II30263), .B(II30264), .Z(WX9958) ) ;
INV     gate7501  (.A(WX9958), .Z(WX10029) ) ;
NAND2   gate7502  (.A(II30294), .B(II30295), .Z(WX9959) ) ;
INV     gate7503  (.A(WX9959), .Z(WX10031) ) ;
NAND2   gate7504  (.A(II30325), .B(II30326), .Z(WX9960) ) ;
INV     gate7505  (.A(WX9960), .Z(WX10033) ) ;
NAND2   gate7506  (.A(II30356), .B(II30357), .Z(WX9961) ) ;
INV     gate7507  (.A(WX9961), .Z(WX10035) ) ;
NAND2   gate7508  (.A(II30387), .B(II30388), .Z(WX9962) ) ;
INV     gate7509  (.A(WX9962), .Z(WX10037) ) ;
NAND2   gate7510  (.A(II30418), .B(II30419), .Z(WX9963) ) ;
INV     gate7511  (.A(WX9963), .Z(WX10039) ) ;
NAND2   gate7512  (.A(II30449), .B(II30450), .Z(WX9964) ) ;
INV     gate7513  (.A(WX9964), .Z(WX10041) ) ;
NAND2   gate7514  (.A(II30480), .B(II30481), .Z(WX9965) ) ;
INV     gate7515  (.A(WX9965), .Z(WX10043) ) ;
NAND2   gate7516  (.A(II30511), .B(II30512), .Z(WX9966) ) ;
INV     gate7517  (.A(WX9966), .Z(WX10045) ) ;
INV     gate7518  (.A(TM0), .Z(WX10047) ) ;
INV     gate7519  (.A(TM0), .Z(WX10048) ) ;
INV     gate7520  (.A(TM0), .Z(WX10049) ) ;
INV     gate7521  (.A(TM1), .Z(WX10050) ) ;
INV     gate7522  (.A(TM1), .Z(WX10051) ) ;
INV     gate7523  (.A(WX10051), .Z(WX10052) ) ;
INV     gate7524  (.A(WX10049), .Z(WX10053) ) ;
INV     gate7525  (.A(WX10047), .Z(WX10056) ) ;
INV     gate7526  (.A(WX10056), .Z(WX10060) ) ;
OR2     gate7527  (.A(WX10059), .B(WX10058), .Z(WX10061) ) ;
INV     gate7528  (.A(WX10061), .Z(WX10062) ) ;
INV     gate7529  (.A(WX10062), .Z(WX10063) ) ;
INV     gate7530  (.A(WX10056), .Z(WX10067) ) ;
OR2     gate7531  (.A(WX10066), .B(WX10065), .Z(WX10068) ) ;
INV     gate7532  (.A(WX10068), .Z(WX10069) ) ;
INV     gate7533  (.A(WX10069), .Z(WX10070) ) ;
INV     gate7534  (.A(WX10056), .Z(WX10074) ) ;
OR2     gate7535  (.A(WX10073), .B(WX10072), .Z(WX10075) ) ;
INV     gate7536  (.A(WX10075), .Z(WX10076) ) ;
INV     gate7537  (.A(WX10076), .Z(WX10077) ) ;
INV     gate7538  (.A(WX10056), .Z(WX10081) ) ;
OR2     gate7539  (.A(WX10080), .B(WX10079), .Z(WX10082) ) ;
INV     gate7540  (.A(WX10082), .Z(WX10083) ) ;
INV     gate7541  (.A(WX10083), .Z(WX10084) ) ;
INV     gate7542  (.A(WX10056), .Z(WX10088) ) ;
OR2     gate7543  (.A(WX10087), .B(WX10086), .Z(WX10089) ) ;
INV     gate7544  (.A(WX10089), .Z(WX10090) ) ;
INV     gate7545  (.A(WX10090), .Z(WX10091) ) ;
INV     gate7546  (.A(WX10056), .Z(WX10095) ) ;
OR2     gate7547  (.A(WX10094), .B(WX10093), .Z(WX10096) ) ;
INV     gate7548  (.A(WX10096), .Z(WX10097) ) ;
INV     gate7549  (.A(WX10097), .Z(WX10098) ) ;
INV     gate7550  (.A(WX10056), .Z(WX10102) ) ;
OR2     gate7551  (.A(WX10101), .B(WX10100), .Z(WX10103) ) ;
INV     gate7552  (.A(WX10103), .Z(WX10104) ) ;
INV     gate7553  (.A(WX10104), .Z(WX10105) ) ;
INV     gate7554  (.A(WX10056), .Z(WX10109) ) ;
OR2     gate7555  (.A(WX10108), .B(WX10107), .Z(WX10110) ) ;
INV     gate7556  (.A(WX10110), .Z(WX10111) ) ;
INV     gate7557  (.A(WX10111), .Z(WX10112) ) ;
INV     gate7558  (.A(WX10056), .Z(WX10116) ) ;
OR2     gate7559  (.A(WX10115), .B(WX10114), .Z(WX10117) ) ;
INV     gate7560  (.A(WX10117), .Z(WX10118) ) ;
INV     gate7561  (.A(WX10118), .Z(WX10119) ) ;
INV     gate7562  (.A(WX10056), .Z(WX10123) ) ;
OR2     gate7563  (.A(WX10122), .B(WX10121), .Z(WX10124) ) ;
INV     gate7564  (.A(WX10124), .Z(WX10125) ) ;
INV     gate7565  (.A(WX10125), .Z(WX10126) ) ;
INV     gate7566  (.A(WX10056), .Z(WX10130) ) ;
OR2     gate7567  (.A(WX10129), .B(WX10128), .Z(WX10131) ) ;
INV     gate7568  (.A(WX10131), .Z(WX10132) ) ;
INV     gate7569  (.A(WX10132), .Z(WX10133) ) ;
INV     gate7570  (.A(WX10056), .Z(WX10137) ) ;
OR2     gate7571  (.A(WX10136), .B(WX10135), .Z(WX10138) ) ;
INV     gate7572  (.A(WX10138), .Z(WX10139) ) ;
INV     gate7573  (.A(WX10139), .Z(WX10140) ) ;
INV     gate7574  (.A(WX10056), .Z(WX10144) ) ;
OR2     gate7575  (.A(WX10143), .B(WX10142), .Z(WX10145) ) ;
INV     gate7576  (.A(WX10145), .Z(WX10146) ) ;
INV     gate7577  (.A(WX10146), .Z(WX10147) ) ;
INV     gate7578  (.A(WX10056), .Z(WX10151) ) ;
OR2     gate7579  (.A(WX10150), .B(WX10149), .Z(WX10152) ) ;
INV     gate7580  (.A(WX10152), .Z(WX10153) ) ;
INV     gate7581  (.A(WX10153), .Z(WX10154) ) ;
INV     gate7582  (.A(WX10056), .Z(WX10158) ) ;
OR2     gate7583  (.A(WX10157), .B(WX10156), .Z(WX10159) ) ;
INV     gate7584  (.A(WX10159), .Z(WX10160) ) ;
INV     gate7585  (.A(WX10160), .Z(WX10161) ) ;
INV     gate7586  (.A(WX10056), .Z(WX10165) ) ;
OR2     gate7587  (.A(WX10164), .B(WX10163), .Z(WX10166) ) ;
INV     gate7588  (.A(WX10166), .Z(WX10167) ) ;
INV     gate7589  (.A(WX10167), .Z(WX10168) ) ;
INV     gate7590  (.A(WX10056), .Z(WX10172) ) ;
OR2     gate7591  (.A(WX10171), .B(WX10170), .Z(WX10173) ) ;
INV     gate7592  (.A(WX10173), .Z(WX10174) ) ;
INV     gate7593  (.A(WX10174), .Z(WX10175) ) ;
INV     gate7594  (.A(WX10056), .Z(WX10179) ) ;
OR2     gate7595  (.A(WX10178), .B(WX10177), .Z(WX10180) ) ;
INV     gate7596  (.A(WX10180), .Z(WX10181) ) ;
INV     gate7597  (.A(WX10181), .Z(WX10182) ) ;
INV     gate7598  (.A(WX10056), .Z(WX10186) ) ;
OR2     gate7599  (.A(WX10185), .B(WX10184), .Z(WX10187) ) ;
INV     gate7600  (.A(WX10187), .Z(WX10188) ) ;
INV     gate7601  (.A(WX10188), .Z(WX10189) ) ;
INV     gate7602  (.A(WX10056), .Z(WX10193) ) ;
OR2     gate7603  (.A(WX10192), .B(WX10191), .Z(WX10194) ) ;
INV     gate7604  (.A(WX10194), .Z(WX10195) ) ;
INV     gate7605  (.A(WX10195), .Z(WX10196) ) ;
INV     gate7606  (.A(WX10056), .Z(WX10200) ) ;
OR2     gate7607  (.A(WX10199), .B(WX10198), .Z(WX10201) ) ;
INV     gate7608  (.A(WX10201), .Z(WX10202) ) ;
INV     gate7609  (.A(WX10202), .Z(WX10203) ) ;
INV     gate7610  (.A(WX10056), .Z(WX10207) ) ;
OR2     gate7611  (.A(WX10206), .B(WX10205), .Z(WX10208) ) ;
INV     gate7612  (.A(WX10208), .Z(WX10209) ) ;
INV     gate7613  (.A(WX10209), .Z(WX10210) ) ;
INV     gate7614  (.A(WX10056), .Z(WX10214) ) ;
OR2     gate7615  (.A(WX10213), .B(WX10212), .Z(WX10215) ) ;
INV     gate7616  (.A(WX10215), .Z(WX10216) ) ;
INV     gate7617  (.A(WX10216), .Z(WX10217) ) ;
INV     gate7618  (.A(WX10056), .Z(WX10221) ) ;
OR2     gate7619  (.A(WX10220), .B(WX10219), .Z(WX10222) ) ;
INV     gate7620  (.A(WX10222), .Z(WX10223) ) ;
INV     gate7621  (.A(WX10223), .Z(WX10224) ) ;
INV     gate7622  (.A(WX10056), .Z(WX10228) ) ;
OR2     gate7623  (.A(WX10227), .B(WX10226), .Z(WX10229) ) ;
INV     gate7624  (.A(WX10229), .Z(WX10230) ) ;
INV     gate7625  (.A(WX10230), .Z(WX10231) ) ;
INV     gate7626  (.A(WX10056), .Z(WX10235) ) ;
OR2     gate7627  (.A(WX10234), .B(WX10233), .Z(WX10236) ) ;
INV     gate7628  (.A(WX10236), .Z(WX10237) ) ;
INV     gate7629  (.A(WX10237), .Z(WX10238) ) ;
INV     gate7630  (.A(WX10056), .Z(WX10242) ) ;
OR2     gate7631  (.A(WX10241), .B(WX10240), .Z(WX10243) ) ;
INV     gate7632  (.A(WX10243), .Z(WX10244) ) ;
INV     gate7633  (.A(WX10244), .Z(WX10245) ) ;
INV     gate7634  (.A(WX10056), .Z(WX10249) ) ;
OR2     gate7635  (.A(WX10248), .B(WX10247), .Z(WX10250) ) ;
INV     gate7636  (.A(WX10250), .Z(WX10251) ) ;
INV     gate7637  (.A(WX10251), .Z(WX10252) ) ;
INV     gate7638  (.A(WX10056), .Z(WX10256) ) ;
OR2     gate7639  (.A(WX10255), .B(WX10254), .Z(WX10257) ) ;
INV     gate7640  (.A(WX10257), .Z(WX10258) ) ;
INV     gate7641  (.A(WX10258), .Z(WX10259) ) ;
INV     gate7642  (.A(WX10056), .Z(WX10263) ) ;
OR2     gate7643  (.A(WX10262), .B(WX10261), .Z(WX10264) ) ;
INV     gate7644  (.A(WX10264), .Z(WX10265) ) ;
INV     gate7645  (.A(WX10265), .Z(WX10266) ) ;
INV     gate7646  (.A(WX10056), .Z(WX10270) ) ;
OR2     gate7647  (.A(WX10269), .B(WX10268), .Z(WX10271) ) ;
INV     gate7648  (.A(WX10271), .Z(WX10272) ) ;
INV     gate7649  (.A(WX10272), .Z(WX10273) ) ;
INV     gate7650  (.A(WX10056), .Z(WX10277) ) ;
OR2     gate7651  (.A(WX10276), .B(WX10275), .Z(WX10278) ) ;
INV     gate7652  (.A(WX10278), .Z(WX10279) ) ;
INV     gate7653  (.A(WX10279), .Z(WX10280) ) ;
INV     gate7654  (.A(RESET), .Z(WX10281) ) ;
INV     gate7655  (.A(WX10281), .Z(WX10314) ) ;
INV     gate7656  (.A(WX11343), .Z(WX11347) ) ;
INV     gate7657  (.A(WX11347), .Z(WX10381) ) ;
INV     gate7658  (.A(WX11341), .Z(WX11348) ) ;
INV     gate7659  (.A(WX11348), .Z(WX10385) ) ;
INV     gate7660  (.A(WX11348), .Z(WX10389) ) ;
OR2     gate7661  (.A(WX10380), .B(WX10379), .Z(WX10382) ) ;
INV     gate7662  (.A(WX10382), .Z(WX10391) ) ;
INV     gate7663  (.A(WX10391), .Z(WX10392) ) ;
INV     gate7664  (.A(WX11347), .Z(WX10395) ) ;
INV     gate7665  (.A(WX11348), .Z(WX10399) ) ;
INV     gate7666  (.A(WX11348), .Z(WX10403) ) ;
OR2     gate7667  (.A(WX10394), .B(WX10393), .Z(WX10396) ) ;
INV     gate7668  (.A(WX10396), .Z(WX10405) ) ;
INV     gate7669  (.A(WX10405), .Z(WX10406) ) ;
INV     gate7670  (.A(WX11347), .Z(WX10409) ) ;
INV     gate7671  (.A(WX11348), .Z(WX10413) ) ;
INV     gate7672  (.A(WX11348), .Z(WX10417) ) ;
OR2     gate7673  (.A(WX10408), .B(WX10407), .Z(WX10410) ) ;
INV     gate7674  (.A(WX10410), .Z(WX10419) ) ;
INV     gate7675  (.A(WX10419), .Z(WX10420) ) ;
INV     gate7676  (.A(WX11347), .Z(WX10423) ) ;
INV     gate7677  (.A(WX11348), .Z(WX10427) ) ;
INV     gate7678  (.A(WX11348), .Z(WX10431) ) ;
OR2     gate7679  (.A(WX10422), .B(WX10421), .Z(WX10424) ) ;
INV     gate7680  (.A(WX10424), .Z(WX10433) ) ;
INV     gate7681  (.A(WX10433), .Z(WX10434) ) ;
INV     gate7682  (.A(WX11347), .Z(WX10437) ) ;
INV     gate7683  (.A(WX11348), .Z(WX10441) ) ;
INV     gate7684  (.A(WX11348), .Z(WX10445) ) ;
OR2     gate7685  (.A(WX10436), .B(WX10435), .Z(WX10438) ) ;
INV     gate7686  (.A(WX10438), .Z(WX10447) ) ;
INV     gate7687  (.A(WX10447), .Z(WX10448) ) ;
INV     gate7688  (.A(WX11347), .Z(WX10451) ) ;
INV     gate7689  (.A(WX11348), .Z(WX10455) ) ;
INV     gate7690  (.A(WX11348), .Z(WX10459) ) ;
OR2     gate7691  (.A(WX10450), .B(WX10449), .Z(WX10452) ) ;
INV     gate7692  (.A(WX10452), .Z(WX10461) ) ;
INV     gate7693  (.A(WX10461), .Z(WX10462) ) ;
INV     gate7694  (.A(WX11347), .Z(WX10465) ) ;
INV     gate7695  (.A(WX11348), .Z(WX10469) ) ;
INV     gate7696  (.A(WX11348), .Z(WX10473) ) ;
OR2     gate7697  (.A(WX10464), .B(WX10463), .Z(WX10466) ) ;
INV     gate7698  (.A(WX10466), .Z(WX10475) ) ;
INV     gate7699  (.A(WX10475), .Z(WX10476) ) ;
INV     gate7700  (.A(WX11347), .Z(WX10479) ) ;
INV     gate7701  (.A(WX11348), .Z(WX10483) ) ;
INV     gate7702  (.A(WX11348), .Z(WX10487) ) ;
OR2     gate7703  (.A(WX10478), .B(WX10477), .Z(WX10480) ) ;
INV     gate7704  (.A(WX10480), .Z(WX10489) ) ;
INV     gate7705  (.A(WX10489), .Z(WX10490) ) ;
INV     gate7706  (.A(WX11347), .Z(WX10493) ) ;
INV     gate7707  (.A(WX11348), .Z(WX10497) ) ;
INV     gate7708  (.A(WX11348), .Z(WX10501) ) ;
OR2     gate7709  (.A(WX10492), .B(WX10491), .Z(WX10494) ) ;
INV     gate7710  (.A(WX10494), .Z(WX10503) ) ;
INV     gate7711  (.A(WX10503), .Z(WX10504) ) ;
INV     gate7712  (.A(WX11347), .Z(WX10507) ) ;
INV     gate7713  (.A(WX11348), .Z(WX10511) ) ;
INV     gate7714  (.A(WX11348), .Z(WX10515) ) ;
OR2     gate7715  (.A(WX10506), .B(WX10505), .Z(WX10508) ) ;
INV     gate7716  (.A(WX10508), .Z(WX10517) ) ;
INV     gate7717  (.A(WX10517), .Z(WX10518) ) ;
INV     gate7718  (.A(WX11347), .Z(WX10521) ) ;
INV     gate7719  (.A(WX11348), .Z(WX10525) ) ;
INV     gate7720  (.A(WX11348), .Z(WX10529) ) ;
OR2     gate7721  (.A(WX10520), .B(WX10519), .Z(WX10522) ) ;
INV     gate7722  (.A(WX10522), .Z(WX10531) ) ;
INV     gate7723  (.A(WX10531), .Z(WX10532) ) ;
INV     gate7724  (.A(WX11347), .Z(WX10535) ) ;
INV     gate7725  (.A(WX11348), .Z(WX10539) ) ;
INV     gate7726  (.A(WX11348), .Z(WX10543) ) ;
OR2     gate7727  (.A(WX10534), .B(WX10533), .Z(WX10536) ) ;
INV     gate7728  (.A(WX10536), .Z(WX10545) ) ;
INV     gate7729  (.A(WX10545), .Z(WX10546) ) ;
INV     gate7730  (.A(WX11347), .Z(WX10549) ) ;
INV     gate7731  (.A(WX11348), .Z(WX10553) ) ;
INV     gate7732  (.A(WX11348), .Z(WX10557) ) ;
OR2     gate7733  (.A(WX10548), .B(WX10547), .Z(WX10550) ) ;
INV     gate7734  (.A(WX10550), .Z(WX10559) ) ;
INV     gate7735  (.A(WX10559), .Z(WX10560) ) ;
INV     gate7736  (.A(WX11347), .Z(WX10563) ) ;
INV     gate7737  (.A(WX11348), .Z(WX10567) ) ;
INV     gate7738  (.A(WX11348), .Z(WX10571) ) ;
OR2     gate7739  (.A(WX10562), .B(WX10561), .Z(WX10564) ) ;
INV     gate7740  (.A(WX10564), .Z(WX10573) ) ;
INV     gate7741  (.A(WX10573), .Z(WX10574) ) ;
INV     gate7742  (.A(WX11347), .Z(WX10577) ) ;
INV     gate7743  (.A(WX11348), .Z(WX10581) ) ;
INV     gate7744  (.A(WX11348), .Z(WX10585) ) ;
OR2     gate7745  (.A(WX10576), .B(WX10575), .Z(WX10578) ) ;
INV     gate7746  (.A(WX10578), .Z(WX10587) ) ;
INV     gate7747  (.A(WX10587), .Z(WX10588) ) ;
INV     gate7748  (.A(WX11347), .Z(WX10591) ) ;
INV     gate7749  (.A(WX11348), .Z(WX10595) ) ;
INV     gate7750  (.A(WX11348), .Z(WX10599) ) ;
OR2     gate7751  (.A(WX10590), .B(WX10589), .Z(WX10592) ) ;
INV     gate7752  (.A(WX10592), .Z(WX10601) ) ;
INV     gate7753  (.A(WX10601), .Z(WX10602) ) ;
INV     gate7754  (.A(WX11347), .Z(WX10605) ) ;
INV     gate7755  (.A(WX11348), .Z(WX10609) ) ;
INV     gate7756  (.A(WX11348), .Z(WX10613) ) ;
OR2     gate7757  (.A(WX10604), .B(WX10603), .Z(WX10606) ) ;
INV     gate7758  (.A(WX10606), .Z(WX10615) ) ;
INV     gate7759  (.A(WX10615), .Z(WX10616) ) ;
INV     gate7760  (.A(WX11347), .Z(WX10619) ) ;
INV     gate7761  (.A(WX11348), .Z(WX10623) ) ;
INV     gate7762  (.A(WX11348), .Z(WX10627) ) ;
OR2     gate7763  (.A(WX10618), .B(WX10617), .Z(WX10620) ) ;
INV     gate7764  (.A(WX10620), .Z(WX10629) ) ;
INV     gate7765  (.A(WX10629), .Z(WX10630) ) ;
INV     gate7766  (.A(WX11347), .Z(WX10633) ) ;
INV     gate7767  (.A(WX11348), .Z(WX10637) ) ;
INV     gate7768  (.A(WX11348), .Z(WX10641) ) ;
OR2     gate7769  (.A(WX10632), .B(WX10631), .Z(WX10634) ) ;
INV     gate7770  (.A(WX10634), .Z(WX10643) ) ;
INV     gate7771  (.A(WX10643), .Z(WX10644) ) ;
INV     gate7772  (.A(WX11347), .Z(WX10647) ) ;
INV     gate7773  (.A(WX11348), .Z(WX10651) ) ;
INV     gate7774  (.A(WX11348), .Z(WX10655) ) ;
OR2     gate7775  (.A(WX10646), .B(WX10645), .Z(WX10648) ) ;
INV     gate7776  (.A(WX10648), .Z(WX10657) ) ;
INV     gate7777  (.A(WX10657), .Z(WX10658) ) ;
INV     gate7778  (.A(WX11347), .Z(WX10661) ) ;
INV     gate7779  (.A(WX11348), .Z(WX10665) ) ;
INV     gate7780  (.A(WX11348), .Z(WX10669) ) ;
OR2     gate7781  (.A(WX10660), .B(WX10659), .Z(WX10662) ) ;
INV     gate7782  (.A(WX10662), .Z(WX10671) ) ;
INV     gate7783  (.A(WX10671), .Z(WX10672) ) ;
INV     gate7784  (.A(WX11347), .Z(WX10675) ) ;
INV     gate7785  (.A(WX11348), .Z(WX10679) ) ;
INV     gate7786  (.A(WX11348), .Z(WX10683) ) ;
OR2     gate7787  (.A(WX10674), .B(WX10673), .Z(WX10676) ) ;
INV     gate7788  (.A(WX10676), .Z(WX10685) ) ;
INV     gate7789  (.A(WX10685), .Z(WX10686) ) ;
INV     gate7790  (.A(WX11347), .Z(WX10689) ) ;
INV     gate7791  (.A(WX11348), .Z(WX10693) ) ;
INV     gate7792  (.A(WX11348), .Z(WX10697) ) ;
OR2     gate7793  (.A(WX10688), .B(WX10687), .Z(WX10690) ) ;
INV     gate7794  (.A(WX10690), .Z(WX10699) ) ;
INV     gate7795  (.A(WX10699), .Z(WX10700) ) ;
INV     gate7796  (.A(WX11347), .Z(WX10703) ) ;
INV     gate7797  (.A(WX11348), .Z(WX10707) ) ;
INV     gate7798  (.A(WX11348), .Z(WX10711) ) ;
OR2     gate7799  (.A(WX10702), .B(WX10701), .Z(WX10704) ) ;
INV     gate7800  (.A(WX10704), .Z(WX10713) ) ;
INV     gate7801  (.A(WX10713), .Z(WX10714) ) ;
INV     gate7802  (.A(WX11347), .Z(WX10717) ) ;
INV     gate7803  (.A(WX11348), .Z(WX10721) ) ;
INV     gate7804  (.A(WX11348), .Z(WX10725) ) ;
OR2     gate7805  (.A(WX10716), .B(WX10715), .Z(WX10718) ) ;
INV     gate7806  (.A(WX10718), .Z(WX10727) ) ;
INV     gate7807  (.A(WX10727), .Z(WX10728) ) ;
INV     gate7808  (.A(WX11347), .Z(WX10731) ) ;
INV     gate7809  (.A(WX11348), .Z(WX10735) ) ;
INV     gate7810  (.A(WX11348), .Z(WX10739) ) ;
OR2     gate7811  (.A(WX10730), .B(WX10729), .Z(WX10732) ) ;
INV     gate7812  (.A(WX10732), .Z(WX10741) ) ;
INV     gate7813  (.A(WX10741), .Z(WX10742) ) ;
INV     gate7814  (.A(WX11347), .Z(WX10745) ) ;
INV     gate7815  (.A(WX11348), .Z(WX10749) ) ;
INV     gate7816  (.A(WX11348), .Z(WX10753) ) ;
OR2     gate7817  (.A(WX10744), .B(WX10743), .Z(WX10746) ) ;
INV     gate7818  (.A(WX10746), .Z(WX10755) ) ;
INV     gate7819  (.A(WX10755), .Z(WX10756) ) ;
INV     gate7820  (.A(WX11347), .Z(WX10759) ) ;
INV     gate7821  (.A(WX11348), .Z(WX10763) ) ;
INV     gate7822  (.A(WX11348), .Z(WX10767) ) ;
OR2     gate7823  (.A(WX10758), .B(WX10757), .Z(WX10760) ) ;
INV     gate7824  (.A(WX10760), .Z(WX10769) ) ;
INV     gate7825  (.A(WX10769), .Z(WX10770) ) ;
INV     gate7826  (.A(WX11347), .Z(WX10773) ) ;
INV     gate7827  (.A(WX11348), .Z(WX10777) ) ;
INV     gate7828  (.A(WX11348), .Z(WX10781) ) ;
OR2     gate7829  (.A(WX10772), .B(WX10771), .Z(WX10774) ) ;
INV     gate7830  (.A(WX10774), .Z(WX10783) ) ;
INV     gate7831  (.A(WX10783), .Z(WX10784) ) ;
INV     gate7832  (.A(WX11347), .Z(WX10787) ) ;
INV     gate7833  (.A(WX11348), .Z(WX10791) ) ;
INV     gate7834  (.A(WX11348), .Z(WX10795) ) ;
OR2     gate7835  (.A(WX10786), .B(WX10785), .Z(WX10788) ) ;
INV     gate7836  (.A(WX10788), .Z(WX10797) ) ;
INV     gate7837  (.A(WX10797), .Z(WX10798) ) ;
INV     gate7838  (.A(WX11347), .Z(WX10801) ) ;
INV     gate7839  (.A(WX11348), .Z(WX10805) ) ;
INV     gate7840  (.A(WX11348), .Z(WX10809) ) ;
OR2     gate7841  (.A(WX10800), .B(WX10799), .Z(WX10802) ) ;
INV     gate7842  (.A(WX10802), .Z(WX10811) ) ;
INV     gate7843  (.A(WX10811), .Z(WX10812) ) ;
INV     gate7844  (.A(WX11347), .Z(WX10815) ) ;
INV     gate7845  (.A(WX11348), .Z(WX10819) ) ;
INV     gate7846  (.A(WX11348), .Z(WX10823) ) ;
OR2     gate7847  (.A(WX10814), .B(WX10813), .Z(WX10816) ) ;
INV     gate7848  (.A(WX10816), .Z(WX10825) ) ;
INV     gate7849  (.A(WX10825), .Z(WX10826) ) ;
INV     gate7850  (.A(WX10829), .Z(WX10827) ) ;
INV     gate7851  (.A(WX11308), .Z(WX11309) ) ;
INV     gate7852  (.A(WX11309), .Z(WX10892) ) ;
INV     gate7853  (.A(WX11310), .Z(WX11311) ) ;
INV     gate7854  (.A(WX11311), .Z(WX10893) ) ;
INV     gate7855  (.A(WX11312), .Z(WX11313) ) ;
INV     gate7856  (.A(WX11313), .Z(WX10894) ) ;
INV     gate7857  (.A(WX11314), .Z(WX11315) ) ;
INV     gate7858  (.A(WX11315), .Z(WX10895) ) ;
INV     gate7859  (.A(WX11316), .Z(WX11317) ) ;
INV     gate7860  (.A(WX11317), .Z(WX10896) ) ;
INV     gate7861  (.A(WX11318), .Z(WX11319) ) ;
INV     gate7862  (.A(WX11319), .Z(WX10897) ) ;
INV     gate7863  (.A(WX11320), .Z(WX11321) ) ;
INV     gate7864  (.A(WX11321), .Z(WX10898) ) ;
INV     gate7865  (.A(WX11322), .Z(WX11323) ) ;
INV     gate7866  (.A(WX11323), .Z(WX10899) ) ;
INV     gate7867  (.A(WX11324), .Z(WX11325) ) ;
INV     gate7868  (.A(WX11325), .Z(WX10900) ) ;
INV     gate7869  (.A(WX11326), .Z(WX11327) ) ;
INV     gate7870  (.A(WX11327), .Z(WX10901) ) ;
INV     gate7871  (.A(WX11328), .Z(WX11329) ) ;
INV     gate7872  (.A(WX11329), .Z(WX10902) ) ;
INV     gate7873  (.A(WX11330), .Z(WX11331) ) ;
INV     gate7874  (.A(WX11331), .Z(WX10903) ) ;
INV     gate7875  (.A(WX11332), .Z(WX11333) ) ;
INV     gate7876  (.A(WX11333), .Z(WX10904) ) ;
INV     gate7877  (.A(WX11334), .Z(WX11335) ) ;
INV     gate7878  (.A(WX11335), .Z(WX10905) ) ;
INV     gate7879  (.A(WX11336), .Z(WX11337) ) ;
INV     gate7880  (.A(WX11337), .Z(WX10906) ) ;
INV     gate7881  (.A(WX11338), .Z(WX11339) ) ;
INV     gate7882  (.A(WX11339), .Z(WX10907) ) ;
INV     gate7883  (.A(WX11276), .Z(WX11277) ) ;
INV     gate7884  (.A(WX11277), .Z(WX10908) ) ;
INV     gate7885  (.A(WX11278), .Z(WX11279) ) ;
INV     gate7886  (.A(WX11279), .Z(WX10909) ) ;
INV     gate7887  (.A(WX11280), .Z(WX11281) ) ;
INV     gate7888  (.A(WX11281), .Z(WX10910) ) ;
INV     gate7889  (.A(WX11282), .Z(WX11283) ) ;
INV     gate7890  (.A(WX11283), .Z(WX10911) ) ;
INV     gate7891  (.A(WX11284), .Z(WX11285) ) ;
INV     gate7892  (.A(WX11285), .Z(WX10912) ) ;
INV     gate7893  (.A(WX11286), .Z(WX11287) ) ;
INV     gate7894  (.A(WX11287), .Z(WX10913) ) ;
INV     gate7895  (.A(WX11288), .Z(WX11289) ) ;
INV     gate7896  (.A(WX11289), .Z(WX10914) ) ;
INV     gate7897  (.A(WX11290), .Z(WX11291) ) ;
INV     gate7898  (.A(WX11291), .Z(WX10915) ) ;
INV     gate7899  (.A(WX11292), .Z(WX11293) ) ;
INV     gate7900  (.A(WX11293), .Z(WX10916) ) ;
INV     gate7901  (.A(WX11294), .Z(WX11295) ) ;
INV     gate7902  (.A(WX11295), .Z(WX10917) ) ;
INV     gate7903  (.A(WX11296), .Z(WX11297) ) ;
INV     gate7904  (.A(WX11297), .Z(WX10918) ) ;
INV     gate7905  (.A(WX11298), .Z(WX11299) ) ;
INV     gate7906  (.A(WX11299), .Z(WX10919) ) ;
INV     gate7907  (.A(WX11300), .Z(WX11301) ) ;
INV     gate7908  (.A(WX11301), .Z(WX10920) ) ;
INV     gate7909  (.A(WX11302), .Z(WX11303) ) ;
INV     gate7910  (.A(WX11303), .Z(WX10921) ) ;
INV     gate7911  (.A(WX11304), .Z(WX11305) ) ;
INV     gate7912  (.A(WX11305), .Z(WX10922) ) ;
INV     gate7913  (.A(WX11306), .Z(WX11307) ) ;
INV     gate7914  (.A(WX11307), .Z(WX10923) ) ;
INV     gate7915  (.A(WX10892), .Z(WX10924) ) ;
INV     gate7916  (.A(WX10893), .Z(WX10925) ) ;
INV     gate7917  (.A(WX10894), .Z(WX10926) ) ;
INV     gate7918  (.A(WX10895), .Z(WX10927) ) ;
INV     gate7919  (.A(WX10896), .Z(WX10928) ) ;
INV     gate7920  (.A(WX10897), .Z(WX10929) ) ;
INV     gate7921  (.A(WX10898), .Z(WX10930) ) ;
INV     gate7922  (.A(WX10899), .Z(WX10931) ) ;
INV     gate7923  (.A(WX10900), .Z(WX10932) ) ;
INV     gate7924  (.A(WX10901), .Z(WX10933) ) ;
INV     gate7925  (.A(WX10902), .Z(WX10934) ) ;
INV     gate7926  (.A(WX10903), .Z(WX10935) ) ;
INV     gate7927  (.A(WX10904), .Z(WX10936) ) ;
INV     gate7928  (.A(WX10905), .Z(WX10937) ) ;
INV     gate7929  (.A(WX10906), .Z(WX10938) ) ;
INV     gate7930  (.A(WX10907), .Z(WX10939) ) ;
INV     gate7931  (.A(WX10908), .Z(WX10940) ) ;
INV     gate7932  (.A(WX10909), .Z(WX10941) ) ;
INV     gate7933  (.A(WX10910), .Z(WX10942) ) ;
INV     gate7934  (.A(WX10911), .Z(WX10943) ) ;
INV     gate7935  (.A(WX10912), .Z(WX10944) ) ;
INV     gate7936  (.A(WX10913), .Z(WX10945) ) ;
INV     gate7937  (.A(WX10914), .Z(WX10946) ) ;
INV     gate7938  (.A(WX10915), .Z(WX10947) ) ;
INV     gate7939  (.A(WX10916), .Z(WX10948) ) ;
INV     gate7940  (.A(WX10917), .Z(WX10949) ) ;
INV     gate7941  (.A(WX10918), .Z(WX10950) ) ;
INV     gate7942  (.A(WX10919), .Z(WX10951) ) ;
INV     gate7943  (.A(WX10920), .Z(WX10952) ) ;
INV     gate7944  (.A(WX10921), .Z(WX10953) ) ;
INV     gate7945  (.A(WX10922), .Z(WX10954) ) ;
INV     gate7946  (.A(WX10923), .Z(WX10955) ) ;
INV     gate7947  (.A(WX11181), .Z(WX10956) ) ;
INV     gate7948  (.A(WX11183), .Z(WX10957) ) ;
INV     gate7949  (.A(WX11185), .Z(WX10958) ) ;
INV     gate7950  (.A(WX11187), .Z(WX10959) ) ;
INV     gate7951  (.A(WX11189), .Z(WX10960) ) ;
INV     gate7952  (.A(WX11191), .Z(WX10961) ) ;
INV     gate7953  (.A(WX11193), .Z(WX10962) ) ;
INV     gate7954  (.A(WX11195), .Z(WX10963) ) ;
INV     gate7955  (.A(WX11197), .Z(WX10964) ) ;
INV     gate7956  (.A(WX11199), .Z(WX10965) ) ;
INV     gate7957  (.A(WX11201), .Z(WX10966) ) ;
INV     gate7958  (.A(WX11203), .Z(WX10967) ) ;
INV     gate7959  (.A(WX11205), .Z(WX10968) ) ;
INV     gate7960  (.A(WX11207), .Z(WX10969) ) ;
INV     gate7961  (.A(WX11209), .Z(WX10970) ) ;
INV     gate7962  (.A(WX11211), .Z(WX10971) ) ;
INV     gate7963  (.A(WX11213), .Z(WX10972) ) ;
INV     gate7964  (.A(WX11215), .Z(WX10973) ) ;
INV     gate7965  (.A(WX11217), .Z(WX10974) ) ;
INV     gate7966  (.A(WX11219), .Z(WX10975) ) ;
INV     gate7967  (.A(WX11221), .Z(WX10976) ) ;
INV     gate7968  (.A(WX11223), .Z(WX10977) ) ;
INV     gate7969  (.A(WX11225), .Z(WX10978) ) ;
INV     gate7970  (.A(WX11227), .Z(WX10979) ) ;
INV     gate7971  (.A(WX11229), .Z(WX10980) ) ;
INV     gate7972  (.A(WX11231), .Z(WX10981) ) ;
INV     gate7973  (.A(WX11233), .Z(WX10982) ) ;
INV     gate7974  (.A(WX11235), .Z(WX10983) ) ;
INV     gate7975  (.A(WX11237), .Z(WX10984) ) ;
INV     gate7976  (.A(WX11239), .Z(WX10985) ) ;
INV     gate7977  (.A(WX11241), .Z(WX10986) ) ;
INV     gate7978  (.A(WX11243), .Z(WX10987) ) ;
NAND2   gate7979  (.A(II34547), .B(II34548), .Z(WX11260) ) ;
INV     gate7980  (.A(WX11260), .Z(WX11276) ) ;
NAND2   gate7981  (.A(II34578), .B(II34579), .Z(WX11261) ) ;
INV     gate7982  (.A(WX11261), .Z(WX11278) ) ;
NAND2   gate7983  (.A(II34609), .B(II34610), .Z(WX11262) ) ;
INV     gate7984  (.A(WX11262), .Z(WX11280) ) ;
NAND2   gate7985  (.A(II34640), .B(II34641), .Z(WX11263) ) ;
INV     gate7986  (.A(WX11263), .Z(WX11282) ) ;
NAND2   gate7987  (.A(II34671), .B(II34672), .Z(WX11264) ) ;
INV     gate7988  (.A(WX11264), .Z(WX11284) ) ;
NAND2   gate7989  (.A(II34702), .B(II34703), .Z(WX11265) ) ;
INV     gate7990  (.A(WX11265), .Z(WX11286) ) ;
NAND2   gate7991  (.A(II34733), .B(II34734), .Z(WX11266) ) ;
INV     gate7992  (.A(WX11266), .Z(WX11288) ) ;
NAND2   gate7993  (.A(II34764), .B(II34765), .Z(WX11267) ) ;
INV     gate7994  (.A(WX11267), .Z(WX11290) ) ;
NAND2   gate7995  (.A(II34795), .B(II34796), .Z(WX11268) ) ;
INV     gate7996  (.A(WX11268), .Z(WX11292) ) ;
NAND2   gate7997  (.A(II34826), .B(II34827), .Z(WX11269) ) ;
INV     gate7998  (.A(WX11269), .Z(WX11294) ) ;
NAND2   gate7999  (.A(II34857), .B(II34858), .Z(WX11270) ) ;
INV     gate8000  (.A(WX11270), .Z(WX11296) ) ;
NAND2   gate8001  (.A(II34888), .B(II34889), .Z(WX11271) ) ;
INV     gate8002  (.A(WX11271), .Z(WX11298) ) ;
NAND2   gate8003  (.A(II34919), .B(II34920), .Z(WX11272) ) ;
INV     gate8004  (.A(WX11272), .Z(WX11300) ) ;
NAND2   gate8005  (.A(II34950), .B(II34951), .Z(WX11273) ) ;
INV     gate8006  (.A(WX11273), .Z(WX11302) ) ;
NAND2   gate8007  (.A(II34981), .B(II34982), .Z(WX11274) ) ;
INV     gate8008  (.A(WX11274), .Z(WX11304) ) ;
NAND2   gate8009  (.A(II35012), .B(II35013), .Z(WX11275) ) ;
INV     gate8010  (.A(WX11275), .Z(WX11306) ) ;
NAND2   gate8011  (.A(II34051), .B(II34052), .Z(WX11244) ) ;
INV     gate8012  (.A(WX11244), .Z(WX11308) ) ;
NAND2   gate8013  (.A(II34082), .B(II34083), .Z(WX11245) ) ;
INV     gate8014  (.A(WX11245), .Z(WX11310) ) ;
NAND2   gate8015  (.A(II34113), .B(II34114), .Z(WX11246) ) ;
INV     gate8016  (.A(WX11246), .Z(WX11312) ) ;
NAND2   gate8017  (.A(II34144), .B(II34145), .Z(WX11247) ) ;
INV     gate8018  (.A(WX11247), .Z(WX11314) ) ;
NAND2   gate8019  (.A(II34175), .B(II34176), .Z(WX11248) ) ;
INV     gate8020  (.A(WX11248), .Z(WX11316) ) ;
NAND2   gate8021  (.A(II34206), .B(II34207), .Z(WX11249) ) ;
INV     gate8022  (.A(WX11249), .Z(WX11318) ) ;
NAND2   gate8023  (.A(II34237), .B(II34238), .Z(WX11250) ) ;
INV     gate8024  (.A(WX11250), .Z(WX11320) ) ;
NAND2   gate8025  (.A(II34268), .B(II34269), .Z(WX11251) ) ;
INV     gate8026  (.A(WX11251), .Z(WX11322) ) ;
NAND2   gate8027  (.A(II34299), .B(II34300), .Z(WX11252) ) ;
INV     gate8028  (.A(WX11252), .Z(WX11324) ) ;
NAND2   gate8029  (.A(II34330), .B(II34331), .Z(WX11253) ) ;
INV     gate8030  (.A(WX11253), .Z(WX11326) ) ;
NAND2   gate8031  (.A(II34361), .B(II34362), .Z(WX11254) ) ;
INV     gate8032  (.A(WX11254), .Z(WX11328) ) ;
NAND2   gate8033  (.A(II34392), .B(II34393), .Z(WX11255) ) ;
INV     gate8034  (.A(WX11255), .Z(WX11330) ) ;
NAND2   gate8035  (.A(II34423), .B(II34424), .Z(WX11256) ) ;
INV     gate8036  (.A(WX11256), .Z(WX11332) ) ;
NAND2   gate8037  (.A(II34454), .B(II34455), .Z(WX11257) ) ;
INV     gate8038  (.A(WX11257), .Z(WX11334) ) ;
NAND2   gate8039  (.A(II34485), .B(II34486), .Z(WX11258) ) ;
INV     gate8040  (.A(WX11258), .Z(WX11336) ) ;
NAND2   gate8041  (.A(II34516), .B(II34517), .Z(WX11259) ) ;
INV     gate8042  (.A(WX11259), .Z(WX11338) ) ;
INV     gate8043  (.A(TM0), .Z(WX11340) ) ;
INV     gate8044  (.A(TM0), .Z(WX11341) ) ;
INV     gate8045  (.A(TM0), .Z(WX11342) ) ;
INV     gate8046  (.A(TM1), .Z(WX11343) ) ;
INV     gate8047  (.A(TM1), .Z(WX11344) ) ;
INV     gate8048  (.A(WX11344), .Z(WX11345) ) ;
INV     gate8049  (.A(WX11342), .Z(WX11346) ) ;
INV     gate8050  (.A(WX11340), .Z(WX11349) ) ;
INV     gate8051  (.A(WX11349), .Z(WX11353) ) ;
OR2     gate8052  (.A(WX11352), .B(WX11351), .Z(WX11354) ) ;
INV     gate8053  (.A(WX11354), .Z(WX11355) ) ;
INV     gate8054  (.A(WX11355), .Z(WX11356) ) ;
INV     gate8055  (.A(WX11349), .Z(WX11360) ) ;
OR2     gate8056  (.A(WX11359), .B(WX11358), .Z(WX11361) ) ;
INV     gate8057  (.A(WX11361), .Z(WX11362) ) ;
INV     gate8058  (.A(WX11362), .Z(WX11363) ) ;
INV     gate8059  (.A(WX11349), .Z(WX11367) ) ;
OR2     gate8060  (.A(WX11366), .B(WX11365), .Z(WX11368) ) ;
INV     gate8061  (.A(WX11368), .Z(WX11369) ) ;
INV     gate8062  (.A(WX11369), .Z(WX11370) ) ;
INV     gate8063  (.A(WX11349), .Z(WX11374) ) ;
OR2     gate8064  (.A(WX11373), .B(WX11372), .Z(WX11375) ) ;
INV     gate8065  (.A(WX11375), .Z(WX11376) ) ;
INV     gate8066  (.A(WX11376), .Z(WX11377) ) ;
INV     gate8067  (.A(WX11349), .Z(WX11381) ) ;
OR2     gate8068  (.A(WX11380), .B(WX11379), .Z(WX11382) ) ;
INV     gate8069  (.A(WX11382), .Z(WX11383) ) ;
INV     gate8070  (.A(WX11383), .Z(WX11384) ) ;
INV     gate8071  (.A(WX11349), .Z(WX11388) ) ;
OR2     gate8072  (.A(WX11387), .B(WX11386), .Z(WX11389) ) ;
INV     gate8073  (.A(WX11389), .Z(WX11390) ) ;
INV     gate8074  (.A(WX11390), .Z(WX11391) ) ;
INV     gate8075  (.A(WX11349), .Z(WX11395) ) ;
OR2     gate8076  (.A(WX11394), .B(WX11393), .Z(WX11396) ) ;
INV     gate8077  (.A(WX11396), .Z(WX11397) ) ;
INV     gate8078  (.A(WX11397), .Z(WX11398) ) ;
INV     gate8079  (.A(WX11349), .Z(WX11402) ) ;
OR2     gate8080  (.A(WX11401), .B(WX11400), .Z(WX11403) ) ;
INV     gate8081  (.A(WX11403), .Z(WX11404) ) ;
INV     gate8082  (.A(WX11404), .Z(WX11405) ) ;
INV     gate8083  (.A(WX11349), .Z(WX11409) ) ;
OR2     gate8084  (.A(WX11408), .B(WX11407), .Z(WX11410) ) ;
INV     gate8085  (.A(WX11410), .Z(WX11411) ) ;
INV     gate8086  (.A(WX11411), .Z(WX11412) ) ;
INV     gate8087  (.A(WX11349), .Z(WX11416) ) ;
OR2     gate8088  (.A(WX11415), .B(WX11414), .Z(WX11417) ) ;
INV     gate8089  (.A(WX11417), .Z(WX11418) ) ;
INV     gate8090  (.A(WX11418), .Z(WX11419) ) ;
INV     gate8091  (.A(WX11349), .Z(WX11423) ) ;
OR2     gate8092  (.A(WX11422), .B(WX11421), .Z(WX11424) ) ;
INV     gate8093  (.A(WX11424), .Z(WX11425) ) ;
INV     gate8094  (.A(WX11425), .Z(WX11426) ) ;
INV     gate8095  (.A(WX11349), .Z(WX11430) ) ;
OR2     gate8096  (.A(WX11429), .B(WX11428), .Z(WX11431) ) ;
INV     gate8097  (.A(WX11431), .Z(WX11432) ) ;
INV     gate8098  (.A(WX11432), .Z(WX11433) ) ;
INV     gate8099  (.A(WX11349), .Z(WX11437) ) ;
OR2     gate8100  (.A(WX11436), .B(WX11435), .Z(WX11438) ) ;
INV     gate8101  (.A(WX11438), .Z(WX11439) ) ;
INV     gate8102  (.A(WX11439), .Z(WX11440) ) ;
INV     gate8103  (.A(WX11349), .Z(WX11444) ) ;
OR2     gate8104  (.A(WX11443), .B(WX11442), .Z(WX11445) ) ;
INV     gate8105  (.A(WX11445), .Z(WX11446) ) ;
INV     gate8106  (.A(WX11446), .Z(WX11447) ) ;
INV     gate8107  (.A(WX11349), .Z(WX11451) ) ;
OR2     gate8108  (.A(WX11450), .B(WX11449), .Z(WX11452) ) ;
INV     gate8109  (.A(WX11452), .Z(WX11453) ) ;
INV     gate8110  (.A(WX11453), .Z(WX11454) ) ;
INV     gate8111  (.A(WX11349), .Z(WX11458) ) ;
OR2     gate8112  (.A(WX11457), .B(WX11456), .Z(WX11459) ) ;
INV     gate8113  (.A(WX11459), .Z(WX11460) ) ;
INV     gate8114  (.A(WX11460), .Z(WX11461) ) ;
INV     gate8115  (.A(WX11349), .Z(WX11465) ) ;
OR2     gate8116  (.A(WX11464), .B(WX11463), .Z(WX11466) ) ;
INV     gate8117  (.A(WX11466), .Z(WX11467) ) ;
INV     gate8118  (.A(WX11467), .Z(WX11468) ) ;
INV     gate8119  (.A(WX11349), .Z(WX11472) ) ;
OR2     gate8120  (.A(WX11471), .B(WX11470), .Z(WX11473) ) ;
INV     gate8121  (.A(WX11473), .Z(WX11474) ) ;
INV     gate8122  (.A(WX11474), .Z(WX11475) ) ;
INV     gate8123  (.A(WX11349), .Z(WX11479) ) ;
OR2     gate8124  (.A(WX11478), .B(WX11477), .Z(WX11480) ) ;
INV     gate8125  (.A(WX11480), .Z(WX11481) ) ;
INV     gate8126  (.A(WX11481), .Z(WX11482) ) ;
INV     gate8127  (.A(WX11349), .Z(WX11486) ) ;
OR2     gate8128  (.A(WX11485), .B(WX11484), .Z(WX11487) ) ;
INV     gate8129  (.A(WX11487), .Z(WX11488) ) ;
INV     gate8130  (.A(WX11488), .Z(WX11489) ) ;
INV     gate8131  (.A(WX11349), .Z(WX11493) ) ;
OR2     gate8132  (.A(WX11492), .B(WX11491), .Z(WX11494) ) ;
INV     gate8133  (.A(WX11494), .Z(WX11495) ) ;
INV     gate8134  (.A(WX11495), .Z(WX11496) ) ;
INV     gate8135  (.A(WX11349), .Z(WX11500) ) ;
OR2     gate8136  (.A(WX11499), .B(WX11498), .Z(WX11501) ) ;
INV     gate8137  (.A(WX11501), .Z(WX11502) ) ;
INV     gate8138  (.A(WX11502), .Z(WX11503) ) ;
INV     gate8139  (.A(WX11349), .Z(WX11507) ) ;
OR2     gate8140  (.A(WX11506), .B(WX11505), .Z(WX11508) ) ;
INV     gate8141  (.A(WX11508), .Z(WX11509) ) ;
INV     gate8142  (.A(WX11509), .Z(WX11510) ) ;
INV     gate8143  (.A(WX11349), .Z(WX11514) ) ;
OR2     gate8144  (.A(WX11513), .B(WX11512), .Z(WX11515) ) ;
INV     gate8145  (.A(WX11515), .Z(WX11516) ) ;
INV     gate8146  (.A(WX11516), .Z(WX11517) ) ;
INV     gate8147  (.A(WX11349), .Z(WX11521) ) ;
OR2     gate8148  (.A(WX11520), .B(WX11519), .Z(WX11522) ) ;
INV     gate8149  (.A(WX11522), .Z(WX11523) ) ;
INV     gate8150  (.A(WX11523), .Z(WX11524) ) ;
INV     gate8151  (.A(WX11349), .Z(WX11528) ) ;
OR2     gate8152  (.A(WX11527), .B(WX11526), .Z(WX11529) ) ;
INV     gate8153  (.A(WX11529), .Z(WX11530) ) ;
INV     gate8154  (.A(WX11530), .Z(WX11531) ) ;
INV     gate8155  (.A(WX11349), .Z(WX11535) ) ;
OR2     gate8156  (.A(WX11534), .B(WX11533), .Z(WX11536) ) ;
INV     gate8157  (.A(WX11536), .Z(WX11537) ) ;
INV     gate8158  (.A(WX11537), .Z(WX11538) ) ;
INV     gate8159  (.A(WX11349), .Z(WX11542) ) ;
OR2     gate8160  (.A(WX11541), .B(WX11540), .Z(WX11543) ) ;
INV     gate8161  (.A(WX11543), .Z(WX11544) ) ;
INV     gate8162  (.A(WX11544), .Z(WX11545) ) ;
INV     gate8163  (.A(WX11349), .Z(WX11549) ) ;
OR2     gate8164  (.A(WX11548), .B(WX11547), .Z(WX11550) ) ;
INV     gate8165  (.A(WX11550), .Z(WX11551) ) ;
INV     gate8166  (.A(WX11551), .Z(WX11552) ) ;
INV     gate8167  (.A(WX11349), .Z(WX11556) ) ;
OR2     gate8168  (.A(WX11555), .B(WX11554), .Z(WX11557) ) ;
INV     gate8169  (.A(WX11557), .Z(WX11558) ) ;
INV     gate8170  (.A(WX11558), .Z(WX11559) ) ;
INV     gate8171  (.A(WX11349), .Z(WX11563) ) ;
OR2     gate8172  (.A(WX11562), .B(WX11561), .Z(WX11564) ) ;
INV     gate8173  (.A(WX11564), .Z(WX11565) ) ;
INV     gate8174  (.A(WX11565), .Z(WX11566) ) ;
INV     gate8175  (.A(WX11349), .Z(WX11570) ) ;
OR2     gate8176  (.A(WX11569), .B(WX11568), .Z(WX11571) ) ;
INV     gate8177  (.A(WX11571), .Z(WX11572) ) ;
INV     gate8178  (.A(WX11572), .Z(WX11573) ) ;
INV     gate8179  (.A(RESET), .Z(WX11574) ) ;
INV     gate8180  (.A(WX11574), .Z(WX11607) ) ;
OR2     gate8181  (.A(WX44), .B(WX43), .Z(WX46) ) ;
AND2    gate8182  (.A(WX46), .B(WX1003), .Z(WX35) ) ;
OR2     gate8183  (.A(WX40), .B(WX39), .Z(WX42) ) ;
AND2    gate8184  (.A(WX42), .B(WX37), .Z(WX36) ) ;
AND2    gate8185  (.A(CRC_OUT_9_31), .B(WX1004), .Z(WX39) ) ;
AND2    gate8186  (.A(WX2305), .B(WX41), .Z(WX40) ) ;
AND2    gate8187  (.A(WX485), .B(WX1004), .Z(WX43) ) ;
AND2    gate8188  (.A(DATA_9_31), .B(WX45), .Z(WX44) ) ;
OR2     gate8189  (.A(WX58), .B(WX57), .Z(WX60) ) ;
AND2    gate8190  (.A(WX60), .B(WX1003), .Z(WX49) ) ;
OR2     gate8191  (.A(WX54), .B(WX53), .Z(WX56) ) ;
AND2    gate8192  (.A(WX56), .B(WX51), .Z(WX50) ) ;
AND2    gate8193  (.A(CRC_OUT_9_30), .B(WX1004), .Z(WX53) ) ;
AND2    gate8194  (.A(WX2312), .B(WX55), .Z(WX54) ) ;
AND2    gate8195  (.A(WX487), .B(WX1004), .Z(WX57) ) ;
AND2    gate8196  (.A(DATA_9_30), .B(WX59), .Z(WX58) ) ;
OR2     gate8197  (.A(WX72), .B(WX71), .Z(WX74) ) ;
AND2    gate8198  (.A(WX74), .B(WX1003), .Z(WX63) ) ;
OR2     gate8199  (.A(WX68), .B(WX67), .Z(WX70) ) ;
AND2    gate8200  (.A(WX70), .B(WX65), .Z(WX64) ) ;
AND2    gate8201  (.A(CRC_OUT_9_29), .B(WX1004), .Z(WX67) ) ;
AND2    gate8202  (.A(WX2319), .B(WX69), .Z(WX68) ) ;
AND2    gate8203  (.A(WX489), .B(WX1004), .Z(WX71) ) ;
AND2    gate8204  (.A(DATA_9_29), .B(WX73), .Z(WX72) ) ;
OR2     gate8205  (.A(WX86), .B(WX85), .Z(WX88) ) ;
AND2    gate8206  (.A(WX88), .B(WX1003), .Z(WX77) ) ;
OR2     gate8207  (.A(WX82), .B(WX81), .Z(WX84) ) ;
AND2    gate8208  (.A(WX84), .B(WX79), .Z(WX78) ) ;
AND2    gate8209  (.A(CRC_OUT_9_28), .B(WX1004), .Z(WX81) ) ;
AND2    gate8210  (.A(WX2326), .B(WX83), .Z(WX82) ) ;
AND2    gate8211  (.A(WX491), .B(WX1004), .Z(WX85) ) ;
AND2    gate8212  (.A(DATA_9_28), .B(WX87), .Z(WX86) ) ;
OR2     gate8213  (.A(WX100), .B(WX99), .Z(WX102) ) ;
AND2    gate8214  (.A(WX102), .B(WX1003), .Z(WX91) ) ;
OR2     gate8215  (.A(WX96), .B(WX95), .Z(WX98) ) ;
AND2    gate8216  (.A(WX98), .B(WX93), .Z(WX92) ) ;
AND2    gate8217  (.A(CRC_OUT_9_27), .B(WX1004), .Z(WX95) ) ;
AND2    gate8218  (.A(WX2333), .B(WX97), .Z(WX96) ) ;
AND2    gate8219  (.A(WX493), .B(WX1004), .Z(WX99) ) ;
AND2    gate8220  (.A(DATA_9_27), .B(WX101), .Z(WX100) ) ;
OR2     gate8221  (.A(WX114), .B(WX113), .Z(WX116) ) ;
AND2    gate8222  (.A(WX116), .B(WX1003), .Z(WX105) ) ;
OR2     gate8223  (.A(WX110), .B(WX109), .Z(WX112) ) ;
AND2    gate8224  (.A(WX112), .B(WX107), .Z(WX106) ) ;
AND2    gate8225  (.A(CRC_OUT_9_26), .B(WX1004), .Z(WX109) ) ;
AND2    gate8226  (.A(WX2340), .B(WX111), .Z(WX110) ) ;
AND2    gate8227  (.A(WX495), .B(WX1004), .Z(WX113) ) ;
AND2    gate8228  (.A(DATA_9_26), .B(WX115), .Z(WX114) ) ;
OR2     gate8229  (.A(WX128), .B(WX127), .Z(WX130) ) ;
AND2    gate8230  (.A(WX130), .B(WX1003), .Z(WX119) ) ;
OR2     gate8231  (.A(WX124), .B(WX123), .Z(WX126) ) ;
AND2    gate8232  (.A(WX126), .B(WX121), .Z(WX120) ) ;
AND2    gate8233  (.A(CRC_OUT_9_25), .B(WX1004), .Z(WX123) ) ;
AND2    gate8234  (.A(WX2347), .B(WX125), .Z(WX124) ) ;
AND2    gate8235  (.A(WX497), .B(WX1004), .Z(WX127) ) ;
AND2    gate8236  (.A(DATA_9_25), .B(WX129), .Z(WX128) ) ;
OR2     gate8237  (.A(WX142), .B(WX141), .Z(WX144) ) ;
AND2    gate8238  (.A(WX144), .B(WX1003), .Z(WX133) ) ;
OR2     gate8239  (.A(WX138), .B(WX137), .Z(WX140) ) ;
AND2    gate8240  (.A(WX140), .B(WX135), .Z(WX134) ) ;
AND2    gate8241  (.A(CRC_OUT_9_24), .B(WX1004), .Z(WX137) ) ;
AND2    gate8242  (.A(WX2354), .B(WX139), .Z(WX138) ) ;
AND2    gate8243  (.A(WX499), .B(WX1004), .Z(WX141) ) ;
AND2    gate8244  (.A(DATA_9_24), .B(WX143), .Z(WX142) ) ;
OR2     gate8245  (.A(WX156), .B(WX155), .Z(WX158) ) ;
AND2    gate8246  (.A(WX158), .B(WX1003), .Z(WX147) ) ;
OR2     gate8247  (.A(WX152), .B(WX151), .Z(WX154) ) ;
AND2    gate8248  (.A(WX154), .B(WX149), .Z(WX148) ) ;
AND2    gate8249  (.A(CRC_OUT_9_23), .B(WX1004), .Z(WX151) ) ;
AND2    gate8250  (.A(WX2361), .B(WX153), .Z(WX152) ) ;
AND2    gate8251  (.A(WX501), .B(WX1004), .Z(WX155) ) ;
AND2    gate8252  (.A(DATA_9_23), .B(WX157), .Z(WX156) ) ;
OR2     gate8253  (.A(WX170), .B(WX169), .Z(WX172) ) ;
AND2    gate8254  (.A(WX172), .B(WX1003), .Z(WX161) ) ;
OR2     gate8255  (.A(WX166), .B(WX165), .Z(WX168) ) ;
AND2    gate8256  (.A(WX168), .B(WX163), .Z(WX162) ) ;
AND2    gate8257  (.A(CRC_OUT_9_22), .B(WX1004), .Z(WX165) ) ;
AND2    gate8258  (.A(WX2368), .B(WX167), .Z(WX166) ) ;
AND2    gate8259  (.A(WX503), .B(WX1004), .Z(WX169) ) ;
AND2    gate8260  (.A(DATA_9_22), .B(WX171), .Z(WX170) ) ;
OR2     gate8261  (.A(WX184), .B(WX183), .Z(WX186) ) ;
AND2    gate8262  (.A(WX186), .B(WX1003), .Z(WX175) ) ;
OR2     gate8263  (.A(WX180), .B(WX179), .Z(WX182) ) ;
AND2    gate8264  (.A(WX182), .B(WX177), .Z(WX176) ) ;
AND2    gate8265  (.A(CRC_OUT_9_21), .B(WX1004), .Z(WX179) ) ;
AND2    gate8266  (.A(WX2375), .B(WX181), .Z(WX180) ) ;
AND2    gate8267  (.A(WX505), .B(WX1004), .Z(WX183) ) ;
AND2    gate8268  (.A(DATA_9_21), .B(WX185), .Z(WX184) ) ;
OR2     gate8269  (.A(WX198), .B(WX197), .Z(WX200) ) ;
AND2    gate8270  (.A(WX200), .B(WX1003), .Z(WX189) ) ;
OR2     gate8271  (.A(WX194), .B(WX193), .Z(WX196) ) ;
AND2    gate8272  (.A(WX196), .B(WX191), .Z(WX190) ) ;
AND2    gate8273  (.A(CRC_OUT_9_20), .B(WX1004), .Z(WX193) ) ;
AND2    gate8274  (.A(WX2382), .B(WX195), .Z(WX194) ) ;
AND2    gate8275  (.A(WX507), .B(WX1004), .Z(WX197) ) ;
AND2    gate8276  (.A(DATA_9_20), .B(WX199), .Z(WX198) ) ;
OR2     gate8277  (.A(WX212), .B(WX211), .Z(WX214) ) ;
AND2    gate8278  (.A(WX214), .B(WX1003), .Z(WX203) ) ;
OR2     gate8279  (.A(WX208), .B(WX207), .Z(WX210) ) ;
AND2    gate8280  (.A(WX210), .B(WX205), .Z(WX204) ) ;
AND2    gate8281  (.A(CRC_OUT_9_19), .B(WX1004), .Z(WX207) ) ;
AND2    gate8282  (.A(WX2389), .B(WX209), .Z(WX208) ) ;
AND2    gate8283  (.A(WX509), .B(WX1004), .Z(WX211) ) ;
AND2    gate8284  (.A(DATA_9_19), .B(WX213), .Z(WX212) ) ;
OR2     gate8285  (.A(WX226), .B(WX225), .Z(WX228) ) ;
AND2    gate8286  (.A(WX228), .B(WX1003), .Z(WX217) ) ;
OR2     gate8287  (.A(WX222), .B(WX221), .Z(WX224) ) ;
AND2    gate8288  (.A(WX224), .B(WX219), .Z(WX218) ) ;
AND2    gate8289  (.A(CRC_OUT_9_18), .B(WX1004), .Z(WX221) ) ;
AND2    gate8290  (.A(WX2396), .B(WX223), .Z(WX222) ) ;
AND2    gate8291  (.A(WX511), .B(WX1004), .Z(WX225) ) ;
AND2    gate8292  (.A(DATA_9_18), .B(WX227), .Z(WX226) ) ;
OR2     gate8293  (.A(WX240), .B(WX239), .Z(WX242) ) ;
AND2    gate8294  (.A(WX242), .B(WX1003), .Z(WX231) ) ;
OR2     gate8295  (.A(WX236), .B(WX235), .Z(WX238) ) ;
AND2    gate8296  (.A(WX238), .B(WX233), .Z(WX232) ) ;
AND2    gate8297  (.A(CRC_OUT_9_17), .B(WX1004), .Z(WX235) ) ;
AND2    gate8298  (.A(WX2403), .B(WX237), .Z(WX236) ) ;
AND2    gate8299  (.A(WX513), .B(WX1004), .Z(WX239) ) ;
AND2    gate8300  (.A(DATA_9_17), .B(WX241), .Z(WX240) ) ;
OR2     gate8301  (.A(WX254), .B(WX253), .Z(WX256) ) ;
AND2    gate8302  (.A(WX256), .B(WX1003), .Z(WX245) ) ;
OR2     gate8303  (.A(WX250), .B(WX249), .Z(WX252) ) ;
AND2    gate8304  (.A(WX252), .B(WX247), .Z(WX246) ) ;
AND2    gate8305  (.A(CRC_OUT_9_16), .B(WX1004), .Z(WX249) ) ;
AND2    gate8306  (.A(WX2410), .B(WX251), .Z(WX250) ) ;
AND2    gate8307  (.A(WX515), .B(WX1004), .Z(WX253) ) ;
AND2    gate8308  (.A(DATA_9_16), .B(WX255), .Z(WX254) ) ;
OR2     gate8309  (.A(WX268), .B(WX267), .Z(WX270) ) ;
AND2    gate8310  (.A(WX270), .B(WX1003), .Z(WX259) ) ;
OR2     gate8311  (.A(WX264), .B(WX263), .Z(WX266) ) ;
AND2    gate8312  (.A(WX266), .B(WX261), .Z(WX260) ) ;
AND2    gate8313  (.A(CRC_OUT_9_15), .B(WX1004), .Z(WX263) ) ;
AND2    gate8314  (.A(WX2417), .B(WX265), .Z(WX264) ) ;
AND2    gate8315  (.A(WX517), .B(WX1004), .Z(WX267) ) ;
AND2    gate8316  (.A(DATA_9_15), .B(WX269), .Z(WX268) ) ;
OR2     gate8317  (.A(WX282), .B(WX281), .Z(WX284) ) ;
AND2    gate8318  (.A(WX284), .B(WX1003), .Z(WX273) ) ;
OR2     gate8319  (.A(WX278), .B(WX277), .Z(WX280) ) ;
AND2    gate8320  (.A(WX280), .B(WX275), .Z(WX274) ) ;
AND2    gate8321  (.A(CRC_OUT_9_14), .B(WX1004), .Z(WX277) ) ;
AND2    gate8322  (.A(WX2424), .B(WX279), .Z(WX278) ) ;
AND2    gate8323  (.A(WX519), .B(WX1004), .Z(WX281) ) ;
AND2    gate8324  (.A(DATA_9_14), .B(WX283), .Z(WX282) ) ;
OR2     gate8325  (.A(WX296), .B(WX295), .Z(WX298) ) ;
AND2    gate8326  (.A(WX298), .B(WX1003), .Z(WX287) ) ;
OR2     gate8327  (.A(WX292), .B(WX291), .Z(WX294) ) ;
AND2    gate8328  (.A(WX294), .B(WX289), .Z(WX288) ) ;
AND2    gate8329  (.A(CRC_OUT_9_13), .B(WX1004), .Z(WX291) ) ;
AND2    gate8330  (.A(WX2431), .B(WX293), .Z(WX292) ) ;
AND2    gate8331  (.A(WX521), .B(WX1004), .Z(WX295) ) ;
AND2    gate8332  (.A(DATA_9_13), .B(WX297), .Z(WX296) ) ;
OR2     gate8333  (.A(WX310), .B(WX309), .Z(WX312) ) ;
AND2    gate8334  (.A(WX312), .B(WX1003), .Z(WX301) ) ;
OR2     gate8335  (.A(WX306), .B(WX305), .Z(WX308) ) ;
AND2    gate8336  (.A(WX308), .B(WX303), .Z(WX302) ) ;
AND2    gate8337  (.A(CRC_OUT_9_12), .B(WX1004), .Z(WX305) ) ;
AND2    gate8338  (.A(WX2438), .B(WX307), .Z(WX306) ) ;
AND2    gate8339  (.A(WX523), .B(WX1004), .Z(WX309) ) ;
AND2    gate8340  (.A(DATA_9_12), .B(WX311), .Z(WX310) ) ;
OR2     gate8341  (.A(WX324), .B(WX323), .Z(WX326) ) ;
AND2    gate8342  (.A(WX326), .B(WX1003), .Z(WX315) ) ;
OR2     gate8343  (.A(WX320), .B(WX319), .Z(WX322) ) ;
AND2    gate8344  (.A(WX322), .B(WX317), .Z(WX316) ) ;
AND2    gate8345  (.A(CRC_OUT_9_11), .B(WX1004), .Z(WX319) ) ;
AND2    gate8346  (.A(WX2445), .B(WX321), .Z(WX320) ) ;
AND2    gate8347  (.A(WX525), .B(WX1004), .Z(WX323) ) ;
AND2    gate8348  (.A(DATA_9_11), .B(WX325), .Z(WX324) ) ;
OR2     gate8349  (.A(WX338), .B(WX337), .Z(WX340) ) ;
AND2    gate8350  (.A(WX340), .B(WX1003), .Z(WX329) ) ;
OR2     gate8351  (.A(WX334), .B(WX333), .Z(WX336) ) ;
AND2    gate8352  (.A(WX336), .B(WX331), .Z(WX330) ) ;
AND2    gate8353  (.A(CRC_OUT_9_10), .B(WX1004), .Z(WX333) ) ;
AND2    gate8354  (.A(WX2452), .B(WX335), .Z(WX334) ) ;
AND2    gate8355  (.A(WX527), .B(WX1004), .Z(WX337) ) ;
AND2    gate8356  (.A(DATA_9_10), .B(WX339), .Z(WX338) ) ;
OR2     gate8357  (.A(WX352), .B(WX351), .Z(WX354) ) ;
AND2    gate8358  (.A(WX354), .B(WX1003), .Z(WX343) ) ;
OR2     gate8359  (.A(WX348), .B(WX347), .Z(WX350) ) ;
AND2    gate8360  (.A(WX350), .B(WX345), .Z(WX344) ) ;
AND2    gate8361  (.A(CRC_OUT_9_9), .B(WX1004), .Z(WX347) ) ;
AND2    gate8362  (.A(WX2459), .B(WX349), .Z(WX348) ) ;
AND2    gate8363  (.A(WX529), .B(WX1004), .Z(WX351) ) ;
AND2    gate8364  (.A(DATA_9_9), .B(WX353), .Z(WX352) ) ;
OR2     gate8365  (.A(WX366), .B(WX365), .Z(WX368) ) ;
AND2    gate8366  (.A(WX368), .B(WX1003), .Z(WX357) ) ;
OR2     gate8367  (.A(WX362), .B(WX361), .Z(WX364) ) ;
AND2    gate8368  (.A(WX364), .B(WX359), .Z(WX358) ) ;
AND2    gate8369  (.A(CRC_OUT_9_8), .B(WX1004), .Z(WX361) ) ;
AND2    gate8370  (.A(WX2466), .B(WX363), .Z(WX362) ) ;
AND2    gate8371  (.A(WX531), .B(WX1004), .Z(WX365) ) ;
AND2    gate8372  (.A(DATA_9_8), .B(WX367), .Z(WX366) ) ;
OR2     gate8373  (.A(WX380), .B(WX379), .Z(WX382) ) ;
AND2    gate8374  (.A(WX382), .B(WX1003), .Z(WX371) ) ;
OR2     gate8375  (.A(WX376), .B(WX375), .Z(WX378) ) ;
AND2    gate8376  (.A(WX378), .B(WX373), .Z(WX372) ) ;
AND2    gate8377  (.A(CRC_OUT_9_7), .B(WX1004), .Z(WX375) ) ;
AND2    gate8378  (.A(WX2473), .B(WX377), .Z(WX376) ) ;
AND2    gate8379  (.A(WX533), .B(WX1004), .Z(WX379) ) ;
AND2    gate8380  (.A(DATA_9_7), .B(WX381), .Z(WX380) ) ;
OR2     gate8381  (.A(WX394), .B(WX393), .Z(WX396) ) ;
AND2    gate8382  (.A(WX396), .B(WX1003), .Z(WX385) ) ;
OR2     gate8383  (.A(WX390), .B(WX389), .Z(WX392) ) ;
AND2    gate8384  (.A(WX392), .B(WX387), .Z(WX386) ) ;
AND2    gate8385  (.A(CRC_OUT_9_6), .B(WX1004), .Z(WX389) ) ;
AND2    gate8386  (.A(WX2480), .B(WX391), .Z(WX390) ) ;
AND2    gate8387  (.A(WX535), .B(WX1004), .Z(WX393) ) ;
AND2    gate8388  (.A(DATA_9_6), .B(WX395), .Z(WX394) ) ;
OR2     gate8389  (.A(WX408), .B(WX407), .Z(WX410) ) ;
AND2    gate8390  (.A(WX410), .B(WX1003), .Z(WX399) ) ;
OR2     gate8391  (.A(WX404), .B(WX403), .Z(WX406) ) ;
AND2    gate8392  (.A(WX406), .B(WX401), .Z(WX400) ) ;
AND2    gate8393  (.A(CRC_OUT_9_5), .B(WX1004), .Z(WX403) ) ;
AND2    gate8394  (.A(WX2487), .B(WX405), .Z(WX404) ) ;
AND2    gate8395  (.A(WX537), .B(WX1004), .Z(WX407) ) ;
AND2    gate8396  (.A(DATA_9_5), .B(WX409), .Z(WX408) ) ;
OR2     gate8397  (.A(WX422), .B(WX421), .Z(WX424) ) ;
AND2    gate8398  (.A(WX424), .B(WX1003), .Z(WX413) ) ;
OR2     gate8399  (.A(WX418), .B(WX417), .Z(WX420) ) ;
AND2    gate8400  (.A(WX420), .B(WX415), .Z(WX414) ) ;
AND2    gate8401  (.A(CRC_OUT_9_4), .B(WX1004), .Z(WX417) ) ;
AND2    gate8402  (.A(WX2494), .B(WX419), .Z(WX418) ) ;
AND2    gate8403  (.A(WX539), .B(WX1004), .Z(WX421) ) ;
AND2    gate8404  (.A(DATA_9_4), .B(WX423), .Z(WX422) ) ;
OR2     gate8405  (.A(WX436), .B(WX435), .Z(WX438) ) ;
AND2    gate8406  (.A(WX438), .B(WX1003), .Z(WX427) ) ;
OR2     gate8407  (.A(WX432), .B(WX431), .Z(WX434) ) ;
AND2    gate8408  (.A(WX434), .B(WX429), .Z(WX428) ) ;
AND2    gate8409  (.A(CRC_OUT_9_3), .B(WX1004), .Z(WX431) ) ;
AND2    gate8410  (.A(WX2501), .B(WX433), .Z(WX432) ) ;
AND2    gate8411  (.A(WX541), .B(WX1004), .Z(WX435) ) ;
AND2    gate8412  (.A(DATA_9_3), .B(WX437), .Z(WX436) ) ;
OR2     gate8413  (.A(WX450), .B(WX449), .Z(WX452) ) ;
AND2    gate8414  (.A(WX452), .B(WX1003), .Z(WX441) ) ;
OR2     gate8415  (.A(WX446), .B(WX445), .Z(WX448) ) ;
AND2    gate8416  (.A(WX448), .B(WX443), .Z(WX442) ) ;
AND2    gate8417  (.A(CRC_OUT_9_2), .B(WX1004), .Z(WX445) ) ;
AND2    gate8418  (.A(WX2508), .B(WX447), .Z(WX446) ) ;
AND2    gate8419  (.A(WX543), .B(WX1004), .Z(WX449) ) ;
AND2    gate8420  (.A(DATA_9_2), .B(WX451), .Z(WX450) ) ;
OR2     gate8421  (.A(WX464), .B(WX463), .Z(WX466) ) ;
AND2    gate8422  (.A(WX466), .B(WX1003), .Z(WX455) ) ;
OR2     gate8423  (.A(WX460), .B(WX459), .Z(WX462) ) ;
AND2    gate8424  (.A(WX462), .B(WX457), .Z(WX456) ) ;
AND2    gate8425  (.A(CRC_OUT_9_1), .B(WX1004), .Z(WX459) ) ;
AND2    gate8426  (.A(WX2515), .B(WX461), .Z(WX460) ) ;
AND2    gate8427  (.A(WX545), .B(WX1004), .Z(WX463) ) ;
AND2    gate8428  (.A(DATA_9_1), .B(WX465), .Z(WX464) ) ;
OR2     gate8429  (.A(WX478), .B(WX477), .Z(WX480) ) ;
AND2    gate8430  (.A(WX480), .B(WX1003), .Z(WX469) ) ;
OR2     gate8431  (.A(WX474), .B(WX473), .Z(WX476) ) ;
AND2    gate8432  (.A(WX476), .B(WX471), .Z(WX470) ) ;
AND2    gate8433  (.A(CRC_OUT_9_0), .B(WX1004), .Z(WX473) ) ;
AND2    gate8434  (.A(WX2522), .B(WX475), .Z(WX474) ) ;
AND2    gate8435  (.A(WX547), .B(WX1004), .Z(WX477) ) ;
AND2    gate8436  (.A(DATA_9_0), .B(WX479), .Z(WX478) ) ;
NAND2   gate8437  (.A(II3053), .B(II3054), .Z(WX1006) ) ;
AND2    gate8438  (.A(WX1006), .B(WX1005), .Z(WX1007) ) ;
AND2    gate8439  (.A(WX580), .B(WX1009), .Z(WX1008) ) ;
NAND2   gate8440  (.A(II3066), .B(II3067), .Z(WX1013) ) ;
AND2    gate8441  (.A(WX1013), .B(WX1005), .Z(WX1014) ) ;
AND2    gate8442  (.A(WX581), .B(WX1016), .Z(WX1015) ) ;
NAND2   gate8443  (.A(II3079), .B(II3080), .Z(WX1020) ) ;
AND2    gate8444  (.A(WX1020), .B(WX1005), .Z(WX1021) ) ;
AND2    gate8445  (.A(WX582), .B(WX1023), .Z(WX1022) ) ;
NAND2   gate8446  (.A(II3092), .B(II3093), .Z(WX1027) ) ;
AND2    gate8447  (.A(WX1027), .B(WX1005), .Z(WX1028) ) ;
AND2    gate8448  (.A(WX583), .B(WX1030), .Z(WX1029) ) ;
NAND2   gate8449  (.A(II3105), .B(II3106), .Z(WX1034) ) ;
AND2    gate8450  (.A(WX1034), .B(WX1005), .Z(WX1035) ) ;
AND2    gate8451  (.A(WX584), .B(WX1037), .Z(WX1036) ) ;
NAND2   gate8452  (.A(II3118), .B(II3119), .Z(WX1041) ) ;
AND2    gate8453  (.A(WX1041), .B(WX1005), .Z(WX1042) ) ;
AND2    gate8454  (.A(WX585), .B(WX1044), .Z(WX1043) ) ;
NAND2   gate8455  (.A(II3131), .B(II3132), .Z(WX1048) ) ;
AND2    gate8456  (.A(WX1048), .B(WX1005), .Z(WX1049) ) ;
AND2    gate8457  (.A(WX586), .B(WX1051), .Z(WX1050) ) ;
NAND2   gate8458  (.A(II3144), .B(II3145), .Z(WX1055) ) ;
AND2    gate8459  (.A(WX1055), .B(WX1005), .Z(WX1056) ) ;
AND2    gate8460  (.A(WX587), .B(WX1058), .Z(WX1057) ) ;
NAND2   gate8461  (.A(II3157), .B(II3158), .Z(WX1062) ) ;
AND2    gate8462  (.A(WX1062), .B(WX1005), .Z(WX1063) ) ;
AND2    gate8463  (.A(WX588), .B(WX1065), .Z(WX1064) ) ;
NAND2   gate8464  (.A(II3170), .B(II3171), .Z(WX1069) ) ;
AND2    gate8465  (.A(WX1069), .B(WX1005), .Z(WX1070) ) ;
AND2    gate8466  (.A(WX589), .B(WX1072), .Z(WX1071) ) ;
NAND2   gate8467  (.A(II3183), .B(II3184), .Z(WX1076) ) ;
AND2    gate8468  (.A(WX1076), .B(WX1005), .Z(WX1077) ) ;
AND2    gate8469  (.A(WX590), .B(WX1079), .Z(WX1078) ) ;
NAND2   gate8470  (.A(II3196), .B(II3197), .Z(WX1083) ) ;
AND2    gate8471  (.A(WX1083), .B(WX1005), .Z(WX1084) ) ;
AND2    gate8472  (.A(WX591), .B(WX1086), .Z(WX1085) ) ;
NAND2   gate8473  (.A(II3209), .B(II3210), .Z(WX1090) ) ;
AND2    gate8474  (.A(WX1090), .B(WX1005), .Z(WX1091) ) ;
AND2    gate8475  (.A(WX592), .B(WX1093), .Z(WX1092) ) ;
NAND2   gate8476  (.A(II3222), .B(II3223), .Z(WX1097) ) ;
AND2    gate8477  (.A(WX1097), .B(WX1005), .Z(WX1098) ) ;
AND2    gate8478  (.A(WX593), .B(WX1100), .Z(WX1099) ) ;
NAND2   gate8479  (.A(II3235), .B(II3236), .Z(WX1104) ) ;
AND2    gate8480  (.A(WX1104), .B(WX1005), .Z(WX1105) ) ;
AND2    gate8481  (.A(WX594), .B(WX1107), .Z(WX1106) ) ;
NAND2   gate8482  (.A(II3248), .B(II3249), .Z(WX1111) ) ;
AND2    gate8483  (.A(WX1111), .B(WX1005), .Z(WX1112) ) ;
AND2    gate8484  (.A(WX595), .B(WX1114), .Z(WX1113) ) ;
NAND2   gate8485  (.A(II3261), .B(II3262), .Z(WX1118) ) ;
AND2    gate8486  (.A(WX1118), .B(WX1005), .Z(WX1119) ) ;
AND2    gate8487  (.A(WX596), .B(WX1121), .Z(WX1120) ) ;
NAND2   gate8488  (.A(II3274), .B(II3275), .Z(WX1125) ) ;
AND2    gate8489  (.A(WX1125), .B(WX1005), .Z(WX1126) ) ;
AND2    gate8490  (.A(WX597), .B(WX1128), .Z(WX1127) ) ;
NAND2   gate8491  (.A(II3287), .B(II3288), .Z(WX1132) ) ;
AND2    gate8492  (.A(WX1132), .B(WX1005), .Z(WX1133) ) ;
AND2    gate8493  (.A(WX598), .B(WX1135), .Z(WX1134) ) ;
NAND2   gate8494  (.A(II3300), .B(II3301), .Z(WX1139) ) ;
AND2    gate8495  (.A(WX1139), .B(WX1005), .Z(WX1140) ) ;
AND2    gate8496  (.A(WX599), .B(WX1142), .Z(WX1141) ) ;
NAND2   gate8497  (.A(II3313), .B(II3314), .Z(WX1146) ) ;
AND2    gate8498  (.A(WX1146), .B(WX1005), .Z(WX1147) ) ;
AND2    gate8499  (.A(WX600), .B(WX1149), .Z(WX1148) ) ;
NAND2   gate8500  (.A(II3326), .B(II3327), .Z(WX1153) ) ;
AND2    gate8501  (.A(WX1153), .B(WX1005), .Z(WX1154) ) ;
AND2    gate8502  (.A(WX601), .B(WX1156), .Z(WX1155) ) ;
NAND2   gate8503  (.A(II3339), .B(II3340), .Z(WX1160) ) ;
AND2    gate8504  (.A(WX1160), .B(WX1005), .Z(WX1161) ) ;
AND2    gate8505  (.A(WX602), .B(WX1163), .Z(WX1162) ) ;
NAND2   gate8506  (.A(II3352), .B(II3353), .Z(WX1167) ) ;
AND2    gate8507  (.A(WX1167), .B(WX1005), .Z(WX1168) ) ;
AND2    gate8508  (.A(WX603), .B(WX1170), .Z(WX1169) ) ;
NAND2   gate8509  (.A(II3365), .B(II3366), .Z(WX1174) ) ;
AND2    gate8510  (.A(WX1174), .B(WX1005), .Z(WX1175) ) ;
AND2    gate8511  (.A(WX604), .B(WX1177), .Z(WX1176) ) ;
NAND2   gate8512  (.A(II3378), .B(II3379), .Z(WX1181) ) ;
AND2    gate8513  (.A(WX1181), .B(WX1005), .Z(WX1182) ) ;
AND2    gate8514  (.A(WX605), .B(WX1184), .Z(WX1183) ) ;
NAND2   gate8515  (.A(II3391), .B(II3392), .Z(WX1188) ) ;
AND2    gate8516  (.A(WX1188), .B(WX1005), .Z(WX1189) ) ;
AND2    gate8517  (.A(WX606), .B(WX1191), .Z(WX1190) ) ;
NAND2   gate8518  (.A(II3404), .B(II3405), .Z(WX1195) ) ;
AND2    gate8519  (.A(WX1195), .B(WX1005), .Z(WX1196) ) ;
AND2    gate8520  (.A(WX607), .B(WX1198), .Z(WX1197) ) ;
NAND2   gate8521  (.A(II3417), .B(II3418), .Z(WX1202) ) ;
AND2    gate8522  (.A(WX1202), .B(WX1005), .Z(WX1203) ) ;
AND2    gate8523  (.A(WX608), .B(WX1205), .Z(WX1204) ) ;
NAND2   gate8524  (.A(II3430), .B(II3431), .Z(WX1209) ) ;
AND2    gate8525  (.A(WX1209), .B(WX1005), .Z(WX1210) ) ;
AND2    gate8526  (.A(WX609), .B(WX1212), .Z(WX1211) ) ;
NAND2   gate8527  (.A(II3443), .B(II3444), .Z(WX1216) ) ;
AND2    gate8528  (.A(WX1216), .B(WX1005), .Z(WX1217) ) ;
AND2    gate8529  (.A(WX610), .B(WX1219), .Z(WX1218) ) ;
NAND2   gate8530  (.A(II3456), .B(II3457), .Z(WX1223) ) ;
AND2    gate8531  (.A(WX1223), .B(WX1005), .Z(WX1224) ) ;
AND2    gate8532  (.A(WX611), .B(WX1226), .Z(WX1225) ) ;
NAND2   gate8533  (.A(II3515), .B(II3516), .Z(WX1234) ) ;
NAND2   gate8534  (.A(II3711), .B(II3712), .Z(WX1262) ) ;
NAND2   gate8535  (.A(II3704), .B(II3705), .Z(WX1261) ) ;
NAND2   gate8536  (.A(II3697), .B(II3698), .Z(WX1260) ) ;
NAND2   gate8537  (.A(II3508), .B(II3509), .Z(WX1233) ) ;
NAND2   gate8538  (.A(II3690), .B(II3691), .Z(WX1259) ) ;
NAND2   gate8539  (.A(II3683), .B(II3684), .Z(WX1258) ) ;
NAND2   gate8540  (.A(II3676), .B(II3677), .Z(WX1257) ) ;
NAND2   gate8541  (.A(II3669), .B(II3670), .Z(WX1256) ) ;
NAND2   gate8542  (.A(II3662), .B(II3663), .Z(WX1255) ) ;
NAND2   gate8543  (.A(II3655), .B(II3656), .Z(WX1254) ) ;
NAND2   gate8544  (.A(II3493), .B(II3494), .Z(WX1232) ) ;
NAND2   gate8545  (.A(II3648), .B(II3649), .Z(WX1253) ) ;
NAND2   gate8546  (.A(II3641), .B(II3642), .Z(WX1252) ) ;
NAND2   gate8547  (.A(II3634), .B(II3635), .Z(WX1251) ) ;
NAND2   gate8548  (.A(II3627), .B(II3628), .Z(WX1250) ) ;
NAND2   gate8549  (.A(II3478), .B(II3479), .Z(WX1231) ) ;
NAND2   gate8550  (.A(II3620), .B(II3621), .Z(WX1249) ) ;
NAND2   gate8551  (.A(II3613), .B(II3614), .Z(WX1248) ) ;
NAND2   gate8552  (.A(II3606), .B(II3607), .Z(WX1247) ) ;
NAND2   gate8553  (.A(II3599), .B(II3600), .Z(WX1246) ) ;
NAND2   gate8554  (.A(II3592), .B(II3593), .Z(WX1245) ) ;
NAND2   gate8555  (.A(II3585), .B(II3586), .Z(WX1244) ) ;
NAND2   gate8556  (.A(II3578), .B(II3579), .Z(WX1243) ) ;
NAND2   gate8557  (.A(II3571), .B(II3572), .Z(WX1242) ) ;
NAND2   gate8558  (.A(II3564), .B(II3565), .Z(WX1241) ) ;
NAND2   gate8559  (.A(II3557), .B(II3558), .Z(WX1240) ) ;
NAND2   gate8560  (.A(II3550), .B(II3551), .Z(WX1239) ) ;
NAND2   gate8561  (.A(II3543), .B(II3544), .Z(WX1238) ) ;
NAND2   gate8562  (.A(II3536), .B(II3537), .Z(WX1237) ) ;
NAND2   gate8563  (.A(II3529), .B(II3530), .Z(WX1236) ) ;
NAND2   gate8564  (.A(II3522), .B(II3523), .Z(WX1235) ) ;
OR2     gate8565  (.A(WX1337), .B(WX1336), .Z(WX1339) ) ;
AND2    gate8566  (.A(WX1339), .B(WX2296), .Z(WX1328) ) ;
OR2     gate8567  (.A(WX1333), .B(WX1332), .Z(WX1335) ) ;
AND2    gate8568  (.A(WX1335), .B(WX1330), .Z(WX1329) ) ;
AND2    gate8569  (.A(CRC_OUT_8_31), .B(WX2297), .Z(WX1332) ) ;
AND2    gate8570  (.A(WX3598), .B(WX1334), .Z(WX1333) ) ;
AND2    gate8571  (.A(WX1778), .B(WX2297), .Z(WX1336) ) ;
AND2    gate8572  (.A(WX2305), .B(WX1338), .Z(WX1337) ) ;
OR2     gate8573  (.A(WX1351), .B(WX1350), .Z(WX1353) ) ;
AND2    gate8574  (.A(WX1353), .B(WX2296), .Z(WX1342) ) ;
OR2     gate8575  (.A(WX1347), .B(WX1346), .Z(WX1349) ) ;
AND2    gate8576  (.A(WX1349), .B(WX1344), .Z(WX1343) ) ;
AND2    gate8577  (.A(CRC_OUT_8_30), .B(WX2297), .Z(WX1346) ) ;
AND2    gate8578  (.A(WX3605), .B(WX1348), .Z(WX1347) ) ;
AND2    gate8579  (.A(WX1780), .B(WX2297), .Z(WX1350) ) ;
AND2    gate8580  (.A(WX2312), .B(WX1352), .Z(WX1351) ) ;
OR2     gate8581  (.A(WX1365), .B(WX1364), .Z(WX1367) ) ;
AND2    gate8582  (.A(WX1367), .B(WX2296), .Z(WX1356) ) ;
OR2     gate8583  (.A(WX1361), .B(WX1360), .Z(WX1363) ) ;
AND2    gate8584  (.A(WX1363), .B(WX1358), .Z(WX1357) ) ;
AND2    gate8585  (.A(CRC_OUT_8_29), .B(WX2297), .Z(WX1360) ) ;
AND2    gate8586  (.A(WX3612), .B(WX1362), .Z(WX1361) ) ;
AND2    gate8587  (.A(WX1782), .B(WX2297), .Z(WX1364) ) ;
AND2    gate8588  (.A(WX2319), .B(WX1366), .Z(WX1365) ) ;
OR2     gate8589  (.A(WX1379), .B(WX1378), .Z(WX1381) ) ;
AND2    gate8590  (.A(WX1381), .B(WX2296), .Z(WX1370) ) ;
OR2     gate8591  (.A(WX1375), .B(WX1374), .Z(WX1377) ) ;
AND2    gate8592  (.A(WX1377), .B(WX1372), .Z(WX1371) ) ;
AND2    gate8593  (.A(CRC_OUT_8_28), .B(WX2297), .Z(WX1374) ) ;
AND2    gate8594  (.A(WX3619), .B(WX1376), .Z(WX1375) ) ;
AND2    gate8595  (.A(WX1784), .B(WX2297), .Z(WX1378) ) ;
AND2    gate8596  (.A(WX2326), .B(WX1380), .Z(WX1379) ) ;
OR2     gate8597  (.A(WX1393), .B(WX1392), .Z(WX1395) ) ;
AND2    gate8598  (.A(WX1395), .B(WX2296), .Z(WX1384) ) ;
OR2     gate8599  (.A(WX1389), .B(WX1388), .Z(WX1391) ) ;
AND2    gate8600  (.A(WX1391), .B(WX1386), .Z(WX1385) ) ;
AND2    gate8601  (.A(CRC_OUT_8_27), .B(WX2297), .Z(WX1388) ) ;
AND2    gate8602  (.A(WX3626), .B(WX1390), .Z(WX1389) ) ;
AND2    gate8603  (.A(WX1786), .B(WX2297), .Z(WX1392) ) ;
AND2    gate8604  (.A(WX2333), .B(WX1394), .Z(WX1393) ) ;
OR2     gate8605  (.A(WX1407), .B(WX1406), .Z(WX1409) ) ;
AND2    gate8606  (.A(WX1409), .B(WX2296), .Z(WX1398) ) ;
OR2     gate8607  (.A(WX1403), .B(WX1402), .Z(WX1405) ) ;
AND2    gate8608  (.A(WX1405), .B(WX1400), .Z(WX1399) ) ;
AND2    gate8609  (.A(CRC_OUT_8_26), .B(WX2297), .Z(WX1402) ) ;
AND2    gate8610  (.A(WX3633), .B(WX1404), .Z(WX1403) ) ;
AND2    gate8611  (.A(WX1788), .B(WX2297), .Z(WX1406) ) ;
AND2    gate8612  (.A(WX2340), .B(WX1408), .Z(WX1407) ) ;
OR2     gate8613  (.A(WX1421), .B(WX1420), .Z(WX1423) ) ;
AND2    gate8614  (.A(WX1423), .B(WX2296), .Z(WX1412) ) ;
OR2     gate8615  (.A(WX1417), .B(WX1416), .Z(WX1419) ) ;
AND2    gate8616  (.A(WX1419), .B(WX1414), .Z(WX1413) ) ;
AND2    gate8617  (.A(CRC_OUT_8_25), .B(WX2297), .Z(WX1416) ) ;
AND2    gate8618  (.A(WX3640), .B(WX1418), .Z(WX1417) ) ;
AND2    gate8619  (.A(WX1790), .B(WX2297), .Z(WX1420) ) ;
AND2    gate8620  (.A(WX2347), .B(WX1422), .Z(WX1421) ) ;
OR2     gate8621  (.A(WX1435), .B(WX1434), .Z(WX1437) ) ;
AND2    gate8622  (.A(WX1437), .B(WX2296), .Z(WX1426) ) ;
OR2     gate8623  (.A(WX1431), .B(WX1430), .Z(WX1433) ) ;
AND2    gate8624  (.A(WX1433), .B(WX1428), .Z(WX1427) ) ;
AND2    gate8625  (.A(CRC_OUT_8_24), .B(WX2297), .Z(WX1430) ) ;
AND2    gate8626  (.A(WX3647), .B(WX1432), .Z(WX1431) ) ;
AND2    gate8627  (.A(WX1792), .B(WX2297), .Z(WX1434) ) ;
AND2    gate8628  (.A(WX2354), .B(WX1436), .Z(WX1435) ) ;
OR2     gate8629  (.A(WX1449), .B(WX1448), .Z(WX1451) ) ;
AND2    gate8630  (.A(WX1451), .B(WX2296), .Z(WX1440) ) ;
OR2     gate8631  (.A(WX1445), .B(WX1444), .Z(WX1447) ) ;
AND2    gate8632  (.A(WX1447), .B(WX1442), .Z(WX1441) ) ;
AND2    gate8633  (.A(CRC_OUT_8_23), .B(WX2297), .Z(WX1444) ) ;
AND2    gate8634  (.A(WX3654), .B(WX1446), .Z(WX1445) ) ;
AND2    gate8635  (.A(WX1794), .B(WX2297), .Z(WX1448) ) ;
AND2    gate8636  (.A(WX2361), .B(WX1450), .Z(WX1449) ) ;
OR2     gate8637  (.A(WX1463), .B(WX1462), .Z(WX1465) ) ;
AND2    gate8638  (.A(WX1465), .B(WX2296), .Z(WX1454) ) ;
OR2     gate8639  (.A(WX1459), .B(WX1458), .Z(WX1461) ) ;
AND2    gate8640  (.A(WX1461), .B(WX1456), .Z(WX1455) ) ;
AND2    gate8641  (.A(CRC_OUT_8_22), .B(WX2297), .Z(WX1458) ) ;
AND2    gate8642  (.A(WX3661), .B(WX1460), .Z(WX1459) ) ;
AND2    gate8643  (.A(WX1796), .B(WX2297), .Z(WX1462) ) ;
AND2    gate8644  (.A(WX2368), .B(WX1464), .Z(WX1463) ) ;
OR2     gate8645  (.A(WX1477), .B(WX1476), .Z(WX1479) ) ;
AND2    gate8646  (.A(WX1479), .B(WX2296), .Z(WX1468) ) ;
OR2     gate8647  (.A(WX1473), .B(WX1472), .Z(WX1475) ) ;
AND2    gate8648  (.A(WX1475), .B(WX1470), .Z(WX1469) ) ;
AND2    gate8649  (.A(CRC_OUT_8_21), .B(WX2297), .Z(WX1472) ) ;
AND2    gate8650  (.A(WX3668), .B(WX1474), .Z(WX1473) ) ;
AND2    gate8651  (.A(WX1798), .B(WX2297), .Z(WX1476) ) ;
AND2    gate8652  (.A(WX2375), .B(WX1478), .Z(WX1477) ) ;
OR2     gate8653  (.A(WX1491), .B(WX1490), .Z(WX1493) ) ;
AND2    gate8654  (.A(WX1493), .B(WX2296), .Z(WX1482) ) ;
OR2     gate8655  (.A(WX1487), .B(WX1486), .Z(WX1489) ) ;
AND2    gate8656  (.A(WX1489), .B(WX1484), .Z(WX1483) ) ;
AND2    gate8657  (.A(CRC_OUT_8_20), .B(WX2297), .Z(WX1486) ) ;
AND2    gate8658  (.A(WX3675), .B(WX1488), .Z(WX1487) ) ;
AND2    gate8659  (.A(WX1800), .B(WX2297), .Z(WX1490) ) ;
AND2    gate8660  (.A(WX2382), .B(WX1492), .Z(WX1491) ) ;
OR2     gate8661  (.A(WX1505), .B(WX1504), .Z(WX1507) ) ;
AND2    gate8662  (.A(WX1507), .B(WX2296), .Z(WX1496) ) ;
OR2     gate8663  (.A(WX1501), .B(WX1500), .Z(WX1503) ) ;
AND2    gate8664  (.A(WX1503), .B(WX1498), .Z(WX1497) ) ;
AND2    gate8665  (.A(CRC_OUT_8_19), .B(WX2297), .Z(WX1500) ) ;
AND2    gate8666  (.A(WX3682), .B(WX1502), .Z(WX1501) ) ;
AND2    gate8667  (.A(WX1802), .B(WX2297), .Z(WX1504) ) ;
AND2    gate8668  (.A(WX2389), .B(WX1506), .Z(WX1505) ) ;
OR2     gate8669  (.A(WX1519), .B(WX1518), .Z(WX1521) ) ;
AND2    gate8670  (.A(WX1521), .B(WX2296), .Z(WX1510) ) ;
OR2     gate8671  (.A(WX1515), .B(WX1514), .Z(WX1517) ) ;
AND2    gate8672  (.A(WX1517), .B(WX1512), .Z(WX1511) ) ;
AND2    gate8673  (.A(CRC_OUT_8_18), .B(WX2297), .Z(WX1514) ) ;
AND2    gate8674  (.A(WX3689), .B(WX1516), .Z(WX1515) ) ;
AND2    gate8675  (.A(WX1804), .B(WX2297), .Z(WX1518) ) ;
AND2    gate8676  (.A(WX2396), .B(WX1520), .Z(WX1519) ) ;
OR2     gate8677  (.A(WX1533), .B(WX1532), .Z(WX1535) ) ;
AND2    gate8678  (.A(WX1535), .B(WX2296), .Z(WX1524) ) ;
OR2     gate8679  (.A(WX1529), .B(WX1528), .Z(WX1531) ) ;
AND2    gate8680  (.A(WX1531), .B(WX1526), .Z(WX1525) ) ;
AND2    gate8681  (.A(CRC_OUT_8_17), .B(WX2297), .Z(WX1528) ) ;
AND2    gate8682  (.A(WX3696), .B(WX1530), .Z(WX1529) ) ;
AND2    gate8683  (.A(WX1806), .B(WX2297), .Z(WX1532) ) ;
AND2    gate8684  (.A(WX2403), .B(WX1534), .Z(WX1533) ) ;
OR2     gate8685  (.A(WX1547), .B(WX1546), .Z(WX1549) ) ;
AND2    gate8686  (.A(WX1549), .B(WX2296), .Z(WX1538) ) ;
OR2     gate8687  (.A(WX1543), .B(WX1542), .Z(WX1545) ) ;
AND2    gate8688  (.A(WX1545), .B(WX1540), .Z(WX1539) ) ;
AND2    gate8689  (.A(CRC_OUT_8_16), .B(WX2297), .Z(WX1542) ) ;
AND2    gate8690  (.A(WX3703), .B(WX1544), .Z(WX1543) ) ;
AND2    gate8691  (.A(WX1808), .B(WX2297), .Z(WX1546) ) ;
AND2    gate8692  (.A(WX2410), .B(WX1548), .Z(WX1547) ) ;
OR2     gate8693  (.A(WX1561), .B(WX1560), .Z(WX1563) ) ;
AND2    gate8694  (.A(WX1563), .B(WX2296), .Z(WX1552) ) ;
OR2     gate8695  (.A(WX1557), .B(WX1556), .Z(WX1559) ) ;
AND2    gate8696  (.A(WX1559), .B(WX1554), .Z(WX1553) ) ;
AND2    gate8697  (.A(CRC_OUT_8_15), .B(WX2297), .Z(WX1556) ) ;
AND2    gate8698  (.A(WX3710), .B(WX1558), .Z(WX1557) ) ;
AND2    gate8699  (.A(WX1810), .B(WX2297), .Z(WX1560) ) ;
AND2    gate8700  (.A(WX2417), .B(WX1562), .Z(WX1561) ) ;
OR2     gate8701  (.A(WX1575), .B(WX1574), .Z(WX1577) ) ;
AND2    gate8702  (.A(WX1577), .B(WX2296), .Z(WX1566) ) ;
OR2     gate8703  (.A(WX1571), .B(WX1570), .Z(WX1573) ) ;
AND2    gate8704  (.A(WX1573), .B(WX1568), .Z(WX1567) ) ;
AND2    gate8705  (.A(CRC_OUT_8_14), .B(WX2297), .Z(WX1570) ) ;
AND2    gate8706  (.A(WX3717), .B(WX1572), .Z(WX1571) ) ;
AND2    gate8707  (.A(WX1812), .B(WX2297), .Z(WX1574) ) ;
AND2    gate8708  (.A(WX2424), .B(WX1576), .Z(WX1575) ) ;
OR2     gate8709  (.A(WX1589), .B(WX1588), .Z(WX1591) ) ;
AND2    gate8710  (.A(WX1591), .B(WX2296), .Z(WX1580) ) ;
OR2     gate8711  (.A(WX1585), .B(WX1584), .Z(WX1587) ) ;
AND2    gate8712  (.A(WX1587), .B(WX1582), .Z(WX1581) ) ;
AND2    gate8713  (.A(CRC_OUT_8_13), .B(WX2297), .Z(WX1584) ) ;
AND2    gate8714  (.A(WX3724), .B(WX1586), .Z(WX1585) ) ;
AND2    gate8715  (.A(WX1814), .B(WX2297), .Z(WX1588) ) ;
AND2    gate8716  (.A(WX2431), .B(WX1590), .Z(WX1589) ) ;
OR2     gate8717  (.A(WX1603), .B(WX1602), .Z(WX1605) ) ;
AND2    gate8718  (.A(WX1605), .B(WX2296), .Z(WX1594) ) ;
OR2     gate8719  (.A(WX1599), .B(WX1598), .Z(WX1601) ) ;
AND2    gate8720  (.A(WX1601), .B(WX1596), .Z(WX1595) ) ;
AND2    gate8721  (.A(CRC_OUT_8_12), .B(WX2297), .Z(WX1598) ) ;
AND2    gate8722  (.A(WX3731), .B(WX1600), .Z(WX1599) ) ;
AND2    gate8723  (.A(WX1816), .B(WX2297), .Z(WX1602) ) ;
AND2    gate8724  (.A(WX2438), .B(WX1604), .Z(WX1603) ) ;
OR2     gate8725  (.A(WX1617), .B(WX1616), .Z(WX1619) ) ;
AND2    gate8726  (.A(WX1619), .B(WX2296), .Z(WX1608) ) ;
OR2     gate8727  (.A(WX1613), .B(WX1612), .Z(WX1615) ) ;
AND2    gate8728  (.A(WX1615), .B(WX1610), .Z(WX1609) ) ;
AND2    gate8729  (.A(CRC_OUT_8_11), .B(WX2297), .Z(WX1612) ) ;
AND2    gate8730  (.A(WX3738), .B(WX1614), .Z(WX1613) ) ;
AND2    gate8731  (.A(WX1818), .B(WX2297), .Z(WX1616) ) ;
AND2    gate8732  (.A(WX2445), .B(WX1618), .Z(WX1617) ) ;
OR2     gate8733  (.A(WX1631), .B(WX1630), .Z(WX1633) ) ;
AND2    gate8734  (.A(WX1633), .B(WX2296), .Z(WX1622) ) ;
OR2     gate8735  (.A(WX1627), .B(WX1626), .Z(WX1629) ) ;
AND2    gate8736  (.A(WX1629), .B(WX1624), .Z(WX1623) ) ;
AND2    gate8737  (.A(CRC_OUT_8_10), .B(WX2297), .Z(WX1626) ) ;
AND2    gate8738  (.A(WX3745), .B(WX1628), .Z(WX1627) ) ;
AND2    gate8739  (.A(WX1820), .B(WX2297), .Z(WX1630) ) ;
AND2    gate8740  (.A(WX2452), .B(WX1632), .Z(WX1631) ) ;
OR2     gate8741  (.A(WX1645), .B(WX1644), .Z(WX1647) ) ;
AND2    gate8742  (.A(WX1647), .B(WX2296), .Z(WX1636) ) ;
OR2     gate8743  (.A(WX1641), .B(WX1640), .Z(WX1643) ) ;
AND2    gate8744  (.A(WX1643), .B(WX1638), .Z(WX1637) ) ;
AND2    gate8745  (.A(CRC_OUT_8_9), .B(WX2297), .Z(WX1640) ) ;
AND2    gate8746  (.A(WX3752), .B(WX1642), .Z(WX1641) ) ;
AND2    gate8747  (.A(WX1822), .B(WX2297), .Z(WX1644) ) ;
AND2    gate8748  (.A(WX2459), .B(WX1646), .Z(WX1645) ) ;
OR2     gate8749  (.A(WX1659), .B(WX1658), .Z(WX1661) ) ;
AND2    gate8750  (.A(WX1661), .B(WX2296), .Z(WX1650) ) ;
OR2     gate8751  (.A(WX1655), .B(WX1654), .Z(WX1657) ) ;
AND2    gate8752  (.A(WX1657), .B(WX1652), .Z(WX1651) ) ;
AND2    gate8753  (.A(CRC_OUT_8_8), .B(WX2297), .Z(WX1654) ) ;
AND2    gate8754  (.A(WX3759), .B(WX1656), .Z(WX1655) ) ;
AND2    gate8755  (.A(WX1824), .B(WX2297), .Z(WX1658) ) ;
AND2    gate8756  (.A(WX2466), .B(WX1660), .Z(WX1659) ) ;
OR2     gate8757  (.A(WX1673), .B(WX1672), .Z(WX1675) ) ;
AND2    gate8758  (.A(WX1675), .B(WX2296), .Z(WX1664) ) ;
OR2     gate8759  (.A(WX1669), .B(WX1668), .Z(WX1671) ) ;
AND2    gate8760  (.A(WX1671), .B(WX1666), .Z(WX1665) ) ;
AND2    gate8761  (.A(CRC_OUT_8_7), .B(WX2297), .Z(WX1668) ) ;
AND2    gate8762  (.A(WX3766), .B(WX1670), .Z(WX1669) ) ;
AND2    gate8763  (.A(WX1826), .B(WX2297), .Z(WX1672) ) ;
AND2    gate8764  (.A(WX2473), .B(WX1674), .Z(WX1673) ) ;
OR2     gate8765  (.A(WX1687), .B(WX1686), .Z(WX1689) ) ;
AND2    gate8766  (.A(WX1689), .B(WX2296), .Z(WX1678) ) ;
OR2     gate8767  (.A(WX1683), .B(WX1682), .Z(WX1685) ) ;
AND2    gate8768  (.A(WX1685), .B(WX1680), .Z(WX1679) ) ;
AND2    gate8769  (.A(CRC_OUT_8_6), .B(WX2297), .Z(WX1682) ) ;
AND2    gate8770  (.A(WX3773), .B(WX1684), .Z(WX1683) ) ;
AND2    gate8771  (.A(WX1828), .B(WX2297), .Z(WX1686) ) ;
AND2    gate8772  (.A(WX2480), .B(WX1688), .Z(WX1687) ) ;
OR2     gate8773  (.A(WX1701), .B(WX1700), .Z(WX1703) ) ;
AND2    gate8774  (.A(WX1703), .B(WX2296), .Z(WX1692) ) ;
OR2     gate8775  (.A(WX1697), .B(WX1696), .Z(WX1699) ) ;
AND2    gate8776  (.A(WX1699), .B(WX1694), .Z(WX1693) ) ;
AND2    gate8777  (.A(CRC_OUT_8_5), .B(WX2297), .Z(WX1696) ) ;
AND2    gate8778  (.A(WX3780), .B(WX1698), .Z(WX1697) ) ;
AND2    gate8779  (.A(WX1830), .B(WX2297), .Z(WX1700) ) ;
AND2    gate8780  (.A(WX2487), .B(WX1702), .Z(WX1701) ) ;
OR2     gate8781  (.A(WX1715), .B(WX1714), .Z(WX1717) ) ;
AND2    gate8782  (.A(WX1717), .B(WX2296), .Z(WX1706) ) ;
OR2     gate8783  (.A(WX1711), .B(WX1710), .Z(WX1713) ) ;
AND2    gate8784  (.A(WX1713), .B(WX1708), .Z(WX1707) ) ;
AND2    gate8785  (.A(CRC_OUT_8_4), .B(WX2297), .Z(WX1710) ) ;
AND2    gate8786  (.A(WX3787), .B(WX1712), .Z(WX1711) ) ;
AND2    gate8787  (.A(WX1832), .B(WX2297), .Z(WX1714) ) ;
AND2    gate8788  (.A(WX2494), .B(WX1716), .Z(WX1715) ) ;
OR2     gate8789  (.A(WX1729), .B(WX1728), .Z(WX1731) ) ;
AND2    gate8790  (.A(WX1731), .B(WX2296), .Z(WX1720) ) ;
OR2     gate8791  (.A(WX1725), .B(WX1724), .Z(WX1727) ) ;
AND2    gate8792  (.A(WX1727), .B(WX1722), .Z(WX1721) ) ;
AND2    gate8793  (.A(CRC_OUT_8_3), .B(WX2297), .Z(WX1724) ) ;
AND2    gate8794  (.A(WX3794), .B(WX1726), .Z(WX1725) ) ;
AND2    gate8795  (.A(WX1834), .B(WX2297), .Z(WX1728) ) ;
AND2    gate8796  (.A(WX2501), .B(WX1730), .Z(WX1729) ) ;
OR2     gate8797  (.A(WX1743), .B(WX1742), .Z(WX1745) ) ;
AND2    gate8798  (.A(WX1745), .B(WX2296), .Z(WX1734) ) ;
OR2     gate8799  (.A(WX1739), .B(WX1738), .Z(WX1741) ) ;
AND2    gate8800  (.A(WX1741), .B(WX1736), .Z(WX1735) ) ;
AND2    gate8801  (.A(CRC_OUT_8_2), .B(WX2297), .Z(WX1738) ) ;
AND2    gate8802  (.A(WX3801), .B(WX1740), .Z(WX1739) ) ;
AND2    gate8803  (.A(WX1836), .B(WX2297), .Z(WX1742) ) ;
AND2    gate8804  (.A(WX2508), .B(WX1744), .Z(WX1743) ) ;
OR2     gate8805  (.A(WX1757), .B(WX1756), .Z(WX1759) ) ;
AND2    gate8806  (.A(WX1759), .B(WX2296), .Z(WX1748) ) ;
OR2     gate8807  (.A(WX1753), .B(WX1752), .Z(WX1755) ) ;
AND2    gate8808  (.A(WX1755), .B(WX1750), .Z(WX1749) ) ;
AND2    gate8809  (.A(CRC_OUT_8_1), .B(WX2297), .Z(WX1752) ) ;
AND2    gate8810  (.A(WX3808), .B(WX1754), .Z(WX1753) ) ;
AND2    gate8811  (.A(WX1838), .B(WX2297), .Z(WX1756) ) ;
AND2    gate8812  (.A(WX2515), .B(WX1758), .Z(WX1757) ) ;
OR2     gate8813  (.A(WX1771), .B(WX1770), .Z(WX1773) ) ;
AND2    gate8814  (.A(WX1773), .B(WX2296), .Z(WX1762) ) ;
OR2     gate8815  (.A(WX1767), .B(WX1766), .Z(WX1769) ) ;
AND2    gate8816  (.A(WX1769), .B(WX1764), .Z(WX1763) ) ;
AND2    gate8817  (.A(CRC_OUT_8_0), .B(WX2297), .Z(WX1766) ) ;
AND2    gate8818  (.A(WX3815), .B(WX1768), .Z(WX1767) ) ;
AND2    gate8819  (.A(WX1840), .B(WX2297), .Z(WX1770) ) ;
AND2    gate8820  (.A(WX2522), .B(WX1772), .Z(WX1771) ) ;
NAND2   gate8821  (.A(II7058), .B(II7059), .Z(WX2299) ) ;
AND2    gate8822  (.A(WX2299), .B(WX2298), .Z(WX2300) ) ;
AND2    gate8823  (.A(WX1873), .B(WX2302), .Z(WX2301) ) ;
NAND2   gate8824  (.A(II7071), .B(II7072), .Z(WX2306) ) ;
AND2    gate8825  (.A(WX2306), .B(WX2298), .Z(WX2307) ) ;
AND2    gate8826  (.A(WX1874), .B(WX2309), .Z(WX2308) ) ;
NAND2   gate8827  (.A(II7084), .B(II7085), .Z(WX2313) ) ;
AND2    gate8828  (.A(WX2313), .B(WX2298), .Z(WX2314) ) ;
AND2    gate8829  (.A(WX1875), .B(WX2316), .Z(WX2315) ) ;
NAND2   gate8830  (.A(II7097), .B(II7098), .Z(WX2320) ) ;
AND2    gate8831  (.A(WX2320), .B(WX2298), .Z(WX2321) ) ;
AND2    gate8832  (.A(WX1876), .B(WX2323), .Z(WX2322) ) ;
NAND2   gate8833  (.A(II7110), .B(II7111), .Z(WX2327) ) ;
AND2    gate8834  (.A(WX2327), .B(WX2298), .Z(WX2328) ) ;
AND2    gate8835  (.A(WX1877), .B(WX2330), .Z(WX2329) ) ;
NAND2   gate8836  (.A(II7123), .B(II7124), .Z(WX2334) ) ;
AND2    gate8837  (.A(WX2334), .B(WX2298), .Z(WX2335) ) ;
AND2    gate8838  (.A(WX1878), .B(WX2337), .Z(WX2336) ) ;
NAND2   gate8839  (.A(II7136), .B(II7137), .Z(WX2341) ) ;
AND2    gate8840  (.A(WX2341), .B(WX2298), .Z(WX2342) ) ;
AND2    gate8841  (.A(WX1879), .B(WX2344), .Z(WX2343) ) ;
NAND2   gate8842  (.A(II7149), .B(II7150), .Z(WX2348) ) ;
AND2    gate8843  (.A(WX2348), .B(WX2298), .Z(WX2349) ) ;
AND2    gate8844  (.A(WX1880), .B(WX2351), .Z(WX2350) ) ;
NAND2   gate8845  (.A(II7162), .B(II7163), .Z(WX2355) ) ;
AND2    gate8846  (.A(WX2355), .B(WX2298), .Z(WX2356) ) ;
AND2    gate8847  (.A(WX1881), .B(WX2358), .Z(WX2357) ) ;
NAND2   gate8848  (.A(II7175), .B(II7176), .Z(WX2362) ) ;
AND2    gate8849  (.A(WX2362), .B(WX2298), .Z(WX2363) ) ;
AND2    gate8850  (.A(WX1882), .B(WX2365), .Z(WX2364) ) ;
NAND2   gate8851  (.A(II7188), .B(II7189), .Z(WX2369) ) ;
AND2    gate8852  (.A(WX2369), .B(WX2298), .Z(WX2370) ) ;
AND2    gate8853  (.A(WX1883), .B(WX2372), .Z(WX2371) ) ;
NAND2   gate8854  (.A(II7201), .B(II7202), .Z(WX2376) ) ;
AND2    gate8855  (.A(WX2376), .B(WX2298), .Z(WX2377) ) ;
AND2    gate8856  (.A(WX1884), .B(WX2379), .Z(WX2378) ) ;
NAND2   gate8857  (.A(II7214), .B(II7215), .Z(WX2383) ) ;
AND2    gate8858  (.A(WX2383), .B(WX2298), .Z(WX2384) ) ;
AND2    gate8859  (.A(WX1885), .B(WX2386), .Z(WX2385) ) ;
NAND2   gate8860  (.A(II7227), .B(II7228), .Z(WX2390) ) ;
AND2    gate8861  (.A(WX2390), .B(WX2298), .Z(WX2391) ) ;
AND2    gate8862  (.A(WX1886), .B(WX2393), .Z(WX2392) ) ;
NAND2   gate8863  (.A(II7240), .B(II7241), .Z(WX2397) ) ;
AND2    gate8864  (.A(WX2397), .B(WX2298), .Z(WX2398) ) ;
AND2    gate8865  (.A(WX1887), .B(WX2400), .Z(WX2399) ) ;
NAND2   gate8866  (.A(II7253), .B(II7254), .Z(WX2404) ) ;
AND2    gate8867  (.A(WX2404), .B(WX2298), .Z(WX2405) ) ;
AND2    gate8868  (.A(WX1888), .B(WX2407), .Z(WX2406) ) ;
NAND2   gate8869  (.A(II7266), .B(II7267), .Z(WX2411) ) ;
AND2    gate8870  (.A(WX2411), .B(WX2298), .Z(WX2412) ) ;
AND2    gate8871  (.A(WX1889), .B(WX2414), .Z(WX2413) ) ;
NAND2   gate8872  (.A(II7279), .B(II7280), .Z(WX2418) ) ;
AND2    gate8873  (.A(WX2418), .B(WX2298), .Z(WX2419) ) ;
AND2    gate8874  (.A(WX1890), .B(WX2421), .Z(WX2420) ) ;
NAND2   gate8875  (.A(II7292), .B(II7293), .Z(WX2425) ) ;
AND2    gate8876  (.A(WX2425), .B(WX2298), .Z(WX2426) ) ;
AND2    gate8877  (.A(WX1891), .B(WX2428), .Z(WX2427) ) ;
NAND2   gate8878  (.A(II7305), .B(II7306), .Z(WX2432) ) ;
AND2    gate8879  (.A(WX2432), .B(WX2298), .Z(WX2433) ) ;
AND2    gate8880  (.A(WX1892), .B(WX2435), .Z(WX2434) ) ;
NAND2   gate8881  (.A(II7318), .B(II7319), .Z(WX2439) ) ;
AND2    gate8882  (.A(WX2439), .B(WX2298), .Z(WX2440) ) ;
AND2    gate8883  (.A(WX1893), .B(WX2442), .Z(WX2441) ) ;
NAND2   gate8884  (.A(II7331), .B(II7332), .Z(WX2446) ) ;
AND2    gate8885  (.A(WX2446), .B(WX2298), .Z(WX2447) ) ;
AND2    gate8886  (.A(WX1894), .B(WX2449), .Z(WX2448) ) ;
NAND2   gate8887  (.A(II7344), .B(II7345), .Z(WX2453) ) ;
AND2    gate8888  (.A(WX2453), .B(WX2298), .Z(WX2454) ) ;
AND2    gate8889  (.A(WX1895), .B(WX2456), .Z(WX2455) ) ;
NAND2   gate8890  (.A(II7357), .B(II7358), .Z(WX2460) ) ;
AND2    gate8891  (.A(WX2460), .B(WX2298), .Z(WX2461) ) ;
AND2    gate8892  (.A(WX1896), .B(WX2463), .Z(WX2462) ) ;
NAND2   gate8893  (.A(II7370), .B(II7371), .Z(WX2467) ) ;
AND2    gate8894  (.A(WX2467), .B(WX2298), .Z(WX2468) ) ;
AND2    gate8895  (.A(WX1897), .B(WX2470), .Z(WX2469) ) ;
NAND2   gate8896  (.A(II7383), .B(II7384), .Z(WX2474) ) ;
AND2    gate8897  (.A(WX2474), .B(WX2298), .Z(WX2475) ) ;
AND2    gate8898  (.A(WX1898), .B(WX2477), .Z(WX2476) ) ;
NAND2   gate8899  (.A(II7396), .B(II7397), .Z(WX2481) ) ;
AND2    gate8900  (.A(WX2481), .B(WX2298), .Z(WX2482) ) ;
AND2    gate8901  (.A(WX1899), .B(WX2484), .Z(WX2483) ) ;
NAND2   gate8902  (.A(II7409), .B(II7410), .Z(WX2488) ) ;
AND2    gate8903  (.A(WX2488), .B(WX2298), .Z(WX2489) ) ;
AND2    gate8904  (.A(WX1900), .B(WX2491), .Z(WX2490) ) ;
NAND2   gate8905  (.A(II7422), .B(II7423), .Z(WX2495) ) ;
AND2    gate8906  (.A(WX2495), .B(WX2298), .Z(WX2496) ) ;
AND2    gate8907  (.A(WX1901), .B(WX2498), .Z(WX2497) ) ;
NAND2   gate8908  (.A(II7435), .B(II7436), .Z(WX2502) ) ;
AND2    gate8909  (.A(WX2502), .B(WX2298), .Z(WX2503) ) ;
AND2    gate8910  (.A(WX1902), .B(WX2505), .Z(WX2504) ) ;
NAND2   gate8911  (.A(II7448), .B(II7449), .Z(WX2509) ) ;
AND2    gate8912  (.A(WX2509), .B(WX2298), .Z(WX2510) ) ;
AND2    gate8913  (.A(WX1903), .B(WX2512), .Z(WX2511) ) ;
NAND2   gate8914  (.A(II7461), .B(II7462), .Z(WX2516) ) ;
AND2    gate8915  (.A(WX2516), .B(WX2298), .Z(WX2517) ) ;
AND2    gate8916  (.A(WX1904), .B(WX2519), .Z(WX2518) ) ;
NAND2   gate8917  (.A(II7520), .B(II7521), .Z(WX2527) ) ;
NAND2   gate8918  (.A(II7716), .B(II7717), .Z(WX2555) ) ;
NAND2   gate8919  (.A(II7709), .B(II7710), .Z(WX2554) ) ;
NAND2   gate8920  (.A(II7702), .B(II7703), .Z(WX2553) ) ;
NAND2   gate8921  (.A(II7513), .B(II7514), .Z(WX2526) ) ;
NAND2   gate8922  (.A(II7695), .B(II7696), .Z(WX2552) ) ;
NAND2   gate8923  (.A(II7688), .B(II7689), .Z(WX2551) ) ;
NAND2   gate8924  (.A(II7681), .B(II7682), .Z(WX2550) ) ;
NAND2   gate8925  (.A(II7674), .B(II7675), .Z(WX2549) ) ;
NAND2   gate8926  (.A(II7667), .B(II7668), .Z(WX2548) ) ;
NAND2   gate8927  (.A(II7660), .B(II7661), .Z(WX2547) ) ;
NAND2   gate8928  (.A(II7498), .B(II7499), .Z(WX2525) ) ;
NAND2   gate8929  (.A(II7653), .B(II7654), .Z(WX2546) ) ;
NAND2   gate8930  (.A(II7646), .B(II7647), .Z(WX2545) ) ;
NAND2   gate8931  (.A(II7639), .B(II7640), .Z(WX2544) ) ;
NAND2   gate8932  (.A(II7632), .B(II7633), .Z(WX2543) ) ;
NAND2   gate8933  (.A(II7483), .B(II7484), .Z(WX2524) ) ;
NAND2   gate8934  (.A(II7625), .B(II7626), .Z(WX2542) ) ;
NAND2   gate8935  (.A(II7618), .B(II7619), .Z(WX2541) ) ;
NAND2   gate8936  (.A(II7611), .B(II7612), .Z(WX2540) ) ;
NAND2   gate8937  (.A(II7604), .B(II7605), .Z(WX2539) ) ;
NAND2   gate8938  (.A(II7597), .B(II7598), .Z(WX2538) ) ;
NAND2   gate8939  (.A(II7590), .B(II7591), .Z(WX2537) ) ;
NAND2   gate8940  (.A(II7583), .B(II7584), .Z(WX2536) ) ;
NAND2   gate8941  (.A(II7576), .B(II7577), .Z(WX2535) ) ;
NAND2   gate8942  (.A(II7569), .B(II7570), .Z(WX2534) ) ;
NAND2   gate8943  (.A(II7562), .B(II7563), .Z(WX2533) ) ;
NAND2   gate8944  (.A(II7555), .B(II7556), .Z(WX2532) ) ;
NAND2   gate8945  (.A(II7548), .B(II7549), .Z(WX2531) ) ;
NAND2   gate8946  (.A(II7541), .B(II7542), .Z(WX2530) ) ;
NAND2   gate8947  (.A(II7534), .B(II7535), .Z(WX2529) ) ;
NAND2   gate8948  (.A(II7527), .B(II7528), .Z(WX2528) ) ;
OR2     gate8949  (.A(WX2630), .B(WX2629), .Z(WX2632) ) ;
AND2    gate8950  (.A(WX2632), .B(WX3589), .Z(WX2621) ) ;
OR2     gate8951  (.A(WX2626), .B(WX2625), .Z(WX2628) ) ;
AND2    gate8952  (.A(WX2628), .B(WX2623), .Z(WX2622) ) ;
AND2    gate8953  (.A(CRC_OUT_7_31), .B(WX3590), .Z(WX2625) ) ;
AND2    gate8954  (.A(WX4891), .B(WX2627), .Z(WX2626) ) ;
AND2    gate8955  (.A(WX3071), .B(WX3590), .Z(WX2629) ) ;
AND2    gate8956  (.A(WX3598), .B(WX2631), .Z(WX2630) ) ;
OR2     gate8957  (.A(WX2644), .B(WX2643), .Z(WX2646) ) ;
AND2    gate8958  (.A(WX2646), .B(WX3589), .Z(WX2635) ) ;
OR2     gate8959  (.A(WX2640), .B(WX2639), .Z(WX2642) ) ;
AND2    gate8960  (.A(WX2642), .B(WX2637), .Z(WX2636) ) ;
AND2    gate8961  (.A(CRC_OUT_7_30), .B(WX3590), .Z(WX2639) ) ;
AND2    gate8962  (.A(WX4898), .B(WX2641), .Z(WX2640) ) ;
AND2    gate8963  (.A(WX3073), .B(WX3590), .Z(WX2643) ) ;
AND2    gate8964  (.A(WX3605), .B(WX2645), .Z(WX2644) ) ;
OR2     gate8965  (.A(WX2658), .B(WX2657), .Z(WX2660) ) ;
AND2    gate8966  (.A(WX2660), .B(WX3589), .Z(WX2649) ) ;
OR2     gate8967  (.A(WX2654), .B(WX2653), .Z(WX2656) ) ;
AND2    gate8968  (.A(WX2656), .B(WX2651), .Z(WX2650) ) ;
AND2    gate8969  (.A(CRC_OUT_7_29), .B(WX3590), .Z(WX2653) ) ;
AND2    gate8970  (.A(WX4905), .B(WX2655), .Z(WX2654) ) ;
AND2    gate8971  (.A(WX3075), .B(WX3590), .Z(WX2657) ) ;
AND2    gate8972  (.A(WX3612), .B(WX2659), .Z(WX2658) ) ;
OR2     gate8973  (.A(WX2672), .B(WX2671), .Z(WX2674) ) ;
AND2    gate8974  (.A(WX2674), .B(WX3589), .Z(WX2663) ) ;
OR2     gate8975  (.A(WX2668), .B(WX2667), .Z(WX2670) ) ;
AND2    gate8976  (.A(WX2670), .B(WX2665), .Z(WX2664) ) ;
AND2    gate8977  (.A(CRC_OUT_7_28), .B(WX3590), .Z(WX2667) ) ;
AND2    gate8978  (.A(WX4912), .B(WX2669), .Z(WX2668) ) ;
AND2    gate8979  (.A(WX3077), .B(WX3590), .Z(WX2671) ) ;
AND2    gate8980  (.A(WX3619), .B(WX2673), .Z(WX2672) ) ;
OR2     gate8981  (.A(WX2686), .B(WX2685), .Z(WX2688) ) ;
AND2    gate8982  (.A(WX2688), .B(WX3589), .Z(WX2677) ) ;
OR2     gate8983  (.A(WX2682), .B(WX2681), .Z(WX2684) ) ;
AND2    gate8984  (.A(WX2684), .B(WX2679), .Z(WX2678) ) ;
AND2    gate8985  (.A(CRC_OUT_7_27), .B(WX3590), .Z(WX2681) ) ;
AND2    gate8986  (.A(WX4919), .B(WX2683), .Z(WX2682) ) ;
AND2    gate8987  (.A(WX3079), .B(WX3590), .Z(WX2685) ) ;
AND2    gate8988  (.A(WX3626), .B(WX2687), .Z(WX2686) ) ;
OR2     gate8989  (.A(WX2700), .B(WX2699), .Z(WX2702) ) ;
AND2    gate8990  (.A(WX2702), .B(WX3589), .Z(WX2691) ) ;
OR2     gate8991  (.A(WX2696), .B(WX2695), .Z(WX2698) ) ;
AND2    gate8992  (.A(WX2698), .B(WX2693), .Z(WX2692) ) ;
AND2    gate8993  (.A(CRC_OUT_7_26), .B(WX3590), .Z(WX2695) ) ;
AND2    gate8994  (.A(WX4926), .B(WX2697), .Z(WX2696) ) ;
AND2    gate8995  (.A(WX3081), .B(WX3590), .Z(WX2699) ) ;
AND2    gate8996  (.A(WX3633), .B(WX2701), .Z(WX2700) ) ;
OR2     gate8997  (.A(WX2714), .B(WX2713), .Z(WX2716) ) ;
AND2    gate8998  (.A(WX2716), .B(WX3589), .Z(WX2705) ) ;
OR2     gate8999  (.A(WX2710), .B(WX2709), .Z(WX2712) ) ;
AND2    gate9000  (.A(WX2712), .B(WX2707), .Z(WX2706) ) ;
AND2    gate9001  (.A(CRC_OUT_7_25), .B(WX3590), .Z(WX2709) ) ;
AND2    gate9002  (.A(WX4933), .B(WX2711), .Z(WX2710) ) ;
AND2    gate9003  (.A(WX3083), .B(WX3590), .Z(WX2713) ) ;
AND2    gate9004  (.A(WX3640), .B(WX2715), .Z(WX2714) ) ;
OR2     gate9005  (.A(WX2728), .B(WX2727), .Z(WX2730) ) ;
AND2    gate9006  (.A(WX2730), .B(WX3589), .Z(WX2719) ) ;
OR2     gate9007  (.A(WX2724), .B(WX2723), .Z(WX2726) ) ;
AND2    gate9008  (.A(WX2726), .B(WX2721), .Z(WX2720) ) ;
AND2    gate9009  (.A(CRC_OUT_7_24), .B(WX3590), .Z(WX2723) ) ;
AND2    gate9010  (.A(WX4940), .B(WX2725), .Z(WX2724) ) ;
AND2    gate9011  (.A(WX3085), .B(WX3590), .Z(WX2727) ) ;
AND2    gate9012  (.A(WX3647), .B(WX2729), .Z(WX2728) ) ;
OR2     gate9013  (.A(WX2742), .B(WX2741), .Z(WX2744) ) ;
AND2    gate9014  (.A(WX2744), .B(WX3589), .Z(WX2733) ) ;
OR2     gate9015  (.A(WX2738), .B(WX2737), .Z(WX2740) ) ;
AND2    gate9016  (.A(WX2740), .B(WX2735), .Z(WX2734) ) ;
AND2    gate9017  (.A(CRC_OUT_7_23), .B(WX3590), .Z(WX2737) ) ;
AND2    gate9018  (.A(WX4947), .B(WX2739), .Z(WX2738) ) ;
AND2    gate9019  (.A(WX3087), .B(WX3590), .Z(WX2741) ) ;
AND2    gate9020  (.A(WX3654), .B(WX2743), .Z(WX2742) ) ;
OR2     gate9021  (.A(WX2756), .B(WX2755), .Z(WX2758) ) ;
AND2    gate9022  (.A(WX2758), .B(WX3589), .Z(WX2747) ) ;
OR2     gate9023  (.A(WX2752), .B(WX2751), .Z(WX2754) ) ;
AND2    gate9024  (.A(WX2754), .B(WX2749), .Z(WX2748) ) ;
AND2    gate9025  (.A(CRC_OUT_7_22), .B(WX3590), .Z(WX2751) ) ;
AND2    gate9026  (.A(WX4954), .B(WX2753), .Z(WX2752) ) ;
AND2    gate9027  (.A(WX3089), .B(WX3590), .Z(WX2755) ) ;
AND2    gate9028  (.A(WX3661), .B(WX2757), .Z(WX2756) ) ;
OR2     gate9029  (.A(WX2770), .B(WX2769), .Z(WX2772) ) ;
AND2    gate9030  (.A(WX2772), .B(WX3589), .Z(WX2761) ) ;
OR2     gate9031  (.A(WX2766), .B(WX2765), .Z(WX2768) ) ;
AND2    gate9032  (.A(WX2768), .B(WX2763), .Z(WX2762) ) ;
AND2    gate9033  (.A(CRC_OUT_7_21), .B(WX3590), .Z(WX2765) ) ;
AND2    gate9034  (.A(WX4961), .B(WX2767), .Z(WX2766) ) ;
AND2    gate9035  (.A(WX3091), .B(WX3590), .Z(WX2769) ) ;
AND2    gate9036  (.A(WX3668), .B(WX2771), .Z(WX2770) ) ;
OR2     gate9037  (.A(WX2784), .B(WX2783), .Z(WX2786) ) ;
AND2    gate9038  (.A(WX2786), .B(WX3589), .Z(WX2775) ) ;
OR2     gate9039  (.A(WX2780), .B(WX2779), .Z(WX2782) ) ;
AND2    gate9040  (.A(WX2782), .B(WX2777), .Z(WX2776) ) ;
AND2    gate9041  (.A(CRC_OUT_7_20), .B(WX3590), .Z(WX2779) ) ;
AND2    gate9042  (.A(WX4968), .B(WX2781), .Z(WX2780) ) ;
AND2    gate9043  (.A(WX3093), .B(WX3590), .Z(WX2783) ) ;
AND2    gate9044  (.A(WX3675), .B(WX2785), .Z(WX2784) ) ;
OR2     gate9045  (.A(WX2798), .B(WX2797), .Z(WX2800) ) ;
AND2    gate9046  (.A(WX2800), .B(WX3589), .Z(WX2789) ) ;
OR2     gate9047  (.A(WX2794), .B(WX2793), .Z(WX2796) ) ;
AND2    gate9048  (.A(WX2796), .B(WX2791), .Z(WX2790) ) ;
AND2    gate9049  (.A(CRC_OUT_7_19), .B(WX3590), .Z(WX2793) ) ;
AND2    gate9050  (.A(WX4975), .B(WX2795), .Z(WX2794) ) ;
AND2    gate9051  (.A(WX3095), .B(WX3590), .Z(WX2797) ) ;
AND2    gate9052  (.A(WX3682), .B(WX2799), .Z(WX2798) ) ;
OR2     gate9053  (.A(WX2812), .B(WX2811), .Z(WX2814) ) ;
AND2    gate9054  (.A(WX2814), .B(WX3589), .Z(WX2803) ) ;
OR2     gate9055  (.A(WX2808), .B(WX2807), .Z(WX2810) ) ;
AND2    gate9056  (.A(WX2810), .B(WX2805), .Z(WX2804) ) ;
AND2    gate9057  (.A(CRC_OUT_7_18), .B(WX3590), .Z(WX2807) ) ;
AND2    gate9058  (.A(WX4982), .B(WX2809), .Z(WX2808) ) ;
AND2    gate9059  (.A(WX3097), .B(WX3590), .Z(WX2811) ) ;
AND2    gate9060  (.A(WX3689), .B(WX2813), .Z(WX2812) ) ;
OR2     gate9061  (.A(WX2826), .B(WX2825), .Z(WX2828) ) ;
AND2    gate9062  (.A(WX2828), .B(WX3589), .Z(WX2817) ) ;
OR2     gate9063  (.A(WX2822), .B(WX2821), .Z(WX2824) ) ;
AND2    gate9064  (.A(WX2824), .B(WX2819), .Z(WX2818) ) ;
AND2    gate9065  (.A(CRC_OUT_7_17), .B(WX3590), .Z(WX2821) ) ;
AND2    gate9066  (.A(WX4989), .B(WX2823), .Z(WX2822) ) ;
AND2    gate9067  (.A(WX3099), .B(WX3590), .Z(WX2825) ) ;
AND2    gate9068  (.A(WX3696), .B(WX2827), .Z(WX2826) ) ;
OR2     gate9069  (.A(WX2840), .B(WX2839), .Z(WX2842) ) ;
AND2    gate9070  (.A(WX2842), .B(WX3589), .Z(WX2831) ) ;
OR2     gate9071  (.A(WX2836), .B(WX2835), .Z(WX2838) ) ;
AND2    gate9072  (.A(WX2838), .B(WX2833), .Z(WX2832) ) ;
AND2    gate9073  (.A(CRC_OUT_7_16), .B(WX3590), .Z(WX2835) ) ;
AND2    gate9074  (.A(WX4996), .B(WX2837), .Z(WX2836) ) ;
AND2    gate9075  (.A(WX3101), .B(WX3590), .Z(WX2839) ) ;
AND2    gate9076  (.A(WX3703), .B(WX2841), .Z(WX2840) ) ;
OR2     gate9077  (.A(WX2854), .B(WX2853), .Z(WX2856) ) ;
AND2    gate9078  (.A(WX2856), .B(WX3589), .Z(WX2845) ) ;
OR2     gate9079  (.A(WX2850), .B(WX2849), .Z(WX2852) ) ;
AND2    gate9080  (.A(WX2852), .B(WX2847), .Z(WX2846) ) ;
AND2    gate9081  (.A(CRC_OUT_7_15), .B(WX3590), .Z(WX2849) ) ;
AND2    gate9082  (.A(WX5003), .B(WX2851), .Z(WX2850) ) ;
AND2    gate9083  (.A(WX3103), .B(WX3590), .Z(WX2853) ) ;
AND2    gate9084  (.A(WX3710), .B(WX2855), .Z(WX2854) ) ;
OR2     gate9085  (.A(WX2868), .B(WX2867), .Z(WX2870) ) ;
AND2    gate9086  (.A(WX2870), .B(WX3589), .Z(WX2859) ) ;
OR2     gate9087  (.A(WX2864), .B(WX2863), .Z(WX2866) ) ;
AND2    gate9088  (.A(WX2866), .B(WX2861), .Z(WX2860) ) ;
AND2    gate9089  (.A(CRC_OUT_7_14), .B(WX3590), .Z(WX2863) ) ;
AND2    gate9090  (.A(WX5010), .B(WX2865), .Z(WX2864) ) ;
AND2    gate9091  (.A(WX3105), .B(WX3590), .Z(WX2867) ) ;
AND2    gate9092  (.A(WX3717), .B(WX2869), .Z(WX2868) ) ;
OR2     gate9093  (.A(WX2882), .B(WX2881), .Z(WX2884) ) ;
AND2    gate9094  (.A(WX2884), .B(WX3589), .Z(WX2873) ) ;
OR2     gate9095  (.A(WX2878), .B(WX2877), .Z(WX2880) ) ;
AND2    gate9096  (.A(WX2880), .B(WX2875), .Z(WX2874) ) ;
AND2    gate9097  (.A(CRC_OUT_7_13), .B(WX3590), .Z(WX2877) ) ;
AND2    gate9098  (.A(WX5017), .B(WX2879), .Z(WX2878) ) ;
AND2    gate9099  (.A(WX3107), .B(WX3590), .Z(WX2881) ) ;
AND2    gate9100  (.A(WX3724), .B(WX2883), .Z(WX2882) ) ;
OR2     gate9101  (.A(WX2896), .B(WX2895), .Z(WX2898) ) ;
AND2    gate9102  (.A(WX2898), .B(WX3589), .Z(WX2887) ) ;
OR2     gate9103  (.A(WX2892), .B(WX2891), .Z(WX2894) ) ;
AND2    gate9104  (.A(WX2894), .B(WX2889), .Z(WX2888) ) ;
AND2    gate9105  (.A(CRC_OUT_7_12), .B(WX3590), .Z(WX2891) ) ;
AND2    gate9106  (.A(WX5024), .B(WX2893), .Z(WX2892) ) ;
AND2    gate9107  (.A(WX3109), .B(WX3590), .Z(WX2895) ) ;
AND2    gate9108  (.A(WX3731), .B(WX2897), .Z(WX2896) ) ;
OR2     gate9109  (.A(WX2910), .B(WX2909), .Z(WX2912) ) ;
AND2    gate9110  (.A(WX2912), .B(WX3589), .Z(WX2901) ) ;
OR2     gate9111  (.A(WX2906), .B(WX2905), .Z(WX2908) ) ;
AND2    gate9112  (.A(WX2908), .B(WX2903), .Z(WX2902) ) ;
AND2    gate9113  (.A(CRC_OUT_7_11), .B(WX3590), .Z(WX2905) ) ;
AND2    gate9114  (.A(WX5031), .B(WX2907), .Z(WX2906) ) ;
AND2    gate9115  (.A(WX3111), .B(WX3590), .Z(WX2909) ) ;
AND2    gate9116  (.A(WX3738), .B(WX2911), .Z(WX2910) ) ;
OR2     gate9117  (.A(WX2924), .B(WX2923), .Z(WX2926) ) ;
AND2    gate9118  (.A(WX2926), .B(WX3589), .Z(WX2915) ) ;
OR2     gate9119  (.A(WX2920), .B(WX2919), .Z(WX2922) ) ;
AND2    gate9120  (.A(WX2922), .B(WX2917), .Z(WX2916) ) ;
AND2    gate9121  (.A(CRC_OUT_7_10), .B(WX3590), .Z(WX2919) ) ;
AND2    gate9122  (.A(WX5038), .B(WX2921), .Z(WX2920) ) ;
AND2    gate9123  (.A(WX3113), .B(WX3590), .Z(WX2923) ) ;
AND2    gate9124  (.A(WX3745), .B(WX2925), .Z(WX2924) ) ;
OR2     gate9125  (.A(WX2938), .B(WX2937), .Z(WX2940) ) ;
AND2    gate9126  (.A(WX2940), .B(WX3589), .Z(WX2929) ) ;
OR2     gate9127  (.A(WX2934), .B(WX2933), .Z(WX2936) ) ;
AND2    gate9128  (.A(WX2936), .B(WX2931), .Z(WX2930) ) ;
AND2    gate9129  (.A(CRC_OUT_7_9), .B(WX3590), .Z(WX2933) ) ;
AND2    gate9130  (.A(WX5045), .B(WX2935), .Z(WX2934) ) ;
AND2    gate9131  (.A(WX3115), .B(WX3590), .Z(WX2937) ) ;
AND2    gate9132  (.A(WX3752), .B(WX2939), .Z(WX2938) ) ;
OR2     gate9133  (.A(WX2952), .B(WX2951), .Z(WX2954) ) ;
AND2    gate9134  (.A(WX2954), .B(WX3589), .Z(WX2943) ) ;
OR2     gate9135  (.A(WX2948), .B(WX2947), .Z(WX2950) ) ;
AND2    gate9136  (.A(WX2950), .B(WX2945), .Z(WX2944) ) ;
AND2    gate9137  (.A(CRC_OUT_7_8), .B(WX3590), .Z(WX2947) ) ;
AND2    gate9138  (.A(WX5052), .B(WX2949), .Z(WX2948) ) ;
AND2    gate9139  (.A(WX3117), .B(WX3590), .Z(WX2951) ) ;
AND2    gate9140  (.A(WX3759), .B(WX2953), .Z(WX2952) ) ;
OR2     gate9141  (.A(WX2966), .B(WX2965), .Z(WX2968) ) ;
AND2    gate9142  (.A(WX2968), .B(WX3589), .Z(WX2957) ) ;
OR2     gate9143  (.A(WX2962), .B(WX2961), .Z(WX2964) ) ;
AND2    gate9144  (.A(WX2964), .B(WX2959), .Z(WX2958) ) ;
AND2    gate9145  (.A(CRC_OUT_7_7), .B(WX3590), .Z(WX2961) ) ;
AND2    gate9146  (.A(WX5059), .B(WX2963), .Z(WX2962) ) ;
AND2    gate9147  (.A(WX3119), .B(WX3590), .Z(WX2965) ) ;
AND2    gate9148  (.A(WX3766), .B(WX2967), .Z(WX2966) ) ;
OR2     gate9149  (.A(WX2980), .B(WX2979), .Z(WX2982) ) ;
AND2    gate9150  (.A(WX2982), .B(WX3589), .Z(WX2971) ) ;
OR2     gate9151  (.A(WX2976), .B(WX2975), .Z(WX2978) ) ;
AND2    gate9152  (.A(WX2978), .B(WX2973), .Z(WX2972) ) ;
AND2    gate9153  (.A(CRC_OUT_7_6), .B(WX3590), .Z(WX2975) ) ;
AND2    gate9154  (.A(WX5066), .B(WX2977), .Z(WX2976) ) ;
AND2    gate9155  (.A(WX3121), .B(WX3590), .Z(WX2979) ) ;
AND2    gate9156  (.A(WX3773), .B(WX2981), .Z(WX2980) ) ;
OR2     gate9157  (.A(WX2994), .B(WX2993), .Z(WX2996) ) ;
AND2    gate9158  (.A(WX2996), .B(WX3589), .Z(WX2985) ) ;
OR2     gate9159  (.A(WX2990), .B(WX2989), .Z(WX2992) ) ;
AND2    gate9160  (.A(WX2992), .B(WX2987), .Z(WX2986) ) ;
AND2    gate9161  (.A(CRC_OUT_7_5), .B(WX3590), .Z(WX2989) ) ;
AND2    gate9162  (.A(WX5073), .B(WX2991), .Z(WX2990) ) ;
AND2    gate9163  (.A(WX3123), .B(WX3590), .Z(WX2993) ) ;
AND2    gate9164  (.A(WX3780), .B(WX2995), .Z(WX2994) ) ;
OR2     gate9165  (.A(WX3008), .B(WX3007), .Z(WX3010) ) ;
AND2    gate9166  (.A(WX3010), .B(WX3589), .Z(WX2999) ) ;
OR2     gate9167  (.A(WX3004), .B(WX3003), .Z(WX3006) ) ;
AND2    gate9168  (.A(WX3006), .B(WX3001), .Z(WX3000) ) ;
AND2    gate9169  (.A(CRC_OUT_7_4), .B(WX3590), .Z(WX3003) ) ;
AND2    gate9170  (.A(WX5080), .B(WX3005), .Z(WX3004) ) ;
AND2    gate9171  (.A(WX3125), .B(WX3590), .Z(WX3007) ) ;
AND2    gate9172  (.A(WX3787), .B(WX3009), .Z(WX3008) ) ;
OR2     gate9173  (.A(WX3022), .B(WX3021), .Z(WX3024) ) ;
AND2    gate9174  (.A(WX3024), .B(WX3589), .Z(WX3013) ) ;
OR2     gate9175  (.A(WX3018), .B(WX3017), .Z(WX3020) ) ;
AND2    gate9176  (.A(WX3020), .B(WX3015), .Z(WX3014) ) ;
AND2    gate9177  (.A(CRC_OUT_7_3), .B(WX3590), .Z(WX3017) ) ;
AND2    gate9178  (.A(WX5087), .B(WX3019), .Z(WX3018) ) ;
AND2    gate9179  (.A(WX3127), .B(WX3590), .Z(WX3021) ) ;
AND2    gate9180  (.A(WX3794), .B(WX3023), .Z(WX3022) ) ;
OR2     gate9181  (.A(WX3036), .B(WX3035), .Z(WX3038) ) ;
AND2    gate9182  (.A(WX3038), .B(WX3589), .Z(WX3027) ) ;
OR2     gate9183  (.A(WX3032), .B(WX3031), .Z(WX3034) ) ;
AND2    gate9184  (.A(WX3034), .B(WX3029), .Z(WX3028) ) ;
AND2    gate9185  (.A(CRC_OUT_7_2), .B(WX3590), .Z(WX3031) ) ;
AND2    gate9186  (.A(WX5094), .B(WX3033), .Z(WX3032) ) ;
AND2    gate9187  (.A(WX3129), .B(WX3590), .Z(WX3035) ) ;
AND2    gate9188  (.A(WX3801), .B(WX3037), .Z(WX3036) ) ;
OR2     gate9189  (.A(WX3050), .B(WX3049), .Z(WX3052) ) ;
AND2    gate9190  (.A(WX3052), .B(WX3589), .Z(WX3041) ) ;
OR2     gate9191  (.A(WX3046), .B(WX3045), .Z(WX3048) ) ;
AND2    gate9192  (.A(WX3048), .B(WX3043), .Z(WX3042) ) ;
AND2    gate9193  (.A(CRC_OUT_7_1), .B(WX3590), .Z(WX3045) ) ;
AND2    gate9194  (.A(WX5101), .B(WX3047), .Z(WX3046) ) ;
AND2    gate9195  (.A(WX3131), .B(WX3590), .Z(WX3049) ) ;
AND2    gate9196  (.A(WX3808), .B(WX3051), .Z(WX3050) ) ;
OR2     gate9197  (.A(WX3064), .B(WX3063), .Z(WX3066) ) ;
AND2    gate9198  (.A(WX3066), .B(WX3589), .Z(WX3055) ) ;
OR2     gate9199  (.A(WX3060), .B(WX3059), .Z(WX3062) ) ;
AND2    gate9200  (.A(WX3062), .B(WX3057), .Z(WX3056) ) ;
AND2    gate9201  (.A(CRC_OUT_7_0), .B(WX3590), .Z(WX3059) ) ;
AND2    gate9202  (.A(WX5108), .B(WX3061), .Z(WX3060) ) ;
AND2    gate9203  (.A(WX3133), .B(WX3590), .Z(WX3063) ) ;
AND2    gate9204  (.A(WX3815), .B(WX3065), .Z(WX3064) ) ;
NAND2   gate9205  (.A(II11063), .B(II11064), .Z(WX3592) ) ;
AND2    gate9206  (.A(WX3592), .B(WX3591), .Z(WX3593) ) ;
AND2    gate9207  (.A(WX3166), .B(WX3595), .Z(WX3594) ) ;
NAND2   gate9208  (.A(II11076), .B(II11077), .Z(WX3599) ) ;
AND2    gate9209  (.A(WX3599), .B(WX3591), .Z(WX3600) ) ;
AND2    gate9210  (.A(WX3167), .B(WX3602), .Z(WX3601) ) ;
NAND2   gate9211  (.A(II11089), .B(II11090), .Z(WX3606) ) ;
AND2    gate9212  (.A(WX3606), .B(WX3591), .Z(WX3607) ) ;
AND2    gate9213  (.A(WX3168), .B(WX3609), .Z(WX3608) ) ;
NAND2   gate9214  (.A(II11102), .B(II11103), .Z(WX3613) ) ;
AND2    gate9215  (.A(WX3613), .B(WX3591), .Z(WX3614) ) ;
AND2    gate9216  (.A(WX3169), .B(WX3616), .Z(WX3615) ) ;
NAND2   gate9217  (.A(II11115), .B(II11116), .Z(WX3620) ) ;
AND2    gate9218  (.A(WX3620), .B(WX3591), .Z(WX3621) ) ;
AND2    gate9219  (.A(WX3170), .B(WX3623), .Z(WX3622) ) ;
NAND2   gate9220  (.A(II11128), .B(II11129), .Z(WX3627) ) ;
AND2    gate9221  (.A(WX3627), .B(WX3591), .Z(WX3628) ) ;
AND2    gate9222  (.A(WX3171), .B(WX3630), .Z(WX3629) ) ;
NAND2   gate9223  (.A(II11141), .B(II11142), .Z(WX3634) ) ;
AND2    gate9224  (.A(WX3634), .B(WX3591), .Z(WX3635) ) ;
AND2    gate9225  (.A(WX3172), .B(WX3637), .Z(WX3636) ) ;
NAND2   gate9226  (.A(II11154), .B(II11155), .Z(WX3641) ) ;
AND2    gate9227  (.A(WX3641), .B(WX3591), .Z(WX3642) ) ;
AND2    gate9228  (.A(WX3173), .B(WX3644), .Z(WX3643) ) ;
NAND2   gate9229  (.A(II11167), .B(II11168), .Z(WX3648) ) ;
AND2    gate9230  (.A(WX3648), .B(WX3591), .Z(WX3649) ) ;
AND2    gate9231  (.A(WX3174), .B(WX3651), .Z(WX3650) ) ;
NAND2   gate9232  (.A(II11180), .B(II11181), .Z(WX3655) ) ;
AND2    gate9233  (.A(WX3655), .B(WX3591), .Z(WX3656) ) ;
AND2    gate9234  (.A(WX3175), .B(WX3658), .Z(WX3657) ) ;
NAND2   gate9235  (.A(II11193), .B(II11194), .Z(WX3662) ) ;
AND2    gate9236  (.A(WX3662), .B(WX3591), .Z(WX3663) ) ;
AND2    gate9237  (.A(WX3176), .B(WX3665), .Z(WX3664) ) ;
NAND2   gate9238  (.A(II11206), .B(II11207), .Z(WX3669) ) ;
AND2    gate9239  (.A(WX3669), .B(WX3591), .Z(WX3670) ) ;
AND2    gate9240  (.A(WX3177), .B(WX3672), .Z(WX3671) ) ;
NAND2   gate9241  (.A(II11219), .B(II11220), .Z(WX3676) ) ;
AND2    gate9242  (.A(WX3676), .B(WX3591), .Z(WX3677) ) ;
AND2    gate9243  (.A(WX3178), .B(WX3679), .Z(WX3678) ) ;
NAND2   gate9244  (.A(II11232), .B(II11233), .Z(WX3683) ) ;
AND2    gate9245  (.A(WX3683), .B(WX3591), .Z(WX3684) ) ;
AND2    gate9246  (.A(WX3179), .B(WX3686), .Z(WX3685) ) ;
NAND2   gate9247  (.A(II11245), .B(II11246), .Z(WX3690) ) ;
AND2    gate9248  (.A(WX3690), .B(WX3591), .Z(WX3691) ) ;
AND2    gate9249  (.A(WX3180), .B(WX3693), .Z(WX3692) ) ;
NAND2   gate9250  (.A(II11258), .B(II11259), .Z(WX3697) ) ;
AND2    gate9251  (.A(WX3697), .B(WX3591), .Z(WX3698) ) ;
AND2    gate9252  (.A(WX3181), .B(WX3700), .Z(WX3699) ) ;
NAND2   gate9253  (.A(II11271), .B(II11272), .Z(WX3704) ) ;
AND2    gate9254  (.A(WX3704), .B(WX3591), .Z(WX3705) ) ;
AND2    gate9255  (.A(WX3182), .B(WX3707), .Z(WX3706) ) ;
NAND2   gate9256  (.A(II11284), .B(II11285), .Z(WX3711) ) ;
AND2    gate9257  (.A(WX3711), .B(WX3591), .Z(WX3712) ) ;
AND2    gate9258  (.A(WX3183), .B(WX3714), .Z(WX3713) ) ;
NAND2   gate9259  (.A(II11297), .B(II11298), .Z(WX3718) ) ;
AND2    gate9260  (.A(WX3718), .B(WX3591), .Z(WX3719) ) ;
AND2    gate9261  (.A(WX3184), .B(WX3721), .Z(WX3720) ) ;
NAND2   gate9262  (.A(II11310), .B(II11311), .Z(WX3725) ) ;
AND2    gate9263  (.A(WX3725), .B(WX3591), .Z(WX3726) ) ;
AND2    gate9264  (.A(WX3185), .B(WX3728), .Z(WX3727) ) ;
NAND2   gate9265  (.A(II11323), .B(II11324), .Z(WX3732) ) ;
AND2    gate9266  (.A(WX3732), .B(WX3591), .Z(WX3733) ) ;
AND2    gate9267  (.A(WX3186), .B(WX3735), .Z(WX3734) ) ;
NAND2   gate9268  (.A(II11336), .B(II11337), .Z(WX3739) ) ;
AND2    gate9269  (.A(WX3739), .B(WX3591), .Z(WX3740) ) ;
AND2    gate9270  (.A(WX3187), .B(WX3742), .Z(WX3741) ) ;
NAND2   gate9271  (.A(II11349), .B(II11350), .Z(WX3746) ) ;
AND2    gate9272  (.A(WX3746), .B(WX3591), .Z(WX3747) ) ;
AND2    gate9273  (.A(WX3188), .B(WX3749), .Z(WX3748) ) ;
NAND2   gate9274  (.A(II11362), .B(II11363), .Z(WX3753) ) ;
AND2    gate9275  (.A(WX3753), .B(WX3591), .Z(WX3754) ) ;
AND2    gate9276  (.A(WX3189), .B(WX3756), .Z(WX3755) ) ;
NAND2   gate9277  (.A(II11375), .B(II11376), .Z(WX3760) ) ;
AND2    gate9278  (.A(WX3760), .B(WX3591), .Z(WX3761) ) ;
AND2    gate9279  (.A(WX3190), .B(WX3763), .Z(WX3762) ) ;
NAND2   gate9280  (.A(II11388), .B(II11389), .Z(WX3767) ) ;
AND2    gate9281  (.A(WX3767), .B(WX3591), .Z(WX3768) ) ;
AND2    gate9282  (.A(WX3191), .B(WX3770), .Z(WX3769) ) ;
NAND2   gate9283  (.A(II11401), .B(II11402), .Z(WX3774) ) ;
AND2    gate9284  (.A(WX3774), .B(WX3591), .Z(WX3775) ) ;
AND2    gate9285  (.A(WX3192), .B(WX3777), .Z(WX3776) ) ;
NAND2   gate9286  (.A(II11414), .B(II11415), .Z(WX3781) ) ;
AND2    gate9287  (.A(WX3781), .B(WX3591), .Z(WX3782) ) ;
AND2    gate9288  (.A(WX3193), .B(WX3784), .Z(WX3783) ) ;
NAND2   gate9289  (.A(II11427), .B(II11428), .Z(WX3788) ) ;
AND2    gate9290  (.A(WX3788), .B(WX3591), .Z(WX3789) ) ;
AND2    gate9291  (.A(WX3194), .B(WX3791), .Z(WX3790) ) ;
NAND2   gate9292  (.A(II11440), .B(II11441), .Z(WX3795) ) ;
AND2    gate9293  (.A(WX3795), .B(WX3591), .Z(WX3796) ) ;
AND2    gate9294  (.A(WX3195), .B(WX3798), .Z(WX3797) ) ;
NAND2   gate9295  (.A(II11453), .B(II11454), .Z(WX3802) ) ;
AND2    gate9296  (.A(WX3802), .B(WX3591), .Z(WX3803) ) ;
AND2    gate9297  (.A(WX3196), .B(WX3805), .Z(WX3804) ) ;
NAND2   gate9298  (.A(II11466), .B(II11467), .Z(WX3809) ) ;
AND2    gate9299  (.A(WX3809), .B(WX3591), .Z(WX3810) ) ;
AND2    gate9300  (.A(WX3197), .B(WX3812), .Z(WX3811) ) ;
NAND2   gate9301  (.A(II11525), .B(II11526), .Z(WX3820) ) ;
NAND2   gate9302  (.A(II11721), .B(II11722), .Z(WX3848) ) ;
NAND2   gate9303  (.A(II11714), .B(II11715), .Z(WX3847) ) ;
NAND2   gate9304  (.A(II11707), .B(II11708), .Z(WX3846) ) ;
NAND2   gate9305  (.A(II11518), .B(II11519), .Z(WX3819) ) ;
NAND2   gate9306  (.A(II11700), .B(II11701), .Z(WX3845) ) ;
NAND2   gate9307  (.A(II11693), .B(II11694), .Z(WX3844) ) ;
NAND2   gate9308  (.A(II11686), .B(II11687), .Z(WX3843) ) ;
NAND2   gate9309  (.A(II11679), .B(II11680), .Z(WX3842) ) ;
NAND2   gate9310  (.A(II11672), .B(II11673), .Z(WX3841) ) ;
NAND2   gate9311  (.A(II11665), .B(II11666), .Z(WX3840) ) ;
NAND2   gate9312  (.A(II11503), .B(II11504), .Z(WX3818) ) ;
NAND2   gate9313  (.A(II11658), .B(II11659), .Z(WX3839) ) ;
NAND2   gate9314  (.A(II11651), .B(II11652), .Z(WX3838) ) ;
NAND2   gate9315  (.A(II11644), .B(II11645), .Z(WX3837) ) ;
NAND2   gate9316  (.A(II11637), .B(II11638), .Z(WX3836) ) ;
NAND2   gate9317  (.A(II11488), .B(II11489), .Z(WX3817) ) ;
NAND2   gate9318  (.A(II11630), .B(II11631), .Z(WX3835) ) ;
NAND2   gate9319  (.A(II11623), .B(II11624), .Z(WX3834) ) ;
NAND2   gate9320  (.A(II11616), .B(II11617), .Z(WX3833) ) ;
NAND2   gate9321  (.A(II11609), .B(II11610), .Z(WX3832) ) ;
NAND2   gate9322  (.A(II11602), .B(II11603), .Z(WX3831) ) ;
NAND2   gate9323  (.A(II11595), .B(II11596), .Z(WX3830) ) ;
NAND2   gate9324  (.A(II11588), .B(II11589), .Z(WX3829) ) ;
NAND2   gate9325  (.A(II11581), .B(II11582), .Z(WX3828) ) ;
NAND2   gate9326  (.A(II11574), .B(II11575), .Z(WX3827) ) ;
NAND2   gate9327  (.A(II11567), .B(II11568), .Z(WX3826) ) ;
NAND2   gate9328  (.A(II11560), .B(II11561), .Z(WX3825) ) ;
NAND2   gate9329  (.A(II11553), .B(II11554), .Z(WX3824) ) ;
NAND2   gate9330  (.A(II11546), .B(II11547), .Z(WX3823) ) ;
NAND2   gate9331  (.A(II11539), .B(II11540), .Z(WX3822) ) ;
NAND2   gate9332  (.A(II11532), .B(II11533), .Z(WX3821) ) ;
OR2     gate9333  (.A(WX3923), .B(WX3922), .Z(WX3925) ) ;
AND2    gate9334  (.A(WX3925), .B(WX4882), .Z(WX3914) ) ;
OR2     gate9335  (.A(WX3919), .B(WX3918), .Z(WX3921) ) ;
AND2    gate9336  (.A(WX3921), .B(WX3916), .Z(WX3915) ) ;
AND2    gate9337  (.A(CRC_OUT_6_31), .B(WX4883), .Z(WX3918) ) ;
AND2    gate9338  (.A(WX6184), .B(WX3920), .Z(WX3919) ) ;
AND2    gate9339  (.A(WX4364), .B(WX4883), .Z(WX3922) ) ;
AND2    gate9340  (.A(WX4891), .B(WX3924), .Z(WX3923) ) ;
OR2     gate9341  (.A(WX3937), .B(WX3936), .Z(WX3939) ) ;
AND2    gate9342  (.A(WX3939), .B(WX4882), .Z(WX3928) ) ;
OR2     gate9343  (.A(WX3933), .B(WX3932), .Z(WX3935) ) ;
AND2    gate9344  (.A(WX3935), .B(WX3930), .Z(WX3929) ) ;
AND2    gate9345  (.A(CRC_OUT_6_30), .B(WX4883), .Z(WX3932) ) ;
AND2    gate9346  (.A(WX6191), .B(WX3934), .Z(WX3933) ) ;
AND2    gate9347  (.A(WX4366), .B(WX4883), .Z(WX3936) ) ;
AND2    gate9348  (.A(WX4898), .B(WX3938), .Z(WX3937) ) ;
OR2     gate9349  (.A(WX3951), .B(WX3950), .Z(WX3953) ) ;
AND2    gate9350  (.A(WX3953), .B(WX4882), .Z(WX3942) ) ;
OR2     gate9351  (.A(WX3947), .B(WX3946), .Z(WX3949) ) ;
AND2    gate9352  (.A(WX3949), .B(WX3944), .Z(WX3943) ) ;
AND2    gate9353  (.A(CRC_OUT_6_29), .B(WX4883), .Z(WX3946) ) ;
AND2    gate9354  (.A(WX6198), .B(WX3948), .Z(WX3947) ) ;
AND2    gate9355  (.A(WX4368), .B(WX4883), .Z(WX3950) ) ;
AND2    gate9356  (.A(WX4905), .B(WX3952), .Z(WX3951) ) ;
OR2     gate9357  (.A(WX3965), .B(WX3964), .Z(WX3967) ) ;
AND2    gate9358  (.A(WX3967), .B(WX4882), .Z(WX3956) ) ;
OR2     gate9359  (.A(WX3961), .B(WX3960), .Z(WX3963) ) ;
AND2    gate9360  (.A(WX3963), .B(WX3958), .Z(WX3957) ) ;
AND2    gate9361  (.A(CRC_OUT_6_28), .B(WX4883), .Z(WX3960) ) ;
AND2    gate9362  (.A(WX6205), .B(WX3962), .Z(WX3961) ) ;
AND2    gate9363  (.A(WX4370), .B(WX4883), .Z(WX3964) ) ;
AND2    gate9364  (.A(WX4912), .B(WX3966), .Z(WX3965) ) ;
OR2     gate9365  (.A(WX3979), .B(WX3978), .Z(WX3981) ) ;
AND2    gate9366  (.A(WX3981), .B(WX4882), .Z(WX3970) ) ;
OR2     gate9367  (.A(WX3975), .B(WX3974), .Z(WX3977) ) ;
AND2    gate9368  (.A(WX3977), .B(WX3972), .Z(WX3971) ) ;
AND2    gate9369  (.A(CRC_OUT_6_27), .B(WX4883), .Z(WX3974) ) ;
AND2    gate9370  (.A(WX6212), .B(WX3976), .Z(WX3975) ) ;
AND2    gate9371  (.A(WX4372), .B(WX4883), .Z(WX3978) ) ;
AND2    gate9372  (.A(WX4919), .B(WX3980), .Z(WX3979) ) ;
OR2     gate9373  (.A(WX3993), .B(WX3992), .Z(WX3995) ) ;
AND2    gate9374  (.A(WX3995), .B(WX4882), .Z(WX3984) ) ;
OR2     gate9375  (.A(WX3989), .B(WX3988), .Z(WX3991) ) ;
AND2    gate9376  (.A(WX3991), .B(WX3986), .Z(WX3985) ) ;
AND2    gate9377  (.A(CRC_OUT_6_26), .B(WX4883), .Z(WX3988) ) ;
AND2    gate9378  (.A(WX6219), .B(WX3990), .Z(WX3989) ) ;
AND2    gate9379  (.A(WX4374), .B(WX4883), .Z(WX3992) ) ;
AND2    gate9380  (.A(WX4926), .B(WX3994), .Z(WX3993) ) ;
OR2     gate9381  (.A(WX4007), .B(WX4006), .Z(WX4009) ) ;
AND2    gate9382  (.A(WX4009), .B(WX4882), .Z(WX3998) ) ;
OR2     gate9383  (.A(WX4003), .B(WX4002), .Z(WX4005) ) ;
AND2    gate9384  (.A(WX4005), .B(WX4000), .Z(WX3999) ) ;
AND2    gate9385  (.A(CRC_OUT_6_25), .B(WX4883), .Z(WX4002) ) ;
AND2    gate9386  (.A(WX6226), .B(WX4004), .Z(WX4003) ) ;
AND2    gate9387  (.A(WX4376), .B(WX4883), .Z(WX4006) ) ;
AND2    gate9388  (.A(WX4933), .B(WX4008), .Z(WX4007) ) ;
OR2     gate9389  (.A(WX4021), .B(WX4020), .Z(WX4023) ) ;
AND2    gate9390  (.A(WX4023), .B(WX4882), .Z(WX4012) ) ;
OR2     gate9391  (.A(WX4017), .B(WX4016), .Z(WX4019) ) ;
AND2    gate9392  (.A(WX4019), .B(WX4014), .Z(WX4013) ) ;
AND2    gate9393  (.A(CRC_OUT_6_24), .B(WX4883), .Z(WX4016) ) ;
AND2    gate9394  (.A(WX6233), .B(WX4018), .Z(WX4017) ) ;
AND2    gate9395  (.A(WX4378), .B(WX4883), .Z(WX4020) ) ;
AND2    gate9396  (.A(WX4940), .B(WX4022), .Z(WX4021) ) ;
OR2     gate9397  (.A(WX4035), .B(WX4034), .Z(WX4037) ) ;
AND2    gate9398  (.A(WX4037), .B(WX4882), .Z(WX4026) ) ;
OR2     gate9399  (.A(WX4031), .B(WX4030), .Z(WX4033) ) ;
AND2    gate9400  (.A(WX4033), .B(WX4028), .Z(WX4027) ) ;
AND2    gate9401  (.A(CRC_OUT_6_23), .B(WX4883), .Z(WX4030) ) ;
AND2    gate9402  (.A(WX6240), .B(WX4032), .Z(WX4031) ) ;
AND2    gate9403  (.A(WX4380), .B(WX4883), .Z(WX4034) ) ;
AND2    gate9404  (.A(WX4947), .B(WX4036), .Z(WX4035) ) ;
OR2     gate9405  (.A(WX4049), .B(WX4048), .Z(WX4051) ) ;
AND2    gate9406  (.A(WX4051), .B(WX4882), .Z(WX4040) ) ;
OR2     gate9407  (.A(WX4045), .B(WX4044), .Z(WX4047) ) ;
AND2    gate9408  (.A(WX4047), .B(WX4042), .Z(WX4041) ) ;
AND2    gate9409  (.A(CRC_OUT_6_22), .B(WX4883), .Z(WX4044) ) ;
AND2    gate9410  (.A(WX6247), .B(WX4046), .Z(WX4045) ) ;
AND2    gate9411  (.A(WX4382), .B(WX4883), .Z(WX4048) ) ;
AND2    gate9412  (.A(WX4954), .B(WX4050), .Z(WX4049) ) ;
OR2     gate9413  (.A(WX4063), .B(WX4062), .Z(WX4065) ) ;
AND2    gate9414  (.A(WX4065), .B(WX4882), .Z(WX4054) ) ;
OR2     gate9415  (.A(WX4059), .B(WX4058), .Z(WX4061) ) ;
AND2    gate9416  (.A(WX4061), .B(WX4056), .Z(WX4055) ) ;
AND2    gate9417  (.A(CRC_OUT_6_21), .B(WX4883), .Z(WX4058) ) ;
AND2    gate9418  (.A(WX6254), .B(WX4060), .Z(WX4059) ) ;
AND2    gate9419  (.A(WX4384), .B(WX4883), .Z(WX4062) ) ;
AND2    gate9420  (.A(WX4961), .B(WX4064), .Z(WX4063) ) ;
OR2     gate9421  (.A(WX4077), .B(WX4076), .Z(WX4079) ) ;
AND2    gate9422  (.A(WX4079), .B(WX4882), .Z(WX4068) ) ;
OR2     gate9423  (.A(WX4073), .B(WX4072), .Z(WX4075) ) ;
AND2    gate9424  (.A(WX4075), .B(WX4070), .Z(WX4069) ) ;
AND2    gate9425  (.A(CRC_OUT_6_20), .B(WX4883), .Z(WX4072) ) ;
AND2    gate9426  (.A(WX6261), .B(WX4074), .Z(WX4073) ) ;
AND2    gate9427  (.A(WX4386), .B(WX4883), .Z(WX4076) ) ;
AND2    gate9428  (.A(WX4968), .B(WX4078), .Z(WX4077) ) ;
OR2     gate9429  (.A(WX4091), .B(WX4090), .Z(WX4093) ) ;
AND2    gate9430  (.A(WX4093), .B(WX4882), .Z(WX4082) ) ;
OR2     gate9431  (.A(WX4087), .B(WX4086), .Z(WX4089) ) ;
AND2    gate9432  (.A(WX4089), .B(WX4084), .Z(WX4083) ) ;
AND2    gate9433  (.A(CRC_OUT_6_19), .B(WX4883), .Z(WX4086) ) ;
AND2    gate9434  (.A(WX6268), .B(WX4088), .Z(WX4087) ) ;
AND2    gate9435  (.A(WX4388), .B(WX4883), .Z(WX4090) ) ;
AND2    gate9436  (.A(WX4975), .B(WX4092), .Z(WX4091) ) ;
OR2     gate9437  (.A(WX4105), .B(WX4104), .Z(WX4107) ) ;
AND2    gate9438  (.A(WX4107), .B(WX4882), .Z(WX4096) ) ;
OR2     gate9439  (.A(WX4101), .B(WX4100), .Z(WX4103) ) ;
AND2    gate9440  (.A(WX4103), .B(WX4098), .Z(WX4097) ) ;
AND2    gate9441  (.A(CRC_OUT_6_18), .B(WX4883), .Z(WX4100) ) ;
AND2    gate9442  (.A(WX6275), .B(WX4102), .Z(WX4101) ) ;
AND2    gate9443  (.A(WX4390), .B(WX4883), .Z(WX4104) ) ;
AND2    gate9444  (.A(WX4982), .B(WX4106), .Z(WX4105) ) ;
OR2     gate9445  (.A(WX4119), .B(WX4118), .Z(WX4121) ) ;
AND2    gate9446  (.A(WX4121), .B(WX4882), .Z(WX4110) ) ;
OR2     gate9447  (.A(WX4115), .B(WX4114), .Z(WX4117) ) ;
AND2    gate9448  (.A(WX4117), .B(WX4112), .Z(WX4111) ) ;
AND2    gate9449  (.A(CRC_OUT_6_17), .B(WX4883), .Z(WX4114) ) ;
AND2    gate9450  (.A(WX6282), .B(WX4116), .Z(WX4115) ) ;
AND2    gate9451  (.A(WX4392), .B(WX4883), .Z(WX4118) ) ;
AND2    gate9452  (.A(WX4989), .B(WX4120), .Z(WX4119) ) ;
OR2     gate9453  (.A(WX4133), .B(WX4132), .Z(WX4135) ) ;
AND2    gate9454  (.A(WX4135), .B(WX4882), .Z(WX4124) ) ;
OR2     gate9455  (.A(WX4129), .B(WX4128), .Z(WX4131) ) ;
AND2    gate9456  (.A(WX4131), .B(WX4126), .Z(WX4125) ) ;
AND2    gate9457  (.A(CRC_OUT_6_16), .B(WX4883), .Z(WX4128) ) ;
AND2    gate9458  (.A(WX6289), .B(WX4130), .Z(WX4129) ) ;
AND2    gate9459  (.A(WX4394), .B(WX4883), .Z(WX4132) ) ;
AND2    gate9460  (.A(WX4996), .B(WX4134), .Z(WX4133) ) ;
OR2     gate9461  (.A(WX4147), .B(WX4146), .Z(WX4149) ) ;
AND2    gate9462  (.A(WX4149), .B(WX4882), .Z(WX4138) ) ;
OR2     gate9463  (.A(WX4143), .B(WX4142), .Z(WX4145) ) ;
AND2    gate9464  (.A(WX4145), .B(WX4140), .Z(WX4139) ) ;
AND2    gate9465  (.A(CRC_OUT_6_15), .B(WX4883), .Z(WX4142) ) ;
AND2    gate9466  (.A(WX6296), .B(WX4144), .Z(WX4143) ) ;
AND2    gate9467  (.A(WX4396), .B(WX4883), .Z(WX4146) ) ;
AND2    gate9468  (.A(WX5003), .B(WX4148), .Z(WX4147) ) ;
OR2     gate9469  (.A(WX4161), .B(WX4160), .Z(WX4163) ) ;
AND2    gate9470  (.A(WX4163), .B(WX4882), .Z(WX4152) ) ;
OR2     gate9471  (.A(WX4157), .B(WX4156), .Z(WX4159) ) ;
AND2    gate9472  (.A(WX4159), .B(WX4154), .Z(WX4153) ) ;
AND2    gate9473  (.A(CRC_OUT_6_14), .B(WX4883), .Z(WX4156) ) ;
AND2    gate9474  (.A(WX6303), .B(WX4158), .Z(WX4157) ) ;
AND2    gate9475  (.A(WX4398), .B(WX4883), .Z(WX4160) ) ;
AND2    gate9476  (.A(WX5010), .B(WX4162), .Z(WX4161) ) ;
OR2     gate9477  (.A(WX4175), .B(WX4174), .Z(WX4177) ) ;
AND2    gate9478  (.A(WX4177), .B(WX4882), .Z(WX4166) ) ;
OR2     gate9479  (.A(WX4171), .B(WX4170), .Z(WX4173) ) ;
AND2    gate9480  (.A(WX4173), .B(WX4168), .Z(WX4167) ) ;
AND2    gate9481  (.A(CRC_OUT_6_13), .B(WX4883), .Z(WX4170) ) ;
AND2    gate9482  (.A(WX6310), .B(WX4172), .Z(WX4171) ) ;
AND2    gate9483  (.A(WX4400), .B(WX4883), .Z(WX4174) ) ;
AND2    gate9484  (.A(WX5017), .B(WX4176), .Z(WX4175) ) ;
OR2     gate9485  (.A(WX4189), .B(WX4188), .Z(WX4191) ) ;
AND2    gate9486  (.A(WX4191), .B(WX4882), .Z(WX4180) ) ;
OR2     gate9487  (.A(WX4185), .B(WX4184), .Z(WX4187) ) ;
AND2    gate9488  (.A(WX4187), .B(WX4182), .Z(WX4181) ) ;
AND2    gate9489  (.A(CRC_OUT_6_12), .B(WX4883), .Z(WX4184) ) ;
AND2    gate9490  (.A(WX6317), .B(WX4186), .Z(WX4185) ) ;
AND2    gate9491  (.A(WX4402), .B(WX4883), .Z(WX4188) ) ;
AND2    gate9492  (.A(WX5024), .B(WX4190), .Z(WX4189) ) ;
OR2     gate9493  (.A(WX4203), .B(WX4202), .Z(WX4205) ) ;
AND2    gate9494  (.A(WX4205), .B(WX4882), .Z(WX4194) ) ;
OR2     gate9495  (.A(WX4199), .B(WX4198), .Z(WX4201) ) ;
AND2    gate9496  (.A(WX4201), .B(WX4196), .Z(WX4195) ) ;
AND2    gate9497  (.A(CRC_OUT_6_11), .B(WX4883), .Z(WX4198) ) ;
AND2    gate9498  (.A(WX6324), .B(WX4200), .Z(WX4199) ) ;
AND2    gate9499  (.A(WX4404), .B(WX4883), .Z(WX4202) ) ;
AND2    gate9500  (.A(WX5031), .B(WX4204), .Z(WX4203) ) ;
OR2     gate9501  (.A(WX4217), .B(WX4216), .Z(WX4219) ) ;
AND2    gate9502  (.A(WX4219), .B(WX4882), .Z(WX4208) ) ;
OR2     gate9503  (.A(WX4213), .B(WX4212), .Z(WX4215) ) ;
AND2    gate9504  (.A(WX4215), .B(WX4210), .Z(WX4209) ) ;
AND2    gate9505  (.A(CRC_OUT_6_10), .B(WX4883), .Z(WX4212) ) ;
AND2    gate9506  (.A(WX6331), .B(WX4214), .Z(WX4213) ) ;
AND2    gate9507  (.A(WX4406), .B(WX4883), .Z(WX4216) ) ;
AND2    gate9508  (.A(WX5038), .B(WX4218), .Z(WX4217) ) ;
OR2     gate9509  (.A(WX4231), .B(WX4230), .Z(WX4233) ) ;
AND2    gate9510  (.A(WX4233), .B(WX4882), .Z(WX4222) ) ;
OR2     gate9511  (.A(WX4227), .B(WX4226), .Z(WX4229) ) ;
AND2    gate9512  (.A(WX4229), .B(WX4224), .Z(WX4223) ) ;
AND2    gate9513  (.A(CRC_OUT_6_9), .B(WX4883), .Z(WX4226) ) ;
AND2    gate9514  (.A(WX6338), .B(WX4228), .Z(WX4227) ) ;
AND2    gate9515  (.A(WX4408), .B(WX4883), .Z(WX4230) ) ;
AND2    gate9516  (.A(WX5045), .B(WX4232), .Z(WX4231) ) ;
OR2     gate9517  (.A(WX4245), .B(WX4244), .Z(WX4247) ) ;
AND2    gate9518  (.A(WX4247), .B(WX4882), .Z(WX4236) ) ;
OR2     gate9519  (.A(WX4241), .B(WX4240), .Z(WX4243) ) ;
AND2    gate9520  (.A(WX4243), .B(WX4238), .Z(WX4237) ) ;
AND2    gate9521  (.A(CRC_OUT_6_8), .B(WX4883), .Z(WX4240) ) ;
AND2    gate9522  (.A(WX6345), .B(WX4242), .Z(WX4241) ) ;
AND2    gate9523  (.A(WX4410), .B(WX4883), .Z(WX4244) ) ;
AND2    gate9524  (.A(WX5052), .B(WX4246), .Z(WX4245) ) ;
OR2     gate9525  (.A(WX4259), .B(WX4258), .Z(WX4261) ) ;
AND2    gate9526  (.A(WX4261), .B(WX4882), .Z(WX4250) ) ;
OR2     gate9527  (.A(WX4255), .B(WX4254), .Z(WX4257) ) ;
AND2    gate9528  (.A(WX4257), .B(WX4252), .Z(WX4251) ) ;
AND2    gate9529  (.A(CRC_OUT_6_7), .B(WX4883), .Z(WX4254) ) ;
AND2    gate9530  (.A(WX6352), .B(WX4256), .Z(WX4255) ) ;
AND2    gate9531  (.A(WX4412), .B(WX4883), .Z(WX4258) ) ;
AND2    gate9532  (.A(WX5059), .B(WX4260), .Z(WX4259) ) ;
OR2     gate9533  (.A(WX4273), .B(WX4272), .Z(WX4275) ) ;
AND2    gate9534  (.A(WX4275), .B(WX4882), .Z(WX4264) ) ;
OR2     gate9535  (.A(WX4269), .B(WX4268), .Z(WX4271) ) ;
AND2    gate9536  (.A(WX4271), .B(WX4266), .Z(WX4265) ) ;
AND2    gate9537  (.A(CRC_OUT_6_6), .B(WX4883), .Z(WX4268) ) ;
AND2    gate9538  (.A(WX6359), .B(WX4270), .Z(WX4269) ) ;
AND2    gate9539  (.A(WX4414), .B(WX4883), .Z(WX4272) ) ;
AND2    gate9540  (.A(WX5066), .B(WX4274), .Z(WX4273) ) ;
OR2     gate9541  (.A(WX4287), .B(WX4286), .Z(WX4289) ) ;
AND2    gate9542  (.A(WX4289), .B(WX4882), .Z(WX4278) ) ;
OR2     gate9543  (.A(WX4283), .B(WX4282), .Z(WX4285) ) ;
AND2    gate9544  (.A(WX4285), .B(WX4280), .Z(WX4279) ) ;
AND2    gate9545  (.A(CRC_OUT_6_5), .B(WX4883), .Z(WX4282) ) ;
AND2    gate9546  (.A(WX6366), .B(WX4284), .Z(WX4283) ) ;
AND2    gate9547  (.A(WX4416), .B(WX4883), .Z(WX4286) ) ;
AND2    gate9548  (.A(WX5073), .B(WX4288), .Z(WX4287) ) ;
OR2     gate9549  (.A(WX4301), .B(WX4300), .Z(WX4303) ) ;
AND2    gate9550  (.A(WX4303), .B(WX4882), .Z(WX4292) ) ;
OR2     gate9551  (.A(WX4297), .B(WX4296), .Z(WX4299) ) ;
AND2    gate9552  (.A(WX4299), .B(WX4294), .Z(WX4293) ) ;
AND2    gate9553  (.A(CRC_OUT_6_4), .B(WX4883), .Z(WX4296) ) ;
AND2    gate9554  (.A(WX6373), .B(WX4298), .Z(WX4297) ) ;
AND2    gate9555  (.A(WX4418), .B(WX4883), .Z(WX4300) ) ;
AND2    gate9556  (.A(WX5080), .B(WX4302), .Z(WX4301) ) ;
OR2     gate9557  (.A(WX4315), .B(WX4314), .Z(WX4317) ) ;
AND2    gate9558  (.A(WX4317), .B(WX4882), .Z(WX4306) ) ;
OR2     gate9559  (.A(WX4311), .B(WX4310), .Z(WX4313) ) ;
AND2    gate9560  (.A(WX4313), .B(WX4308), .Z(WX4307) ) ;
AND2    gate9561  (.A(CRC_OUT_6_3), .B(WX4883), .Z(WX4310) ) ;
AND2    gate9562  (.A(WX6380), .B(WX4312), .Z(WX4311) ) ;
AND2    gate9563  (.A(WX4420), .B(WX4883), .Z(WX4314) ) ;
AND2    gate9564  (.A(WX5087), .B(WX4316), .Z(WX4315) ) ;
OR2     gate9565  (.A(WX4329), .B(WX4328), .Z(WX4331) ) ;
AND2    gate9566  (.A(WX4331), .B(WX4882), .Z(WX4320) ) ;
OR2     gate9567  (.A(WX4325), .B(WX4324), .Z(WX4327) ) ;
AND2    gate9568  (.A(WX4327), .B(WX4322), .Z(WX4321) ) ;
AND2    gate9569  (.A(CRC_OUT_6_2), .B(WX4883), .Z(WX4324) ) ;
AND2    gate9570  (.A(WX6387), .B(WX4326), .Z(WX4325) ) ;
AND2    gate9571  (.A(WX4422), .B(WX4883), .Z(WX4328) ) ;
AND2    gate9572  (.A(WX5094), .B(WX4330), .Z(WX4329) ) ;
OR2     gate9573  (.A(WX4343), .B(WX4342), .Z(WX4345) ) ;
AND2    gate9574  (.A(WX4345), .B(WX4882), .Z(WX4334) ) ;
OR2     gate9575  (.A(WX4339), .B(WX4338), .Z(WX4341) ) ;
AND2    gate9576  (.A(WX4341), .B(WX4336), .Z(WX4335) ) ;
AND2    gate9577  (.A(CRC_OUT_6_1), .B(WX4883), .Z(WX4338) ) ;
AND2    gate9578  (.A(WX6394), .B(WX4340), .Z(WX4339) ) ;
AND2    gate9579  (.A(WX4424), .B(WX4883), .Z(WX4342) ) ;
AND2    gate9580  (.A(WX5101), .B(WX4344), .Z(WX4343) ) ;
OR2     gate9581  (.A(WX4357), .B(WX4356), .Z(WX4359) ) ;
AND2    gate9582  (.A(WX4359), .B(WX4882), .Z(WX4348) ) ;
OR2     gate9583  (.A(WX4353), .B(WX4352), .Z(WX4355) ) ;
AND2    gate9584  (.A(WX4355), .B(WX4350), .Z(WX4349) ) ;
AND2    gate9585  (.A(CRC_OUT_6_0), .B(WX4883), .Z(WX4352) ) ;
AND2    gate9586  (.A(WX6401), .B(WX4354), .Z(WX4353) ) ;
AND2    gate9587  (.A(WX4426), .B(WX4883), .Z(WX4356) ) ;
AND2    gate9588  (.A(WX5108), .B(WX4358), .Z(WX4357) ) ;
NAND2   gate9589  (.A(II15068), .B(II15069), .Z(WX4885) ) ;
AND2    gate9590  (.A(WX4885), .B(WX4884), .Z(WX4886) ) ;
AND2    gate9591  (.A(WX4459), .B(WX4888), .Z(WX4887) ) ;
NAND2   gate9592  (.A(II15081), .B(II15082), .Z(WX4892) ) ;
AND2    gate9593  (.A(WX4892), .B(WX4884), .Z(WX4893) ) ;
AND2    gate9594  (.A(WX4460), .B(WX4895), .Z(WX4894) ) ;
NAND2   gate9595  (.A(II15094), .B(II15095), .Z(WX4899) ) ;
AND2    gate9596  (.A(WX4899), .B(WX4884), .Z(WX4900) ) ;
AND2    gate9597  (.A(WX4461), .B(WX4902), .Z(WX4901) ) ;
NAND2   gate9598  (.A(II15107), .B(II15108), .Z(WX4906) ) ;
AND2    gate9599  (.A(WX4906), .B(WX4884), .Z(WX4907) ) ;
AND2    gate9600  (.A(WX4462), .B(WX4909), .Z(WX4908) ) ;
NAND2   gate9601  (.A(II15120), .B(II15121), .Z(WX4913) ) ;
AND2    gate9602  (.A(WX4913), .B(WX4884), .Z(WX4914) ) ;
AND2    gate9603  (.A(WX4463), .B(WX4916), .Z(WX4915) ) ;
NAND2   gate9604  (.A(II15133), .B(II15134), .Z(WX4920) ) ;
AND2    gate9605  (.A(WX4920), .B(WX4884), .Z(WX4921) ) ;
AND2    gate9606  (.A(WX4464), .B(WX4923), .Z(WX4922) ) ;
NAND2   gate9607  (.A(II15146), .B(II15147), .Z(WX4927) ) ;
AND2    gate9608  (.A(WX4927), .B(WX4884), .Z(WX4928) ) ;
AND2    gate9609  (.A(WX4465), .B(WX4930), .Z(WX4929) ) ;
NAND2   gate9610  (.A(II15159), .B(II15160), .Z(WX4934) ) ;
AND2    gate9611  (.A(WX4934), .B(WX4884), .Z(WX4935) ) ;
AND2    gate9612  (.A(WX4466), .B(WX4937), .Z(WX4936) ) ;
NAND2   gate9613  (.A(II15172), .B(II15173), .Z(WX4941) ) ;
AND2    gate9614  (.A(WX4941), .B(WX4884), .Z(WX4942) ) ;
AND2    gate9615  (.A(WX4467), .B(WX4944), .Z(WX4943) ) ;
NAND2   gate9616  (.A(II15185), .B(II15186), .Z(WX4948) ) ;
AND2    gate9617  (.A(WX4948), .B(WX4884), .Z(WX4949) ) ;
AND2    gate9618  (.A(WX4468), .B(WX4951), .Z(WX4950) ) ;
NAND2   gate9619  (.A(II15198), .B(II15199), .Z(WX4955) ) ;
AND2    gate9620  (.A(WX4955), .B(WX4884), .Z(WX4956) ) ;
AND2    gate9621  (.A(WX4469), .B(WX4958), .Z(WX4957) ) ;
NAND2   gate9622  (.A(II15211), .B(II15212), .Z(WX4962) ) ;
AND2    gate9623  (.A(WX4962), .B(WX4884), .Z(WX4963) ) ;
AND2    gate9624  (.A(WX4470), .B(WX4965), .Z(WX4964) ) ;
NAND2   gate9625  (.A(II15224), .B(II15225), .Z(WX4969) ) ;
AND2    gate9626  (.A(WX4969), .B(WX4884), .Z(WX4970) ) ;
AND2    gate9627  (.A(WX4471), .B(WX4972), .Z(WX4971) ) ;
NAND2   gate9628  (.A(II15237), .B(II15238), .Z(WX4976) ) ;
AND2    gate9629  (.A(WX4976), .B(WX4884), .Z(WX4977) ) ;
AND2    gate9630  (.A(WX4472), .B(WX4979), .Z(WX4978) ) ;
NAND2   gate9631  (.A(II15250), .B(II15251), .Z(WX4983) ) ;
AND2    gate9632  (.A(WX4983), .B(WX4884), .Z(WX4984) ) ;
AND2    gate9633  (.A(WX4473), .B(WX4986), .Z(WX4985) ) ;
NAND2   gate9634  (.A(II15263), .B(II15264), .Z(WX4990) ) ;
AND2    gate9635  (.A(WX4990), .B(WX4884), .Z(WX4991) ) ;
AND2    gate9636  (.A(WX4474), .B(WX4993), .Z(WX4992) ) ;
NAND2   gate9637  (.A(II15276), .B(II15277), .Z(WX4997) ) ;
AND2    gate9638  (.A(WX4997), .B(WX4884), .Z(WX4998) ) ;
AND2    gate9639  (.A(WX4475), .B(WX5000), .Z(WX4999) ) ;
NAND2   gate9640  (.A(II15289), .B(II15290), .Z(WX5004) ) ;
AND2    gate9641  (.A(WX5004), .B(WX4884), .Z(WX5005) ) ;
AND2    gate9642  (.A(WX4476), .B(WX5007), .Z(WX5006) ) ;
NAND2   gate9643  (.A(II15302), .B(II15303), .Z(WX5011) ) ;
AND2    gate9644  (.A(WX5011), .B(WX4884), .Z(WX5012) ) ;
AND2    gate9645  (.A(WX4477), .B(WX5014), .Z(WX5013) ) ;
NAND2   gate9646  (.A(II15315), .B(II15316), .Z(WX5018) ) ;
AND2    gate9647  (.A(WX5018), .B(WX4884), .Z(WX5019) ) ;
AND2    gate9648  (.A(WX4478), .B(WX5021), .Z(WX5020) ) ;
NAND2   gate9649  (.A(II15328), .B(II15329), .Z(WX5025) ) ;
AND2    gate9650  (.A(WX5025), .B(WX4884), .Z(WX5026) ) ;
AND2    gate9651  (.A(WX4479), .B(WX5028), .Z(WX5027) ) ;
NAND2   gate9652  (.A(II15341), .B(II15342), .Z(WX5032) ) ;
AND2    gate9653  (.A(WX5032), .B(WX4884), .Z(WX5033) ) ;
AND2    gate9654  (.A(WX4480), .B(WX5035), .Z(WX5034) ) ;
NAND2   gate9655  (.A(II15354), .B(II15355), .Z(WX5039) ) ;
AND2    gate9656  (.A(WX5039), .B(WX4884), .Z(WX5040) ) ;
AND2    gate9657  (.A(WX4481), .B(WX5042), .Z(WX5041) ) ;
NAND2   gate9658  (.A(II15367), .B(II15368), .Z(WX5046) ) ;
AND2    gate9659  (.A(WX5046), .B(WX4884), .Z(WX5047) ) ;
AND2    gate9660  (.A(WX4482), .B(WX5049), .Z(WX5048) ) ;
NAND2   gate9661  (.A(II15380), .B(II15381), .Z(WX5053) ) ;
AND2    gate9662  (.A(WX5053), .B(WX4884), .Z(WX5054) ) ;
AND2    gate9663  (.A(WX4483), .B(WX5056), .Z(WX5055) ) ;
NAND2   gate9664  (.A(II15393), .B(II15394), .Z(WX5060) ) ;
AND2    gate9665  (.A(WX5060), .B(WX4884), .Z(WX5061) ) ;
AND2    gate9666  (.A(WX4484), .B(WX5063), .Z(WX5062) ) ;
NAND2   gate9667  (.A(II15406), .B(II15407), .Z(WX5067) ) ;
AND2    gate9668  (.A(WX5067), .B(WX4884), .Z(WX5068) ) ;
AND2    gate9669  (.A(WX4485), .B(WX5070), .Z(WX5069) ) ;
NAND2   gate9670  (.A(II15419), .B(II15420), .Z(WX5074) ) ;
AND2    gate9671  (.A(WX5074), .B(WX4884), .Z(WX5075) ) ;
AND2    gate9672  (.A(WX4486), .B(WX5077), .Z(WX5076) ) ;
NAND2   gate9673  (.A(II15432), .B(II15433), .Z(WX5081) ) ;
AND2    gate9674  (.A(WX5081), .B(WX4884), .Z(WX5082) ) ;
AND2    gate9675  (.A(WX4487), .B(WX5084), .Z(WX5083) ) ;
NAND2   gate9676  (.A(II15445), .B(II15446), .Z(WX5088) ) ;
AND2    gate9677  (.A(WX5088), .B(WX4884), .Z(WX5089) ) ;
AND2    gate9678  (.A(WX4488), .B(WX5091), .Z(WX5090) ) ;
NAND2   gate9679  (.A(II15458), .B(II15459), .Z(WX5095) ) ;
AND2    gate9680  (.A(WX5095), .B(WX4884), .Z(WX5096) ) ;
AND2    gate9681  (.A(WX4489), .B(WX5098), .Z(WX5097) ) ;
NAND2   gate9682  (.A(II15471), .B(II15472), .Z(WX5102) ) ;
AND2    gate9683  (.A(WX5102), .B(WX4884), .Z(WX5103) ) ;
AND2    gate9684  (.A(WX4490), .B(WX5105), .Z(WX5104) ) ;
NAND2   gate9685  (.A(II15530), .B(II15531), .Z(WX5113) ) ;
NAND2   gate9686  (.A(II15726), .B(II15727), .Z(WX5141) ) ;
NAND2   gate9687  (.A(II15719), .B(II15720), .Z(WX5140) ) ;
NAND2   gate9688  (.A(II15712), .B(II15713), .Z(WX5139) ) ;
NAND2   gate9689  (.A(II15523), .B(II15524), .Z(WX5112) ) ;
NAND2   gate9690  (.A(II15705), .B(II15706), .Z(WX5138) ) ;
NAND2   gate9691  (.A(II15698), .B(II15699), .Z(WX5137) ) ;
NAND2   gate9692  (.A(II15691), .B(II15692), .Z(WX5136) ) ;
NAND2   gate9693  (.A(II15684), .B(II15685), .Z(WX5135) ) ;
NAND2   gate9694  (.A(II15677), .B(II15678), .Z(WX5134) ) ;
NAND2   gate9695  (.A(II15670), .B(II15671), .Z(WX5133) ) ;
NAND2   gate9696  (.A(II15508), .B(II15509), .Z(WX5111) ) ;
NAND2   gate9697  (.A(II15663), .B(II15664), .Z(WX5132) ) ;
NAND2   gate9698  (.A(II15656), .B(II15657), .Z(WX5131) ) ;
NAND2   gate9699  (.A(II15649), .B(II15650), .Z(WX5130) ) ;
NAND2   gate9700  (.A(II15642), .B(II15643), .Z(WX5129) ) ;
NAND2   gate9701  (.A(II15493), .B(II15494), .Z(WX5110) ) ;
NAND2   gate9702  (.A(II15635), .B(II15636), .Z(WX5128) ) ;
NAND2   gate9703  (.A(II15628), .B(II15629), .Z(WX5127) ) ;
NAND2   gate9704  (.A(II15621), .B(II15622), .Z(WX5126) ) ;
NAND2   gate9705  (.A(II15614), .B(II15615), .Z(WX5125) ) ;
NAND2   gate9706  (.A(II15607), .B(II15608), .Z(WX5124) ) ;
NAND2   gate9707  (.A(II15600), .B(II15601), .Z(WX5123) ) ;
NAND2   gate9708  (.A(II15593), .B(II15594), .Z(WX5122) ) ;
NAND2   gate9709  (.A(II15586), .B(II15587), .Z(WX5121) ) ;
NAND2   gate9710  (.A(II15579), .B(II15580), .Z(WX5120) ) ;
NAND2   gate9711  (.A(II15572), .B(II15573), .Z(WX5119) ) ;
NAND2   gate9712  (.A(II15565), .B(II15566), .Z(WX5118) ) ;
NAND2   gate9713  (.A(II15558), .B(II15559), .Z(WX5117) ) ;
NAND2   gate9714  (.A(II15551), .B(II15552), .Z(WX5116) ) ;
NAND2   gate9715  (.A(II15544), .B(II15545), .Z(WX5115) ) ;
NAND2   gate9716  (.A(II15537), .B(II15538), .Z(WX5114) ) ;
OR2     gate9717  (.A(WX5216), .B(WX5215), .Z(WX5218) ) ;
AND2    gate9718  (.A(WX5218), .B(WX6175), .Z(WX5207) ) ;
OR2     gate9719  (.A(WX5212), .B(WX5211), .Z(WX5214) ) ;
AND2    gate9720  (.A(WX5214), .B(WX5209), .Z(WX5208) ) ;
AND2    gate9721  (.A(CRC_OUT_5_31), .B(WX6176), .Z(WX5211) ) ;
AND2    gate9722  (.A(WX7477), .B(WX5213), .Z(WX5212) ) ;
AND2    gate9723  (.A(WX5657), .B(WX6176), .Z(WX5215) ) ;
AND2    gate9724  (.A(WX6184), .B(WX5217), .Z(WX5216) ) ;
OR2     gate9725  (.A(WX5230), .B(WX5229), .Z(WX5232) ) ;
AND2    gate9726  (.A(WX5232), .B(WX6175), .Z(WX5221) ) ;
OR2     gate9727  (.A(WX5226), .B(WX5225), .Z(WX5228) ) ;
AND2    gate9728  (.A(WX5228), .B(WX5223), .Z(WX5222) ) ;
AND2    gate9729  (.A(CRC_OUT_5_30), .B(WX6176), .Z(WX5225) ) ;
AND2    gate9730  (.A(WX7484), .B(WX5227), .Z(WX5226) ) ;
AND2    gate9731  (.A(WX5659), .B(WX6176), .Z(WX5229) ) ;
AND2    gate9732  (.A(WX6191), .B(WX5231), .Z(WX5230) ) ;
OR2     gate9733  (.A(WX5244), .B(WX5243), .Z(WX5246) ) ;
AND2    gate9734  (.A(WX5246), .B(WX6175), .Z(WX5235) ) ;
OR2     gate9735  (.A(WX5240), .B(WX5239), .Z(WX5242) ) ;
AND2    gate9736  (.A(WX5242), .B(WX5237), .Z(WX5236) ) ;
AND2    gate9737  (.A(CRC_OUT_5_29), .B(WX6176), .Z(WX5239) ) ;
AND2    gate9738  (.A(WX7491), .B(WX5241), .Z(WX5240) ) ;
AND2    gate9739  (.A(WX5661), .B(WX6176), .Z(WX5243) ) ;
AND2    gate9740  (.A(WX6198), .B(WX5245), .Z(WX5244) ) ;
OR2     gate9741  (.A(WX5258), .B(WX5257), .Z(WX5260) ) ;
AND2    gate9742  (.A(WX5260), .B(WX6175), .Z(WX5249) ) ;
OR2     gate9743  (.A(WX5254), .B(WX5253), .Z(WX5256) ) ;
AND2    gate9744  (.A(WX5256), .B(WX5251), .Z(WX5250) ) ;
AND2    gate9745  (.A(CRC_OUT_5_28), .B(WX6176), .Z(WX5253) ) ;
AND2    gate9746  (.A(WX7498), .B(WX5255), .Z(WX5254) ) ;
AND2    gate9747  (.A(WX5663), .B(WX6176), .Z(WX5257) ) ;
AND2    gate9748  (.A(WX6205), .B(WX5259), .Z(WX5258) ) ;
OR2     gate9749  (.A(WX5272), .B(WX5271), .Z(WX5274) ) ;
AND2    gate9750  (.A(WX5274), .B(WX6175), .Z(WX5263) ) ;
OR2     gate9751  (.A(WX5268), .B(WX5267), .Z(WX5270) ) ;
AND2    gate9752  (.A(WX5270), .B(WX5265), .Z(WX5264) ) ;
AND2    gate9753  (.A(CRC_OUT_5_27), .B(WX6176), .Z(WX5267) ) ;
AND2    gate9754  (.A(WX7505), .B(WX5269), .Z(WX5268) ) ;
AND2    gate9755  (.A(WX5665), .B(WX6176), .Z(WX5271) ) ;
AND2    gate9756  (.A(WX6212), .B(WX5273), .Z(WX5272) ) ;
OR2     gate9757  (.A(WX5286), .B(WX5285), .Z(WX5288) ) ;
AND2    gate9758  (.A(WX5288), .B(WX6175), .Z(WX5277) ) ;
OR2     gate9759  (.A(WX5282), .B(WX5281), .Z(WX5284) ) ;
AND2    gate9760  (.A(WX5284), .B(WX5279), .Z(WX5278) ) ;
AND2    gate9761  (.A(CRC_OUT_5_26), .B(WX6176), .Z(WX5281) ) ;
AND2    gate9762  (.A(WX7512), .B(WX5283), .Z(WX5282) ) ;
AND2    gate9763  (.A(WX5667), .B(WX6176), .Z(WX5285) ) ;
AND2    gate9764  (.A(WX6219), .B(WX5287), .Z(WX5286) ) ;
OR2     gate9765  (.A(WX5300), .B(WX5299), .Z(WX5302) ) ;
AND2    gate9766  (.A(WX5302), .B(WX6175), .Z(WX5291) ) ;
OR2     gate9767  (.A(WX5296), .B(WX5295), .Z(WX5298) ) ;
AND2    gate9768  (.A(WX5298), .B(WX5293), .Z(WX5292) ) ;
AND2    gate9769  (.A(CRC_OUT_5_25), .B(WX6176), .Z(WX5295) ) ;
AND2    gate9770  (.A(WX7519), .B(WX5297), .Z(WX5296) ) ;
AND2    gate9771  (.A(WX5669), .B(WX6176), .Z(WX5299) ) ;
AND2    gate9772  (.A(WX6226), .B(WX5301), .Z(WX5300) ) ;
OR2     gate9773  (.A(WX5314), .B(WX5313), .Z(WX5316) ) ;
AND2    gate9774  (.A(WX5316), .B(WX6175), .Z(WX5305) ) ;
OR2     gate9775  (.A(WX5310), .B(WX5309), .Z(WX5312) ) ;
AND2    gate9776  (.A(WX5312), .B(WX5307), .Z(WX5306) ) ;
AND2    gate9777  (.A(CRC_OUT_5_24), .B(WX6176), .Z(WX5309) ) ;
AND2    gate9778  (.A(WX7526), .B(WX5311), .Z(WX5310) ) ;
AND2    gate9779  (.A(WX5671), .B(WX6176), .Z(WX5313) ) ;
AND2    gate9780  (.A(WX6233), .B(WX5315), .Z(WX5314) ) ;
OR2     gate9781  (.A(WX5328), .B(WX5327), .Z(WX5330) ) ;
AND2    gate9782  (.A(WX5330), .B(WX6175), .Z(WX5319) ) ;
OR2     gate9783  (.A(WX5324), .B(WX5323), .Z(WX5326) ) ;
AND2    gate9784  (.A(WX5326), .B(WX5321), .Z(WX5320) ) ;
AND2    gate9785  (.A(CRC_OUT_5_23), .B(WX6176), .Z(WX5323) ) ;
AND2    gate9786  (.A(WX7533), .B(WX5325), .Z(WX5324) ) ;
AND2    gate9787  (.A(WX5673), .B(WX6176), .Z(WX5327) ) ;
AND2    gate9788  (.A(WX6240), .B(WX5329), .Z(WX5328) ) ;
OR2     gate9789  (.A(WX5342), .B(WX5341), .Z(WX5344) ) ;
AND2    gate9790  (.A(WX5344), .B(WX6175), .Z(WX5333) ) ;
OR2     gate9791  (.A(WX5338), .B(WX5337), .Z(WX5340) ) ;
AND2    gate9792  (.A(WX5340), .B(WX5335), .Z(WX5334) ) ;
AND2    gate9793  (.A(CRC_OUT_5_22), .B(WX6176), .Z(WX5337) ) ;
AND2    gate9794  (.A(WX7540), .B(WX5339), .Z(WX5338) ) ;
AND2    gate9795  (.A(WX5675), .B(WX6176), .Z(WX5341) ) ;
AND2    gate9796  (.A(WX6247), .B(WX5343), .Z(WX5342) ) ;
OR2     gate9797  (.A(WX5356), .B(WX5355), .Z(WX5358) ) ;
AND2    gate9798  (.A(WX5358), .B(WX6175), .Z(WX5347) ) ;
OR2     gate9799  (.A(WX5352), .B(WX5351), .Z(WX5354) ) ;
AND2    gate9800  (.A(WX5354), .B(WX5349), .Z(WX5348) ) ;
AND2    gate9801  (.A(CRC_OUT_5_21), .B(WX6176), .Z(WX5351) ) ;
AND2    gate9802  (.A(WX7547), .B(WX5353), .Z(WX5352) ) ;
AND2    gate9803  (.A(WX5677), .B(WX6176), .Z(WX5355) ) ;
AND2    gate9804  (.A(WX6254), .B(WX5357), .Z(WX5356) ) ;
OR2     gate9805  (.A(WX5370), .B(WX5369), .Z(WX5372) ) ;
AND2    gate9806  (.A(WX5372), .B(WX6175), .Z(WX5361) ) ;
OR2     gate9807  (.A(WX5366), .B(WX5365), .Z(WX5368) ) ;
AND2    gate9808  (.A(WX5368), .B(WX5363), .Z(WX5362) ) ;
AND2    gate9809  (.A(CRC_OUT_5_20), .B(WX6176), .Z(WX5365) ) ;
AND2    gate9810  (.A(WX7554), .B(WX5367), .Z(WX5366) ) ;
AND2    gate9811  (.A(WX5679), .B(WX6176), .Z(WX5369) ) ;
AND2    gate9812  (.A(WX6261), .B(WX5371), .Z(WX5370) ) ;
OR2     gate9813  (.A(WX5384), .B(WX5383), .Z(WX5386) ) ;
AND2    gate9814  (.A(WX5386), .B(WX6175), .Z(WX5375) ) ;
OR2     gate9815  (.A(WX5380), .B(WX5379), .Z(WX5382) ) ;
AND2    gate9816  (.A(WX5382), .B(WX5377), .Z(WX5376) ) ;
AND2    gate9817  (.A(CRC_OUT_5_19), .B(WX6176), .Z(WX5379) ) ;
AND2    gate9818  (.A(WX7561), .B(WX5381), .Z(WX5380) ) ;
AND2    gate9819  (.A(WX5681), .B(WX6176), .Z(WX5383) ) ;
AND2    gate9820  (.A(WX6268), .B(WX5385), .Z(WX5384) ) ;
OR2     gate9821  (.A(WX5398), .B(WX5397), .Z(WX5400) ) ;
AND2    gate9822  (.A(WX5400), .B(WX6175), .Z(WX5389) ) ;
OR2     gate9823  (.A(WX5394), .B(WX5393), .Z(WX5396) ) ;
AND2    gate9824  (.A(WX5396), .B(WX5391), .Z(WX5390) ) ;
AND2    gate9825  (.A(CRC_OUT_5_18), .B(WX6176), .Z(WX5393) ) ;
AND2    gate9826  (.A(WX7568), .B(WX5395), .Z(WX5394) ) ;
AND2    gate9827  (.A(WX5683), .B(WX6176), .Z(WX5397) ) ;
AND2    gate9828  (.A(WX6275), .B(WX5399), .Z(WX5398) ) ;
OR2     gate9829  (.A(WX5412), .B(WX5411), .Z(WX5414) ) ;
AND2    gate9830  (.A(WX5414), .B(WX6175), .Z(WX5403) ) ;
OR2     gate9831  (.A(WX5408), .B(WX5407), .Z(WX5410) ) ;
AND2    gate9832  (.A(WX5410), .B(WX5405), .Z(WX5404) ) ;
AND2    gate9833  (.A(CRC_OUT_5_17), .B(WX6176), .Z(WX5407) ) ;
AND2    gate9834  (.A(WX7575), .B(WX5409), .Z(WX5408) ) ;
AND2    gate9835  (.A(WX5685), .B(WX6176), .Z(WX5411) ) ;
AND2    gate9836  (.A(WX6282), .B(WX5413), .Z(WX5412) ) ;
OR2     gate9837  (.A(WX5426), .B(WX5425), .Z(WX5428) ) ;
AND2    gate9838  (.A(WX5428), .B(WX6175), .Z(WX5417) ) ;
OR2     gate9839  (.A(WX5422), .B(WX5421), .Z(WX5424) ) ;
AND2    gate9840  (.A(WX5424), .B(WX5419), .Z(WX5418) ) ;
AND2    gate9841  (.A(CRC_OUT_5_16), .B(WX6176), .Z(WX5421) ) ;
AND2    gate9842  (.A(WX7582), .B(WX5423), .Z(WX5422) ) ;
AND2    gate9843  (.A(WX5687), .B(WX6176), .Z(WX5425) ) ;
AND2    gate9844  (.A(WX6289), .B(WX5427), .Z(WX5426) ) ;
OR2     gate9845  (.A(WX5440), .B(WX5439), .Z(WX5442) ) ;
AND2    gate9846  (.A(WX5442), .B(WX6175), .Z(WX5431) ) ;
OR2     gate9847  (.A(WX5436), .B(WX5435), .Z(WX5438) ) ;
AND2    gate9848  (.A(WX5438), .B(WX5433), .Z(WX5432) ) ;
AND2    gate9849  (.A(CRC_OUT_5_15), .B(WX6176), .Z(WX5435) ) ;
AND2    gate9850  (.A(WX7589), .B(WX5437), .Z(WX5436) ) ;
AND2    gate9851  (.A(WX5689), .B(WX6176), .Z(WX5439) ) ;
AND2    gate9852  (.A(WX6296), .B(WX5441), .Z(WX5440) ) ;
OR2     gate9853  (.A(WX5454), .B(WX5453), .Z(WX5456) ) ;
AND2    gate9854  (.A(WX5456), .B(WX6175), .Z(WX5445) ) ;
OR2     gate9855  (.A(WX5450), .B(WX5449), .Z(WX5452) ) ;
AND2    gate9856  (.A(WX5452), .B(WX5447), .Z(WX5446) ) ;
AND2    gate9857  (.A(CRC_OUT_5_14), .B(WX6176), .Z(WX5449) ) ;
AND2    gate9858  (.A(WX7596), .B(WX5451), .Z(WX5450) ) ;
AND2    gate9859  (.A(WX5691), .B(WX6176), .Z(WX5453) ) ;
AND2    gate9860  (.A(WX6303), .B(WX5455), .Z(WX5454) ) ;
OR2     gate9861  (.A(WX5468), .B(WX5467), .Z(WX5470) ) ;
AND2    gate9862  (.A(WX5470), .B(WX6175), .Z(WX5459) ) ;
OR2     gate9863  (.A(WX5464), .B(WX5463), .Z(WX5466) ) ;
AND2    gate9864  (.A(WX5466), .B(WX5461), .Z(WX5460) ) ;
AND2    gate9865  (.A(CRC_OUT_5_13), .B(WX6176), .Z(WX5463) ) ;
AND2    gate9866  (.A(WX7603), .B(WX5465), .Z(WX5464) ) ;
AND2    gate9867  (.A(WX5693), .B(WX6176), .Z(WX5467) ) ;
AND2    gate9868  (.A(WX6310), .B(WX5469), .Z(WX5468) ) ;
OR2     gate9869  (.A(WX5482), .B(WX5481), .Z(WX5484) ) ;
AND2    gate9870  (.A(WX5484), .B(WX6175), .Z(WX5473) ) ;
OR2     gate9871  (.A(WX5478), .B(WX5477), .Z(WX5480) ) ;
AND2    gate9872  (.A(WX5480), .B(WX5475), .Z(WX5474) ) ;
AND2    gate9873  (.A(CRC_OUT_5_12), .B(WX6176), .Z(WX5477) ) ;
AND2    gate9874  (.A(WX7610), .B(WX5479), .Z(WX5478) ) ;
AND2    gate9875  (.A(WX5695), .B(WX6176), .Z(WX5481) ) ;
AND2    gate9876  (.A(WX6317), .B(WX5483), .Z(WX5482) ) ;
OR2     gate9877  (.A(WX5496), .B(WX5495), .Z(WX5498) ) ;
AND2    gate9878  (.A(WX5498), .B(WX6175), .Z(WX5487) ) ;
OR2     gate9879  (.A(WX5492), .B(WX5491), .Z(WX5494) ) ;
AND2    gate9880  (.A(WX5494), .B(WX5489), .Z(WX5488) ) ;
AND2    gate9881  (.A(CRC_OUT_5_11), .B(WX6176), .Z(WX5491) ) ;
AND2    gate9882  (.A(WX7617), .B(WX5493), .Z(WX5492) ) ;
AND2    gate9883  (.A(WX5697), .B(WX6176), .Z(WX5495) ) ;
AND2    gate9884  (.A(WX6324), .B(WX5497), .Z(WX5496) ) ;
OR2     gate9885  (.A(WX5510), .B(WX5509), .Z(WX5512) ) ;
AND2    gate9886  (.A(WX5512), .B(WX6175), .Z(WX5501) ) ;
OR2     gate9887  (.A(WX5506), .B(WX5505), .Z(WX5508) ) ;
AND2    gate9888  (.A(WX5508), .B(WX5503), .Z(WX5502) ) ;
AND2    gate9889  (.A(CRC_OUT_5_10), .B(WX6176), .Z(WX5505) ) ;
AND2    gate9890  (.A(WX7624), .B(WX5507), .Z(WX5506) ) ;
AND2    gate9891  (.A(WX5699), .B(WX6176), .Z(WX5509) ) ;
AND2    gate9892  (.A(WX6331), .B(WX5511), .Z(WX5510) ) ;
OR2     gate9893  (.A(WX5524), .B(WX5523), .Z(WX5526) ) ;
AND2    gate9894  (.A(WX5526), .B(WX6175), .Z(WX5515) ) ;
OR2     gate9895  (.A(WX5520), .B(WX5519), .Z(WX5522) ) ;
AND2    gate9896  (.A(WX5522), .B(WX5517), .Z(WX5516) ) ;
AND2    gate9897  (.A(CRC_OUT_5_9), .B(WX6176), .Z(WX5519) ) ;
AND2    gate9898  (.A(WX7631), .B(WX5521), .Z(WX5520) ) ;
AND2    gate9899  (.A(WX5701), .B(WX6176), .Z(WX5523) ) ;
AND2    gate9900  (.A(WX6338), .B(WX5525), .Z(WX5524) ) ;
OR2     gate9901  (.A(WX5538), .B(WX5537), .Z(WX5540) ) ;
AND2    gate9902  (.A(WX5540), .B(WX6175), .Z(WX5529) ) ;
OR2     gate9903  (.A(WX5534), .B(WX5533), .Z(WX5536) ) ;
AND2    gate9904  (.A(WX5536), .B(WX5531), .Z(WX5530) ) ;
AND2    gate9905  (.A(CRC_OUT_5_8), .B(WX6176), .Z(WX5533) ) ;
AND2    gate9906  (.A(WX7638), .B(WX5535), .Z(WX5534) ) ;
AND2    gate9907  (.A(WX5703), .B(WX6176), .Z(WX5537) ) ;
AND2    gate9908  (.A(WX6345), .B(WX5539), .Z(WX5538) ) ;
OR2     gate9909  (.A(WX5552), .B(WX5551), .Z(WX5554) ) ;
AND2    gate9910  (.A(WX5554), .B(WX6175), .Z(WX5543) ) ;
OR2     gate9911  (.A(WX5548), .B(WX5547), .Z(WX5550) ) ;
AND2    gate9912  (.A(WX5550), .B(WX5545), .Z(WX5544) ) ;
AND2    gate9913  (.A(CRC_OUT_5_7), .B(WX6176), .Z(WX5547) ) ;
AND2    gate9914  (.A(WX7645), .B(WX5549), .Z(WX5548) ) ;
AND2    gate9915  (.A(WX5705), .B(WX6176), .Z(WX5551) ) ;
AND2    gate9916  (.A(WX6352), .B(WX5553), .Z(WX5552) ) ;
OR2     gate9917  (.A(WX5566), .B(WX5565), .Z(WX5568) ) ;
AND2    gate9918  (.A(WX5568), .B(WX6175), .Z(WX5557) ) ;
OR2     gate9919  (.A(WX5562), .B(WX5561), .Z(WX5564) ) ;
AND2    gate9920  (.A(WX5564), .B(WX5559), .Z(WX5558) ) ;
AND2    gate9921  (.A(CRC_OUT_5_6), .B(WX6176), .Z(WX5561) ) ;
AND2    gate9922  (.A(WX7652), .B(WX5563), .Z(WX5562) ) ;
AND2    gate9923  (.A(WX5707), .B(WX6176), .Z(WX5565) ) ;
AND2    gate9924  (.A(WX6359), .B(WX5567), .Z(WX5566) ) ;
OR2     gate9925  (.A(WX5580), .B(WX5579), .Z(WX5582) ) ;
AND2    gate9926  (.A(WX5582), .B(WX6175), .Z(WX5571) ) ;
OR2     gate9927  (.A(WX5576), .B(WX5575), .Z(WX5578) ) ;
AND2    gate9928  (.A(WX5578), .B(WX5573), .Z(WX5572) ) ;
AND2    gate9929  (.A(CRC_OUT_5_5), .B(WX6176), .Z(WX5575) ) ;
AND2    gate9930  (.A(WX7659), .B(WX5577), .Z(WX5576) ) ;
AND2    gate9931  (.A(WX5709), .B(WX6176), .Z(WX5579) ) ;
AND2    gate9932  (.A(WX6366), .B(WX5581), .Z(WX5580) ) ;
OR2     gate9933  (.A(WX5594), .B(WX5593), .Z(WX5596) ) ;
AND2    gate9934  (.A(WX5596), .B(WX6175), .Z(WX5585) ) ;
OR2     gate9935  (.A(WX5590), .B(WX5589), .Z(WX5592) ) ;
AND2    gate9936  (.A(WX5592), .B(WX5587), .Z(WX5586) ) ;
AND2    gate9937  (.A(CRC_OUT_5_4), .B(WX6176), .Z(WX5589) ) ;
AND2    gate9938  (.A(WX7666), .B(WX5591), .Z(WX5590) ) ;
AND2    gate9939  (.A(WX5711), .B(WX6176), .Z(WX5593) ) ;
AND2    gate9940  (.A(WX6373), .B(WX5595), .Z(WX5594) ) ;
OR2     gate9941  (.A(WX5608), .B(WX5607), .Z(WX5610) ) ;
AND2    gate9942  (.A(WX5610), .B(WX6175), .Z(WX5599) ) ;
OR2     gate9943  (.A(WX5604), .B(WX5603), .Z(WX5606) ) ;
AND2    gate9944  (.A(WX5606), .B(WX5601), .Z(WX5600) ) ;
AND2    gate9945  (.A(CRC_OUT_5_3), .B(WX6176), .Z(WX5603) ) ;
AND2    gate9946  (.A(WX7673), .B(WX5605), .Z(WX5604) ) ;
AND2    gate9947  (.A(WX5713), .B(WX6176), .Z(WX5607) ) ;
AND2    gate9948  (.A(WX6380), .B(WX5609), .Z(WX5608) ) ;
OR2     gate9949  (.A(WX5622), .B(WX5621), .Z(WX5624) ) ;
AND2    gate9950  (.A(WX5624), .B(WX6175), .Z(WX5613) ) ;
OR2     gate9951  (.A(WX5618), .B(WX5617), .Z(WX5620) ) ;
AND2    gate9952  (.A(WX5620), .B(WX5615), .Z(WX5614) ) ;
AND2    gate9953  (.A(CRC_OUT_5_2), .B(WX6176), .Z(WX5617) ) ;
AND2    gate9954  (.A(WX7680), .B(WX5619), .Z(WX5618) ) ;
AND2    gate9955  (.A(WX5715), .B(WX6176), .Z(WX5621) ) ;
AND2    gate9956  (.A(WX6387), .B(WX5623), .Z(WX5622) ) ;
OR2     gate9957  (.A(WX5636), .B(WX5635), .Z(WX5638) ) ;
AND2    gate9958  (.A(WX5638), .B(WX6175), .Z(WX5627) ) ;
OR2     gate9959  (.A(WX5632), .B(WX5631), .Z(WX5634) ) ;
AND2    gate9960  (.A(WX5634), .B(WX5629), .Z(WX5628) ) ;
AND2    gate9961  (.A(CRC_OUT_5_1), .B(WX6176), .Z(WX5631) ) ;
AND2    gate9962  (.A(WX7687), .B(WX5633), .Z(WX5632) ) ;
AND2    gate9963  (.A(WX5717), .B(WX6176), .Z(WX5635) ) ;
AND2    gate9964  (.A(WX6394), .B(WX5637), .Z(WX5636) ) ;
OR2     gate9965  (.A(WX5650), .B(WX5649), .Z(WX5652) ) ;
AND2    gate9966  (.A(WX5652), .B(WX6175), .Z(WX5641) ) ;
OR2     gate9967  (.A(WX5646), .B(WX5645), .Z(WX5648) ) ;
AND2    gate9968  (.A(WX5648), .B(WX5643), .Z(WX5642) ) ;
AND2    gate9969  (.A(CRC_OUT_5_0), .B(WX6176), .Z(WX5645) ) ;
AND2    gate9970  (.A(WX7694), .B(WX5647), .Z(WX5646) ) ;
AND2    gate9971  (.A(WX5719), .B(WX6176), .Z(WX5649) ) ;
AND2    gate9972  (.A(WX6401), .B(WX5651), .Z(WX5650) ) ;
NAND2   gate9973  (.A(II19073), .B(II19074), .Z(WX6178) ) ;
AND2    gate9974  (.A(WX6178), .B(WX6177), .Z(WX6179) ) ;
AND2    gate9975  (.A(WX5752), .B(WX6181), .Z(WX6180) ) ;
NAND2   gate9976  (.A(II19086), .B(II19087), .Z(WX6185) ) ;
AND2    gate9977  (.A(WX6185), .B(WX6177), .Z(WX6186) ) ;
AND2    gate9978  (.A(WX5753), .B(WX6188), .Z(WX6187) ) ;
NAND2   gate9979  (.A(II19099), .B(II19100), .Z(WX6192) ) ;
AND2    gate9980  (.A(WX6192), .B(WX6177), .Z(WX6193) ) ;
AND2    gate9981  (.A(WX5754), .B(WX6195), .Z(WX6194) ) ;
NAND2   gate9982  (.A(II19112), .B(II19113), .Z(WX6199) ) ;
AND2    gate9983  (.A(WX6199), .B(WX6177), .Z(WX6200) ) ;
AND2    gate9984  (.A(WX5755), .B(WX6202), .Z(WX6201) ) ;
NAND2   gate9985  (.A(II19125), .B(II19126), .Z(WX6206) ) ;
AND2    gate9986  (.A(WX6206), .B(WX6177), .Z(WX6207) ) ;
AND2    gate9987  (.A(WX5756), .B(WX6209), .Z(WX6208) ) ;
NAND2   gate9988  (.A(II19138), .B(II19139), .Z(WX6213) ) ;
AND2    gate9989  (.A(WX6213), .B(WX6177), .Z(WX6214) ) ;
AND2    gate9990  (.A(WX5757), .B(WX6216), .Z(WX6215) ) ;
NAND2   gate9991  (.A(II19151), .B(II19152), .Z(WX6220) ) ;
AND2    gate9992  (.A(WX6220), .B(WX6177), .Z(WX6221) ) ;
AND2    gate9993  (.A(WX5758), .B(WX6223), .Z(WX6222) ) ;
NAND2   gate9994  (.A(II19164), .B(II19165), .Z(WX6227) ) ;
AND2    gate9995  (.A(WX6227), .B(WX6177), .Z(WX6228) ) ;
AND2    gate9996  (.A(WX5759), .B(WX6230), .Z(WX6229) ) ;
NAND2   gate9997  (.A(II19177), .B(II19178), .Z(WX6234) ) ;
AND2    gate9998  (.A(WX6234), .B(WX6177), .Z(WX6235) ) ;
AND2    gate9999  (.A(WX5760), .B(WX6237), .Z(WX6236) ) ;
NAND2   gate10000  (.A(II19190), .B(II19191), .Z(WX6241) ) ;
AND2    gate10001  (.A(WX6241), .B(WX6177), .Z(WX6242) ) ;
AND2    gate10002  (.A(WX5761), .B(WX6244), .Z(WX6243) ) ;
NAND2   gate10003  (.A(II19203), .B(II19204), .Z(WX6248) ) ;
AND2    gate10004  (.A(WX6248), .B(WX6177), .Z(WX6249) ) ;
AND2    gate10005  (.A(WX5762), .B(WX6251), .Z(WX6250) ) ;
NAND2   gate10006  (.A(II19216), .B(II19217), .Z(WX6255) ) ;
AND2    gate10007  (.A(WX6255), .B(WX6177), .Z(WX6256) ) ;
AND2    gate10008  (.A(WX5763), .B(WX6258), .Z(WX6257) ) ;
NAND2   gate10009  (.A(II19229), .B(II19230), .Z(WX6262) ) ;
AND2    gate10010  (.A(WX6262), .B(WX6177), .Z(WX6263) ) ;
AND2    gate10011  (.A(WX5764), .B(WX6265), .Z(WX6264) ) ;
NAND2   gate10012  (.A(II19242), .B(II19243), .Z(WX6269) ) ;
AND2    gate10013  (.A(WX6269), .B(WX6177), .Z(WX6270) ) ;
AND2    gate10014  (.A(WX5765), .B(WX6272), .Z(WX6271) ) ;
NAND2   gate10015  (.A(II19255), .B(II19256), .Z(WX6276) ) ;
AND2    gate10016  (.A(WX6276), .B(WX6177), .Z(WX6277) ) ;
AND2    gate10017  (.A(WX5766), .B(WX6279), .Z(WX6278) ) ;
NAND2   gate10018  (.A(II19268), .B(II19269), .Z(WX6283) ) ;
AND2    gate10019  (.A(WX6283), .B(WX6177), .Z(WX6284) ) ;
AND2    gate10020  (.A(WX5767), .B(WX6286), .Z(WX6285) ) ;
NAND2   gate10021  (.A(II19281), .B(II19282), .Z(WX6290) ) ;
AND2    gate10022  (.A(WX6290), .B(WX6177), .Z(WX6291) ) ;
AND2    gate10023  (.A(WX5768), .B(WX6293), .Z(WX6292) ) ;
NAND2   gate10024  (.A(II19294), .B(II19295), .Z(WX6297) ) ;
AND2    gate10025  (.A(WX6297), .B(WX6177), .Z(WX6298) ) ;
AND2    gate10026  (.A(WX5769), .B(WX6300), .Z(WX6299) ) ;
NAND2   gate10027  (.A(II19307), .B(II19308), .Z(WX6304) ) ;
AND2    gate10028  (.A(WX6304), .B(WX6177), .Z(WX6305) ) ;
AND2    gate10029  (.A(WX5770), .B(WX6307), .Z(WX6306) ) ;
NAND2   gate10030  (.A(II19320), .B(II19321), .Z(WX6311) ) ;
AND2    gate10031  (.A(WX6311), .B(WX6177), .Z(WX6312) ) ;
AND2    gate10032  (.A(WX5771), .B(WX6314), .Z(WX6313) ) ;
NAND2   gate10033  (.A(II19333), .B(II19334), .Z(WX6318) ) ;
AND2    gate10034  (.A(WX6318), .B(WX6177), .Z(WX6319) ) ;
AND2    gate10035  (.A(WX5772), .B(WX6321), .Z(WX6320) ) ;
NAND2   gate10036  (.A(II19346), .B(II19347), .Z(WX6325) ) ;
AND2    gate10037  (.A(WX6325), .B(WX6177), .Z(WX6326) ) ;
AND2    gate10038  (.A(WX5773), .B(WX6328), .Z(WX6327) ) ;
NAND2   gate10039  (.A(II19359), .B(II19360), .Z(WX6332) ) ;
AND2    gate10040  (.A(WX6332), .B(WX6177), .Z(WX6333) ) ;
AND2    gate10041  (.A(WX5774), .B(WX6335), .Z(WX6334) ) ;
NAND2   gate10042  (.A(II19372), .B(II19373), .Z(WX6339) ) ;
AND2    gate10043  (.A(WX6339), .B(WX6177), .Z(WX6340) ) ;
AND2    gate10044  (.A(WX5775), .B(WX6342), .Z(WX6341) ) ;
NAND2   gate10045  (.A(II19385), .B(II19386), .Z(WX6346) ) ;
AND2    gate10046  (.A(WX6346), .B(WX6177), .Z(WX6347) ) ;
AND2    gate10047  (.A(WX5776), .B(WX6349), .Z(WX6348) ) ;
NAND2   gate10048  (.A(II19398), .B(II19399), .Z(WX6353) ) ;
AND2    gate10049  (.A(WX6353), .B(WX6177), .Z(WX6354) ) ;
AND2    gate10050  (.A(WX5777), .B(WX6356), .Z(WX6355) ) ;
NAND2   gate10051  (.A(II19411), .B(II19412), .Z(WX6360) ) ;
AND2    gate10052  (.A(WX6360), .B(WX6177), .Z(WX6361) ) ;
AND2    gate10053  (.A(WX5778), .B(WX6363), .Z(WX6362) ) ;
NAND2   gate10054  (.A(II19424), .B(II19425), .Z(WX6367) ) ;
AND2    gate10055  (.A(WX6367), .B(WX6177), .Z(WX6368) ) ;
AND2    gate10056  (.A(WX5779), .B(WX6370), .Z(WX6369) ) ;
NAND2   gate10057  (.A(II19437), .B(II19438), .Z(WX6374) ) ;
AND2    gate10058  (.A(WX6374), .B(WX6177), .Z(WX6375) ) ;
AND2    gate10059  (.A(WX5780), .B(WX6377), .Z(WX6376) ) ;
NAND2   gate10060  (.A(II19450), .B(II19451), .Z(WX6381) ) ;
AND2    gate10061  (.A(WX6381), .B(WX6177), .Z(WX6382) ) ;
AND2    gate10062  (.A(WX5781), .B(WX6384), .Z(WX6383) ) ;
NAND2   gate10063  (.A(II19463), .B(II19464), .Z(WX6388) ) ;
AND2    gate10064  (.A(WX6388), .B(WX6177), .Z(WX6389) ) ;
AND2    gate10065  (.A(WX5782), .B(WX6391), .Z(WX6390) ) ;
NAND2   gate10066  (.A(II19476), .B(II19477), .Z(WX6395) ) ;
AND2    gate10067  (.A(WX6395), .B(WX6177), .Z(WX6396) ) ;
AND2    gate10068  (.A(WX5783), .B(WX6398), .Z(WX6397) ) ;
NAND2   gate10069  (.A(II19535), .B(II19536), .Z(WX6406) ) ;
NAND2   gate10070  (.A(II19731), .B(II19732), .Z(WX6434) ) ;
NAND2   gate10071  (.A(II19724), .B(II19725), .Z(WX6433) ) ;
NAND2   gate10072  (.A(II19717), .B(II19718), .Z(WX6432) ) ;
NAND2   gate10073  (.A(II19528), .B(II19529), .Z(WX6405) ) ;
NAND2   gate10074  (.A(II19710), .B(II19711), .Z(WX6431) ) ;
NAND2   gate10075  (.A(II19703), .B(II19704), .Z(WX6430) ) ;
NAND2   gate10076  (.A(II19696), .B(II19697), .Z(WX6429) ) ;
NAND2   gate10077  (.A(II19689), .B(II19690), .Z(WX6428) ) ;
NAND2   gate10078  (.A(II19682), .B(II19683), .Z(WX6427) ) ;
NAND2   gate10079  (.A(II19675), .B(II19676), .Z(WX6426) ) ;
NAND2   gate10080  (.A(II19513), .B(II19514), .Z(WX6404) ) ;
NAND2   gate10081  (.A(II19668), .B(II19669), .Z(WX6425) ) ;
NAND2   gate10082  (.A(II19661), .B(II19662), .Z(WX6424) ) ;
NAND2   gate10083  (.A(II19654), .B(II19655), .Z(WX6423) ) ;
NAND2   gate10084  (.A(II19647), .B(II19648), .Z(WX6422) ) ;
NAND2   gate10085  (.A(II19498), .B(II19499), .Z(WX6403) ) ;
NAND2   gate10086  (.A(II19640), .B(II19641), .Z(WX6421) ) ;
NAND2   gate10087  (.A(II19633), .B(II19634), .Z(WX6420) ) ;
NAND2   gate10088  (.A(II19626), .B(II19627), .Z(WX6419) ) ;
NAND2   gate10089  (.A(II19619), .B(II19620), .Z(WX6418) ) ;
NAND2   gate10090  (.A(II19612), .B(II19613), .Z(WX6417) ) ;
NAND2   gate10091  (.A(II19605), .B(II19606), .Z(WX6416) ) ;
NAND2   gate10092  (.A(II19598), .B(II19599), .Z(WX6415) ) ;
NAND2   gate10093  (.A(II19591), .B(II19592), .Z(WX6414) ) ;
NAND2   gate10094  (.A(II19584), .B(II19585), .Z(WX6413) ) ;
NAND2   gate10095  (.A(II19577), .B(II19578), .Z(WX6412) ) ;
NAND2   gate10096  (.A(II19570), .B(II19571), .Z(WX6411) ) ;
NAND2   gate10097  (.A(II19563), .B(II19564), .Z(WX6410) ) ;
NAND2   gate10098  (.A(II19556), .B(II19557), .Z(WX6409) ) ;
NAND2   gate10099  (.A(II19549), .B(II19550), .Z(WX6408) ) ;
NAND2   gate10100  (.A(II19542), .B(II19543), .Z(WX6407) ) ;
OR2     gate10101  (.A(WX6509), .B(WX6508), .Z(WX6511) ) ;
AND2    gate10102  (.A(WX6511), .B(WX7468), .Z(WX6500) ) ;
OR2     gate10103  (.A(WX6505), .B(WX6504), .Z(WX6507) ) ;
AND2    gate10104  (.A(WX6507), .B(WX6502), .Z(WX6501) ) ;
AND2    gate10105  (.A(CRC_OUT_4_31), .B(WX7469), .Z(WX6504) ) ;
AND2    gate10106  (.A(WX8770), .B(WX6506), .Z(WX6505) ) ;
AND2    gate10107  (.A(WX6950), .B(WX7469), .Z(WX6508) ) ;
AND2    gate10108  (.A(WX7477), .B(WX6510), .Z(WX6509) ) ;
OR2     gate10109  (.A(WX6523), .B(WX6522), .Z(WX6525) ) ;
AND2    gate10110  (.A(WX6525), .B(WX7468), .Z(WX6514) ) ;
OR2     gate10111  (.A(WX6519), .B(WX6518), .Z(WX6521) ) ;
AND2    gate10112  (.A(WX6521), .B(WX6516), .Z(WX6515) ) ;
AND2    gate10113  (.A(CRC_OUT_4_30), .B(WX7469), .Z(WX6518) ) ;
AND2    gate10114  (.A(WX8777), .B(WX6520), .Z(WX6519) ) ;
AND2    gate10115  (.A(WX6952), .B(WX7469), .Z(WX6522) ) ;
AND2    gate10116  (.A(WX7484), .B(WX6524), .Z(WX6523) ) ;
OR2     gate10117  (.A(WX6537), .B(WX6536), .Z(WX6539) ) ;
AND2    gate10118  (.A(WX6539), .B(WX7468), .Z(WX6528) ) ;
OR2     gate10119  (.A(WX6533), .B(WX6532), .Z(WX6535) ) ;
AND2    gate10120  (.A(WX6535), .B(WX6530), .Z(WX6529) ) ;
AND2    gate10121  (.A(CRC_OUT_4_29), .B(WX7469), .Z(WX6532) ) ;
AND2    gate10122  (.A(WX8784), .B(WX6534), .Z(WX6533) ) ;
AND2    gate10123  (.A(WX6954), .B(WX7469), .Z(WX6536) ) ;
AND2    gate10124  (.A(WX7491), .B(WX6538), .Z(WX6537) ) ;
OR2     gate10125  (.A(WX6551), .B(WX6550), .Z(WX6553) ) ;
AND2    gate10126  (.A(WX6553), .B(WX7468), .Z(WX6542) ) ;
OR2     gate10127  (.A(WX6547), .B(WX6546), .Z(WX6549) ) ;
AND2    gate10128  (.A(WX6549), .B(WX6544), .Z(WX6543) ) ;
AND2    gate10129  (.A(CRC_OUT_4_28), .B(WX7469), .Z(WX6546) ) ;
AND2    gate10130  (.A(WX8791), .B(WX6548), .Z(WX6547) ) ;
AND2    gate10131  (.A(WX6956), .B(WX7469), .Z(WX6550) ) ;
AND2    gate10132  (.A(WX7498), .B(WX6552), .Z(WX6551) ) ;
OR2     gate10133  (.A(WX6565), .B(WX6564), .Z(WX6567) ) ;
AND2    gate10134  (.A(WX6567), .B(WX7468), .Z(WX6556) ) ;
OR2     gate10135  (.A(WX6561), .B(WX6560), .Z(WX6563) ) ;
AND2    gate10136  (.A(WX6563), .B(WX6558), .Z(WX6557) ) ;
AND2    gate10137  (.A(CRC_OUT_4_27), .B(WX7469), .Z(WX6560) ) ;
AND2    gate10138  (.A(WX8798), .B(WX6562), .Z(WX6561) ) ;
AND2    gate10139  (.A(WX6958), .B(WX7469), .Z(WX6564) ) ;
AND2    gate10140  (.A(WX7505), .B(WX6566), .Z(WX6565) ) ;
OR2     gate10141  (.A(WX6579), .B(WX6578), .Z(WX6581) ) ;
AND2    gate10142  (.A(WX6581), .B(WX7468), .Z(WX6570) ) ;
OR2     gate10143  (.A(WX6575), .B(WX6574), .Z(WX6577) ) ;
AND2    gate10144  (.A(WX6577), .B(WX6572), .Z(WX6571) ) ;
AND2    gate10145  (.A(CRC_OUT_4_26), .B(WX7469), .Z(WX6574) ) ;
AND2    gate10146  (.A(WX8805), .B(WX6576), .Z(WX6575) ) ;
AND2    gate10147  (.A(WX6960), .B(WX7469), .Z(WX6578) ) ;
AND2    gate10148  (.A(WX7512), .B(WX6580), .Z(WX6579) ) ;
OR2     gate10149  (.A(WX6593), .B(WX6592), .Z(WX6595) ) ;
AND2    gate10150  (.A(WX6595), .B(WX7468), .Z(WX6584) ) ;
OR2     gate10151  (.A(WX6589), .B(WX6588), .Z(WX6591) ) ;
AND2    gate10152  (.A(WX6591), .B(WX6586), .Z(WX6585) ) ;
AND2    gate10153  (.A(CRC_OUT_4_25), .B(WX7469), .Z(WX6588) ) ;
AND2    gate10154  (.A(WX8812), .B(WX6590), .Z(WX6589) ) ;
AND2    gate10155  (.A(WX6962), .B(WX7469), .Z(WX6592) ) ;
AND2    gate10156  (.A(WX7519), .B(WX6594), .Z(WX6593) ) ;
OR2     gate10157  (.A(WX6607), .B(WX6606), .Z(WX6609) ) ;
AND2    gate10158  (.A(WX6609), .B(WX7468), .Z(WX6598) ) ;
OR2     gate10159  (.A(WX6603), .B(WX6602), .Z(WX6605) ) ;
AND2    gate10160  (.A(WX6605), .B(WX6600), .Z(WX6599) ) ;
AND2    gate10161  (.A(CRC_OUT_4_24), .B(WX7469), .Z(WX6602) ) ;
AND2    gate10162  (.A(WX8819), .B(WX6604), .Z(WX6603) ) ;
AND2    gate10163  (.A(WX6964), .B(WX7469), .Z(WX6606) ) ;
AND2    gate10164  (.A(WX7526), .B(WX6608), .Z(WX6607) ) ;
OR2     gate10165  (.A(WX6621), .B(WX6620), .Z(WX6623) ) ;
AND2    gate10166  (.A(WX6623), .B(WX7468), .Z(WX6612) ) ;
OR2     gate10167  (.A(WX6617), .B(WX6616), .Z(WX6619) ) ;
AND2    gate10168  (.A(WX6619), .B(WX6614), .Z(WX6613) ) ;
AND2    gate10169  (.A(CRC_OUT_4_23), .B(WX7469), .Z(WX6616) ) ;
AND2    gate10170  (.A(WX8826), .B(WX6618), .Z(WX6617) ) ;
AND2    gate10171  (.A(WX6966), .B(WX7469), .Z(WX6620) ) ;
AND2    gate10172  (.A(WX7533), .B(WX6622), .Z(WX6621) ) ;
OR2     gate10173  (.A(WX6635), .B(WX6634), .Z(WX6637) ) ;
AND2    gate10174  (.A(WX6637), .B(WX7468), .Z(WX6626) ) ;
OR2     gate10175  (.A(WX6631), .B(WX6630), .Z(WX6633) ) ;
AND2    gate10176  (.A(WX6633), .B(WX6628), .Z(WX6627) ) ;
AND2    gate10177  (.A(CRC_OUT_4_22), .B(WX7469), .Z(WX6630) ) ;
AND2    gate10178  (.A(WX8833), .B(WX6632), .Z(WX6631) ) ;
AND2    gate10179  (.A(WX6968), .B(WX7469), .Z(WX6634) ) ;
AND2    gate10180  (.A(WX7540), .B(WX6636), .Z(WX6635) ) ;
OR2     gate10181  (.A(WX6649), .B(WX6648), .Z(WX6651) ) ;
AND2    gate10182  (.A(WX6651), .B(WX7468), .Z(WX6640) ) ;
OR2     gate10183  (.A(WX6645), .B(WX6644), .Z(WX6647) ) ;
AND2    gate10184  (.A(WX6647), .B(WX6642), .Z(WX6641) ) ;
AND2    gate10185  (.A(CRC_OUT_4_21), .B(WX7469), .Z(WX6644) ) ;
AND2    gate10186  (.A(WX8840), .B(WX6646), .Z(WX6645) ) ;
AND2    gate10187  (.A(WX6970), .B(WX7469), .Z(WX6648) ) ;
AND2    gate10188  (.A(WX7547), .B(WX6650), .Z(WX6649) ) ;
OR2     gate10189  (.A(WX6663), .B(WX6662), .Z(WX6665) ) ;
AND2    gate10190  (.A(WX6665), .B(WX7468), .Z(WX6654) ) ;
OR2     gate10191  (.A(WX6659), .B(WX6658), .Z(WX6661) ) ;
AND2    gate10192  (.A(WX6661), .B(WX6656), .Z(WX6655) ) ;
AND2    gate10193  (.A(CRC_OUT_4_20), .B(WX7469), .Z(WX6658) ) ;
AND2    gate10194  (.A(WX8847), .B(WX6660), .Z(WX6659) ) ;
AND2    gate10195  (.A(WX6972), .B(WX7469), .Z(WX6662) ) ;
AND2    gate10196  (.A(WX7554), .B(WX6664), .Z(WX6663) ) ;
OR2     gate10197  (.A(WX6677), .B(WX6676), .Z(WX6679) ) ;
AND2    gate10198  (.A(WX6679), .B(WX7468), .Z(WX6668) ) ;
OR2     gate10199  (.A(WX6673), .B(WX6672), .Z(WX6675) ) ;
AND2    gate10200  (.A(WX6675), .B(WX6670), .Z(WX6669) ) ;
AND2    gate10201  (.A(CRC_OUT_4_19), .B(WX7469), .Z(WX6672) ) ;
AND2    gate10202  (.A(WX8854), .B(WX6674), .Z(WX6673) ) ;
AND2    gate10203  (.A(WX6974), .B(WX7469), .Z(WX6676) ) ;
AND2    gate10204  (.A(WX7561), .B(WX6678), .Z(WX6677) ) ;
OR2     gate10205  (.A(WX6691), .B(WX6690), .Z(WX6693) ) ;
AND2    gate10206  (.A(WX6693), .B(WX7468), .Z(WX6682) ) ;
OR2     gate10207  (.A(WX6687), .B(WX6686), .Z(WX6689) ) ;
AND2    gate10208  (.A(WX6689), .B(WX6684), .Z(WX6683) ) ;
AND2    gate10209  (.A(CRC_OUT_4_18), .B(WX7469), .Z(WX6686) ) ;
AND2    gate10210  (.A(WX8861), .B(WX6688), .Z(WX6687) ) ;
AND2    gate10211  (.A(WX6976), .B(WX7469), .Z(WX6690) ) ;
AND2    gate10212  (.A(WX7568), .B(WX6692), .Z(WX6691) ) ;
OR2     gate10213  (.A(WX6705), .B(WX6704), .Z(WX6707) ) ;
AND2    gate10214  (.A(WX6707), .B(WX7468), .Z(WX6696) ) ;
OR2     gate10215  (.A(WX6701), .B(WX6700), .Z(WX6703) ) ;
AND2    gate10216  (.A(WX6703), .B(WX6698), .Z(WX6697) ) ;
AND2    gate10217  (.A(CRC_OUT_4_17), .B(WX7469), .Z(WX6700) ) ;
AND2    gate10218  (.A(WX8868), .B(WX6702), .Z(WX6701) ) ;
AND2    gate10219  (.A(WX6978), .B(WX7469), .Z(WX6704) ) ;
AND2    gate10220  (.A(WX7575), .B(WX6706), .Z(WX6705) ) ;
OR2     gate10221  (.A(WX6719), .B(WX6718), .Z(WX6721) ) ;
AND2    gate10222  (.A(WX6721), .B(WX7468), .Z(WX6710) ) ;
OR2     gate10223  (.A(WX6715), .B(WX6714), .Z(WX6717) ) ;
AND2    gate10224  (.A(WX6717), .B(WX6712), .Z(WX6711) ) ;
AND2    gate10225  (.A(CRC_OUT_4_16), .B(WX7469), .Z(WX6714) ) ;
AND2    gate10226  (.A(WX8875), .B(WX6716), .Z(WX6715) ) ;
AND2    gate10227  (.A(WX6980), .B(WX7469), .Z(WX6718) ) ;
AND2    gate10228  (.A(WX7582), .B(WX6720), .Z(WX6719) ) ;
OR2     gate10229  (.A(WX6733), .B(WX6732), .Z(WX6735) ) ;
AND2    gate10230  (.A(WX6735), .B(WX7468), .Z(WX6724) ) ;
OR2     gate10231  (.A(WX6729), .B(WX6728), .Z(WX6731) ) ;
AND2    gate10232  (.A(WX6731), .B(WX6726), .Z(WX6725) ) ;
AND2    gate10233  (.A(CRC_OUT_4_15), .B(WX7469), .Z(WX6728) ) ;
AND2    gate10234  (.A(WX8882), .B(WX6730), .Z(WX6729) ) ;
AND2    gate10235  (.A(WX6982), .B(WX7469), .Z(WX6732) ) ;
AND2    gate10236  (.A(WX7589), .B(WX6734), .Z(WX6733) ) ;
OR2     gate10237  (.A(WX6747), .B(WX6746), .Z(WX6749) ) ;
AND2    gate10238  (.A(WX6749), .B(WX7468), .Z(WX6738) ) ;
OR2     gate10239  (.A(WX6743), .B(WX6742), .Z(WX6745) ) ;
AND2    gate10240  (.A(WX6745), .B(WX6740), .Z(WX6739) ) ;
AND2    gate10241  (.A(CRC_OUT_4_14), .B(WX7469), .Z(WX6742) ) ;
AND2    gate10242  (.A(WX8889), .B(WX6744), .Z(WX6743) ) ;
AND2    gate10243  (.A(WX6984), .B(WX7469), .Z(WX6746) ) ;
AND2    gate10244  (.A(WX7596), .B(WX6748), .Z(WX6747) ) ;
OR2     gate10245  (.A(WX6761), .B(WX6760), .Z(WX6763) ) ;
AND2    gate10246  (.A(WX6763), .B(WX7468), .Z(WX6752) ) ;
OR2     gate10247  (.A(WX6757), .B(WX6756), .Z(WX6759) ) ;
AND2    gate10248  (.A(WX6759), .B(WX6754), .Z(WX6753) ) ;
AND2    gate10249  (.A(CRC_OUT_4_13), .B(WX7469), .Z(WX6756) ) ;
AND2    gate10250  (.A(WX8896), .B(WX6758), .Z(WX6757) ) ;
AND2    gate10251  (.A(WX6986), .B(WX7469), .Z(WX6760) ) ;
AND2    gate10252  (.A(WX7603), .B(WX6762), .Z(WX6761) ) ;
OR2     gate10253  (.A(WX6775), .B(WX6774), .Z(WX6777) ) ;
AND2    gate10254  (.A(WX6777), .B(WX7468), .Z(WX6766) ) ;
OR2     gate10255  (.A(WX6771), .B(WX6770), .Z(WX6773) ) ;
AND2    gate10256  (.A(WX6773), .B(WX6768), .Z(WX6767) ) ;
AND2    gate10257  (.A(CRC_OUT_4_12), .B(WX7469), .Z(WX6770) ) ;
AND2    gate10258  (.A(WX8903), .B(WX6772), .Z(WX6771) ) ;
AND2    gate10259  (.A(WX6988), .B(WX7469), .Z(WX6774) ) ;
AND2    gate10260  (.A(WX7610), .B(WX6776), .Z(WX6775) ) ;
OR2     gate10261  (.A(WX6789), .B(WX6788), .Z(WX6791) ) ;
AND2    gate10262  (.A(WX6791), .B(WX7468), .Z(WX6780) ) ;
OR2     gate10263  (.A(WX6785), .B(WX6784), .Z(WX6787) ) ;
AND2    gate10264  (.A(WX6787), .B(WX6782), .Z(WX6781) ) ;
AND2    gate10265  (.A(CRC_OUT_4_11), .B(WX7469), .Z(WX6784) ) ;
AND2    gate10266  (.A(WX8910), .B(WX6786), .Z(WX6785) ) ;
AND2    gate10267  (.A(WX6990), .B(WX7469), .Z(WX6788) ) ;
AND2    gate10268  (.A(WX7617), .B(WX6790), .Z(WX6789) ) ;
OR2     gate10269  (.A(WX6803), .B(WX6802), .Z(WX6805) ) ;
AND2    gate10270  (.A(WX6805), .B(WX7468), .Z(WX6794) ) ;
OR2     gate10271  (.A(WX6799), .B(WX6798), .Z(WX6801) ) ;
AND2    gate10272  (.A(WX6801), .B(WX6796), .Z(WX6795) ) ;
AND2    gate10273  (.A(CRC_OUT_4_10), .B(WX7469), .Z(WX6798) ) ;
AND2    gate10274  (.A(WX8917), .B(WX6800), .Z(WX6799) ) ;
AND2    gate10275  (.A(WX6992), .B(WX7469), .Z(WX6802) ) ;
AND2    gate10276  (.A(WX7624), .B(WX6804), .Z(WX6803) ) ;
OR2     gate10277  (.A(WX6817), .B(WX6816), .Z(WX6819) ) ;
AND2    gate10278  (.A(WX6819), .B(WX7468), .Z(WX6808) ) ;
OR2     gate10279  (.A(WX6813), .B(WX6812), .Z(WX6815) ) ;
AND2    gate10280  (.A(WX6815), .B(WX6810), .Z(WX6809) ) ;
AND2    gate10281  (.A(CRC_OUT_4_9), .B(WX7469), .Z(WX6812) ) ;
AND2    gate10282  (.A(WX8924), .B(WX6814), .Z(WX6813) ) ;
AND2    gate10283  (.A(WX6994), .B(WX7469), .Z(WX6816) ) ;
AND2    gate10284  (.A(WX7631), .B(WX6818), .Z(WX6817) ) ;
OR2     gate10285  (.A(WX6831), .B(WX6830), .Z(WX6833) ) ;
AND2    gate10286  (.A(WX6833), .B(WX7468), .Z(WX6822) ) ;
OR2     gate10287  (.A(WX6827), .B(WX6826), .Z(WX6829) ) ;
AND2    gate10288  (.A(WX6829), .B(WX6824), .Z(WX6823) ) ;
AND2    gate10289  (.A(CRC_OUT_4_8), .B(WX7469), .Z(WX6826) ) ;
AND2    gate10290  (.A(WX8931), .B(WX6828), .Z(WX6827) ) ;
AND2    gate10291  (.A(WX6996), .B(WX7469), .Z(WX6830) ) ;
AND2    gate10292  (.A(WX7638), .B(WX6832), .Z(WX6831) ) ;
OR2     gate10293  (.A(WX6845), .B(WX6844), .Z(WX6847) ) ;
AND2    gate10294  (.A(WX6847), .B(WX7468), .Z(WX6836) ) ;
OR2     gate10295  (.A(WX6841), .B(WX6840), .Z(WX6843) ) ;
AND2    gate10296  (.A(WX6843), .B(WX6838), .Z(WX6837) ) ;
AND2    gate10297  (.A(CRC_OUT_4_7), .B(WX7469), .Z(WX6840) ) ;
AND2    gate10298  (.A(WX8938), .B(WX6842), .Z(WX6841) ) ;
AND2    gate10299  (.A(WX6998), .B(WX7469), .Z(WX6844) ) ;
AND2    gate10300  (.A(WX7645), .B(WX6846), .Z(WX6845) ) ;
OR2     gate10301  (.A(WX6859), .B(WX6858), .Z(WX6861) ) ;
AND2    gate10302  (.A(WX6861), .B(WX7468), .Z(WX6850) ) ;
OR2     gate10303  (.A(WX6855), .B(WX6854), .Z(WX6857) ) ;
AND2    gate10304  (.A(WX6857), .B(WX6852), .Z(WX6851) ) ;
AND2    gate10305  (.A(CRC_OUT_4_6), .B(WX7469), .Z(WX6854) ) ;
AND2    gate10306  (.A(WX8945), .B(WX6856), .Z(WX6855) ) ;
AND2    gate10307  (.A(WX7000), .B(WX7469), .Z(WX6858) ) ;
AND2    gate10308  (.A(WX7652), .B(WX6860), .Z(WX6859) ) ;
OR2     gate10309  (.A(WX6873), .B(WX6872), .Z(WX6875) ) ;
AND2    gate10310  (.A(WX6875), .B(WX7468), .Z(WX6864) ) ;
OR2     gate10311  (.A(WX6869), .B(WX6868), .Z(WX6871) ) ;
AND2    gate10312  (.A(WX6871), .B(WX6866), .Z(WX6865) ) ;
AND2    gate10313  (.A(CRC_OUT_4_5), .B(WX7469), .Z(WX6868) ) ;
AND2    gate10314  (.A(WX8952), .B(WX6870), .Z(WX6869) ) ;
AND2    gate10315  (.A(WX7002), .B(WX7469), .Z(WX6872) ) ;
AND2    gate10316  (.A(WX7659), .B(WX6874), .Z(WX6873) ) ;
OR2     gate10317  (.A(WX6887), .B(WX6886), .Z(WX6889) ) ;
AND2    gate10318  (.A(WX6889), .B(WX7468), .Z(WX6878) ) ;
OR2     gate10319  (.A(WX6883), .B(WX6882), .Z(WX6885) ) ;
AND2    gate10320  (.A(WX6885), .B(WX6880), .Z(WX6879) ) ;
AND2    gate10321  (.A(CRC_OUT_4_4), .B(WX7469), .Z(WX6882) ) ;
AND2    gate10322  (.A(WX8959), .B(WX6884), .Z(WX6883) ) ;
AND2    gate10323  (.A(WX7004), .B(WX7469), .Z(WX6886) ) ;
AND2    gate10324  (.A(WX7666), .B(WX6888), .Z(WX6887) ) ;
OR2     gate10325  (.A(WX6901), .B(WX6900), .Z(WX6903) ) ;
AND2    gate10326  (.A(WX6903), .B(WX7468), .Z(WX6892) ) ;
OR2     gate10327  (.A(WX6897), .B(WX6896), .Z(WX6899) ) ;
AND2    gate10328  (.A(WX6899), .B(WX6894), .Z(WX6893) ) ;
AND2    gate10329  (.A(CRC_OUT_4_3), .B(WX7469), .Z(WX6896) ) ;
AND2    gate10330  (.A(WX8966), .B(WX6898), .Z(WX6897) ) ;
AND2    gate10331  (.A(WX7006), .B(WX7469), .Z(WX6900) ) ;
AND2    gate10332  (.A(WX7673), .B(WX6902), .Z(WX6901) ) ;
OR2     gate10333  (.A(WX6915), .B(WX6914), .Z(WX6917) ) ;
AND2    gate10334  (.A(WX6917), .B(WX7468), .Z(WX6906) ) ;
OR2     gate10335  (.A(WX6911), .B(WX6910), .Z(WX6913) ) ;
AND2    gate10336  (.A(WX6913), .B(WX6908), .Z(WX6907) ) ;
AND2    gate10337  (.A(CRC_OUT_4_2), .B(WX7469), .Z(WX6910) ) ;
AND2    gate10338  (.A(WX8973), .B(WX6912), .Z(WX6911) ) ;
AND2    gate10339  (.A(WX7008), .B(WX7469), .Z(WX6914) ) ;
AND2    gate10340  (.A(WX7680), .B(WX6916), .Z(WX6915) ) ;
OR2     gate10341  (.A(WX6929), .B(WX6928), .Z(WX6931) ) ;
AND2    gate10342  (.A(WX6931), .B(WX7468), .Z(WX6920) ) ;
OR2     gate10343  (.A(WX6925), .B(WX6924), .Z(WX6927) ) ;
AND2    gate10344  (.A(WX6927), .B(WX6922), .Z(WX6921) ) ;
AND2    gate10345  (.A(CRC_OUT_4_1), .B(WX7469), .Z(WX6924) ) ;
AND2    gate10346  (.A(WX8980), .B(WX6926), .Z(WX6925) ) ;
AND2    gate10347  (.A(WX7010), .B(WX7469), .Z(WX6928) ) ;
AND2    gate10348  (.A(WX7687), .B(WX6930), .Z(WX6929) ) ;
OR2     gate10349  (.A(WX6943), .B(WX6942), .Z(WX6945) ) ;
AND2    gate10350  (.A(WX6945), .B(WX7468), .Z(WX6934) ) ;
OR2     gate10351  (.A(WX6939), .B(WX6938), .Z(WX6941) ) ;
AND2    gate10352  (.A(WX6941), .B(WX6936), .Z(WX6935) ) ;
AND2    gate10353  (.A(CRC_OUT_4_0), .B(WX7469), .Z(WX6938) ) ;
AND2    gate10354  (.A(WX8987), .B(WX6940), .Z(WX6939) ) ;
AND2    gate10355  (.A(WX7012), .B(WX7469), .Z(WX6942) ) ;
AND2    gate10356  (.A(WX7694), .B(WX6944), .Z(WX6943) ) ;
NAND2   gate10357  (.A(II23078), .B(II23079), .Z(WX7471) ) ;
AND2    gate10358  (.A(WX7471), .B(WX7470), .Z(WX7472) ) ;
AND2    gate10359  (.A(WX7045), .B(WX7474), .Z(WX7473) ) ;
NAND2   gate10360  (.A(II23091), .B(II23092), .Z(WX7478) ) ;
AND2    gate10361  (.A(WX7478), .B(WX7470), .Z(WX7479) ) ;
AND2    gate10362  (.A(WX7046), .B(WX7481), .Z(WX7480) ) ;
NAND2   gate10363  (.A(II23104), .B(II23105), .Z(WX7485) ) ;
AND2    gate10364  (.A(WX7485), .B(WX7470), .Z(WX7486) ) ;
AND2    gate10365  (.A(WX7047), .B(WX7488), .Z(WX7487) ) ;
NAND2   gate10366  (.A(II23117), .B(II23118), .Z(WX7492) ) ;
AND2    gate10367  (.A(WX7492), .B(WX7470), .Z(WX7493) ) ;
AND2    gate10368  (.A(WX7048), .B(WX7495), .Z(WX7494) ) ;
NAND2   gate10369  (.A(II23130), .B(II23131), .Z(WX7499) ) ;
AND2    gate10370  (.A(WX7499), .B(WX7470), .Z(WX7500) ) ;
AND2    gate10371  (.A(WX7049), .B(WX7502), .Z(WX7501) ) ;
NAND2   gate10372  (.A(II23143), .B(II23144), .Z(WX7506) ) ;
AND2    gate10373  (.A(WX7506), .B(WX7470), .Z(WX7507) ) ;
AND2    gate10374  (.A(WX7050), .B(WX7509), .Z(WX7508) ) ;
NAND2   gate10375  (.A(II23156), .B(II23157), .Z(WX7513) ) ;
AND2    gate10376  (.A(WX7513), .B(WX7470), .Z(WX7514) ) ;
AND2    gate10377  (.A(WX7051), .B(WX7516), .Z(WX7515) ) ;
NAND2   gate10378  (.A(II23169), .B(II23170), .Z(WX7520) ) ;
AND2    gate10379  (.A(WX7520), .B(WX7470), .Z(WX7521) ) ;
AND2    gate10380  (.A(WX7052), .B(WX7523), .Z(WX7522) ) ;
NAND2   gate10381  (.A(II23182), .B(II23183), .Z(WX7527) ) ;
AND2    gate10382  (.A(WX7527), .B(WX7470), .Z(WX7528) ) ;
AND2    gate10383  (.A(WX7053), .B(WX7530), .Z(WX7529) ) ;
NAND2   gate10384  (.A(II23195), .B(II23196), .Z(WX7534) ) ;
AND2    gate10385  (.A(WX7534), .B(WX7470), .Z(WX7535) ) ;
AND2    gate10386  (.A(WX7054), .B(WX7537), .Z(WX7536) ) ;
NAND2   gate10387  (.A(II23208), .B(II23209), .Z(WX7541) ) ;
AND2    gate10388  (.A(WX7541), .B(WX7470), .Z(WX7542) ) ;
AND2    gate10389  (.A(WX7055), .B(WX7544), .Z(WX7543) ) ;
NAND2   gate10390  (.A(II23221), .B(II23222), .Z(WX7548) ) ;
AND2    gate10391  (.A(WX7548), .B(WX7470), .Z(WX7549) ) ;
AND2    gate10392  (.A(WX7056), .B(WX7551), .Z(WX7550) ) ;
NAND2   gate10393  (.A(II23234), .B(II23235), .Z(WX7555) ) ;
AND2    gate10394  (.A(WX7555), .B(WX7470), .Z(WX7556) ) ;
AND2    gate10395  (.A(WX7057), .B(WX7558), .Z(WX7557) ) ;
NAND2   gate10396  (.A(II23247), .B(II23248), .Z(WX7562) ) ;
AND2    gate10397  (.A(WX7562), .B(WX7470), .Z(WX7563) ) ;
AND2    gate10398  (.A(WX7058), .B(WX7565), .Z(WX7564) ) ;
NAND2   gate10399  (.A(II23260), .B(II23261), .Z(WX7569) ) ;
AND2    gate10400  (.A(WX7569), .B(WX7470), .Z(WX7570) ) ;
AND2    gate10401  (.A(WX7059), .B(WX7572), .Z(WX7571) ) ;
NAND2   gate10402  (.A(II23273), .B(II23274), .Z(WX7576) ) ;
AND2    gate10403  (.A(WX7576), .B(WX7470), .Z(WX7577) ) ;
AND2    gate10404  (.A(WX7060), .B(WX7579), .Z(WX7578) ) ;
NAND2   gate10405  (.A(II23286), .B(II23287), .Z(WX7583) ) ;
AND2    gate10406  (.A(WX7583), .B(WX7470), .Z(WX7584) ) ;
AND2    gate10407  (.A(WX7061), .B(WX7586), .Z(WX7585) ) ;
NAND2   gate10408  (.A(II23299), .B(II23300), .Z(WX7590) ) ;
AND2    gate10409  (.A(WX7590), .B(WX7470), .Z(WX7591) ) ;
AND2    gate10410  (.A(WX7062), .B(WX7593), .Z(WX7592) ) ;
NAND2   gate10411  (.A(II23312), .B(II23313), .Z(WX7597) ) ;
AND2    gate10412  (.A(WX7597), .B(WX7470), .Z(WX7598) ) ;
AND2    gate10413  (.A(WX7063), .B(WX7600), .Z(WX7599) ) ;
NAND2   gate10414  (.A(II23325), .B(II23326), .Z(WX7604) ) ;
AND2    gate10415  (.A(WX7604), .B(WX7470), .Z(WX7605) ) ;
AND2    gate10416  (.A(WX7064), .B(WX7607), .Z(WX7606) ) ;
NAND2   gate10417  (.A(II23338), .B(II23339), .Z(WX7611) ) ;
AND2    gate10418  (.A(WX7611), .B(WX7470), .Z(WX7612) ) ;
AND2    gate10419  (.A(WX7065), .B(WX7614), .Z(WX7613) ) ;
NAND2   gate10420  (.A(II23351), .B(II23352), .Z(WX7618) ) ;
AND2    gate10421  (.A(WX7618), .B(WX7470), .Z(WX7619) ) ;
AND2    gate10422  (.A(WX7066), .B(WX7621), .Z(WX7620) ) ;
NAND2   gate10423  (.A(II23364), .B(II23365), .Z(WX7625) ) ;
AND2    gate10424  (.A(WX7625), .B(WX7470), .Z(WX7626) ) ;
AND2    gate10425  (.A(WX7067), .B(WX7628), .Z(WX7627) ) ;
NAND2   gate10426  (.A(II23377), .B(II23378), .Z(WX7632) ) ;
AND2    gate10427  (.A(WX7632), .B(WX7470), .Z(WX7633) ) ;
AND2    gate10428  (.A(WX7068), .B(WX7635), .Z(WX7634) ) ;
NAND2   gate10429  (.A(II23390), .B(II23391), .Z(WX7639) ) ;
AND2    gate10430  (.A(WX7639), .B(WX7470), .Z(WX7640) ) ;
AND2    gate10431  (.A(WX7069), .B(WX7642), .Z(WX7641) ) ;
NAND2   gate10432  (.A(II23403), .B(II23404), .Z(WX7646) ) ;
AND2    gate10433  (.A(WX7646), .B(WX7470), .Z(WX7647) ) ;
AND2    gate10434  (.A(WX7070), .B(WX7649), .Z(WX7648) ) ;
NAND2   gate10435  (.A(II23416), .B(II23417), .Z(WX7653) ) ;
AND2    gate10436  (.A(WX7653), .B(WX7470), .Z(WX7654) ) ;
AND2    gate10437  (.A(WX7071), .B(WX7656), .Z(WX7655) ) ;
NAND2   gate10438  (.A(II23429), .B(II23430), .Z(WX7660) ) ;
AND2    gate10439  (.A(WX7660), .B(WX7470), .Z(WX7661) ) ;
AND2    gate10440  (.A(WX7072), .B(WX7663), .Z(WX7662) ) ;
NAND2   gate10441  (.A(II23442), .B(II23443), .Z(WX7667) ) ;
AND2    gate10442  (.A(WX7667), .B(WX7470), .Z(WX7668) ) ;
AND2    gate10443  (.A(WX7073), .B(WX7670), .Z(WX7669) ) ;
NAND2   gate10444  (.A(II23455), .B(II23456), .Z(WX7674) ) ;
AND2    gate10445  (.A(WX7674), .B(WX7470), .Z(WX7675) ) ;
AND2    gate10446  (.A(WX7074), .B(WX7677), .Z(WX7676) ) ;
NAND2   gate10447  (.A(II23468), .B(II23469), .Z(WX7681) ) ;
AND2    gate10448  (.A(WX7681), .B(WX7470), .Z(WX7682) ) ;
AND2    gate10449  (.A(WX7075), .B(WX7684), .Z(WX7683) ) ;
NAND2   gate10450  (.A(II23481), .B(II23482), .Z(WX7688) ) ;
AND2    gate10451  (.A(WX7688), .B(WX7470), .Z(WX7689) ) ;
AND2    gate10452  (.A(WX7076), .B(WX7691), .Z(WX7690) ) ;
NAND2   gate10453  (.A(II23540), .B(II23541), .Z(WX7699) ) ;
NAND2   gate10454  (.A(II23736), .B(II23737), .Z(WX7727) ) ;
NAND2   gate10455  (.A(II23729), .B(II23730), .Z(WX7726) ) ;
NAND2   gate10456  (.A(II23722), .B(II23723), .Z(WX7725) ) ;
NAND2   gate10457  (.A(II23533), .B(II23534), .Z(WX7698) ) ;
NAND2   gate10458  (.A(II23715), .B(II23716), .Z(WX7724) ) ;
NAND2   gate10459  (.A(II23708), .B(II23709), .Z(WX7723) ) ;
NAND2   gate10460  (.A(II23701), .B(II23702), .Z(WX7722) ) ;
NAND2   gate10461  (.A(II23694), .B(II23695), .Z(WX7721) ) ;
NAND2   gate10462  (.A(II23687), .B(II23688), .Z(WX7720) ) ;
NAND2   gate10463  (.A(II23680), .B(II23681), .Z(WX7719) ) ;
NAND2   gate10464  (.A(II23518), .B(II23519), .Z(WX7697) ) ;
NAND2   gate10465  (.A(II23673), .B(II23674), .Z(WX7718) ) ;
NAND2   gate10466  (.A(II23666), .B(II23667), .Z(WX7717) ) ;
NAND2   gate10467  (.A(II23659), .B(II23660), .Z(WX7716) ) ;
NAND2   gate10468  (.A(II23652), .B(II23653), .Z(WX7715) ) ;
NAND2   gate10469  (.A(II23503), .B(II23504), .Z(WX7696) ) ;
NAND2   gate10470  (.A(II23645), .B(II23646), .Z(WX7714) ) ;
NAND2   gate10471  (.A(II23638), .B(II23639), .Z(WX7713) ) ;
NAND2   gate10472  (.A(II23631), .B(II23632), .Z(WX7712) ) ;
NAND2   gate10473  (.A(II23624), .B(II23625), .Z(WX7711) ) ;
NAND2   gate10474  (.A(II23617), .B(II23618), .Z(WX7710) ) ;
NAND2   gate10475  (.A(II23610), .B(II23611), .Z(WX7709) ) ;
NAND2   gate10476  (.A(II23603), .B(II23604), .Z(WX7708) ) ;
NAND2   gate10477  (.A(II23596), .B(II23597), .Z(WX7707) ) ;
NAND2   gate10478  (.A(II23589), .B(II23590), .Z(WX7706) ) ;
NAND2   gate10479  (.A(II23582), .B(II23583), .Z(WX7705) ) ;
NAND2   gate10480  (.A(II23575), .B(II23576), .Z(WX7704) ) ;
NAND2   gate10481  (.A(II23568), .B(II23569), .Z(WX7703) ) ;
NAND2   gate10482  (.A(II23561), .B(II23562), .Z(WX7702) ) ;
NAND2   gate10483  (.A(II23554), .B(II23555), .Z(WX7701) ) ;
NAND2   gate10484  (.A(II23547), .B(II23548), .Z(WX7700) ) ;
OR2     gate10485  (.A(WX7802), .B(WX7801), .Z(WX7804) ) ;
AND2    gate10486  (.A(WX7804), .B(WX8761), .Z(WX7793) ) ;
OR2     gate10487  (.A(WX7798), .B(WX7797), .Z(WX7800) ) ;
AND2    gate10488  (.A(WX7800), .B(WX7795), .Z(WX7794) ) ;
AND2    gate10489  (.A(CRC_OUT_3_31), .B(WX8762), .Z(WX7797) ) ;
AND2    gate10490  (.A(WX10063), .B(WX7799), .Z(WX7798) ) ;
AND2    gate10491  (.A(WX8243), .B(WX8762), .Z(WX7801) ) ;
AND2    gate10492  (.A(WX8770), .B(WX7803), .Z(WX7802) ) ;
OR2     gate10493  (.A(WX7816), .B(WX7815), .Z(WX7818) ) ;
AND2    gate10494  (.A(WX7818), .B(WX8761), .Z(WX7807) ) ;
OR2     gate10495  (.A(WX7812), .B(WX7811), .Z(WX7814) ) ;
AND2    gate10496  (.A(WX7814), .B(WX7809), .Z(WX7808) ) ;
AND2    gate10497  (.A(CRC_OUT_3_30), .B(WX8762), .Z(WX7811) ) ;
AND2    gate10498  (.A(WX10070), .B(WX7813), .Z(WX7812) ) ;
AND2    gate10499  (.A(WX8245), .B(WX8762), .Z(WX7815) ) ;
AND2    gate10500  (.A(WX8777), .B(WX7817), .Z(WX7816) ) ;
OR2     gate10501  (.A(WX7830), .B(WX7829), .Z(WX7832) ) ;
AND2    gate10502  (.A(WX7832), .B(WX8761), .Z(WX7821) ) ;
OR2     gate10503  (.A(WX7826), .B(WX7825), .Z(WX7828) ) ;
AND2    gate10504  (.A(WX7828), .B(WX7823), .Z(WX7822) ) ;
AND2    gate10505  (.A(CRC_OUT_3_29), .B(WX8762), .Z(WX7825) ) ;
AND2    gate10506  (.A(WX10077), .B(WX7827), .Z(WX7826) ) ;
AND2    gate10507  (.A(WX8247), .B(WX8762), .Z(WX7829) ) ;
AND2    gate10508  (.A(WX8784), .B(WX7831), .Z(WX7830) ) ;
OR2     gate10509  (.A(WX7844), .B(WX7843), .Z(WX7846) ) ;
AND2    gate10510  (.A(WX7846), .B(WX8761), .Z(WX7835) ) ;
OR2     gate10511  (.A(WX7840), .B(WX7839), .Z(WX7842) ) ;
AND2    gate10512  (.A(WX7842), .B(WX7837), .Z(WX7836) ) ;
AND2    gate10513  (.A(CRC_OUT_3_28), .B(WX8762), .Z(WX7839) ) ;
AND2    gate10514  (.A(WX10084), .B(WX7841), .Z(WX7840) ) ;
AND2    gate10515  (.A(WX8249), .B(WX8762), .Z(WX7843) ) ;
AND2    gate10516  (.A(WX8791), .B(WX7845), .Z(WX7844) ) ;
OR2     gate10517  (.A(WX7858), .B(WX7857), .Z(WX7860) ) ;
AND2    gate10518  (.A(WX7860), .B(WX8761), .Z(WX7849) ) ;
OR2     gate10519  (.A(WX7854), .B(WX7853), .Z(WX7856) ) ;
AND2    gate10520  (.A(WX7856), .B(WX7851), .Z(WX7850) ) ;
AND2    gate10521  (.A(CRC_OUT_3_27), .B(WX8762), .Z(WX7853) ) ;
AND2    gate10522  (.A(WX10091), .B(WX7855), .Z(WX7854) ) ;
AND2    gate10523  (.A(WX8251), .B(WX8762), .Z(WX7857) ) ;
AND2    gate10524  (.A(WX8798), .B(WX7859), .Z(WX7858) ) ;
OR2     gate10525  (.A(WX7872), .B(WX7871), .Z(WX7874) ) ;
AND2    gate10526  (.A(WX7874), .B(WX8761), .Z(WX7863) ) ;
OR2     gate10527  (.A(WX7868), .B(WX7867), .Z(WX7870) ) ;
AND2    gate10528  (.A(WX7870), .B(WX7865), .Z(WX7864) ) ;
AND2    gate10529  (.A(CRC_OUT_3_26), .B(WX8762), .Z(WX7867) ) ;
AND2    gate10530  (.A(WX10098), .B(WX7869), .Z(WX7868) ) ;
AND2    gate10531  (.A(WX8253), .B(WX8762), .Z(WX7871) ) ;
AND2    gate10532  (.A(WX8805), .B(WX7873), .Z(WX7872) ) ;
OR2     gate10533  (.A(WX7886), .B(WX7885), .Z(WX7888) ) ;
AND2    gate10534  (.A(WX7888), .B(WX8761), .Z(WX7877) ) ;
OR2     gate10535  (.A(WX7882), .B(WX7881), .Z(WX7884) ) ;
AND2    gate10536  (.A(WX7884), .B(WX7879), .Z(WX7878) ) ;
AND2    gate10537  (.A(CRC_OUT_3_25), .B(WX8762), .Z(WX7881) ) ;
AND2    gate10538  (.A(WX10105), .B(WX7883), .Z(WX7882) ) ;
AND2    gate10539  (.A(WX8255), .B(WX8762), .Z(WX7885) ) ;
AND2    gate10540  (.A(WX8812), .B(WX7887), .Z(WX7886) ) ;
OR2     gate10541  (.A(WX7900), .B(WX7899), .Z(WX7902) ) ;
AND2    gate10542  (.A(WX7902), .B(WX8761), .Z(WX7891) ) ;
OR2     gate10543  (.A(WX7896), .B(WX7895), .Z(WX7898) ) ;
AND2    gate10544  (.A(WX7898), .B(WX7893), .Z(WX7892) ) ;
AND2    gate10545  (.A(CRC_OUT_3_24), .B(WX8762), .Z(WX7895) ) ;
AND2    gate10546  (.A(WX10112), .B(WX7897), .Z(WX7896) ) ;
AND2    gate10547  (.A(WX8257), .B(WX8762), .Z(WX7899) ) ;
AND2    gate10548  (.A(WX8819), .B(WX7901), .Z(WX7900) ) ;
OR2     gate10549  (.A(WX7914), .B(WX7913), .Z(WX7916) ) ;
AND2    gate10550  (.A(WX7916), .B(WX8761), .Z(WX7905) ) ;
OR2     gate10551  (.A(WX7910), .B(WX7909), .Z(WX7912) ) ;
AND2    gate10552  (.A(WX7912), .B(WX7907), .Z(WX7906) ) ;
AND2    gate10553  (.A(CRC_OUT_3_23), .B(WX8762), .Z(WX7909) ) ;
AND2    gate10554  (.A(WX10119), .B(WX7911), .Z(WX7910) ) ;
AND2    gate10555  (.A(WX8259), .B(WX8762), .Z(WX7913) ) ;
AND2    gate10556  (.A(WX8826), .B(WX7915), .Z(WX7914) ) ;
OR2     gate10557  (.A(WX7928), .B(WX7927), .Z(WX7930) ) ;
AND2    gate10558  (.A(WX7930), .B(WX8761), .Z(WX7919) ) ;
OR2     gate10559  (.A(WX7924), .B(WX7923), .Z(WX7926) ) ;
AND2    gate10560  (.A(WX7926), .B(WX7921), .Z(WX7920) ) ;
AND2    gate10561  (.A(CRC_OUT_3_22), .B(WX8762), .Z(WX7923) ) ;
AND2    gate10562  (.A(WX10126), .B(WX7925), .Z(WX7924) ) ;
AND2    gate10563  (.A(WX8261), .B(WX8762), .Z(WX7927) ) ;
AND2    gate10564  (.A(WX8833), .B(WX7929), .Z(WX7928) ) ;
OR2     gate10565  (.A(WX7942), .B(WX7941), .Z(WX7944) ) ;
AND2    gate10566  (.A(WX7944), .B(WX8761), .Z(WX7933) ) ;
OR2     gate10567  (.A(WX7938), .B(WX7937), .Z(WX7940) ) ;
AND2    gate10568  (.A(WX7940), .B(WX7935), .Z(WX7934) ) ;
AND2    gate10569  (.A(CRC_OUT_3_21), .B(WX8762), .Z(WX7937) ) ;
AND2    gate10570  (.A(WX10133), .B(WX7939), .Z(WX7938) ) ;
AND2    gate10571  (.A(WX8263), .B(WX8762), .Z(WX7941) ) ;
AND2    gate10572  (.A(WX8840), .B(WX7943), .Z(WX7942) ) ;
OR2     gate10573  (.A(WX7956), .B(WX7955), .Z(WX7958) ) ;
AND2    gate10574  (.A(WX7958), .B(WX8761), .Z(WX7947) ) ;
OR2     gate10575  (.A(WX7952), .B(WX7951), .Z(WX7954) ) ;
AND2    gate10576  (.A(WX7954), .B(WX7949), .Z(WX7948) ) ;
AND2    gate10577  (.A(CRC_OUT_3_20), .B(WX8762), .Z(WX7951) ) ;
AND2    gate10578  (.A(WX10140), .B(WX7953), .Z(WX7952) ) ;
AND2    gate10579  (.A(WX8265), .B(WX8762), .Z(WX7955) ) ;
AND2    gate10580  (.A(WX8847), .B(WX7957), .Z(WX7956) ) ;
OR2     gate10581  (.A(WX7970), .B(WX7969), .Z(WX7972) ) ;
AND2    gate10582  (.A(WX7972), .B(WX8761), .Z(WX7961) ) ;
OR2     gate10583  (.A(WX7966), .B(WX7965), .Z(WX7968) ) ;
AND2    gate10584  (.A(WX7968), .B(WX7963), .Z(WX7962) ) ;
AND2    gate10585  (.A(CRC_OUT_3_19), .B(WX8762), .Z(WX7965) ) ;
AND2    gate10586  (.A(WX10147), .B(WX7967), .Z(WX7966) ) ;
AND2    gate10587  (.A(WX8267), .B(WX8762), .Z(WX7969) ) ;
AND2    gate10588  (.A(WX8854), .B(WX7971), .Z(WX7970) ) ;
OR2     gate10589  (.A(WX7984), .B(WX7983), .Z(WX7986) ) ;
AND2    gate10590  (.A(WX7986), .B(WX8761), .Z(WX7975) ) ;
OR2     gate10591  (.A(WX7980), .B(WX7979), .Z(WX7982) ) ;
AND2    gate10592  (.A(WX7982), .B(WX7977), .Z(WX7976) ) ;
AND2    gate10593  (.A(CRC_OUT_3_18), .B(WX8762), .Z(WX7979) ) ;
AND2    gate10594  (.A(WX10154), .B(WX7981), .Z(WX7980) ) ;
AND2    gate10595  (.A(WX8269), .B(WX8762), .Z(WX7983) ) ;
AND2    gate10596  (.A(WX8861), .B(WX7985), .Z(WX7984) ) ;
OR2     gate10597  (.A(WX7998), .B(WX7997), .Z(WX8000) ) ;
AND2    gate10598  (.A(WX8000), .B(WX8761), .Z(WX7989) ) ;
OR2     gate10599  (.A(WX7994), .B(WX7993), .Z(WX7996) ) ;
AND2    gate10600  (.A(WX7996), .B(WX7991), .Z(WX7990) ) ;
AND2    gate10601  (.A(CRC_OUT_3_17), .B(WX8762), .Z(WX7993) ) ;
AND2    gate10602  (.A(WX10161), .B(WX7995), .Z(WX7994) ) ;
AND2    gate10603  (.A(WX8271), .B(WX8762), .Z(WX7997) ) ;
AND2    gate10604  (.A(WX8868), .B(WX7999), .Z(WX7998) ) ;
OR2     gate10605  (.A(WX8012), .B(WX8011), .Z(WX8014) ) ;
AND2    gate10606  (.A(WX8014), .B(WX8761), .Z(WX8003) ) ;
OR2     gate10607  (.A(WX8008), .B(WX8007), .Z(WX8010) ) ;
AND2    gate10608  (.A(WX8010), .B(WX8005), .Z(WX8004) ) ;
AND2    gate10609  (.A(CRC_OUT_3_16), .B(WX8762), .Z(WX8007) ) ;
AND2    gate10610  (.A(WX10168), .B(WX8009), .Z(WX8008) ) ;
AND2    gate10611  (.A(WX8273), .B(WX8762), .Z(WX8011) ) ;
AND2    gate10612  (.A(WX8875), .B(WX8013), .Z(WX8012) ) ;
OR2     gate10613  (.A(WX8026), .B(WX8025), .Z(WX8028) ) ;
AND2    gate10614  (.A(WX8028), .B(WX8761), .Z(WX8017) ) ;
OR2     gate10615  (.A(WX8022), .B(WX8021), .Z(WX8024) ) ;
AND2    gate10616  (.A(WX8024), .B(WX8019), .Z(WX8018) ) ;
AND2    gate10617  (.A(CRC_OUT_3_15), .B(WX8762), .Z(WX8021) ) ;
AND2    gate10618  (.A(WX10175), .B(WX8023), .Z(WX8022) ) ;
AND2    gate10619  (.A(WX8275), .B(WX8762), .Z(WX8025) ) ;
AND2    gate10620  (.A(WX8882), .B(WX8027), .Z(WX8026) ) ;
OR2     gate10621  (.A(WX8040), .B(WX8039), .Z(WX8042) ) ;
AND2    gate10622  (.A(WX8042), .B(WX8761), .Z(WX8031) ) ;
OR2     gate10623  (.A(WX8036), .B(WX8035), .Z(WX8038) ) ;
AND2    gate10624  (.A(WX8038), .B(WX8033), .Z(WX8032) ) ;
AND2    gate10625  (.A(CRC_OUT_3_14), .B(WX8762), .Z(WX8035) ) ;
AND2    gate10626  (.A(WX10182), .B(WX8037), .Z(WX8036) ) ;
AND2    gate10627  (.A(WX8277), .B(WX8762), .Z(WX8039) ) ;
AND2    gate10628  (.A(WX8889), .B(WX8041), .Z(WX8040) ) ;
OR2     gate10629  (.A(WX8054), .B(WX8053), .Z(WX8056) ) ;
AND2    gate10630  (.A(WX8056), .B(WX8761), .Z(WX8045) ) ;
OR2     gate10631  (.A(WX8050), .B(WX8049), .Z(WX8052) ) ;
AND2    gate10632  (.A(WX8052), .B(WX8047), .Z(WX8046) ) ;
AND2    gate10633  (.A(CRC_OUT_3_13), .B(WX8762), .Z(WX8049) ) ;
AND2    gate10634  (.A(WX10189), .B(WX8051), .Z(WX8050) ) ;
AND2    gate10635  (.A(WX8279), .B(WX8762), .Z(WX8053) ) ;
AND2    gate10636  (.A(WX8896), .B(WX8055), .Z(WX8054) ) ;
OR2     gate10637  (.A(WX8068), .B(WX8067), .Z(WX8070) ) ;
AND2    gate10638  (.A(WX8070), .B(WX8761), .Z(WX8059) ) ;
OR2     gate10639  (.A(WX8064), .B(WX8063), .Z(WX8066) ) ;
AND2    gate10640  (.A(WX8066), .B(WX8061), .Z(WX8060) ) ;
AND2    gate10641  (.A(CRC_OUT_3_12), .B(WX8762), .Z(WX8063) ) ;
AND2    gate10642  (.A(WX10196), .B(WX8065), .Z(WX8064) ) ;
AND2    gate10643  (.A(WX8281), .B(WX8762), .Z(WX8067) ) ;
AND2    gate10644  (.A(WX8903), .B(WX8069), .Z(WX8068) ) ;
OR2     gate10645  (.A(WX8082), .B(WX8081), .Z(WX8084) ) ;
AND2    gate10646  (.A(WX8084), .B(WX8761), .Z(WX8073) ) ;
OR2     gate10647  (.A(WX8078), .B(WX8077), .Z(WX8080) ) ;
AND2    gate10648  (.A(WX8080), .B(WX8075), .Z(WX8074) ) ;
AND2    gate10649  (.A(CRC_OUT_3_11), .B(WX8762), .Z(WX8077) ) ;
AND2    gate10650  (.A(WX10203), .B(WX8079), .Z(WX8078) ) ;
AND2    gate10651  (.A(WX8283), .B(WX8762), .Z(WX8081) ) ;
AND2    gate10652  (.A(WX8910), .B(WX8083), .Z(WX8082) ) ;
OR2     gate10653  (.A(WX8096), .B(WX8095), .Z(WX8098) ) ;
AND2    gate10654  (.A(WX8098), .B(WX8761), .Z(WX8087) ) ;
OR2     gate10655  (.A(WX8092), .B(WX8091), .Z(WX8094) ) ;
AND2    gate10656  (.A(WX8094), .B(WX8089), .Z(WX8088) ) ;
AND2    gate10657  (.A(CRC_OUT_3_10), .B(WX8762), .Z(WX8091) ) ;
AND2    gate10658  (.A(WX10210), .B(WX8093), .Z(WX8092) ) ;
AND2    gate10659  (.A(WX8285), .B(WX8762), .Z(WX8095) ) ;
AND2    gate10660  (.A(WX8917), .B(WX8097), .Z(WX8096) ) ;
OR2     gate10661  (.A(WX8110), .B(WX8109), .Z(WX8112) ) ;
AND2    gate10662  (.A(WX8112), .B(WX8761), .Z(WX8101) ) ;
OR2     gate10663  (.A(WX8106), .B(WX8105), .Z(WX8108) ) ;
AND2    gate10664  (.A(WX8108), .B(WX8103), .Z(WX8102) ) ;
AND2    gate10665  (.A(CRC_OUT_3_9), .B(WX8762), .Z(WX8105) ) ;
AND2    gate10666  (.A(WX10217), .B(WX8107), .Z(WX8106) ) ;
AND2    gate10667  (.A(WX8287), .B(WX8762), .Z(WX8109) ) ;
AND2    gate10668  (.A(WX8924), .B(WX8111), .Z(WX8110) ) ;
OR2     gate10669  (.A(WX8124), .B(WX8123), .Z(WX8126) ) ;
AND2    gate10670  (.A(WX8126), .B(WX8761), .Z(WX8115) ) ;
OR2     gate10671  (.A(WX8120), .B(WX8119), .Z(WX8122) ) ;
AND2    gate10672  (.A(WX8122), .B(WX8117), .Z(WX8116) ) ;
AND2    gate10673  (.A(CRC_OUT_3_8), .B(WX8762), .Z(WX8119) ) ;
AND2    gate10674  (.A(WX10224), .B(WX8121), .Z(WX8120) ) ;
AND2    gate10675  (.A(WX8289), .B(WX8762), .Z(WX8123) ) ;
AND2    gate10676  (.A(WX8931), .B(WX8125), .Z(WX8124) ) ;
OR2     gate10677  (.A(WX8138), .B(WX8137), .Z(WX8140) ) ;
AND2    gate10678  (.A(WX8140), .B(WX8761), .Z(WX8129) ) ;
OR2     gate10679  (.A(WX8134), .B(WX8133), .Z(WX8136) ) ;
AND2    gate10680  (.A(WX8136), .B(WX8131), .Z(WX8130) ) ;
AND2    gate10681  (.A(CRC_OUT_3_7), .B(WX8762), .Z(WX8133) ) ;
AND2    gate10682  (.A(WX10231), .B(WX8135), .Z(WX8134) ) ;
AND2    gate10683  (.A(WX8291), .B(WX8762), .Z(WX8137) ) ;
AND2    gate10684  (.A(WX8938), .B(WX8139), .Z(WX8138) ) ;
OR2     gate10685  (.A(WX8152), .B(WX8151), .Z(WX8154) ) ;
AND2    gate10686  (.A(WX8154), .B(WX8761), .Z(WX8143) ) ;
OR2     gate10687  (.A(WX8148), .B(WX8147), .Z(WX8150) ) ;
AND2    gate10688  (.A(WX8150), .B(WX8145), .Z(WX8144) ) ;
AND2    gate10689  (.A(CRC_OUT_3_6), .B(WX8762), .Z(WX8147) ) ;
AND2    gate10690  (.A(WX10238), .B(WX8149), .Z(WX8148) ) ;
AND2    gate10691  (.A(WX8293), .B(WX8762), .Z(WX8151) ) ;
AND2    gate10692  (.A(WX8945), .B(WX8153), .Z(WX8152) ) ;
OR2     gate10693  (.A(WX8166), .B(WX8165), .Z(WX8168) ) ;
AND2    gate10694  (.A(WX8168), .B(WX8761), .Z(WX8157) ) ;
OR2     gate10695  (.A(WX8162), .B(WX8161), .Z(WX8164) ) ;
AND2    gate10696  (.A(WX8164), .B(WX8159), .Z(WX8158) ) ;
AND2    gate10697  (.A(CRC_OUT_3_5), .B(WX8762), .Z(WX8161) ) ;
AND2    gate10698  (.A(WX10245), .B(WX8163), .Z(WX8162) ) ;
AND2    gate10699  (.A(WX8295), .B(WX8762), .Z(WX8165) ) ;
AND2    gate10700  (.A(WX8952), .B(WX8167), .Z(WX8166) ) ;
OR2     gate10701  (.A(WX8180), .B(WX8179), .Z(WX8182) ) ;
AND2    gate10702  (.A(WX8182), .B(WX8761), .Z(WX8171) ) ;
OR2     gate10703  (.A(WX8176), .B(WX8175), .Z(WX8178) ) ;
AND2    gate10704  (.A(WX8178), .B(WX8173), .Z(WX8172) ) ;
AND2    gate10705  (.A(CRC_OUT_3_4), .B(WX8762), .Z(WX8175) ) ;
AND2    gate10706  (.A(WX10252), .B(WX8177), .Z(WX8176) ) ;
AND2    gate10707  (.A(WX8297), .B(WX8762), .Z(WX8179) ) ;
AND2    gate10708  (.A(WX8959), .B(WX8181), .Z(WX8180) ) ;
OR2     gate10709  (.A(WX8194), .B(WX8193), .Z(WX8196) ) ;
AND2    gate10710  (.A(WX8196), .B(WX8761), .Z(WX8185) ) ;
OR2     gate10711  (.A(WX8190), .B(WX8189), .Z(WX8192) ) ;
AND2    gate10712  (.A(WX8192), .B(WX8187), .Z(WX8186) ) ;
AND2    gate10713  (.A(CRC_OUT_3_3), .B(WX8762), .Z(WX8189) ) ;
AND2    gate10714  (.A(WX10259), .B(WX8191), .Z(WX8190) ) ;
AND2    gate10715  (.A(WX8299), .B(WX8762), .Z(WX8193) ) ;
AND2    gate10716  (.A(WX8966), .B(WX8195), .Z(WX8194) ) ;
OR2     gate10717  (.A(WX8208), .B(WX8207), .Z(WX8210) ) ;
AND2    gate10718  (.A(WX8210), .B(WX8761), .Z(WX8199) ) ;
OR2     gate10719  (.A(WX8204), .B(WX8203), .Z(WX8206) ) ;
AND2    gate10720  (.A(WX8206), .B(WX8201), .Z(WX8200) ) ;
AND2    gate10721  (.A(CRC_OUT_3_2), .B(WX8762), .Z(WX8203) ) ;
AND2    gate10722  (.A(WX10266), .B(WX8205), .Z(WX8204) ) ;
AND2    gate10723  (.A(WX8301), .B(WX8762), .Z(WX8207) ) ;
AND2    gate10724  (.A(WX8973), .B(WX8209), .Z(WX8208) ) ;
OR2     gate10725  (.A(WX8222), .B(WX8221), .Z(WX8224) ) ;
AND2    gate10726  (.A(WX8224), .B(WX8761), .Z(WX8213) ) ;
OR2     gate10727  (.A(WX8218), .B(WX8217), .Z(WX8220) ) ;
AND2    gate10728  (.A(WX8220), .B(WX8215), .Z(WX8214) ) ;
AND2    gate10729  (.A(CRC_OUT_3_1), .B(WX8762), .Z(WX8217) ) ;
AND2    gate10730  (.A(WX10273), .B(WX8219), .Z(WX8218) ) ;
AND2    gate10731  (.A(WX8303), .B(WX8762), .Z(WX8221) ) ;
AND2    gate10732  (.A(WX8980), .B(WX8223), .Z(WX8222) ) ;
OR2     gate10733  (.A(WX8236), .B(WX8235), .Z(WX8238) ) ;
AND2    gate10734  (.A(WX8238), .B(WX8761), .Z(WX8227) ) ;
OR2     gate10735  (.A(WX8232), .B(WX8231), .Z(WX8234) ) ;
AND2    gate10736  (.A(WX8234), .B(WX8229), .Z(WX8228) ) ;
AND2    gate10737  (.A(CRC_OUT_3_0), .B(WX8762), .Z(WX8231) ) ;
AND2    gate10738  (.A(WX10280), .B(WX8233), .Z(WX8232) ) ;
AND2    gate10739  (.A(WX8305), .B(WX8762), .Z(WX8235) ) ;
AND2    gate10740  (.A(WX8987), .B(WX8237), .Z(WX8236) ) ;
NAND2   gate10741  (.A(II27083), .B(II27084), .Z(WX8764) ) ;
AND2    gate10742  (.A(WX8764), .B(WX8763), .Z(WX8765) ) ;
AND2    gate10743  (.A(WX8338), .B(WX8767), .Z(WX8766) ) ;
NAND2   gate10744  (.A(II27096), .B(II27097), .Z(WX8771) ) ;
AND2    gate10745  (.A(WX8771), .B(WX8763), .Z(WX8772) ) ;
AND2    gate10746  (.A(WX8339), .B(WX8774), .Z(WX8773) ) ;
NAND2   gate10747  (.A(II27109), .B(II27110), .Z(WX8778) ) ;
AND2    gate10748  (.A(WX8778), .B(WX8763), .Z(WX8779) ) ;
AND2    gate10749  (.A(WX8340), .B(WX8781), .Z(WX8780) ) ;
NAND2   gate10750  (.A(II27122), .B(II27123), .Z(WX8785) ) ;
AND2    gate10751  (.A(WX8785), .B(WX8763), .Z(WX8786) ) ;
AND2    gate10752  (.A(WX8341), .B(WX8788), .Z(WX8787) ) ;
NAND2   gate10753  (.A(II27135), .B(II27136), .Z(WX8792) ) ;
AND2    gate10754  (.A(WX8792), .B(WX8763), .Z(WX8793) ) ;
AND2    gate10755  (.A(WX8342), .B(WX8795), .Z(WX8794) ) ;
NAND2   gate10756  (.A(II27148), .B(II27149), .Z(WX8799) ) ;
AND2    gate10757  (.A(WX8799), .B(WX8763), .Z(WX8800) ) ;
AND2    gate10758  (.A(WX8343), .B(WX8802), .Z(WX8801) ) ;
NAND2   gate10759  (.A(II27161), .B(II27162), .Z(WX8806) ) ;
AND2    gate10760  (.A(WX8806), .B(WX8763), .Z(WX8807) ) ;
AND2    gate10761  (.A(WX8344), .B(WX8809), .Z(WX8808) ) ;
NAND2   gate10762  (.A(II27174), .B(II27175), .Z(WX8813) ) ;
AND2    gate10763  (.A(WX8813), .B(WX8763), .Z(WX8814) ) ;
AND2    gate10764  (.A(WX8345), .B(WX8816), .Z(WX8815) ) ;
NAND2   gate10765  (.A(II27187), .B(II27188), .Z(WX8820) ) ;
AND2    gate10766  (.A(WX8820), .B(WX8763), .Z(WX8821) ) ;
AND2    gate10767  (.A(WX8346), .B(WX8823), .Z(WX8822) ) ;
NAND2   gate10768  (.A(II27200), .B(II27201), .Z(WX8827) ) ;
AND2    gate10769  (.A(WX8827), .B(WX8763), .Z(WX8828) ) ;
AND2    gate10770  (.A(WX8347), .B(WX8830), .Z(WX8829) ) ;
NAND2   gate10771  (.A(II27213), .B(II27214), .Z(WX8834) ) ;
AND2    gate10772  (.A(WX8834), .B(WX8763), .Z(WX8835) ) ;
AND2    gate10773  (.A(WX8348), .B(WX8837), .Z(WX8836) ) ;
NAND2   gate10774  (.A(II27226), .B(II27227), .Z(WX8841) ) ;
AND2    gate10775  (.A(WX8841), .B(WX8763), .Z(WX8842) ) ;
AND2    gate10776  (.A(WX8349), .B(WX8844), .Z(WX8843) ) ;
NAND2   gate10777  (.A(II27239), .B(II27240), .Z(WX8848) ) ;
AND2    gate10778  (.A(WX8848), .B(WX8763), .Z(WX8849) ) ;
AND2    gate10779  (.A(WX8350), .B(WX8851), .Z(WX8850) ) ;
NAND2   gate10780  (.A(II27252), .B(II27253), .Z(WX8855) ) ;
AND2    gate10781  (.A(WX8855), .B(WX8763), .Z(WX8856) ) ;
AND2    gate10782  (.A(WX8351), .B(WX8858), .Z(WX8857) ) ;
NAND2   gate10783  (.A(II27265), .B(II27266), .Z(WX8862) ) ;
AND2    gate10784  (.A(WX8862), .B(WX8763), .Z(WX8863) ) ;
AND2    gate10785  (.A(WX8352), .B(WX8865), .Z(WX8864) ) ;
NAND2   gate10786  (.A(II27278), .B(II27279), .Z(WX8869) ) ;
AND2    gate10787  (.A(WX8869), .B(WX8763), .Z(WX8870) ) ;
AND2    gate10788  (.A(WX8353), .B(WX8872), .Z(WX8871) ) ;
NAND2   gate10789  (.A(II27291), .B(II27292), .Z(WX8876) ) ;
AND2    gate10790  (.A(WX8876), .B(WX8763), .Z(WX8877) ) ;
AND2    gate10791  (.A(WX8354), .B(WX8879), .Z(WX8878) ) ;
NAND2   gate10792  (.A(II27304), .B(II27305), .Z(WX8883) ) ;
AND2    gate10793  (.A(WX8883), .B(WX8763), .Z(WX8884) ) ;
AND2    gate10794  (.A(WX8355), .B(WX8886), .Z(WX8885) ) ;
NAND2   gate10795  (.A(II27317), .B(II27318), .Z(WX8890) ) ;
AND2    gate10796  (.A(WX8890), .B(WX8763), .Z(WX8891) ) ;
AND2    gate10797  (.A(WX8356), .B(WX8893), .Z(WX8892) ) ;
NAND2   gate10798  (.A(II27330), .B(II27331), .Z(WX8897) ) ;
AND2    gate10799  (.A(WX8897), .B(WX8763), .Z(WX8898) ) ;
AND2    gate10800  (.A(WX8357), .B(WX8900), .Z(WX8899) ) ;
NAND2   gate10801  (.A(II27343), .B(II27344), .Z(WX8904) ) ;
AND2    gate10802  (.A(WX8904), .B(WX8763), .Z(WX8905) ) ;
AND2    gate10803  (.A(WX8358), .B(WX8907), .Z(WX8906) ) ;
NAND2   gate10804  (.A(II27356), .B(II27357), .Z(WX8911) ) ;
AND2    gate10805  (.A(WX8911), .B(WX8763), .Z(WX8912) ) ;
AND2    gate10806  (.A(WX8359), .B(WX8914), .Z(WX8913) ) ;
NAND2   gate10807  (.A(II27369), .B(II27370), .Z(WX8918) ) ;
AND2    gate10808  (.A(WX8918), .B(WX8763), .Z(WX8919) ) ;
AND2    gate10809  (.A(WX8360), .B(WX8921), .Z(WX8920) ) ;
NAND2   gate10810  (.A(II27382), .B(II27383), .Z(WX8925) ) ;
AND2    gate10811  (.A(WX8925), .B(WX8763), .Z(WX8926) ) ;
AND2    gate10812  (.A(WX8361), .B(WX8928), .Z(WX8927) ) ;
NAND2   gate10813  (.A(II27395), .B(II27396), .Z(WX8932) ) ;
AND2    gate10814  (.A(WX8932), .B(WX8763), .Z(WX8933) ) ;
AND2    gate10815  (.A(WX8362), .B(WX8935), .Z(WX8934) ) ;
NAND2   gate10816  (.A(II27408), .B(II27409), .Z(WX8939) ) ;
AND2    gate10817  (.A(WX8939), .B(WX8763), .Z(WX8940) ) ;
AND2    gate10818  (.A(WX8363), .B(WX8942), .Z(WX8941) ) ;
NAND2   gate10819  (.A(II27421), .B(II27422), .Z(WX8946) ) ;
AND2    gate10820  (.A(WX8946), .B(WX8763), .Z(WX8947) ) ;
AND2    gate10821  (.A(WX8364), .B(WX8949), .Z(WX8948) ) ;
NAND2   gate10822  (.A(II27434), .B(II27435), .Z(WX8953) ) ;
AND2    gate10823  (.A(WX8953), .B(WX8763), .Z(WX8954) ) ;
AND2    gate10824  (.A(WX8365), .B(WX8956), .Z(WX8955) ) ;
NAND2   gate10825  (.A(II27447), .B(II27448), .Z(WX8960) ) ;
AND2    gate10826  (.A(WX8960), .B(WX8763), .Z(WX8961) ) ;
AND2    gate10827  (.A(WX8366), .B(WX8963), .Z(WX8962) ) ;
NAND2   gate10828  (.A(II27460), .B(II27461), .Z(WX8967) ) ;
AND2    gate10829  (.A(WX8967), .B(WX8763), .Z(WX8968) ) ;
AND2    gate10830  (.A(WX8367), .B(WX8970), .Z(WX8969) ) ;
NAND2   gate10831  (.A(II27473), .B(II27474), .Z(WX8974) ) ;
AND2    gate10832  (.A(WX8974), .B(WX8763), .Z(WX8975) ) ;
AND2    gate10833  (.A(WX8368), .B(WX8977), .Z(WX8976) ) ;
NAND2   gate10834  (.A(II27486), .B(II27487), .Z(WX8981) ) ;
AND2    gate10835  (.A(WX8981), .B(WX8763), .Z(WX8982) ) ;
AND2    gate10836  (.A(WX8369), .B(WX8984), .Z(WX8983) ) ;
NAND2   gate10837  (.A(II27545), .B(II27546), .Z(WX8992) ) ;
NAND2   gate10838  (.A(II27741), .B(II27742), .Z(WX9020) ) ;
NAND2   gate10839  (.A(II27734), .B(II27735), .Z(WX9019) ) ;
NAND2   gate10840  (.A(II27727), .B(II27728), .Z(WX9018) ) ;
NAND2   gate10841  (.A(II27538), .B(II27539), .Z(WX8991) ) ;
NAND2   gate10842  (.A(II27720), .B(II27721), .Z(WX9017) ) ;
NAND2   gate10843  (.A(II27713), .B(II27714), .Z(WX9016) ) ;
NAND2   gate10844  (.A(II27706), .B(II27707), .Z(WX9015) ) ;
NAND2   gate10845  (.A(II27699), .B(II27700), .Z(WX9014) ) ;
NAND2   gate10846  (.A(II27692), .B(II27693), .Z(WX9013) ) ;
NAND2   gate10847  (.A(II27685), .B(II27686), .Z(WX9012) ) ;
NAND2   gate10848  (.A(II27523), .B(II27524), .Z(WX8990) ) ;
NAND2   gate10849  (.A(II27678), .B(II27679), .Z(WX9011) ) ;
NAND2   gate10850  (.A(II27671), .B(II27672), .Z(WX9010) ) ;
NAND2   gate10851  (.A(II27664), .B(II27665), .Z(WX9009) ) ;
NAND2   gate10852  (.A(II27657), .B(II27658), .Z(WX9008) ) ;
NAND2   gate10853  (.A(II27508), .B(II27509), .Z(WX8989) ) ;
NAND2   gate10854  (.A(II27650), .B(II27651), .Z(WX9007) ) ;
NAND2   gate10855  (.A(II27643), .B(II27644), .Z(WX9006) ) ;
NAND2   gate10856  (.A(II27636), .B(II27637), .Z(WX9005) ) ;
NAND2   gate10857  (.A(II27629), .B(II27630), .Z(WX9004) ) ;
NAND2   gate10858  (.A(II27622), .B(II27623), .Z(WX9003) ) ;
NAND2   gate10859  (.A(II27615), .B(II27616), .Z(WX9002) ) ;
NAND2   gate10860  (.A(II27608), .B(II27609), .Z(WX9001) ) ;
NAND2   gate10861  (.A(II27601), .B(II27602), .Z(WX9000) ) ;
NAND2   gate10862  (.A(II27594), .B(II27595), .Z(WX8999) ) ;
NAND2   gate10863  (.A(II27587), .B(II27588), .Z(WX8998) ) ;
NAND2   gate10864  (.A(II27580), .B(II27581), .Z(WX8997) ) ;
NAND2   gate10865  (.A(II27573), .B(II27574), .Z(WX8996) ) ;
NAND2   gate10866  (.A(II27566), .B(II27567), .Z(WX8995) ) ;
NAND2   gate10867  (.A(II27559), .B(II27560), .Z(WX8994) ) ;
NAND2   gate10868  (.A(II27552), .B(II27553), .Z(WX8993) ) ;
OR2     gate10869  (.A(WX9095), .B(WX9094), .Z(WX9097) ) ;
AND2    gate10870  (.A(WX9097), .B(WX10054), .Z(WX9086) ) ;
OR2     gate10871  (.A(WX9091), .B(WX9090), .Z(WX9093) ) ;
AND2    gate10872  (.A(WX9093), .B(WX9088), .Z(WX9087) ) ;
AND2    gate10873  (.A(CRC_OUT_2_31), .B(WX10055), .Z(WX9090) ) ;
AND2    gate10874  (.A(WX11356), .B(WX9092), .Z(WX9091) ) ;
AND2    gate10875  (.A(WX9536), .B(WX10055), .Z(WX9094) ) ;
AND2    gate10876  (.A(WX10063), .B(WX9096), .Z(WX9095) ) ;
OR2     gate10877  (.A(WX9109), .B(WX9108), .Z(WX9111) ) ;
AND2    gate10878  (.A(WX9111), .B(WX10054), .Z(WX9100) ) ;
OR2     gate10879  (.A(WX9105), .B(WX9104), .Z(WX9107) ) ;
AND2    gate10880  (.A(WX9107), .B(WX9102), .Z(WX9101) ) ;
AND2    gate10881  (.A(CRC_OUT_2_30), .B(WX10055), .Z(WX9104) ) ;
AND2    gate10882  (.A(WX11363), .B(WX9106), .Z(WX9105) ) ;
AND2    gate10883  (.A(WX9538), .B(WX10055), .Z(WX9108) ) ;
AND2    gate10884  (.A(WX10070), .B(WX9110), .Z(WX9109) ) ;
OR2     gate10885  (.A(WX9123), .B(WX9122), .Z(WX9125) ) ;
AND2    gate10886  (.A(WX9125), .B(WX10054), .Z(WX9114) ) ;
OR2     gate10887  (.A(WX9119), .B(WX9118), .Z(WX9121) ) ;
AND2    gate10888  (.A(WX9121), .B(WX9116), .Z(WX9115) ) ;
AND2    gate10889  (.A(CRC_OUT_2_29), .B(WX10055), .Z(WX9118) ) ;
AND2    gate10890  (.A(WX11370), .B(WX9120), .Z(WX9119) ) ;
AND2    gate10891  (.A(WX9540), .B(WX10055), .Z(WX9122) ) ;
AND2    gate10892  (.A(WX10077), .B(WX9124), .Z(WX9123) ) ;
OR2     gate10893  (.A(WX9137), .B(WX9136), .Z(WX9139) ) ;
AND2    gate10894  (.A(WX9139), .B(WX10054), .Z(WX9128) ) ;
OR2     gate10895  (.A(WX9133), .B(WX9132), .Z(WX9135) ) ;
AND2    gate10896  (.A(WX9135), .B(WX9130), .Z(WX9129) ) ;
AND2    gate10897  (.A(CRC_OUT_2_28), .B(WX10055), .Z(WX9132) ) ;
AND2    gate10898  (.A(WX11377), .B(WX9134), .Z(WX9133) ) ;
AND2    gate10899  (.A(WX9542), .B(WX10055), .Z(WX9136) ) ;
AND2    gate10900  (.A(WX10084), .B(WX9138), .Z(WX9137) ) ;
OR2     gate10901  (.A(WX9151), .B(WX9150), .Z(WX9153) ) ;
AND2    gate10902  (.A(WX9153), .B(WX10054), .Z(WX9142) ) ;
OR2     gate10903  (.A(WX9147), .B(WX9146), .Z(WX9149) ) ;
AND2    gate10904  (.A(WX9149), .B(WX9144), .Z(WX9143) ) ;
AND2    gate10905  (.A(CRC_OUT_2_27), .B(WX10055), .Z(WX9146) ) ;
AND2    gate10906  (.A(WX11384), .B(WX9148), .Z(WX9147) ) ;
AND2    gate10907  (.A(WX9544), .B(WX10055), .Z(WX9150) ) ;
AND2    gate10908  (.A(WX10091), .B(WX9152), .Z(WX9151) ) ;
OR2     gate10909  (.A(WX9165), .B(WX9164), .Z(WX9167) ) ;
AND2    gate10910  (.A(WX9167), .B(WX10054), .Z(WX9156) ) ;
OR2     gate10911  (.A(WX9161), .B(WX9160), .Z(WX9163) ) ;
AND2    gate10912  (.A(WX9163), .B(WX9158), .Z(WX9157) ) ;
AND2    gate10913  (.A(CRC_OUT_2_26), .B(WX10055), .Z(WX9160) ) ;
AND2    gate10914  (.A(WX11391), .B(WX9162), .Z(WX9161) ) ;
AND2    gate10915  (.A(WX9546), .B(WX10055), .Z(WX9164) ) ;
AND2    gate10916  (.A(WX10098), .B(WX9166), .Z(WX9165) ) ;
OR2     gate10917  (.A(WX9179), .B(WX9178), .Z(WX9181) ) ;
AND2    gate10918  (.A(WX9181), .B(WX10054), .Z(WX9170) ) ;
OR2     gate10919  (.A(WX9175), .B(WX9174), .Z(WX9177) ) ;
AND2    gate10920  (.A(WX9177), .B(WX9172), .Z(WX9171) ) ;
AND2    gate10921  (.A(CRC_OUT_2_25), .B(WX10055), .Z(WX9174) ) ;
AND2    gate10922  (.A(WX11398), .B(WX9176), .Z(WX9175) ) ;
AND2    gate10923  (.A(WX9548), .B(WX10055), .Z(WX9178) ) ;
AND2    gate10924  (.A(WX10105), .B(WX9180), .Z(WX9179) ) ;
OR2     gate10925  (.A(WX9193), .B(WX9192), .Z(WX9195) ) ;
AND2    gate10926  (.A(WX9195), .B(WX10054), .Z(WX9184) ) ;
OR2     gate10927  (.A(WX9189), .B(WX9188), .Z(WX9191) ) ;
AND2    gate10928  (.A(WX9191), .B(WX9186), .Z(WX9185) ) ;
AND2    gate10929  (.A(CRC_OUT_2_24), .B(WX10055), .Z(WX9188) ) ;
AND2    gate10930  (.A(WX11405), .B(WX9190), .Z(WX9189) ) ;
AND2    gate10931  (.A(WX9550), .B(WX10055), .Z(WX9192) ) ;
AND2    gate10932  (.A(WX10112), .B(WX9194), .Z(WX9193) ) ;
OR2     gate10933  (.A(WX9207), .B(WX9206), .Z(WX9209) ) ;
AND2    gate10934  (.A(WX9209), .B(WX10054), .Z(WX9198) ) ;
OR2     gate10935  (.A(WX9203), .B(WX9202), .Z(WX9205) ) ;
AND2    gate10936  (.A(WX9205), .B(WX9200), .Z(WX9199) ) ;
AND2    gate10937  (.A(CRC_OUT_2_23), .B(WX10055), .Z(WX9202) ) ;
AND2    gate10938  (.A(WX11412), .B(WX9204), .Z(WX9203) ) ;
AND2    gate10939  (.A(WX9552), .B(WX10055), .Z(WX9206) ) ;
AND2    gate10940  (.A(WX10119), .B(WX9208), .Z(WX9207) ) ;
OR2     gate10941  (.A(WX9221), .B(WX9220), .Z(WX9223) ) ;
AND2    gate10942  (.A(WX9223), .B(WX10054), .Z(WX9212) ) ;
OR2     gate10943  (.A(WX9217), .B(WX9216), .Z(WX9219) ) ;
AND2    gate10944  (.A(WX9219), .B(WX9214), .Z(WX9213) ) ;
AND2    gate10945  (.A(CRC_OUT_2_22), .B(WX10055), .Z(WX9216) ) ;
AND2    gate10946  (.A(WX11419), .B(WX9218), .Z(WX9217) ) ;
AND2    gate10947  (.A(WX9554), .B(WX10055), .Z(WX9220) ) ;
AND2    gate10948  (.A(WX10126), .B(WX9222), .Z(WX9221) ) ;
OR2     gate10949  (.A(WX9235), .B(WX9234), .Z(WX9237) ) ;
AND2    gate10950  (.A(WX9237), .B(WX10054), .Z(WX9226) ) ;
OR2     gate10951  (.A(WX9231), .B(WX9230), .Z(WX9233) ) ;
AND2    gate10952  (.A(WX9233), .B(WX9228), .Z(WX9227) ) ;
AND2    gate10953  (.A(CRC_OUT_2_21), .B(WX10055), .Z(WX9230) ) ;
AND2    gate10954  (.A(WX11426), .B(WX9232), .Z(WX9231) ) ;
AND2    gate10955  (.A(WX9556), .B(WX10055), .Z(WX9234) ) ;
AND2    gate10956  (.A(WX10133), .B(WX9236), .Z(WX9235) ) ;
OR2     gate10957  (.A(WX9249), .B(WX9248), .Z(WX9251) ) ;
AND2    gate10958  (.A(WX9251), .B(WX10054), .Z(WX9240) ) ;
OR2     gate10959  (.A(WX9245), .B(WX9244), .Z(WX9247) ) ;
AND2    gate10960  (.A(WX9247), .B(WX9242), .Z(WX9241) ) ;
AND2    gate10961  (.A(CRC_OUT_2_20), .B(WX10055), .Z(WX9244) ) ;
AND2    gate10962  (.A(WX11433), .B(WX9246), .Z(WX9245) ) ;
AND2    gate10963  (.A(WX9558), .B(WX10055), .Z(WX9248) ) ;
AND2    gate10964  (.A(WX10140), .B(WX9250), .Z(WX9249) ) ;
OR2     gate10965  (.A(WX9263), .B(WX9262), .Z(WX9265) ) ;
AND2    gate10966  (.A(WX9265), .B(WX10054), .Z(WX9254) ) ;
OR2     gate10967  (.A(WX9259), .B(WX9258), .Z(WX9261) ) ;
AND2    gate10968  (.A(WX9261), .B(WX9256), .Z(WX9255) ) ;
AND2    gate10969  (.A(CRC_OUT_2_19), .B(WX10055), .Z(WX9258) ) ;
AND2    gate10970  (.A(WX11440), .B(WX9260), .Z(WX9259) ) ;
AND2    gate10971  (.A(WX9560), .B(WX10055), .Z(WX9262) ) ;
AND2    gate10972  (.A(WX10147), .B(WX9264), .Z(WX9263) ) ;
OR2     gate10973  (.A(WX9277), .B(WX9276), .Z(WX9279) ) ;
AND2    gate10974  (.A(WX9279), .B(WX10054), .Z(WX9268) ) ;
OR2     gate10975  (.A(WX9273), .B(WX9272), .Z(WX9275) ) ;
AND2    gate10976  (.A(WX9275), .B(WX9270), .Z(WX9269) ) ;
AND2    gate10977  (.A(CRC_OUT_2_18), .B(WX10055), .Z(WX9272) ) ;
AND2    gate10978  (.A(WX11447), .B(WX9274), .Z(WX9273) ) ;
AND2    gate10979  (.A(WX9562), .B(WX10055), .Z(WX9276) ) ;
AND2    gate10980  (.A(WX10154), .B(WX9278), .Z(WX9277) ) ;
OR2     gate10981  (.A(WX9291), .B(WX9290), .Z(WX9293) ) ;
AND2    gate10982  (.A(WX9293), .B(WX10054), .Z(WX9282) ) ;
OR2     gate10983  (.A(WX9287), .B(WX9286), .Z(WX9289) ) ;
AND2    gate10984  (.A(WX9289), .B(WX9284), .Z(WX9283) ) ;
AND2    gate10985  (.A(CRC_OUT_2_17), .B(WX10055), .Z(WX9286) ) ;
AND2    gate10986  (.A(WX11454), .B(WX9288), .Z(WX9287) ) ;
AND2    gate10987  (.A(WX9564), .B(WX10055), .Z(WX9290) ) ;
AND2    gate10988  (.A(WX10161), .B(WX9292), .Z(WX9291) ) ;
OR2     gate10989  (.A(WX9305), .B(WX9304), .Z(WX9307) ) ;
AND2    gate10990  (.A(WX9307), .B(WX10054), .Z(WX9296) ) ;
OR2     gate10991  (.A(WX9301), .B(WX9300), .Z(WX9303) ) ;
AND2    gate10992  (.A(WX9303), .B(WX9298), .Z(WX9297) ) ;
AND2    gate10993  (.A(CRC_OUT_2_16), .B(WX10055), .Z(WX9300) ) ;
AND2    gate10994  (.A(WX11461), .B(WX9302), .Z(WX9301) ) ;
AND2    gate10995  (.A(WX9566), .B(WX10055), .Z(WX9304) ) ;
AND2    gate10996  (.A(WX10168), .B(WX9306), .Z(WX9305) ) ;
OR2     gate10997  (.A(WX9319), .B(WX9318), .Z(WX9321) ) ;
AND2    gate10998  (.A(WX9321), .B(WX10054), .Z(WX9310) ) ;
OR2     gate10999  (.A(WX9315), .B(WX9314), .Z(WX9317) ) ;
AND2    gate11000  (.A(WX9317), .B(WX9312), .Z(WX9311) ) ;
AND2    gate11001  (.A(CRC_OUT_2_15), .B(WX10055), .Z(WX9314) ) ;
AND2    gate11002  (.A(WX11468), .B(WX9316), .Z(WX9315) ) ;
AND2    gate11003  (.A(WX9568), .B(WX10055), .Z(WX9318) ) ;
AND2    gate11004  (.A(WX10175), .B(WX9320), .Z(WX9319) ) ;
OR2     gate11005  (.A(WX9333), .B(WX9332), .Z(WX9335) ) ;
AND2    gate11006  (.A(WX9335), .B(WX10054), .Z(WX9324) ) ;
OR2     gate11007  (.A(WX9329), .B(WX9328), .Z(WX9331) ) ;
AND2    gate11008  (.A(WX9331), .B(WX9326), .Z(WX9325) ) ;
AND2    gate11009  (.A(CRC_OUT_2_14), .B(WX10055), .Z(WX9328) ) ;
AND2    gate11010  (.A(WX11475), .B(WX9330), .Z(WX9329) ) ;
AND2    gate11011  (.A(WX9570), .B(WX10055), .Z(WX9332) ) ;
AND2    gate11012  (.A(WX10182), .B(WX9334), .Z(WX9333) ) ;
OR2     gate11013  (.A(WX9347), .B(WX9346), .Z(WX9349) ) ;
AND2    gate11014  (.A(WX9349), .B(WX10054), .Z(WX9338) ) ;
OR2     gate11015  (.A(WX9343), .B(WX9342), .Z(WX9345) ) ;
AND2    gate11016  (.A(WX9345), .B(WX9340), .Z(WX9339) ) ;
AND2    gate11017  (.A(CRC_OUT_2_13), .B(WX10055), .Z(WX9342) ) ;
AND2    gate11018  (.A(WX11482), .B(WX9344), .Z(WX9343) ) ;
AND2    gate11019  (.A(WX9572), .B(WX10055), .Z(WX9346) ) ;
AND2    gate11020  (.A(WX10189), .B(WX9348), .Z(WX9347) ) ;
OR2     gate11021  (.A(WX9361), .B(WX9360), .Z(WX9363) ) ;
AND2    gate11022  (.A(WX9363), .B(WX10054), .Z(WX9352) ) ;
OR2     gate11023  (.A(WX9357), .B(WX9356), .Z(WX9359) ) ;
AND2    gate11024  (.A(WX9359), .B(WX9354), .Z(WX9353) ) ;
AND2    gate11025  (.A(CRC_OUT_2_12), .B(WX10055), .Z(WX9356) ) ;
AND2    gate11026  (.A(WX11489), .B(WX9358), .Z(WX9357) ) ;
AND2    gate11027  (.A(WX9574), .B(WX10055), .Z(WX9360) ) ;
AND2    gate11028  (.A(WX10196), .B(WX9362), .Z(WX9361) ) ;
OR2     gate11029  (.A(WX9375), .B(WX9374), .Z(WX9377) ) ;
AND2    gate11030  (.A(WX9377), .B(WX10054), .Z(WX9366) ) ;
OR2     gate11031  (.A(WX9371), .B(WX9370), .Z(WX9373) ) ;
AND2    gate11032  (.A(WX9373), .B(WX9368), .Z(WX9367) ) ;
AND2    gate11033  (.A(CRC_OUT_2_11), .B(WX10055), .Z(WX9370) ) ;
AND2    gate11034  (.A(WX11496), .B(WX9372), .Z(WX9371) ) ;
AND2    gate11035  (.A(WX9576), .B(WX10055), .Z(WX9374) ) ;
AND2    gate11036  (.A(WX10203), .B(WX9376), .Z(WX9375) ) ;
OR2     gate11037  (.A(WX9389), .B(WX9388), .Z(WX9391) ) ;
AND2    gate11038  (.A(WX9391), .B(WX10054), .Z(WX9380) ) ;
OR2     gate11039  (.A(WX9385), .B(WX9384), .Z(WX9387) ) ;
AND2    gate11040  (.A(WX9387), .B(WX9382), .Z(WX9381) ) ;
AND2    gate11041  (.A(CRC_OUT_2_10), .B(WX10055), .Z(WX9384) ) ;
AND2    gate11042  (.A(WX11503), .B(WX9386), .Z(WX9385) ) ;
AND2    gate11043  (.A(WX9578), .B(WX10055), .Z(WX9388) ) ;
AND2    gate11044  (.A(WX10210), .B(WX9390), .Z(WX9389) ) ;
OR2     gate11045  (.A(WX9403), .B(WX9402), .Z(WX9405) ) ;
AND2    gate11046  (.A(WX9405), .B(WX10054), .Z(WX9394) ) ;
OR2     gate11047  (.A(WX9399), .B(WX9398), .Z(WX9401) ) ;
AND2    gate11048  (.A(WX9401), .B(WX9396), .Z(WX9395) ) ;
AND2    gate11049  (.A(CRC_OUT_2_9), .B(WX10055), .Z(WX9398) ) ;
AND2    gate11050  (.A(WX11510), .B(WX9400), .Z(WX9399) ) ;
AND2    gate11051  (.A(WX9580), .B(WX10055), .Z(WX9402) ) ;
AND2    gate11052  (.A(WX10217), .B(WX9404), .Z(WX9403) ) ;
OR2     gate11053  (.A(WX9417), .B(WX9416), .Z(WX9419) ) ;
AND2    gate11054  (.A(WX9419), .B(WX10054), .Z(WX9408) ) ;
OR2     gate11055  (.A(WX9413), .B(WX9412), .Z(WX9415) ) ;
AND2    gate11056  (.A(WX9415), .B(WX9410), .Z(WX9409) ) ;
AND2    gate11057  (.A(CRC_OUT_2_8), .B(WX10055), .Z(WX9412) ) ;
AND2    gate11058  (.A(WX11517), .B(WX9414), .Z(WX9413) ) ;
AND2    gate11059  (.A(WX9582), .B(WX10055), .Z(WX9416) ) ;
AND2    gate11060  (.A(WX10224), .B(WX9418), .Z(WX9417) ) ;
OR2     gate11061  (.A(WX9431), .B(WX9430), .Z(WX9433) ) ;
AND2    gate11062  (.A(WX9433), .B(WX10054), .Z(WX9422) ) ;
OR2     gate11063  (.A(WX9427), .B(WX9426), .Z(WX9429) ) ;
AND2    gate11064  (.A(WX9429), .B(WX9424), .Z(WX9423) ) ;
AND2    gate11065  (.A(CRC_OUT_2_7), .B(WX10055), .Z(WX9426) ) ;
AND2    gate11066  (.A(WX11524), .B(WX9428), .Z(WX9427) ) ;
AND2    gate11067  (.A(WX9584), .B(WX10055), .Z(WX9430) ) ;
AND2    gate11068  (.A(WX10231), .B(WX9432), .Z(WX9431) ) ;
OR2     gate11069  (.A(WX9445), .B(WX9444), .Z(WX9447) ) ;
AND2    gate11070  (.A(WX9447), .B(WX10054), .Z(WX9436) ) ;
OR2     gate11071  (.A(WX9441), .B(WX9440), .Z(WX9443) ) ;
AND2    gate11072  (.A(WX9443), .B(WX9438), .Z(WX9437) ) ;
AND2    gate11073  (.A(CRC_OUT_2_6), .B(WX10055), .Z(WX9440) ) ;
AND2    gate11074  (.A(WX11531), .B(WX9442), .Z(WX9441) ) ;
AND2    gate11075  (.A(WX9586), .B(WX10055), .Z(WX9444) ) ;
AND2    gate11076  (.A(WX10238), .B(WX9446), .Z(WX9445) ) ;
OR2     gate11077  (.A(WX9459), .B(WX9458), .Z(WX9461) ) ;
AND2    gate11078  (.A(WX9461), .B(WX10054), .Z(WX9450) ) ;
OR2     gate11079  (.A(WX9455), .B(WX9454), .Z(WX9457) ) ;
AND2    gate11080  (.A(WX9457), .B(WX9452), .Z(WX9451) ) ;
AND2    gate11081  (.A(CRC_OUT_2_5), .B(WX10055), .Z(WX9454) ) ;
AND2    gate11082  (.A(WX11538), .B(WX9456), .Z(WX9455) ) ;
AND2    gate11083  (.A(WX9588), .B(WX10055), .Z(WX9458) ) ;
AND2    gate11084  (.A(WX10245), .B(WX9460), .Z(WX9459) ) ;
OR2     gate11085  (.A(WX9473), .B(WX9472), .Z(WX9475) ) ;
AND2    gate11086  (.A(WX9475), .B(WX10054), .Z(WX9464) ) ;
OR2     gate11087  (.A(WX9469), .B(WX9468), .Z(WX9471) ) ;
AND2    gate11088  (.A(WX9471), .B(WX9466), .Z(WX9465) ) ;
AND2    gate11089  (.A(CRC_OUT_2_4), .B(WX10055), .Z(WX9468) ) ;
AND2    gate11090  (.A(WX11545), .B(WX9470), .Z(WX9469) ) ;
AND2    gate11091  (.A(WX9590), .B(WX10055), .Z(WX9472) ) ;
AND2    gate11092  (.A(WX10252), .B(WX9474), .Z(WX9473) ) ;
OR2     gate11093  (.A(WX9487), .B(WX9486), .Z(WX9489) ) ;
AND2    gate11094  (.A(WX9489), .B(WX10054), .Z(WX9478) ) ;
OR2     gate11095  (.A(WX9483), .B(WX9482), .Z(WX9485) ) ;
AND2    gate11096  (.A(WX9485), .B(WX9480), .Z(WX9479) ) ;
AND2    gate11097  (.A(CRC_OUT_2_3), .B(WX10055), .Z(WX9482) ) ;
AND2    gate11098  (.A(WX11552), .B(WX9484), .Z(WX9483) ) ;
AND2    gate11099  (.A(WX9592), .B(WX10055), .Z(WX9486) ) ;
AND2    gate11100  (.A(WX10259), .B(WX9488), .Z(WX9487) ) ;
OR2     gate11101  (.A(WX9501), .B(WX9500), .Z(WX9503) ) ;
AND2    gate11102  (.A(WX9503), .B(WX10054), .Z(WX9492) ) ;
OR2     gate11103  (.A(WX9497), .B(WX9496), .Z(WX9499) ) ;
AND2    gate11104  (.A(WX9499), .B(WX9494), .Z(WX9493) ) ;
AND2    gate11105  (.A(CRC_OUT_2_2), .B(WX10055), .Z(WX9496) ) ;
AND2    gate11106  (.A(WX11559), .B(WX9498), .Z(WX9497) ) ;
AND2    gate11107  (.A(WX9594), .B(WX10055), .Z(WX9500) ) ;
AND2    gate11108  (.A(WX10266), .B(WX9502), .Z(WX9501) ) ;
OR2     gate11109  (.A(WX9515), .B(WX9514), .Z(WX9517) ) ;
AND2    gate11110  (.A(WX9517), .B(WX10054), .Z(WX9506) ) ;
OR2     gate11111  (.A(WX9511), .B(WX9510), .Z(WX9513) ) ;
AND2    gate11112  (.A(WX9513), .B(WX9508), .Z(WX9507) ) ;
AND2    gate11113  (.A(CRC_OUT_2_1), .B(WX10055), .Z(WX9510) ) ;
AND2    gate11114  (.A(WX11566), .B(WX9512), .Z(WX9511) ) ;
AND2    gate11115  (.A(WX9596), .B(WX10055), .Z(WX9514) ) ;
AND2    gate11116  (.A(WX10273), .B(WX9516), .Z(WX9515) ) ;
OR2     gate11117  (.A(WX9529), .B(WX9528), .Z(WX9531) ) ;
AND2    gate11118  (.A(WX9531), .B(WX10054), .Z(WX9520) ) ;
OR2     gate11119  (.A(WX9525), .B(WX9524), .Z(WX9527) ) ;
AND2    gate11120  (.A(WX9527), .B(WX9522), .Z(WX9521) ) ;
AND2    gate11121  (.A(CRC_OUT_2_0), .B(WX10055), .Z(WX9524) ) ;
AND2    gate11122  (.A(WX11573), .B(WX9526), .Z(WX9525) ) ;
AND2    gate11123  (.A(WX9598), .B(WX10055), .Z(WX9528) ) ;
AND2    gate11124  (.A(WX10280), .B(WX9530), .Z(WX9529) ) ;
NAND2   gate11125  (.A(II31088), .B(II31089), .Z(WX10057) ) ;
AND2    gate11126  (.A(WX10057), .B(WX10056), .Z(WX10058) ) ;
AND2    gate11127  (.A(WX9631), .B(WX10060), .Z(WX10059) ) ;
NAND2   gate11128  (.A(II31101), .B(II31102), .Z(WX10064) ) ;
AND2    gate11129  (.A(WX10064), .B(WX10056), .Z(WX10065) ) ;
AND2    gate11130  (.A(WX9632), .B(WX10067), .Z(WX10066) ) ;
NAND2   gate11131  (.A(II31114), .B(II31115), .Z(WX10071) ) ;
AND2    gate11132  (.A(WX10071), .B(WX10056), .Z(WX10072) ) ;
AND2    gate11133  (.A(WX9633), .B(WX10074), .Z(WX10073) ) ;
NAND2   gate11134  (.A(II31127), .B(II31128), .Z(WX10078) ) ;
AND2    gate11135  (.A(WX10078), .B(WX10056), .Z(WX10079) ) ;
AND2    gate11136  (.A(WX9634), .B(WX10081), .Z(WX10080) ) ;
NAND2   gate11137  (.A(II31140), .B(II31141), .Z(WX10085) ) ;
AND2    gate11138  (.A(WX10085), .B(WX10056), .Z(WX10086) ) ;
AND2    gate11139  (.A(WX9635), .B(WX10088), .Z(WX10087) ) ;
NAND2   gate11140  (.A(II31153), .B(II31154), .Z(WX10092) ) ;
AND2    gate11141  (.A(WX10092), .B(WX10056), .Z(WX10093) ) ;
AND2    gate11142  (.A(WX9636), .B(WX10095), .Z(WX10094) ) ;
NAND2   gate11143  (.A(II31166), .B(II31167), .Z(WX10099) ) ;
AND2    gate11144  (.A(WX10099), .B(WX10056), .Z(WX10100) ) ;
AND2    gate11145  (.A(WX9637), .B(WX10102), .Z(WX10101) ) ;
NAND2   gate11146  (.A(II31179), .B(II31180), .Z(WX10106) ) ;
AND2    gate11147  (.A(WX10106), .B(WX10056), .Z(WX10107) ) ;
AND2    gate11148  (.A(WX9638), .B(WX10109), .Z(WX10108) ) ;
NAND2   gate11149  (.A(II31192), .B(II31193), .Z(WX10113) ) ;
AND2    gate11150  (.A(WX10113), .B(WX10056), .Z(WX10114) ) ;
AND2    gate11151  (.A(WX9639), .B(WX10116), .Z(WX10115) ) ;
NAND2   gate11152  (.A(II31205), .B(II31206), .Z(WX10120) ) ;
AND2    gate11153  (.A(WX10120), .B(WX10056), .Z(WX10121) ) ;
AND2    gate11154  (.A(WX9640), .B(WX10123), .Z(WX10122) ) ;
NAND2   gate11155  (.A(II31218), .B(II31219), .Z(WX10127) ) ;
AND2    gate11156  (.A(WX10127), .B(WX10056), .Z(WX10128) ) ;
AND2    gate11157  (.A(WX9641), .B(WX10130), .Z(WX10129) ) ;
NAND2   gate11158  (.A(II31231), .B(II31232), .Z(WX10134) ) ;
AND2    gate11159  (.A(WX10134), .B(WX10056), .Z(WX10135) ) ;
AND2    gate11160  (.A(WX9642), .B(WX10137), .Z(WX10136) ) ;
NAND2   gate11161  (.A(II31244), .B(II31245), .Z(WX10141) ) ;
AND2    gate11162  (.A(WX10141), .B(WX10056), .Z(WX10142) ) ;
AND2    gate11163  (.A(WX9643), .B(WX10144), .Z(WX10143) ) ;
NAND2   gate11164  (.A(II31257), .B(II31258), .Z(WX10148) ) ;
AND2    gate11165  (.A(WX10148), .B(WX10056), .Z(WX10149) ) ;
AND2    gate11166  (.A(WX9644), .B(WX10151), .Z(WX10150) ) ;
NAND2   gate11167  (.A(II31270), .B(II31271), .Z(WX10155) ) ;
AND2    gate11168  (.A(WX10155), .B(WX10056), .Z(WX10156) ) ;
AND2    gate11169  (.A(WX9645), .B(WX10158), .Z(WX10157) ) ;
NAND2   gate11170  (.A(II31283), .B(II31284), .Z(WX10162) ) ;
AND2    gate11171  (.A(WX10162), .B(WX10056), .Z(WX10163) ) ;
AND2    gate11172  (.A(WX9646), .B(WX10165), .Z(WX10164) ) ;
NAND2   gate11173  (.A(II31296), .B(II31297), .Z(WX10169) ) ;
AND2    gate11174  (.A(WX10169), .B(WX10056), .Z(WX10170) ) ;
AND2    gate11175  (.A(WX9647), .B(WX10172), .Z(WX10171) ) ;
NAND2   gate11176  (.A(II31309), .B(II31310), .Z(WX10176) ) ;
AND2    gate11177  (.A(WX10176), .B(WX10056), .Z(WX10177) ) ;
AND2    gate11178  (.A(WX9648), .B(WX10179), .Z(WX10178) ) ;
NAND2   gate11179  (.A(II31322), .B(II31323), .Z(WX10183) ) ;
AND2    gate11180  (.A(WX10183), .B(WX10056), .Z(WX10184) ) ;
AND2    gate11181  (.A(WX9649), .B(WX10186), .Z(WX10185) ) ;
NAND2   gate11182  (.A(II31335), .B(II31336), .Z(WX10190) ) ;
AND2    gate11183  (.A(WX10190), .B(WX10056), .Z(WX10191) ) ;
AND2    gate11184  (.A(WX9650), .B(WX10193), .Z(WX10192) ) ;
NAND2   gate11185  (.A(II31348), .B(II31349), .Z(WX10197) ) ;
AND2    gate11186  (.A(WX10197), .B(WX10056), .Z(WX10198) ) ;
AND2    gate11187  (.A(WX9651), .B(WX10200), .Z(WX10199) ) ;
NAND2   gate11188  (.A(II31361), .B(II31362), .Z(WX10204) ) ;
AND2    gate11189  (.A(WX10204), .B(WX10056), .Z(WX10205) ) ;
AND2    gate11190  (.A(WX9652), .B(WX10207), .Z(WX10206) ) ;
NAND2   gate11191  (.A(II31374), .B(II31375), .Z(WX10211) ) ;
AND2    gate11192  (.A(WX10211), .B(WX10056), .Z(WX10212) ) ;
AND2    gate11193  (.A(WX9653), .B(WX10214), .Z(WX10213) ) ;
NAND2   gate11194  (.A(II31387), .B(II31388), .Z(WX10218) ) ;
AND2    gate11195  (.A(WX10218), .B(WX10056), .Z(WX10219) ) ;
AND2    gate11196  (.A(WX9654), .B(WX10221), .Z(WX10220) ) ;
NAND2   gate11197  (.A(II31400), .B(II31401), .Z(WX10225) ) ;
AND2    gate11198  (.A(WX10225), .B(WX10056), .Z(WX10226) ) ;
AND2    gate11199  (.A(WX9655), .B(WX10228), .Z(WX10227) ) ;
NAND2   gate11200  (.A(II31413), .B(II31414), .Z(WX10232) ) ;
AND2    gate11201  (.A(WX10232), .B(WX10056), .Z(WX10233) ) ;
AND2    gate11202  (.A(WX9656), .B(WX10235), .Z(WX10234) ) ;
NAND2   gate11203  (.A(II31426), .B(II31427), .Z(WX10239) ) ;
AND2    gate11204  (.A(WX10239), .B(WX10056), .Z(WX10240) ) ;
AND2    gate11205  (.A(WX9657), .B(WX10242), .Z(WX10241) ) ;
NAND2   gate11206  (.A(II31439), .B(II31440), .Z(WX10246) ) ;
AND2    gate11207  (.A(WX10246), .B(WX10056), .Z(WX10247) ) ;
AND2    gate11208  (.A(WX9658), .B(WX10249), .Z(WX10248) ) ;
NAND2   gate11209  (.A(II31452), .B(II31453), .Z(WX10253) ) ;
AND2    gate11210  (.A(WX10253), .B(WX10056), .Z(WX10254) ) ;
AND2    gate11211  (.A(WX9659), .B(WX10256), .Z(WX10255) ) ;
NAND2   gate11212  (.A(II31465), .B(II31466), .Z(WX10260) ) ;
AND2    gate11213  (.A(WX10260), .B(WX10056), .Z(WX10261) ) ;
AND2    gate11214  (.A(WX9660), .B(WX10263), .Z(WX10262) ) ;
NAND2   gate11215  (.A(II31478), .B(II31479), .Z(WX10267) ) ;
AND2    gate11216  (.A(WX10267), .B(WX10056), .Z(WX10268) ) ;
AND2    gate11217  (.A(WX9661), .B(WX10270), .Z(WX10269) ) ;
NAND2   gate11218  (.A(II31491), .B(II31492), .Z(WX10274) ) ;
AND2    gate11219  (.A(WX10274), .B(WX10056), .Z(WX10275) ) ;
AND2    gate11220  (.A(WX9662), .B(WX10277), .Z(WX10276) ) ;
NAND2   gate11221  (.A(II31550), .B(II31551), .Z(WX10285) ) ;
NAND2   gate11222  (.A(II31746), .B(II31747), .Z(WX10313) ) ;
NAND2   gate11223  (.A(II31739), .B(II31740), .Z(WX10312) ) ;
NAND2   gate11224  (.A(II31732), .B(II31733), .Z(WX10311) ) ;
NAND2   gate11225  (.A(II31543), .B(II31544), .Z(WX10284) ) ;
NAND2   gate11226  (.A(II31725), .B(II31726), .Z(WX10310) ) ;
NAND2   gate11227  (.A(II31718), .B(II31719), .Z(WX10309) ) ;
NAND2   gate11228  (.A(II31711), .B(II31712), .Z(WX10308) ) ;
NAND2   gate11229  (.A(II31704), .B(II31705), .Z(WX10307) ) ;
NAND2   gate11230  (.A(II31697), .B(II31698), .Z(WX10306) ) ;
NAND2   gate11231  (.A(II31690), .B(II31691), .Z(WX10305) ) ;
NAND2   gate11232  (.A(II31528), .B(II31529), .Z(WX10283) ) ;
NAND2   gate11233  (.A(II31683), .B(II31684), .Z(WX10304) ) ;
NAND2   gate11234  (.A(II31676), .B(II31677), .Z(WX10303) ) ;
NAND2   gate11235  (.A(II31669), .B(II31670), .Z(WX10302) ) ;
NAND2   gate11236  (.A(II31662), .B(II31663), .Z(WX10301) ) ;
NAND2   gate11237  (.A(II31513), .B(II31514), .Z(WX10282) ) ;
NAND2   gate11238  (.A(II31655), .B(II31656), .Z(WX10300) ) ;
NAND2   gate11239  (.A(II31648), .B(II31649), .Z(WX10299) ) ;
NAND2   gate11240  (.A(II31641), .B(II31642), .Z(WX10298) ) ;
NAND2   gate11241  (.A(II31634), .B(II31635), .Z(WX10297) ) ;
NAND2   gate11242  (.A(II31627), .B(II31628), .Z(WX10296) ) ;
NAND2   gate11243  (.A(II31620), .B(II31621), .Z(WX10295) ) ;
NAND2   gate11244  (.A(II31613), .B(II31614), .Z(WX10294) ) ;
NAND2   gate11245  (.A(II31606), .B(II31607), .Z(WX10293) ) ;
NAND2   gate11246  (.A(II31599), .B(II31600), .Z(WX10292) ) ;
NAND2   gate11247  (.A(II31592), .B(II31593), .Z(WX10291) ) ;
NAND2   gate11248  (.A(II31585), .B(II31586), .Z(WX10290) ) ;
NAND2   gate11249  (.A(II31578), .B(II31579), .Z(WX10289) ) ;
NAND2   gate11250  (.A(II31571), .B(II31572), .Z(WX10288) ) ;
NAND2   gate11251  (.A(II31564), .B(II31565), .Z(WX10287) ) ;
NAND2   gate11252  (.A(II31557), .B(II31558), .Z(WX10286) ) ;
OR2     gate11253  (.A(WX10388), .B(WX10387), .Z(WX10390) ) ;
AND2    gate11254  (.A(WX10390), .B(WX11347), .Z(WX10379) ) ;
OR2     gate11255  (.A(WX10384), .B(WX10383), .Z(WX10386) ) ;
AND2    gate11256  (.A(WX10386), .B(WX10381), .Z(WX10380) ) ;
AND2    gate11257  (.A(CRC_OUT_1_31), .B(WX11348), .Z(WX10383) ) ;
AND2    gate11258  (.A(DATA_0_31), .B(WX10385), .Z(WX10384) ) ;
AND2    gate11259  (.A(WX10829), .B(WX11348), .Z(WX10387) ) ;
AND2    gate11260  (.A(WX11356), .B(WX10389), .Z(WX10388) ) ;
OR2     gate11261  (.A(WX10402), .B(WX10401), .Z(WX10404) ) ;
AND2    gate11262  (.A(WX10404), .B(WX11347), .Z(WX10393) ) ;
OR2     gate11263  (.A(WX10398), .B(WX10397), .Z(WX10400) ) ;
AND2    gate11264  (.A(WX10400), .B(WX10395), .Z(WX10394) ) ;
AND2    gate11265  (.A(CRC_OUT_1_30), .B(WX11348), .Z(WX10397) ) ;
AND2    gate11266  (.A(DATA_0_30), .B(WX10399), .Z(WX10398) ) ;
AND2    gate11267  (.A(WX10831), .B(WX11348), .Z(WX10401) ) ;
AND2    gate11268  (.A(WX11363), .B(WX10403), .Z(WX10402) ) ;
OR2     gate11269  (.A(WX10416), .B(WX10415), .Z(WX10418) ) ;
AND2    gate11270  (.A(WX10418), .B(WX11347), .Z(WX10407) ) ;
OR2     gate11271  (.A(WX10412), .B(WX10411), .Z(WX10414) ) ;
AND2    gate11272  (.A(WX10414), .B(WX10409), .Z(WX10408) ) ;
AND2    gate11273  (.A(CRC_OUT_1_29), .B(WX11348), .Z(WX10411) ) ;
AND2    gate11274  (.A(DATA_0_29), .B(WX10413), .Z(WX10412) ) ;
AND2    gate11275  (.A(WX10833), .B(WX11348), .Z(WX10415) ) ;
AND2    gate11276  (.A(WX11370), .B(WX10417), .Z(WX10416) ) ;
OR2     gate11277  (.A(WX10430), .B(WX10429), .Z(WX10432) ) ;
AND2    gate11278  (.A(WX10432), .B(WX11347), .Z(WX10421) ) ;
OR2     gate11279  (.A(WX10426), .B(WX10425), .Z(WX10428) ) ;
AND2    gate11280  (.A(WX10428), .B(WX10423), .Z(WX10422) ) ;
AND2    gate11281  (.A(CRC_OUT_1_28), .B(WX11348), .Z(WX10425) ) ;
AND2    gate11282  (.A(DATA_0_28), .B(WX10427), .Z(WX10426) ) ;
AND2    gate11283  (.A(WX10835), .B(WX11348), .Z(WX10429) ) ;
AND2    gate11284  (.A(WX11377), .B(WX10431), .Z(WX10430) ) ;
OR2     gate11285  (.A(WX10444), .B(WX10443), .Z(WX10446) ) ;
AND2    gate11286  (.A(WX10446), .B(WX11347), .Z(WX10435) ) ;
OR2     gate11287  (.A(WX10440), .B(WX10439), .Z(WX10442) ) ;
AND2    gate11288  (.A(WX10442), .B(WX10437), .Z(WX10436) ) ;
AND2    gate11289  (.A(CRC_OUT_1_27), .B(WX11348), .Z(WX10439) ) ;
AND2    gate11290  (.A(DATA_0_27), .B(WX10441), .Z(WX10440) ) ;
AND2    gate11291  (.A(WX10837), .B(WX11348), .Z(WX10443) ) ;
AND2    gate11292  (.A(WX11384), .B(WX10445), .Z(WX10444) ) ;
OR2     gate11293  (.A(WX10458), .B(WX10457), .Z(WX10460) ) ;
AND2    gate11294  (.A(WX10460), .B(WX11347), .Z(WX10449) ) ;
OR2     gate11295  (.A(WX10454), .B(WX10453), .Z(WX10456) ) ;
AND2    gate11296  (.A(WX10456), .B(WX10451), .Z(WX10450) ) ;
AND2    gate11297  (.A(CRC_OUT_1_26), .B(WX11348), .Z(WX10453) ) ;
AND2    gate11298  (.A(DATA_0_26), .B(WX10455), .Z(WX10454) ) ;
AND2    gate11299  (.A(WX10839), .B(WX11348), .Z(WX10457) ) ;
AND2    gate11300  (.A(WX11391), .B(WX10459), .Z(WX10458) ) ;
OR2     gate11301  (.A(WX10472), .B(WX10471), .Z(WX10474) ) ;
AND2    gate11302  (.A(WX10474), .B(WX11347), .Z(WX10463) ) ;
OR2     gate11303  (.A(WX10468), .B(WX10467), .Z(WX10470) ) ;
AND2    gate11304  (.A(WX10470), .B(WX10465), .Z(WX10464) ) ;
AND2    gate11305  (.A(CRC_OUT_1_25), .B(WX11348), .Z(WX10467) ) ;
AND2    gate11306  (.A(DATA_0_25), .B(WX10469), .Z(WX10468) ) ;
AND2    gate11307  (.A(WX10841), .B(WX11348), .Z(WX10471) ) ;
AND2    gate11308  (.A(WX11398), .B(WX10473), .Z(WX10472) ) ;
OR2     gate11309  (.A(WX10486), .B(WX10485), .Z(WX10488) ) ;
AND2    gate11310  (.A(WX10488), .B(WX11347), .Z(WX10477) ) ;
OR2     gate11311  (.A(WX10482), .B(WX10481), .Z(WX10484) ) ;
AND2    gate11312  (.A(WX10484), .B(WX10479), .Z(WX10478) ) ;
AND2    gate11313  (.A(CRC_OUT_1_24), .B(WX11348), .Z(WX10481) ) ;
AND2    gate11314  (.A(DATA_0_24), .B(WX10483), .Z(WX10482) ) ;
AND2    gate11315  (.A(WX10843), .B(WX11348), .Z(WX10485) ) ;
AND2    gate11316  (.A(WX11405), .B(WX10487), .Z(WX10486) ) ;
OR2     gate11317  (.A(WX10500), .B(WX10499), .Z(WX10502) ) ;
AND2    gate11318  (.A(WX10502), .B(WX11347), .Z(WX10491) ) ;
OR2     gate11319  (.A(WX10496), .B(WX10495), .Z(WX10498) ) ;
AND2    gate11320  (.A(WX10498), .B(WX10493), .Z(WX10492) ) ;
AND2    gate11321  (.A(CRC_OUT_1_23), .B(WX11348), .Z(WX10495) ) ;
AND2    gate11322  (.A(DATA_0_23), .B(WX10497), .Z(WX10496) ) ;
AND2    gate11323  (.A(WX10845), .B(WX11348), .Z(WX10499) ) ;
AND2    gate11324  (.A(WX11412), .B(WX10501), .Z(WX10500) ) ;
OR2     gate11325  (.A(WX10514), .B(WX10513), .Z(WX10516) ) ;
AND2    gate11326  (.A(WX10516), .B(WX11347), .Z(WX10505) ) ;
OR2     gate11327  (.A(WX10510), .B(WX10509), .Z(WX10512) ) ;
AND2    gate11328  (.A(WX10512), .B(WX10507), .Z(WX10506) ) ;
AND2    gate11329  (.A(CRC_OUT_1_22), .B(WX11348), .Z(WX10509) ) ;
AND2    gate11330  (.A(DATA_0_22), .B(WX10511), .Z(WX10510) ) ;
AND2    gate11331  (.A(WX10847), .B(WX11348), .Z(WX10513) ) ;
AND2    gate11332  (.A(WX11419), .B(WX10515), .Z(WX10514) ) ;
OR2     gate11333  (.A(WX10528), .B(WX10527), .Z(WX10530) ) ;
AND2    gate11334  (.A(WX10530), .B(WX11347), .Z(WX10519) ) ;
OR2     gate11335  (.A(WX10524), .B(WX10523), .Z(WX10526) ) ;
AND2    gate11336  (.A(WX10526), .B(WX10521), .Z(WX10520) ) ;
AND2    gate11337  (.A(CRC_OUT_1_21), .B(WX11348), .Z(WX10523) ) ;
AND2    gate11338  (.A(DATA_0_21), .B(WX10525), .Z(WX10524) ) ;
AND2    gate11339  (.A(WX10849), .B(WX11348), .Z(WX10527) ) ;
AND2    gate11340  (.A(WX11426), .B(WX10529), .Z(WX10528) ) ;
OR2     gate11341  (.A(WX10542), .B(WX10541), .Z(WX10544) ) ;
AND2    gate11342  (.A(WX10544), .B(WX11347), .Z(WX10533) ) ;
OR2     gate11343  (.A(WX10538), .B(WX10537), .Z(WX10540) ) ;
AND2    gate11344  (.A(WX10540), .B(WX10535), .Z(WX10534) ) ;
AND2    gate11345  (.A(CRC_OUT_1_20), .B(WX11348), .Z(WX10537) ) ;
AND2    gate11346  (.A(DATA_0_20), .B(WX10539), .Z(WX10538) ) ;
AND2    gate11347  (.A(WX10851), .B(WX11348), .Z(WX10541) ) ;
AND2    gate11348  (.A(WX11433), .B(WX10543), .Z(WX10542) ) ;
OR2     gate11349  (.A(WX10556), .B(WX10555), .Z(WX10558) ) ;
AND2    gate11350  (.A(WX10558), .B(WX11347), .Z(WX10547) ) ;
OR2     gate11351  (.A(WX10552), .B(WX10551), .Z(WX10554) ) ;
AND2    gate11352  (.A(WX10554), .B(WX10549), .Z(WX10548) ) ;
AND2    gate11353  (.A(CRC_OUT_1_19), .B(WX11348), .Z(WX10551) ) ;
AND2    gate11354  (.A(DATA_0_19), .B(WX10553), .Z(WX10552) ) ;
AND2    gate11355  (.A(WX10853), .B(WX11348), .Z(WX10555) ) ;
AND2    gate11356  (.A(WX11440), .B(WX10557), .Z(WX10556) ) ;
OR2     gate11357  (.A(WX10570), .B(WX10569), .Z(WX10572) ) ;
AND2    gate11358  (.A(WX10572), .B(WX11347), .Z(WX10561) ) ;
OR2     gate11359  (.A(WX10566), .B(WX10565), .Z(WX10568) ) ;
AND2    gate11360  (.A(WX10568), .B(WX10563), .Z(WX10562) ) ;
AND2    gate11361  (.A(CRC_OUT_1_18), .B(WX11348), .Z(WX10565) ) ;
AND2    gate11362  (.A(DATA_0_18), .B(WX10567), .Z(WX10566) ) ;
AND2    gate11363  (.A(WX10855), .B(WX11348), .Z(WX10569) ) ;
AND2    gate11364  (.A(WX11447), .B(WX10571), .Z(WX10570) ) ;
OR2     gate11365  (.A(WX10584), .B(WX10583), .Z(WX10586) ) ;
AND2    gate11366  (.A(WX10586), .B(WX11347), .Z(WX10575) ) ;
OR2     gate11367  (.A(WX10580), .B(WX10579), .Z(WX10582) ) ;
AND2    gate11368  (.A(WX10582), .B(WX10577), .Z(WX10576) ) ;
AND2    gate11369  (.A(CRC_OUT_1_17), .B(WX11348), .Z(WX10579) ) ;
AND2    gate11370  (.A(DATA_0_17), .B(WX10581), .Z(WX10580) ) ;
AND2    gate11371  (.A(WX10857), .B(WX11348), .Z(WX10583) ) ;
AND2    gate11372  (.A(WX11454), .B(WX10585), .Z(WX10584) ) ;
OR2     gate11373  (.A(WX10598), .B(WX10597), .Z(WX10600) ) ;
AND2    gate11374  (.A(WX10600), .B(WX11347), .Z(WX10589) ) ;
OR2     gate11375  (.A(WX10594), .B(WX10593), .Z(WX10596) ) ;
AND2    gate11376  (.A(WX10596), .B(WX10591), .Z(WX10590) ) ;
AND2    gate11377  (.A(CRC_OUT_1_16), .B(WX11348), .Z(WX10593) ) ;
AND2    gate11378  (.A(DATA_0_16), .B(WX10595), .Z(WX10594) ) ;
AND2    gate11379  (.A(WX10859), .B(WX11348), .Z(WX10597) ) ;
AND2    gate11380  (.A(WX11461), .B(WX10599), .Z(WX10598) ) ;
OR2     gate11381  (.A(WX10612), .B(WX10611), .Z(WX10614) ) ;
AND2    gate11382  (.A(WX10614), .B(WX11347), .Z(WX10603) ) ;
OR2     gate11383  (.A(WX10608), .B(WX10607), .Z(WX10610) ) ;
AND2    gate11384  (.A(WX10610), .B(WX10605), .Z(WX10604) ) ;
AND2    gate11385  (.A(CRC_OUT_1_15), .B(WX11348), .Z(WX10607) ) ;
AND2    gate11386  (.A(DATA_0_15), .B(WX10609), .Z(WX10608) ) ;
AND2    gate11387  (.A(WX10861), .B(WX11348), .Z(WX10611) ) ;
AND2    gate11388  (.A(WX11468), .B(WX10613), .Z(WX10612) ) ;
OR2     gate11389  (.A(WX10626), .B(WX10625), .Z(WX10628) ) ;
AND2    gate11390  (.A(WX10628), .B(WX11347), .Z(WX10617) ) ;
OR2     gate11391  (.A(WX10622), .B(WX10621), .Z(WX10624) ) ;
AND2    gate11392  (.A(WX10624), .B(WX10619), .Z(WX10618) ) ;
AND2    gate11393  (.A(CRC_OUT_1_14), .B(WX11348), .Z(WX10621) ) ;
AND2    gate11394  (.A(DATA_0_14), .B(WX10623), .Z(WX10622) ) ;
AND2    gate11395  (.A(WX10863), .B(WX11348), .Z(WX10625) ) ;
AND2    gate11396  (.A(WX11475), .B(WX10627), .Z(WX10626) ) ;
OR2     gate11397  (.A(WX10640), .B(WX10639), .Z(WX10642) ) ;
AND2    gate11398  (.A(WX10642), .B(WX11347), .Z(WX10631) ) ;
OR2     gate11399  (.A(WX10636), .B(WX10635), .Z(WX10638) ) ;
AND2    gate11400  (.A(WX10638), .B(WX10633), .Z(WX10632) ) ;
AND2    gate11401  (.A(CRC_OUT_1_13), .B(WX11348), .Z(WX10635) ) ;
AND2    gate11402  (.A(DATA_0_13), .B(WX10637), .Z(WX10636) ) ;
AND2    gate11403  (.A(WX10865), .B(WX11348), .Z(WX10639) ) ;
AND2    gate11404  (.A(WX11482), .B(WX10641), .Z(WX10640) ) ;
OR2     gate11405  (.A(WX10654), .B(WX10653), .Z(WX10656) ) ;
AND2    gate11406  (.A(WX10656), .B(WX11347), .Z(WX10645) ) ;
OR2     gate11407  (.A(WX10650), .B(WX10649), .Z(WX10652) ) ;
AND2    gate11408  (.A(WX10652), .B(WX10647), .Z(WX10646) ) ;
AND2    gate11409  (.A(CRC_OUT_1_12), .B(WX11348), .Z(WX10649) ) ;
AND2    gate11410  (.A(DATA_0_12), .B(WX10651), .Z(WX10650) ) ;
AND2    gate11411  (.A(WX10867), .B(WX11348), .Z(WX10653) ) ;
AND2    gate11412  (.A(WX11489), .B(WX10655), .Z(WX10654) ) ;
OR2     gate11413  (.A(WX10668), .B(WX10667), .Z(WX10670) ) ;
AND2    gate11414  (.A(WX10670), .B(WX11347), .Z(WX10659) ) ;
OR2     gate11415  (.A(WX10664), .B(WX10663), .Z(WX10666) ) ;
AND2    gate11416  (.A(WX10666), .B(WX10661), .Z(WX10660) ) ;
AND2    gate11417  (.A(CRC_OUT_1_11), .B(WX11348), .Z(WX10663) ) ;
AND2    gate11418  (.A(DATA_0_11), .B(WX10665), .Z(WX10664) ) ;
AND2    gate11419  (.A(WX10869), .B(WX11348), .Z(WX10667) ) ;
AND2    gate11420  (.A(WX11496), .B(WX10669), .Z(WX10668) ) ;
OR2     gate11421  (.A(WX10682), .B(WX10681), .Z(WX10684) ) ;
AND2    gate11422  (.A(WX10684), .B(WX11347), .Z(WX10673) ) ;
OR2     gate11423  (.A(WX10678), .B(WX10677), .Z(WX10680) ) ;
AND2    gate11424  (.A(WX10680), .B(WX10675), .Z(WX10674) ) ;
AND2    gate11425  (.A(CRC_OUT_1_10), .B(WX11348), .Z(WX10677) ) ;
AND2    gate11426  (.A(DATA_0_10), .B(WX10679), .Z(WX10678) ) ;
AND2    gate11427  (.A(WX10871), .B(WX11348), .Z(WX10681) ) ;
AND2    gate11428  (.A(WX11503), .B(WX10683), .Z(WX10682) ) ;
OR2     gate11429  (.A(WX10696), .B(WX10695), .Z(WX10698) ) ;
AND2    gate11430  (.A(WX10698), .B(WX11347), .Z(WX10687) ) ;
OR2     gate11431  (.A(WX10692), .B(WX10691), .Z(WX10694) ) ;
AND2    gate11432  (.A(WX10694), .B(WX10689), .Z(WX10688) ) ;
AND2    gate11433  (.A(CRC_OUT_1_9), .B(WX11348), .Z(WX10691) ) ;
AND2    gate11434  (.A(DATA_0_9), .B(WX10693), .Z(WX10692) ) ;
AND2    gate11435  (.A(WX10873), .B(WX11348), .Z(WX10695) ) ;
AND2    gate11436  (.A(WX11510), .B(WX10697), .Z(WX10696) ) ;
OR2     gate11437  (.A(WX10710), .B(WX10709), .Z(WX10712) ) ;
AND2    gate11438  (.A(WX10712), .B(WX11347), .Z(WX10701) ) ;
OR2     gate11439  (.A(WX10706), .B(WX10705), .Z(WX10708) ) ;
AND2    gate11440  (.A(WX10708), .B(WX10703), .Z(WX10702) ) ;
AND2    gate11441  (.A(CRC_OUT_1_8), .B(WX11348), .Z(WX10705) ) ;
AND2    gate11442  (.A(DATA_0_8), .B(WX10707), .Z(WX10706) ) ;
AND2    gate11443  (.A(WX10875), .B(WX11348), .Z(WX10709) ) ;
AND2    gate11444  (.A(WX11517), .B(WX10711), .Z(WX10710) ) ;
OR2     gate11445  (.A(WX10724), .B(WX10723), .Z(WX10726) ) ;
AND2    gate11446  (.A(WX10726), .B(WX11347), .Z(WX10715) ) ;
OR2     gate11447  (.A(WX10720), .B(WX10719), .Z(WX10722) ) ;
AND2    gate11448  (.A(WX10722), .B(WX10717), .Z(WX10716) ) ;
AND2    gate11449  (.A(CRC_OUT_1_7), .B(WX11348), .Z(WX10719) ) ;
AND2    gate11450  (.A(DATA_0_7), .B(WX10721), .Z(WX10720) ) ;
AND2    gate11451  (.A(WX10877), .B(WX11348), .Z(WX10723) ) ;
AND2    gate11452  (.A(WX11524), .B(WX10725), .Z(WX10724) ) ;
OR2     gate11453  (.A(WX10738), .B(WX10737), .Z(WX10740) ) ;
AND2    gate11454  (.A(WX10740), .B(WX11347), .Z(WX10729) ) ;
OR2     gate11455  (.A(WX10734), .B(WX10733), .Z(WX10736) ) ;
AND2    gate11456  (.A(WX10736), .B(WX10731), .Z(WX10730) ) ;
AND2    gate11457  (.A(CRC_OUT_1_6), .B(WX11348), .Z(WX10733) ) ;
AND2    gate11458  (.A(DATA_0_6), .B(WX10735), .Z(WX10734) ) ;
AND2    gate11459  (.A(WX10879), .B(WX11348), .Z(WX10737) ) ;
AND2    gate11460  (.A(WX11531), .B(WX10739), .Z(WX10738) ) ;
OR2     gate11461  (.A(WX10752), .B(WX10751), .Z(WX10754) ) ;
AND2    gate11462  (.A(WX10754), .B(WX11347), .Z(WX10743) ) ;
OR2     gate11463  (.A(WX10748), .B(WX10747), .Z(WX10750) ) ;
AND2    gate11464  (.A(WX10750), .B(WX10745), .Z(WX10744) ) ;
AND2    gate11465  (.A(CRC_OUT_1_5), .B(WX11348), .Z(WX10747) ) ;
AND2    gate11466  (.A(DATA_0_5), .B(WX10749), .Z(WX10748) ) ;
AND2    gate11467  (.A(WX10881), .B(WX11348), .Z(WX10751) ) ;
AND2    gate11468  (.A(WX11538), .B(WX10753), .Z(WX10752) ) ;
OR2     gate11469  (.A(WX10766), .B(WX10765), .Z(WX10768) ) ;
AND2    gate11470  (.A(WX10768), .B(WX11347), .Z(WX10757) ) ;
OR2     gate11471  (.A(WX10762), .B(WX10761), .Z(WX10764) ) ;
AND2    gate11472  (.A(WX10764), .B(WX10759), .Z(WX10758) ) ;
AND2    gate11473  (.A(CRC_OUT_1_4), .B(WX11348), .Z(WX10761) ) ;
AND2    gate11474  (.A(DATA_0_4), .B(WX10763), .Z(WX10762) ) ;
AND2    gate11475  (.A(WX10883), .B(WX11348), .Z(WX10765) ) ;
AND2    gate11476  (.A(WX11545), .B(WX10767), .Z(WX10766) ) ;
OR2     gate11477  (.A(WX10780), .B(WX10779), .Z(WX10782) ) ;
AND2    gate11478  (.A(WX10782), .B(WX11347), .Z(WX10771) ) ;
OR2     gate11479  (.A(WX10776), .B(WX10775), .Z(WX10778) ) ;
AND2    gate11480  (.A(WX10778), .B(WX10773), .Z(WX10772) ) ;
AND2    gate11481  (.A(CRC_OUT_1_3), .B(WX11348), .Z(WX10775) ) ;
AND2    gate11482  (.A(DATA_0_3), .B(WX10777), .Z(WX10776) ) ;
AND2    gate11483  (.A(WX10885), .B(WX11348), .Z(WX10779) ) ;
AND2    gate11484  (.A(WX11552), .B(WX10781), .Z(WX10780) ) ;
OR2     gate11485  (.A(WX10794), .B(WX10793), .Z(WX10796) ) ;
AND2    gate11486  (.A(WX10796), .B(WX11347), .Z(WX10785) ) ;
OR2     gate11487  (.A(WX10790), .B(WX10789), .Z(WX10792) ) ;
AND2    gate11488  (.A(WX10792), .B(WX10787), .Z(WX10786) ) ;
AND2    gate11489  (.A(CRC_OUT_1_2), .B(WX11348), .Z(WX10789) ) ;
AND2    gate11490  (.A(DATA_0_2), .B(WX10791), .Z(WX10790) ) ;
AND2    gate11491  (.A(WX10887), .B(WX11348), .Z(WX10793) ) ;
AND2    gate11492  (.A(WX11559), .B(WX10795), .Z(WX10794) ) ;
OR2     gate11493  (.A(WX10808), .B(WX10807), .Z(WX10810) ) ;
AND2    gate11494  (.A(WX10810), .B(WX11347), .Z(WX10799) ) ;
OR2     gate11495  (.A(WX10804), .B(WX10803), .Z(WX10806) ) ;
AND2    gate11496  (.A(WX10806), .B(WX10801), .Z(WX10800) ) ;
AND2    gate11497  (.A(CRC_OUT_1_1), .B(WX11348), .Z(WX10803) ) ;
AND2    gate11498  (.A(DATA_0_1), .B(WX10805), .Z(WX10804) ) ;
AND2    gate11499  (.A(WX10889), .B(WX11348), .Z(WX10807) ) ;
AND2    gate11500  (.A(WX11566), .B(WX10809), .Z(WX10808) ) ;
OR2     gate11501  (.A(WX10822), .B(WX10821), .Z(WX10824) ) ;
AND2    gate11502  (.A(WX10824), .B(WX11347), .Z(WX10813) ) ;
OR2     gate11503  (.A(WX10818), .B(WX10817), .Z(WX10820) ) ;
AND2    gate11504  (.A(WX10820), .B(WX10815), .Z(WX10814) ) ;
AND2    gate11505  (.A(CRC_OUT_1_0), .B(WX11348), .Z(WX10817) ) ;
AND2    gate11506  (.A(DATA_0_0), .B(WX10819), .Z(WX10818) ) ;
AND2    gate11507  (.A(WX10891), .B(WX11348), .Z(WX10821) ) ;
AND2    gate11508  (.A(WX11573), .B(WX10823), .Z(WX10822) ) ;
NAND2   gate11509  (.A(II35093), .B(II35094), .Z(WX11350) ) ;
AND2    gate11510  (.A(WX11350), .B(WX11349), .Z(WX11351) ) ;
AND2    gate11511  (.A(WX10924), .B(WX11353), .Z(WX11352) ) ;
NAND2   gate11512  (.A(II35106), .B(II35107), .Z(WX11357) ) ;
AND2    gate11513  (.A(WX11357), .B(WX11349), .Z(WX11358) ) ;
AND2    gate11514  (.A(WX10925), .B(WX11360), .Z(WX11359) ) ;
NAND2   gate11515  (.A(II35119), .B(II35120), .Z(WX11364) ) ;
AND2    gate11516  (.A(WX11364), .B(WX11349), .Z(WX11365) ) ;
AND2    gate11517  (.A(WX10926), .B(WX11367), .Z(WX11366) ) ;
NAND2   gate11518  (.A(II35132), .B(II35133), .Z(WX11371) ) ;
AND2    gate11519  (.A(WX11371), .B(WX11349), .Z(WX11372) ) ;
AND2    gate11520  (.A(WX10927), .B(WX11374), .Z(WX11373) ) ;
NAND2   gate11521  (.A(II35145), .B(II35146), .Z(WX11378) ) ;
AND2    gate11522  (.A(WX11378), .B(WX11349), .Z(WX11379) ) ;
AND2    gate11523  (.A(WX10928), .B(WX11381), .Z(WX11380) ) ;
NAND2   gate11524  (.A(II35158), .B(II35159), .Z(WX11385) ) ;
AND2    gate11525  (.A(WX11385), .B(WX11349), .Z(WX11386) ) ;
AND2    gate11526  (.A(WX10929), .B(WX11388), .Z(WX11387) ) ;
NAND2   gate11527  (.A(II35171), .B(II35172), .Z(WX11392) ) ;
AND2    gate11528  (.A(WX11392), .B(WX11349), .Z(WX11393) ) ;
AND2    gate11529  (.A(WX10930), .B(WX11395), .Z(WX11394) ) ;
NAND2   gate11530  (.A(II35184), .B(II35185), .Z(WX11399) ) ;
AND2    gate11531  (.A(WX11399), .B(WX11349), .Z(WX11400) ) ;
AND2    gate11532  (.A(WX10931), .B(WX11402), .Z(WX11401) ) ;
NAND2   gate11533  (.A(II35197), .B(II35198), .Z(WX11406) ) ;
AND2    gate11534  (.A(WX11406), .B(WX11349), .Z(WX11407) ) ;
AND2    gate11535  (.A(WX10932), .B(WX11409), .Z(WX11408) ) ;
NAND2   gate11536  (.A(II35210), .B(II35211), .Z(WX11413) ) ;
AND2    gate11537  (.A(WX11413), .B(WX11349), .Z(WX11414) ) ;
AND2    gate11538  (.A(WX10933), .B(WX11416), .Z(WX11415) ) ;
NAND2   gate11539  (.A(II35223), .B(II35224), .Z(WX11420) ) ;
AND2    gate11540  (.A(WX11420), .B(WX11349), .Z(WX11421) ) ;
AND2    gate11541  (.A(WX10934), .B(WX11423), .Z(WX11422) ) ;
NAND2   gate11542  (.A(II35236), .B(II35237), .Z(WX11427) ) ;
AND2    gate11543  (.A(WX11427), .B(WX11349), .Z(WX11428) ) ;
AND2    gate11544  (.A(WX10935), .B(WX11430), .Z(WX11429) ) ;
NAND2   gate11545  (.A(II35249), .B(II35250), .Z(WX11434) ) ;
AND2    gate11546  (.A(WX11434), .B(WX11349), .Z(WX11435) ) ;
AND2    gate11547  (.A(WX10936), .B(WX11437), .Z(WX11436) ) ;
NAND2   gate11548  (.A(II35262), .B(II35263), .Z(WX11441) ) ;
AND2    gate11549  (.A(WX11441), .B(WX11349), .Z(WX11442) ) ;
AND2    gate11550  (.A(WX10937), .B(WX11444), .Z(WX11443) ) ;
NAND2   gate11551  (.A(II35275), .B(II35276), .Z(WX11448) ) ;
AND2    gate11552  (.A(WX11448), .B(WX11349), .Z(WX11449) ) ;
AND2    gate11553  (.A(WX10938), .B(WX11451), .Z(WX11450) ) ;
NAND2   gate11554  (.A(II35288), .B(II35289), .Z(WX11455) ) ;
AND2    gate11555  (.A(WX11455), .B(WX11349), .Z(WX11456) ) ;
AND2    gate11556  (.A(WX10939), .B(WX11458), .Z(WX11457) ) ;
NAND2   gate11557  (.A(II35301), .B(II35302), .Z(WX11462) ) ;
AND2    gate11558  (.A(WX11462), .B(WX11349), .Z(WX11463) ) ;
AND2    gate11559  (.A(WX10940), .B(WX11465), .Z(WX11464) ) ;
NAND2   gate11560  (.A(II35314), .B(II35315), .Z(WX11469) ) ;
AND2    gate11561  (.A(WX11469), .B(WX11349), .Z(WX11470) ) ;
AND2    gate11562  (.A(WX10941), .B(WX11472), .Z(WX11471) ) ;
NAND2   gate11563  (.A(II35327), .B(II35328), .Z(WX11476) ) ;
AND2    gate11564  (.A(WX11476), .B(WX11349), .Z(WX11477) ) ;
AND2    gate11565  (.A(WX10942), .B(WX11479), .Z(WX11478) ) ;
NAND2   gate11566  (.A(II35340), .B(II35341), .Z(WX11483) ) ;
AND2    gate11567  (.A(WX11483), .B(WX11349), .Z(WX11484) ) ;
AND2    gate11568  (.A(WX10943), .B(WX11486), .Z(WX11485) ) ;
NAND2   gate11569  (.A(II35353), .B(II35354), .Z(WX11490) ) ;
AND2    gate11570  (.A(WX11490), .B(WX11349), .Z(WX11491) ) ;
AND2    gate11571  (.A(WX10944), .B(WX11493), .Z(WX11492) ) ;
NAND2   gate11572  (.A(II35366), .B(II35367), .Z(WX11497) ) ;
AND2    gate11573  (.A(WX11497), .B(WX11349), .Z(WX11498) ) ;
AND2    gate11574  (.A(WX10945), .B(WX11500), .Z(WX11499) ) ;
NAND2   gate11575  (.A(II35379), .B(II35380), .Z(WX11504) ) ;
AND2    gate11576  (.A(WX11504), .B(WX11349), .Z(WX11505) ) ;
AND2    gate11577  (.A(WX10946), .B(WX11507), .Z(WX11506) ) ;
NAND2   gate11578  (.A(II35392), .B(II35393), .Z(WX11511) ) ;
AND2    gate11579  (.A(WX11511), .B(WX11349), .Z(WX11512) ) ;
AND2    gate11580  (.A(WX10947), .B(WX11514), .Z(WX11513) ) ;
NAND2   gate11581  (.A(II35405), .B(II35406), .Z(WX11518) ) ;
AND2    gate11582  (.A(WX11518), .B(WX11349), .Z(WX11519) ) ;
AND2    gate11583  (.A(WX10948), .B(WX11521), .Z(WX11520) ) ;
NAND2   gate11584  (.A(II35418), .B(II35419), .Z(WX11525) ) ;
AND2    gate11585  (.A(WX11525), .B(WX11349), .Z(WX11526) ) ;
AND2    gate11586  (.A(WX10949), .B(WX11528), .Z(WX11527) ) ;
NAND2   gate11587  (.A(II35431), .B(II35432), .Z(WX11532) ) ;
AND2    gate11588  (.A(WX11532), .B(WX11349), .Z(WX11533) ) ;
AND2    gate11589  (.A(WX10950), .B(WX11535), .Z(WX11534) ) ;
NAND2   gate11590  (.A(II35444), .B(II35445), .Z(WX11539) ) ;
AND2    gate11591  (.A(WX11539), .B(WX11349), .Z(WX11540) ) ;
AND2    gate11592  (.A(WX10951), .B(WX11542), .Z(WX11541) ) ;
NAND2   gate11593  (.A(II35457), .B(II35458), .Z(WX11546) ) ;
AND2    gate11594  (.A(WX11546), .B(WX11349), .Z(WX11547) ) ;
AND2    gate11595  (.A(WX10952), .B(WX11549), .Z(WX11548) ) ;
NAND2   gate11596  (.A(II35470), .B(II35471), .Z(WX11553) ) ;
AND2    gate11597  (.A(WX11553), .B(WX11349), .Z(WX11554) ) ;
AND2    gate11598  (.A(WX10953), .B(WX11556), .Z(WX11555) ) ;
NAND2   gate11599  (.A(II35483), .B(II35484), .Z(WX11560) ) ;
AND2    gate11600  (.A(WX11560), .B(WX11349), .Z(WX11561) ) ;
AND2    gate11601  (.A(WX10954), .B(WX11563), .Z(WX11562) ) ;
NAND2   gate11602  (.A(II35496), .B(II35497), .Z(WX11567) ) ;
AND2    gate11603  (.A(WX11567), .B(WX11349), .Z(WX11568) ) ;
AND2    gate11604  (.A(WX10955), .B(WX11570), .Z(WX11569) ) ;
NAND2   gate11605  (.A(II35555), .B(II35556), .Z(WX11578) ) ;
NAND2   gate11606  (.A(II35751), .B(II35752), .Z(WX11606) ) ;
NAND2   gate11607  (.A(II35744), .B(II35745), .Z(WX11605) ) ;
NAND2   gate11608  (.A(II35737), .B(II35738), .Z(WX11604) ) ;
NAND2   gate11609  (.A(II35548), .B(II35549), .Z(WX11577) ) ;
NAND2   gate11610  (.A(II35730), .B(II35731), .Z(WX11603) ) ;
NAND2   gate11611  (.A(II35723), .B(II35724), .Z(WX11602) ) ;
NAND2   gate11612  (.A(II35716), .B(II35717), .Z(WX11601) ) ;
NAND2   gate11613  (.A(II35709), .B(II35710), .Z(WX11600) ) ;
NAND2   gate11614  (.A(II35702), .B(II35703), .Z(WX11599) ) ;
NAND2   gate11615  (.A(II35695), .B(II35696), .Z(WX11598) ) ;
NAND2   gate11616  (.A(II35533), .B(II35534), .Z(WX11576) ) ;
NAND2   gate11617  (.A(II35688), .B(II35689), .Z(WX11597) ) ;
NAND2   gate11618  (.A(II35681), .B(II35682), .Z(WX11596) ) ;
NAND2   gate11619  (.A(II35674), .B(II35675), .Z(WX11595) ) ;
NAND2   gate11620  (.A(II35667), .B(II35668), .Z(WX11594) ) ;
NAND2   gate11621  (.A(II35518), .B(II35519), .Z(WX11575) ) ;
NAND2   gate11622  (.A(II35660), .B(II35661), .Z(WX11593) ) ;
NAND2   gate11623  (.A(II35653), .B(II35654), .Z(WX11592) ) ;
NAND2   gate11624  (.A(II35646), .B(II35647), .Z(WX11591) ) ;
NAND2   gate11625  (.A(II35639), .B(II35640), .Z(WX11590) ) ;
NAND2   gate11626  (.A(II35632), .B(II35633), .Z(WX11589) ) ;
NAND2   gate11627  (.A(II35625), .B(II35626), .Z(WX11588) ) ;
NAND2   gate11628  (.A(II35618), .B(II35619), .Z(WX11587) ) ;
NAND2   gate11629  (.A(II35611), .B(II35612), .Z(WX11586) ) ;
NAND2   gate11630  (.A(II35604), .B(II35605), .Z(WX11585) ) ;
NAND2   gate11631  (.A(II35597), .B(II35598), .Z(WX11584) ) ;
NAND2   gate11632  (.A(II35590), .B(II35591), .Z(WX11583) ) ;
NAND2   gate11633  (.A(II35583), .B(II35584), .Z(WX11582) ) ;
NAND2   gate11634  (.A(II35576), .B(II35577), .Z(WX11581) ) ;
NAND2   gate11635  (.A(II35569), .B(II35570), .Z(WX11580) ) ;
NAND2   gate11636  (.A(II35562), .B(II35563), .Z(WX11579) ) ;
NAND2   gate11637  (.A(WX1001), .B(WX645), .Z(II1988) ) ;
NAND2   gate11638  (.A(WX1001), .B(II1988), .Z(II1989) ) ;
NAND2   gate11639  (.A(WX645), .B(II1988), .Z(II1990) ) ;
NAND2   gate11640  (.A(II1989), .B(II1990), .Z(II1987) ) ;
NAND2   gate11641  (.A(WX709), .B(II1987), .Z(II1995) ) ;
NAND2   gate11642  (.A(WX709), .B(II1995), .Z(II1996) ) ;
NAND2   gate11643  (.A(II1987), .B(II1995), .Z(II1997) ) ;
NAND2   gate11644  (.A(II1996), .B(II1997), .Z(II1986) ) ;
NAND2   gate11645  (.A(WX773), .B(WX837), .Z(II2003) ) ;
NAND2   gate11646  (.A(WX773), .B(II2003), .Z(II2004) ) ;
NAND2   gate11647  (.A(WX837), .B(II2003), .Z(II2005) ) ;
NAND2   gate11648  (.A(II2004), .B(II2005), .Z(II2002) ) ;
NAND2   gate11649  (.A(II1986), .B(II2002), .Z(II2010) ) ;
NAND2   gate11650  (.A(II1986), .B(II2010), .Z(II2011) ) ;
NAND2   gate11651  (.A(II2002), .B(II2010), .Z(II2012) ) ;
NAND2   gate11652  (.A(WX1001), .B(WX647), .Z(II2019) ) ;
NAND2   gate11653  (.A(WX1001), .B(II2019), .Z(II2020) ) ;
NAND2   gate11654  (.A(WX647), .B(II2019), .Z(II2021) ) ;
NAND2   gate11655  (.A(II2020), .B(II2021), .Z(II2018) ) ;
NAND2   gate11656  (.A(WX711), .B(II2018), .Z(II2026) ) ;
NAND2   gate11657  (.A(WX711), .B(II2026), .Z(II2027) ) ;
NAND2   gate11658  (.A(II2018), .B(II2026), .Z(II2028) ) ;
NAND2   gate11659  (.A(II2027), .B(II2028), .Z(II2017) ) ;
NAND2   gate11660  (.A(WX775), .B(WX839), .Z(II2034) ) ;
NAND2   gate11661  (.A(WX775), .B(II2034), .Z(II2035) ) ;
NAND2   gate11662  (.A(WX839), .B(II2034), .Z(II2036) ) ;
NAND2   gate11663  (.A(II2035), .B(II2036), .Z(II2033) ) ;
NAND2   gate11664  (.A(II2017), .B(II2033), .Z(II2041) ) ;
NAND2   gate11665  (.A(II2017), .B(II2041), .Z(II2042) ) ;
NAND2   gate11666  (.A(II2033), .B(II2041), .Z(II2043) ) ;
NAND2   gate11667  (.A(WX1001), .B(WX649), .Z(II2050) ) ;
NAND2   gate11668  (.A(WX1001), .B(II2050), .Z(II2051) ) ;
NAND2   gate11669  (.A(WX649), .B(II2050), .Z(II2052) ) ;
NAND2   gate11670  (.A(II2051), .B(II2052), .Z(II2049) ) ;
NAND2   gate11671  (.A(WX713), .B(II2049), .Z(II2057) ) ;
NAND2   gate11672  (.A(WX713), .B(II2057), .Z(II2058) ) ;
NAND2   gate11673  (.A(II2049), .B(II2057), .Z(II2059) ) ;
NAND2   gate11674  (.A(II2058), .B(II2059), .Z(II2048) ) ;
NAND2   gate11675  (.A(WX777), .B(WX841), .Z(II2065) ) ;
NAND2   gate11676  (.A(WX777), .B(II2065), .Z(II2066) ) ;
NAND2   gate11677  (.A(WX841), .B(II2065), .Z(II2067) ) ;
NAND2   gate11678  (.A(II2066), .B(II2067), .Z(II2064) ) ;
NAND2   gate11679  (.A(II2048), .B(II2064), .Z(II2072) ) ;
NAND2   gate11680  (.A(II2048), .B(II2072), .Z(II2073) ) ;
NAND2   gate11681  (.A(II2064), .B(II2072), .Z(II2074) ) ;
NAND2   gate11682  (.A(WX1001), .B(WX651), .Z(II2081) ) ;
NAND2   gate11683  (.A(WX1001), .B(II2081), .Z(II2082) ) ;
NAND2   gate11684  (.A(WX651), .B(II2081), .Z(II2083) ) ;
NAND2   gate11685  (.A(II2082), .B(II2083), .Z(II2080) ) ;
NAND2   gate11686  (.A(WX715), .B(II2080), .Z(II2088) ) ;
NAND2   gate11687  (.A(WX715), .B(II2088), .Z(II2089) ) ;
NAND2   gate11688  (.A(II2080), .B(II2088), .Z(II2090) ) ;
NAND2   gate11689  (.A(II2089), .B(II2090), .Z(II2079) ) ;
NAND2   gate11690  (.A(WX779), .B(WX843), .Z(II2096) ) ;
NAND2   gate11691  (.A(WX779), .B(II2096), .Z(II2097) ) ;
NAND2   gate11692  (.A(WX843), .B(II2096), .Z(II2098) ) ;
NAND2   gate11693  (.A(II2097), .B(II2098), .Z(II2095) ) ;
NAND2   gate11694  (.A(II2079), .B(II2095), .Z(II2103) ) ;
NAND2   gate11695  (.A(II2079), .B(II2103), .Z(II2104) ) ;
NAND2   gate11696  (.A(II2095), .B(II2103), .Z(II2105) ) ;
NAND2   gate11697  (.A(WX1001), .B(WX653), .Z(II2112) ) ;
NAND2   gate11698  (.A(WX1001), .B(II2112), .Z(II2113) ) ;
NAND2   gate11699  (.A(WX653), .B(II2112), .Z(II2114) ) ;
NAND2   gate11700  (.A(II2113), .B(II2114), .Z(II2111) ) ;
NAND2   gate11701  (.A(WX717), .B(II2111), .Z(II2119) ) ;
NAND2   gate11702  (.A(WX717), .B(II2119), .Z(II2120) ) ;
NAND2   gate11703  (.A(II2111), .B(II2119), .Z(II2121) ) ;
NAND2   gate11704  (.A(II2120), .B(II2121), .Z(II2110) ) ;
NAND2   gate11705  (.A(WX781), .B(WX845), .Z(II2127) ) ;
NAND2   gate11706  (.A(WX781), .B(II2127), .Z(II2128) ) ;
NAND2   gate11707  (.A(WX845), .B(II2127), .Z(II2129) ) ;
NAND2   gate11708  (.A(II2128), .B(II2129), .Z(II2126) ) ;
NAND2   gate11709  (.A(II2110), .B(II2126), .Z(II2134) ) ;
NAND2   gate11710  (.A(II2110), .B(II2134), .Z(II2135) ) ;
NAND2   gate11711  (.A(II2126), .B(II2134), .Z(II2136) ) ;
NAND2   gate11712  (.A(WX1001), .B(WX655), .Z(II2143) ) ;
NAND2   gate11713  (.A(WX1001), .B(II2143), .Z(II2144) ) ;
NAND2   gate11714  (.A(WX655), .B(II2143), .Z(II2145) ) ;
NAND2   gate11715  (.A(II2144), .B(II2145), .Z(II2142) ) ;
NAND2   gate11716  (.A(WX719), .B(II2142), .Z(II2150) ) ;
NAND2   gate11717  (.A(WX719), .B(II2150), .Z(II2151) ) ;
NAND2   gate11718  (.A(II2142), .B(II2150), .Z(II2152) ) ;
NAND2   gate11719  (.A(II2151), .B(II2152), .Z(II2141) ) ;
NAND2   gate11720  (.A(WX783), .B(WX847), .Z(II2158) ) ;
NAND2   gate11721  (.A(WX783), .B(II2158), .Z(II2159) ) ;
NAND2   gate11722  (.A(WX847), .B(II2158), .Z(II2160) ) ;
NAND2   gate11723  (.A(II2159), .B(II2160), .Z(II2157) ) ;
NAND2   gate11724  (.A(II2141), .B(II2157), .Z(II2165) ) ;
NAND2   gate11725  (.A(II2141), .B(II2165), .Z(II2166) ) ;
NAND2   gate11726  (.A(II2157), .B(II2165), .Z(II2167) ) ;
NAND2   gate11727  (.A(WX1001), .B(WX657), .Z(II2174) ) ;
NAND2   gate11728  (.A(WX1001), .B(II2174), .Z(II2175) ) ;
NAND2   gate11729  (.A(WX657), .B(II2174), .Z(II2176) ) ;
NAND2   gate11730  (.A(II2175), .B(II2176), .Z(II2173) ) ;
NAND2   gate11731  (.A(WX721), .B(II2173), .Z(II2181) ) ;
NAND2   gate11732  (.A(WX721), .B(II2181), .Z(II2182) ) ;
NAND2   gate11733  (.A(II2173), .B(II2181), .Z(II2183) ) ;
NAND2   gate11734  (.A(II2182), .B(II2183), .Z(II2172) ) ;
NAND2   gate11735  (.A(WX785), .B(WX849), .Z(II2189) ) ;
NAND2   gate11736  (.A(WX785), .B(II2189), .Z(II2190) ) ;
NAND2   gate11737  (.A(WX849), .B(II2189), .Z(II2191) ) ;
NAND2   gate11738  (.A(II2190), .B(II2191), .Z(II2188) ) ;
NAND2   gate11739  (.A(II2172), .B(II2188), .Z(II2196) ) ;
NAND2   gate11740  (.A(II2172), .B(II2196), .Z(II2197) ) ;
NAND2   gate11741  (.A(II2188), .B(II2196), .Z(II2198) ) ;
NAND2   gate11742  (.A(WX1001), .B(WX659), .Z(II2205) ) ;
NAND2   gate11743  (.A(WX1001), .B(II2205), .Z(II2206) ) ;
NAND2   gate11744  (.A(WX659), .B(II2205), .Z(II2207) ) ;
NAND2   gate11745  (.A(II2206), .B(II2207), .Z(II2204) ) ;
NAND2   gate11746  (.A(WX723), .B(II2204), .Z(II2212) ) ;
NAND2   gate11747  (.A(WX723), .B(II2212), .Z(II2213) ) ;
NAND2   gate11748  (.A(II2204), .B(II2212), .Z(II2214) ) ;
NAND2   gate11749  (.A(II2213), .B(II2214), .Z(II2203) ) ;
NAND2   gate11750  (.A(WX787), .B(WX851), .Z(II2220) ) ;
NAND2   gate11751  (.A(WX787), .B(II2220), .Z(II2221) ) ;
NAND2   gate11752  (.A(WX851), .B(II2220), .Z(II2222) ) ;
NAND2   gate11753  (.A(II2221), .B(II2222), .Z(II2219) ) ;
NAND2   gate11754  (.A(II2203), .B(II2219), .Z(II2227) ) ;
NAND2   gate11755  (.A(II2203), .B(II2227), .Z(II2228) ) ;
NAND2   gate11756  (.A(II2219), .B(II2227), .Z(II2229) ) ;
NAND2   gate11757  (.A(WX1001), .B(WX661), .Z(II2236) ) ;
NAND2   gate11758  (.A(WX1001), .B(II2236), .Z(II2237) ) ;
NAND2   gate11759  (.A(WX661), .B(II2236), .Z(II2238) ) ;
NAND2   gate11760  (.A(II2237), .B(II2238), .Z(II2235) ) ;
NAND2   gate11761  (.A(WX725), .B(II2235), .Z(II2243) ) ;
NAND2   gate11762  (.A(WX725), .B(II2243), .Z(II2244) ) ;
NAND2   gate11763  (.A(II2235), .B(II2243), .Z(II2245) ) ;
NAND2   gate11764  (.A(II2244), .B(II2245), .Z(II2234) ) ;
NAND2   gate11765  (.A(WX789), .B(WX853), .Z(II2251) ) ;
NAND2   gate11766  (.A(WX789), .B(II2251), .Z(II2252) ) ;
NAND2   gate11767  (.A(WX853), .B(II2251), .Z(II2253) ) ;
NAND2   gate11768  (.A(II2252), .B(II2253), .Z(II2250) ) ;
NAND2   gate11769  (.A(II2234), .B(II2250), .Z(II2258) ) ;
NAND2   gate11770  (.A(II2234), .B(II2258), .Z(II2259) ) ;
NAND2   gate11771  (.A(II2250), .B(II2258), .Z(II2260) ) ;
NAND2   gate11772  (.A(WX1001), .B(WX663), .Z(II2267) ) ;
NAND2   gate11773  (.A(WX1001), .B(II2267), .Z(II2268) ) ;
NAND2   gate11774  (.A(WX663), .B(II2267), .Z(II2269) ) ;
NAND2   gate11775  (.A(II2268), .B(II2269), .Z(II2266) ) ;
NAND2   gate11776  (.A(WX727), .B(II2266), .Z(II2274) ) ;
NAND2   gate11777  (.A(WX727), .B(II2274), .Z(II2275) ) ;
NAND2   gate11778  (.A(II2266), .B(II2274), .Z(II2276) ) ;
NAND2   gate11779  (.A(II2275), .B(II2276), .Z(II2265) ) ;
NAND2   gate11780  (.A(WX791), .B(WX855), .Z(II2282) ) ;
NAND2   gate11781  (.A(WX791), .B(II2282), .Z(II2283) ) ;
NAND2   gate11782  (.A(WX855), .B(II2282), .Z(II2284) ) ;
NAND2   gate11783  (.A(II2283), .B(II2284), .Z(II2281) ) ;
NAND2   gate11784  (.A(II2265), .B(II2281), .Z(II2289) ) ;
NAND2   gate11785  (.A(II2265), .B(II2289), .Z(II2290) ) ;
NAND2   gate11786  (.A(II2281), .B(II2289), .Z(II2291) ) ;
NAND2   gate11787  (.A(WX1001), .B(WX665), .Z(II2298) ) ;
NAND2   gate11788  (.A(WX1001), .B(II2298), .Z(II2299) ) ;
NAND2   gate11789  (.A(WX665), .B(II2298), .Z(II2300) ) ;
NAND2   gate11790  (.A(II2299), .B(II2300), .Z(II2297) ) ;
NAND2   gate11791  (.A(WX729), .B(II2297), .Z(II2305) ) ;
NAND2   gate11792  (.A(WX729), .B(II2305), .Z(II2306) ) ;
NAND2   gate11793  (.A(II2297), .B(II2305), .Z(II2307) ) ;
NAND2   gate11794  (.A(II2306), .B(II2307), .Z(II2296) ) ;
NAND2   gate11795  (.A(WX793), .B(WX857), .Z(II2313) ) ;
NAND2   gate11796  (.A(WX793), .B(II2313), .Z(II2314) ) ;
NAND2   gate11797  (.A(WX857), .B(II2313), .Z(II2315) ) ;
NAND2   gate11798  (.A(II2314), .B(II2315), .Z(II2312) ) ;
NAND2   gate11799  (.A(II2296), .B(II2312), .Z(II2320) ) ;
NAND2   gate11800  (.A(II2296), .B(II2320), .Z(II2321) ) ;
NAND2   gate11801  (.A(II2312), .B(II2320), .Z(II2322) ) ;
NAND2   gate11802  (.A(WX1001), .B(WX667), .Z(II2329) ) ;
NAND2   gate11803  (.A(WX1001), .B(II2329), .Z(II2330) ) ;
NAND2   gate11804  (.A(WX667), .B(II2329), .Z(II2331) ) ;
NAND2   gate11805  (.A(II2330), .B(II2331), .Z(II2328) ) ;
NAND2   gate11806  (.A(WX731), .B(II2328), .Z(II2336) ) ;
NAND2   gate11807  (.A(WX731), .B(II2336), .Z(II2337) ) ;
NAND2   gate11808  (.A(II2328), .B(II2336), .Z(II2338) ) ;
NAND2   gate11809  (.A(II2337), .B(II2338), .Z(II2327) ) ;
NAND2   gate11810  (.A(WX795), .B(WX859), .Z(II2344) ) ;
NAND2   gate11811  (.A(WX795), .B(II2344), .Z(II2345) ) ;
NAND2   gate11812  (.A(WX859), .B(II2344), .Z(II2346) ) ;
NAND2   gate11813  (.A(II2345), .B(II2346), .Z(II2343) ) ;
NAND2   gate11814  (.A(II2327), .B(II2343), .Z(II2351) ) ;
NAND2   gate11815  (.A(II2327), .B(II2351), .Z(II2352) ) ;
NAND2   gate11816  (.A(II2343), .B(II2351), .Z(II2353) ) ;
NAND2   gate11817  (.A(WX1001), .B(WX669), .Z(II2360) ) ;
NAND2   gate11818  (.A(WX1001), .B(II2360), .Z(II2361) ) ;
NAND2   gate11819  (.A(WX669), .B(II2360), .Z(II2362) ) ;
NAND2   gate11820  (.A(II2361), .B(II2362), .Z(II2359) ) ;
NAND2   gate11821  (.A(WX733), .B(II2359), .Z(II2367) ) ;
NAND2   gate11822  (.A(WX733), .B(II2367), .Z(II2368) ) ;
NAND2   gate11823  (.A(II2359), .B(II2367), .Z(II2369) ) ;
NAND2   gate11824  (.A(II2368), .B(II2369), .Z(II2358) ) ;
NAND2   gate11825  (.A(WX797), .B(WX861), .Z(II2375) ) ;
NAND2   gate11826  (.A(WX797), .B(II2375), .Z(II2376) ) ;
NAND2   gate11827  (.A(WX861), .B(II2375), .Z(II2377) ) ;
NAND2   gate11828  (.A(II2376), .B(II2377), .Z(II2374) ) ;
NAND2   gate11829  (.A(II2358), .B(II2374), .Z(II2382) ) ;
NAND2   gate11830  (.A(II2358), .B(II2382), .Z(II2383) ) ;
NAND2   gate11831  (.A(II2374), .B(II2382), .Z(II2384) ) ;
NAND2   gate11832  (.A(WX1001), .B(WX671), .Z(II2391) ) ;
NAND2   gate11833  (.A(WX1001), .B(II2391), .Z(II2392) ) ;
NAND2   gate11834  (.A(WX671), .B(II2391), .Z(II2393) ) ;
NAND2   gate11835  (.A(II2392), .B(II2393), .Z(II2390) ) ;
NAND2   gate11836  (.A(WX735), .B(II2390), .Z(II2398) ) ;
NAND2   gate11837  (.A(WX735), .B(II2398), .Z(II2399) ) ;
NAND2   gate11838  (.A(II2390), .B(II2398), .Z(II2400) ) ;
NAND2   gate11839  (.A(II2399), .B(II2400), .Z(II2389) ) ;
NAND2   gate11840  (.A(WX799), .B(WX863), .Z(II2406) ) ;
NAND2   gate11841  (.A(WX799), .B(II2406), .Z(II2407) ) ;
NAND2   gate11842  (.A(WX863), .B(II2406), .Z(II2408) ) ;
NAND2   gate11843  (.A(II2407), .B(II2408), .Z(II2405) ) ;
NAND2   gate11844  (.A(II2389), .B(II2405), .Z(II2413) ) ;
NAND2   gate11845  (.A(II2389), .B(II2413), .Z(II2414) ) ;
NAND2   gate11846  (.A(II2405), .B(II2413), .Z(II2415) ) ;
NAND2   gate11847  (.A(WX1001), .B(WX673), .Z(II2422) ) ;
NAND2   gate11848  (.A(WX1001), .B(II2422), .Z(II2423) ) ;
NAND2   gate11849  (.A(WX673), .B(II2422), .Z(II2424) ) ;
NAND2   gate11850  (.A(II2423), .B(II2424), .Z(II2421) ) ;
NAND2   gate11851  (.A(WX737), .B(II2421), .Z(II2429) ) ;
NAND2   gate11852  (.A(WX737), .B(II2429), .Z(II2430) ) ;
NAND2   gate11853  (.A(II2421), .B(II2429), .Z(II2431) ) ;
NAND2   gate11854  (.A(II2430), .B(II2431), .Z(II2420) ) ;
NAND2   gate11855  (.A(WX801), .B(WX865), .Z(II2437) ) ;
NAND2   gate11856  (.A(WX801), .B(II2437), .Z(II2438) ) ;
NAND2   gate11857  (.A(WX865), .B(II2437), .Z(II2439) ) ;
NAND2   gate11858  (.A(II2438), .B(II2439), .Z(II2436) ) ;
NAND2   gate11859  (.A(II2420), .B(II2436), .Z(II2444) ) ;
NAND2   gate11860  (.A(II2420), .B(II2444), .Z(II2445) ) ;
NAND2   gate11861  (.A(II2436), .B(II2444), .Z(II2446) ) ;
NAND2   gate11862  (.A(WX1001), .B(WX675), .Z(II2453) ) ;
NAND2   gate11863  (.A(WX1001), .B(II2453), .Z(II2454) ) ;
NAND2   gate11864  (.A(WX675), .B(II2453), .Z(II2455) ) ;
NAND2   gate11865  (.A(II2454), .B(II2455), .Z(II2452) ) ;
NAND2   gate11866  (.A(WX739), .B(II2452), .Z(II2460) ) ;
NAND2   gate11867  (.A(WX739), .B(II2460), .Z(II2461) ) ;
NAND2   gate11868  (.A(II2452), .B(II2460), .Z(II2462) ) ;
NAND2   gate11869  (.A(II2461), .B(II2462), .Z(II2451) ) ;
NAND2   gate11870  (.A(WX803), .B(WX867), .Z(II2468) ) ;
NAND2   gate11871  (.A(WX803), .B(II2468), .Z(II2469) ) ;
NAND2   gate11872  (.A(WX867), .B(II2468), .Z(II2470) ) ;
NAND2   gate11873  (.A(II2469), .B(II2470), .Z(II2467) ) ;
NAND2   gate11874  (.A(II2451), .B(II2467), .Z(II2475) ) ;
NAND2   gate11875  (.A(II2451), .B(II2475), .Z(II2476) ) ;
NAND2   gate11876  (.A(II2467), .B(II2475), .Z(II2477) ) ;
NAND2   gate11877  (.A(WX1002), .B(WX677), .Z(II2484) ) ;
NAND2   gate11878  (.A(WX1002), .B(II2484), .Z(II2485) ) ;
NAND2   gate11879  (.A(WX677), .B(II2484), .Z(II2486) ) ;
NAND2   gate11880  (.A(II2485), .B(II2486), .Z(II2483) ) ;
NAND2   gate11881  (.A(WX741), .B(II2483), .Z(II2491) ) ;
NAND2   gate11882  (.A(WX741), .B(II2491), .Z(II2492) ) ;
NAND2   gate11883  (.A(II2483), .B(II2491), .Z(II2493) ) ;
NAND2   gate11884  (.A(II2492), .B(II2493), .Z(II2482) ) ;
NAND2   gate11885  (.A(WX805), .B(WX869), .Z(II2499) ) ;
NAND2   gate11886  (.A(WX805), .B(II2499), .Z(II2500) ) ;
NAND2   gate11887  (.A(WX869), .B(II2499), .Z(II2501) ) ;
NAND2   gate11888  (.A(II2500), .B(II2501), .Z(II2498) ) ;
NAND2   gate11889  (.A(II2482), .B(II2498), .Z(II2506) ) ;
NAND2   gate11890  (.A(II2482), .B(II2506), .Z(II2507) ) ;
NAND2   gate11891  (.A(II2498), .B(II2506), .Z(II2508) ) ;
NAND2   gate11892  (.A(WX1002), .B(WX679), .Z(II2515) ) ;
NAND2   gate11893  (.A(WX1002), .B(II2515), .Z(II2516) ) ;
NAND2   gate11894  (.A(WX679), .B(II2515), .Z(II2517) ) ;
NAND2   gate11895  (.A(II2516), .B(II2517), .Z(II2514) ) ;
NAND2   gate11896  (.A(WX743), .B(II2514), .Z(II2522) ) ;
NAND2   gate11897  (.A(WX743), .B(II2522), .Z(II2523) ) ;
NAND2   gate11898  (.A(II2514), .B(II2522), .Z(II2524) ) ;
NAND2   gate11899  (.A(II2523), .B(II2524), .Z(II2513) ) ;
NAND2   gate11900  (.A(WX807), .B(WX871), .Z(II2530) ) ;
NAND2   gate11901  (.A(WX807), .B(II2530), .Z(II2531) ) ;
NAND2   gate11902  (.A(WX871), .B(II2530), .Z(II2532) ) ;
NAND2   gate11903  (.A(II2531), .B(II2532), .Z(II2529) ) ;
NAND2   gate11904  (.A(II2513), .B(II2529), .Z(II2537) ) ;
NAND2   gate11905  (.A(II2513), .B(II2537), .Z(II2538) ) ;
NAND2   gate11906  (.A(II2529), .B(II2537), .Z(II2539) ) ;
NAND2   gate11907  (.A(WX1002), .B(WX681), .Z(II2546) ) ;
NAND2   gate11908  (.A(WX1002), .B(II2546), .Z(II2547) ) ;
NAND2   gate11909  (.A(WX681), .B(II2546), .Z(II2548) ) ;
NAND2   gate11910  (.A(II2547), .B(II2548), .Z(II2545) ) ;
NAND2   gate11911  (.A(WX745), .B(II2545), .Z(II2553) ) ;
NAND2   gate11912  (.A(WX745), .B(II2553), .Z(II2554) ) ;
NAND2   gate11913  (.A(II2545), .B(II2553), .Z(II2555) ) ;
NAND2   gate11914  (.A(II2554), .B(II2555), .Z(II2544) ) ;
NAND2   gate11915  (.A(WX809), .B(WX873), .Z(II2561) ) ;
NAND2   gate11916  (.A(WX809), .B(II2561), .Z(II2562) ) ;
NAND2   gate11917  (.A(WX873), .B(II2561), .Z(II2563) ) ;
NAND2   gate11918  (.A(II2562), .B(II2563), .Z(II2560) ) ;
NAND2   gate11919  (.A(II2544), .B(II2560), .Z(II2568) ) ;
NAND2   gate11920  (.A(II2544), .B(II2568), .Z(II2569) ) ;
NAND2   gate11921  (.A(II2560), .B(II2568), .Z(II2570) ) ;
NAND2   gate11922  (.A(WX1002), .B(WX683), .Z(II2577) ) ;
NAND2   gate11923  (.A(WX1002), .B(II2577), .Z(II2578) ) ;
NAND2   gate11924  (.A(WX683), .B(II2577), .Z(II2579) ) ;
NAND2   gate11925  (.A(II2578), .B(II2579), .Z(II2576) ) ;
NAND2   gate11926  (.A(WX747), .B(II2576), .Z(II2584) ) ;
NAND2   gate11927  (.A(WX747), .B(II2584), .Z(II2585) ) ;
NAND2   gate11928  (.A(II2576), .B(II2584), .Z(II2586) ) ;
NAND2   gate11929  (.A(II2585), .B(II2586), .Z(II2575) ) ;
NAND2   gate11930  (.A(WX811), .B(WX875), .Z(II2592) ) ;
NAND2   gate11931  (.A(WX811), .B(II2592), .Z(II2593) ) ;
NAND2   gate11932  (.A(WX875), .B(II2592), .Z(II2594) ) ;
NAND2   gate11933  (.A(II2593), .B(II2594), .Z(II2591) ) ;
NAND2   gate11934  (.A(II2575), .B(II2591), .Z(II2599) ) ;
NAND2   gate11935  (.A(II2575), .B(II2599), .Z(II2600) ) ;
NAND2   gate11936  (.A(II2591), .B(II2599), .Z(II2601) ) ;
NAND2   gate11937  (.A(WX1002), .B(WX685), .Z(II2608) ) ;
NAND2   gate11938  (.A(WX1002), .B(II2608), .Z(II2609) ) ;
NAND2   gate11939  (.A(WX685), .B(II2608), .Z(II2610) ) ;
NAND2   gate11940  (.A(II2609), .B(II2610), .Z(II2607) ) ;
NAND2   gate11941  (.A(WX749), .B(II2607), .Z(II2615) ) ;
NAND2   gate11942  (.A(WX749), .B(II2615), .Z(II2616) ) ;
NAND2   gate11943  (.A(II2607), .B(II2615), .Z(II2617) ) ;
NAND2   gate11944  (.A(II2616), .B(II2617), .Z(II2606) ) ;
NAND2   gate11945  (.A(WX813), .B(WX877), .Z(II2623) ) ;
NAND2   gate11946  (.A(WX813), .B(II2623), .Z(II2624) ) ;
NAND2   gate11947  (.A(WX877), .B(II2623), .Z(II2625) ) ;
NAND2   gate11948  (.A(II2624), .B(II2625), .Z(II2622) ) ;
NAND2   gate11949  (.A(II2606), .B(II2622), .Z(II2630) ) ;
NAND2   gate11950  (.A(II2606), .B(II2630), .Z(II2631) ) ;
NAND2   gate11951  (.A(II2622), .B(II2630), .Z(II2632) ) ;
NAND2   gate11952  (.A(WX1002), .B(WX687), .Z(II2639) ) ;
NAND2   gate11953  (.A(WX1002), .B(II2639), .Z(II2640) ) ;
NAND2   gate11954  (.A(WX687), .B(II2639), .Z(II2641) ) ;
NAND2   gate11955  (.A(II2640), .B(II2641), .Z(II2638) ) ;
NAND2   gate11956  (.A(WX751), .B(II2638), .Z(II2646) ) ;
NAND2   gate11957  (.A(WX751), .B(II2646), .Z(II2647) ) ;
NAND2   gate11958  (.A(II2638), .B(II2646), .Z(II2648) ) ;
NAND2   gate11959  (.A(II2647), .B(II2648), .Z(II2637) ) ;
NAND2   gate11960  (.A(WX815), .B(WX879), .Z(II2654) ) ;
NAND2   gate11961  (.A(WX815), .B(II2654), .Z(II2655) ) ;
NAND2   gate11962  (.A(WX879), .B(II2654), .Z(II2656) ) ;
NAND2   gate11963  (.A(II2655), .B(II2656), .Z(II2653) ) ;
NAND2   gate11964  (.A(II2637), .B(II2653), .Z(II2661) ) ;
NAND2   gate11965  (.A(II2637), .B(II2661), .Z(II2662) ) ;
NAND2   gate11966  (.A(II2653), .B(II2661), .Z(II2663) ) ;
NAND2   gate11967  (.A(WX1002), .B(WX689), .Z(II2670) ) ;
NAND2   gate11968  (.A(WX1002), .B(II2670), .Z(II2671) ) ;
NAND2   gate11969  (.A(WX689), .B(II2670), .Z(II2672) ) ;
NAND2   gate11970  (.A(II2671), .B(II2672), .Z(II2669) ) ;
NAND2   gate11971  (.A(WX753), .B(II2669), .Z(II2677) ) ;
NAND2   gate11972  (.A(WX753), .B(II2677), .Z(II2678) ) ;
NAND2   gate11973  (.A(II2669), .B(II2677), .Z(II2679) ) ;
NAND2   gate11974  (.A(II2678), .B(II2679), .Z(II2668) ) ;
NAND2   gate11975  (.A(WX817), .B(WX881), .Z(II2685) ) ;
NAND2   gate11976  (.A(WX817), .B(II2685), .Z(II2686) ) ;
NAND2   gate11977  (.A(WX881), .B(II2685), .Z(II2687) ) ;
NAND2   gate11978  (.A(II2686), .B(II2687), .Z(II2684) ) ;
NAND2   gate11979  (.A(II2668), .B(II2684), .Z(II2692) ) ;
NAND2   gate11980  (.A(II2668), .B(II2692), .Z(II2693) ) ;
NAND2   gate11981  (.A(II2684), .B(II2692), .Z(II2694) ) ;
NAND2   gate11982  (.A(WX1002), .B(WX691), .Z(II2701) ) ;
NAND2   gate11983  (.A(WX1002), .B(II2701), .Z(II2702) ) ;
NAND2   gate11984  (.A(WX691), .B(II2701), .Z(II2703) ) ;
NAND2   gate11985  (.A(II2702), .B(II2703), .Z(II2700) ) ;
NAND2   gate11986  (.A(WX755), .B(II2700), .Z(II2708) ) ;
NAND2   gate11987  (.A(WX755), .B(II2708), .Z(II2709) ) ;
NAND2   gate11988  (.A(II2700), .B(II2708), .Z(II2710) ) ;
NAND2   gate11989  (.A(II2709), .B(II2710), .Z(II2699) ) ;
NAND2   gate11990  (.A(WX819), .B(WX883), .Z(II2716) ) ;
NAND2   gate11991  (.A(WX819), .B(II2716), .Z(II2717) ) ;
NAND2   gate11992  (.A(WX883), .B(II2716), .Z(II2718) ) ;
NAND2   gate11993  (.A(II2717), .B(II2718), .Z(II2715) ) ;
NAND2   gate11994  (.A(II2699), .B(II2715), .Z(II2723) ) ;
NAND2   gate11995  (.A(II2699), .B(II2723), .Z(II2724) ) ;
NAND2   gate11996  (.A(II2715), .B(II2723), .Z(II2725) ) ;
NAND2   gate11997  (.A(WX1002), .B(WX693), .Z(II2732) ) ;
NAND2   gate11998  (.A(WX1002), .B(II2732), .Z(II2733) ) ;
NAND2   gate11999  (.A(WX693), .B(II2732), .Z(II2734) ) ;
NAND2   gate12000  (.A(II2733), .B(II2734), .Z(II2731) ) ;
NAND2   gate12001  (.A(WX757), .B(II2731), .Z(II2739) ) ;
NAND2   gate12002  (.A(WX757), .B(II2739), .Z(II2740) ) ;
NAND2   gate12003  (.A(II2731), .B(II2739), .Z(II2741) ) ;
NAND2   gate12004  (.A(II2740), .B(II2741), .Z(II2730) ) ;
NAND2   gate12005  (.A(WX821), .B(WX885), .Z(II2747) ) ;
NAND2   gate12006  (.A(WX821), .B(II2747), .Z(II2748) ) ;
NAND2   gate12007  (.A(WX885), .B(II2747), .Z(II2749) ) ;
NAND2   gate12008  (.A(II2748), .B(II2749), .Z(II2746) ) ;
NAND2   gate12009  (.A(II2730), .B(II2746), .Z(II2754) ) ;
NAND2   gate12010  (.A(II2730), .B(II2754), .Z(II2755) ) ;
NAND2   gate12011  (.A(II2746), .B(II2754), .Z(II2756) ) ;
NAND2   gate12012  (.A(WX1002), .B(WX695), .Z(II2763) ) ;
NAND2   gate12013  (.A(WX1002), .B(II2763), .Z(II2764) ) ;
NAND2   gate12014  (.A(WX695), .B(II2763), .Z(II2765) ) ;
NAND2   gate12015  (.A(II2764), .B(II2765), .Z(II2762) ) ;
NAND2   gate12016  (.A(WX759), .B(II2762), .Z(II2770) ) ;
NAND2   gate12017  (.A(WX759), .B(II2770), .Z(II2771) ) ;
NAND2   gate12018  (.A(II2762), .B(II2770), .Z(II2772) ) ;
NAND2   gate12019  (.A(II2771), .B(II2772), .Z(II2761) ) ;
NAND2   gate12020  (.A(WX823), .B(WX887), .Z(II2778) ) ;
NAND2   gate12021  (.A(WX823), .B(II2778), .Z(II2779) ) ;
NAND2   gate12022  (.A(WX887), .B(II2778), .Z(II2780) ) ;
NAND2   gate12023  (.A(II2779), .B(II2780), .Z(II2777) ) ;
NAND2   gate12024  (.A(II2761), .B(II2777), .Z(II2785) ) ;
NAND2   gate12025  (.A(II2761), .B(II2785), .Z(II2786) ) ;
NAND2   gate12026  (.A(II2777), .B(II2785), .Z(II2787) ) ;
NAND2   gate12027  (.A(WX1002), .B(WX697), .Z(II2794) ) ;
NAND2   gate12028  (.A(WX1002), .B(II2794), .Z(II2795) ) ;
NAND2   gate12029  (.A(WX697), .B(II2794), .Z(II2796) ) ;
NAND2   gate12030  (.A(II2795), .B(II2796), .Z(II2793) ) ;
NAND2   gate12031  (.A(WX761), .B(II2793), .Z(II2801) ) ;
NAND2   gate12032  (.A(WX761), .B(II2801), .Z(II2802) ) ;
NAND2   gate12033  (.A(II2793), .B(II2801), .Z(II2803) ) ;
NAND2   gate12034  (.A(II2802), .B(II2803), .Z(II2792) ) ;
NAND2   gate12035  (.A(WX825), .B(WX889), .Z(II2809) ) ;
NAND2   gate12036  (.A(WX825), .B(II2809), .Z(II2810) ) ;
NAND2   gate12037  (.A(WX889), .B(II2809), .Z(II2811) ) ;
NAND2   gate12038  (.A(II2810), .B(II2811), .Z(II2808) ) ;
NAND2   gate12039  (.A(II2792), .B(II2808), .Z(II2816) ) ;
NAND2   gate12040  (.A(II2792), .B(II2816), .Z(II2817) ) ;
NAND2   gate12041  (.A(II2808), .B(II2816), .Z(II2818) ) ;
NAND2   gate12042  (.A(WX1002), .B(WX699), .Z(II2825) ) ;
NAND2   gate12043  (.A(WX1002), .B(II2825), .Z(II2826) ) ;
NAND2   gate12044  (.A(WX699), .B(II2825), .Z(II2827) ) ;
NAND2   gate12045  (.A(II2826), .B(II2827), .Z(II2824) ) ;
NAND2   gate12046  (.A(WX763), .B(II2824), .Z(II2832) ) ;
NAND2   gate12047  (.A(WX763), .B(II2832), .Z(II2833) ) ;
NAND2   gate12048  (.A(II2824), .B(II2832), .Z(II2834) ) ;
NAND2   gate12049  (.A(II2833), .B(II2834), .Z(II2823) ) ;
NAND2   gate12050  (.A(WX827), .B(WX891), .Z(II2840) ) ;
NAND2   gate12051  (.A(WX827), .B(II2840), .Z(II2841) ) ;
NAND2   gate12052  (.A(WX891), .B(II2840), .Z(II2842) ) ;
NAND2   gate12053  (.A(II2841), .B(II2842), .Z(II2839) ) ;
NAND2   gate12054  (.A(II2823), .B(II2839), .Z(II2847) ) ;
NAND2   gate12055  (.A(II2823), .B(II2847), .Z(II2848) ) ;
NAND2   gate12056  (.A(II2839), .B(II2847), .Z(II2849) ) ;
NAND2   gate12057  (.A(WX1002), .B(WX701), .Z(II2856) ) ;
NAND2   gate12058  (.A(WX1002), .B(II2856), .Z(II2857) ) ;
NAND2   gate12059  (.A(WX701), .B(II2856), .Z(II2858) ) ;
NAND2   gate12060  (.A(II2857), .B(II2858), .Z(II2855) ) ;
NAND2   gate12061  (.A(WX765), .B(II2855), .Z(II2863) ) ;
NAND2   gate12062  (.A(WX765), .B(II2863), .Z(II2864) ) ;
NAND2   gate12063  (.A(II2855), .B(II2863), .Z(II2865) ) ;
NAND2   gate12064  (.A(II2864), .B(II2865), .Z(II2854) ) ;
NAND2   gate12065  (.A(WX829), .B(WX893), .Z(II2871) ) ;
NAND2   gate12066  (.A(WX829), .B(II2871), .Z(II2872) ) ;
NAND2   gate12067  (.A(WX893), .B(II2871), .Z(II2873) ) ;
NAND2   gate12068  (.A(II2872), .B(II2873), .Z(II2870) ) ;
NAND2   gate12069  (.A(II2854), .B(II2870), .Z(II2878) ) ;
NAND2   gate12070  (.A(II2854), .B(II2878), .Z(II2879) ) ;
NAND2   gate12071  (.A(II2870), .B(II2878), .Z(II2880) ) ;
NAND2   gate12072  (.A(WX1002), .B(WX703), .Z(II2887) ) ;
NAND2   gate12073  (.A(WX1002), .B(II2887), .Z(II2888) ) ;
NAND2   gate12074  (.A(WX703), .B(II2887), .Z(II2889) ) ;
NAND2   gate12075  (.A(II2888), .B(II2889), .Z(II2886) ) ;
NAND2   gate12076  (.A(WX767), .B(II2886), .Z(II2894) ) ;
NAND2   gate12077  (.A(WX767), .B(II2894), .Z(II2895) ) ;
NAND2   gate12078  (.A(II2886), .B(II2894), .Z(II2896) ) ;
NAND2   gate12079  (.A(II2895), .B(II2896), .Z(II2885) ) ;
NAND2   gate12080  (.A(WX831), .B(WX895), .Z(II2902) ) ;
NAND2   gate12081  (.A(WX831), .B(II2902), .Z(II2903) ) ;
NAND2   gate12082  (.A(WX895), .B(II2902), .Z(II2904) ) ;
NAND2   gate12083  (.A(II2903), .B(II2904), .Z(II2901) ) ;
NAND2   gate12084  (.A(II2885), .B(II2901), .Z(II2909) ) ;
NAND2   gate12085  (.A(II2885), .B(II2909), .Z(II2910) ) ;
NAND2   gate12086  (.A(II2901), .B(II2909), .Z(II2911) ) ;
NAND2   gate12087  (.A(WX1002), .B(WX705), .Z(II2918) ) ;
NAND2   gate12088  (.A(WX1002), .B(II2918), .Z(II2919) ) ;
NAND2   gate12089  (.A(WX705), .B(II2918), .Z(II2920) ) ;
NAND2   gate12090  (.A(II2919), .B(II2920), .Z(II2917) ) ;
NAND2   gate12091  (.A(WX769), .B(II2917), .Z(II2925) ) ;
NAND2   gate12092  (.A(WX769), .B(II2925), .Z(II2926) ) ;
NAND2   gate12093  (.A(II2917), .B(II2925), .Z(II2927) ) ;
NAND2   gate12094  (.A(II2926), .B(II2927), .Z(II2916) ) ;
NAND2   gate12095  (.A(WX833), .B(WX897), .Z(II2933) ) ;
NAND2   gate12096  (.A(WX833), .B(II2933), .Z(II2934) ) ;
NAND2   gate12097  (.A(WX897), .B(II2933), .Z(II2935) ) ;
NAND2   gate12098  (.A(II2934), .B(II2935), .Z(II2932) ) ;
NAND2   gate12099  (.A(II2916), .B(II2932), .Z(II2940) ) ;
NAND2   gate12100  (.A(II2916), .B(II2940), .Z(II2941) ) ;
NAND2   gate12101  (.A(II2932), .B(II2940), .Z(II2942) ) ;
NAND2   gate12102  (.A(WX1002), .B(WX707), .Z(II2949) ) ;
NAND2   gate12103  (.A(WX1002), .B(II2949), .Z(II2950) ) ;
NAND2   gate12104  (.A(WX707), .B(II2949), .Z(II2951) ) ;
NAND2   gate12105  (.A(II2950), .B(II2951), .Z(II2948) ) ;
NAND2   gate12106  (.A(WX771), .B(II2948), .Z(II2956) ) ;
NAND2   gate12107  (.A(WX771), .B(II2956), .Z(II2957) ) ;
NAND2   gate12108  (.A(II2948), .B(II2956), .Z(II2958) ) ;
NAND2   gate12109  (.A(II2957), .B(II2958), .Z(II2947) ) ;
NAND2   gate12110  (.A(WX835), .B(WX899), .Z(II2964) ) ;
NAND2   gate12111  (.A(WX835), .B(II2964), .Z(II2965) ) ;
NAND2   gate12112  (.A(WX899), .B(II2964), .Z(II2966) ) ;
NAND2   gate12113  (.A(II2965), .B(II2966), .Z(II2963) ) ;
NAND2   gate12114  (.A(II2947), .B(II2963), .Z(II2971) ) ;
NAND2   gate12115  (.A(II2947), .B(II2971), .Z(II2972) ) ;
NAND2   gate12116  (.A(II2963), .B(II2971), .Z(II2973) ) ;
NAND2   gate12117  (.A(WX580), .B(WX485), .Z(II3052) ) ;
NAND2   gate12118  (.A(WX580), .B(II3052), .Z(II3053) ) ;
NAND2   gate12119  (.A(WX485), .B(II3052), .Z(II3054) ) ;
NAND2   gate12120  (.A(WX581), .B(WX487), .Z(II3065) ) ;
NAND2   gate12121  (.A(WX581), .B(II3065), .Z(II3066) ) ;
NAND2   gate12122  (.A(WX487), .B(II3065), .Z(II3067) ) ;
NAND2   gate12123  (.A(WX582), .B(WX489), .Z(II3078) ) ;
NAND2   gate12124  (.A(WX582), .B(II3078), .Z(II3079) ) ;
NAND2   gate12125  (.A(WX489), .B(II3078), .Z(II3080) ) ;
NAND2   gate12126  (.A(WX583), .B(WX491), .Z(II3091) ) ;
NAND2   gate12127  (.A(WX583), .B(II3091), .Z(II3092) ) ;
NAND2   gate12128  (.A(WX491), .B(II3091), .Z(II3093) ) ;
NAND2   gate12129  (.A(WX584), .B(WX493), .Z(II3104) ) ;
NAND2   gate12130  (.A(WX584), .B(II3104), .Z(II3105) ) ;
NAND2   gate12131  (.A(WX493), .B(II3104), .Z(II3106) ) ;
NAND2   gate12132  (.A(WX585), .B(WX495), .Z(II3117) ) ;
NAND2   gate12133  (.A(WX585), .B(II3117), .Z(II3118) ) ;
NAND2   gate12134  (.A(WX495), .B(II3117), .Z(II3119) ) ;
NAND2   gate12135  (.A(WX586), .B(WX497), .Z(II3130) ) ;
NAND2   gate12136  (.A(WX586), .B(II3130), .Z(II3131) ) ;
NAND2   gate12137  (.A(WX497), .B(II3130), .Z(II3132) ) ;
NAND2   gate12138  (.A(WX587), .B(WX499), .Z(II3143) ) ;
NAND2   gate12139  (.A(WX587), .B(II3143), .Z(II3144) ) ;
NAND2   gate12140  (.A(WX499), .B(II3143), .Z(II3145) ) ;
NAND2   gate12141  (.A(WX588), .B(WX501), .Z(II3156) ) ;
NAND2   gate12142  (.A(WX588), .B(II3156), .Z(II3157) ) ;
NAND2   gate12143  (.A(WX501), .B(II3156), .Z(II3158) ) ;
NAND2   gate12144  (.A(WX589), .B(WX503), .Z(II3169) ) ;
NAND2   gate12145  (.A(WX589), .B(II3169), .Z(II3170) ) ;
NAND2   gate12146  (.A(WX503), .B(II3169), .Z(II3171) ) ;
NAND2   gate12147  (.A(WX590), .B(WX505), .Z(II3182) ) ;
NAND2   gate12148  (.A(WX590), .B(II3182), .Z(II3183) ) ;
NAND2   gate12149  (.A(WX505), .B(II3182), .Z(II3184) ) ;
NAND2   gate12150  (.A(WX591), .B(WX507), .Z(II3195) ) ;
NAND2   gate12151  (.A(WX591), .B(II3195), .Z(II3196) ) ;
NAND2   gate12152  (.A(WX507), .B(II3195), .Z(II3197) ) ;
NAND2   gate12153  (.A(WX592), .B(WX509), .Z(II3208) ) ;
NAND2   gate12154  (.A(WX592), .B(II3208), .Z(II3209) ) ;
NAND2   gate12155  (.A(WX509), .B(II3208), .Z(II3210) ) ;
NAND2   gate12156  (.A(WX593), .B(WX511), .Z(II3221) ) ;
NAND2   gate12157  (.A(WX593), .B(II3221), .Z(II3222) ) ;
NAND2   gate12158  (.A(WX511), .B(II3221), .Z(II3223) ) ;
NAND2   gate12159  (.A(WX594), .B(WX513), .Z(II3234) ) ;
NAND2   gate12160  (.A(WX594), .B(II3234), .Z(II3235) ) ;
NAND2   gate12161  (.A(WX513), .B(II3234), .Z(II3236) ) ;
NAND2   gate12162  (.A(WX595), .B(WX515), .Z(II3247) ) ;
NAND2   gate12163  (.A(WX595), .B(II3247), .Z(II3248) ) ;
NAND2   gate12164  (.A(WX515), .B(II3247), .Z(II3249) ) ;
NAND2   gate12165  (.A(WX596), .B(WX517), .Z(II3260) ) ;
NAND2   gate12166  (.A(WX596), .B(II3260), .Z(II3261) ) ;
NAND2   gate12167  (.A(WX517), .B(II3260), .Z(II3262) ) ;
NAND2   gate12168  (.A(WX597), .B(WX519), .Z(II3273) ) ;
NAND2   gate12169  (.A(WX597), .B(II3273), .Z(II3274) ) ;
NAND2   gate12170  (.A(WX519), .B(II3273), .Z(II3275) ) ;
NAND2   gate12171  (.A(WX598), .B(WX521), .Z(II3286) ) ;
NAND2   gate12172  (.A(WX598), .B(II3286), .Z(II3287) ) ;
NAND2   gate12173  (.A(WX521), .B(II3286), .Z(II3288) ) ;
NAND2   gate12174  (.A(WX599), .B(WX523), .Z(II3299) ) ;
NAND2   gate12175  (.A(WX599), .B(II3299), .Z(II3300) ) ;
NAND2   gate12176  (.A(WX523), .B(II3299), .Z(II3301) ) ;
NAND2   gate12177  (.A(WX600), .B(WX525), .Z(II3312) ) ;
NAND2   gate12178  (.A(WX600), .B(II3312), .Z(II3313) ) ;
NAND2   gate12179  (.A(WX525), .B(II3312), .Z(II3314) ) ;
NAND2   gate12180  (.A(WX601), .B(WX527), .Z(II3325) ) ;
NAND2   gate12181  (.A(WX601), .B(II3325), .Z(II3326) ) ;
NAND2   gate12182  (.A(WX527), .B(II3325), .Z(II3327) ) ;
NAND2   gate12183  (.A(WX602), .B(WX529), .Z(II3338) ) ;
NAND2   gate12184  (.A(WX602), .B(II3338), .Z(II3339) ) ;
NAND2   gate12185  (.A(WX529), .B(II3338), .Z(II3340) ) ;
NAND2   gate12186  (.A(WX603), .B(WX531), .Z(II3351) ) ;
NAND2   gate12187  (.A(WX603), .B(II3351), .Z(II3352) ) ;
NAND2   gate12188  (.A(WX531), .B(II3351), .Z(II3353) ) ;
NAND2   gate12189  (.A(WX604), .B(WX533), .Z(II3364) ) ;
NAND2   gate12190  (.A(WX604), .B(II3364), .Z(II3365) ) ;
NAND2   gate12191  (.A(WX533), .B(II3364), .Z(II3366) ) ;
NAND2   gate12192  (.A(WX605), .B(WX535), .Z(II3377) ) ;
NAND2   gate12193  (.A(WX605), .B(II3377), .Z(II3378) ) ;
NAND2   gate12194  (.A(WX535), .B(II3377), .Z(II3379) ) ;
NAND2   gate12195  (.A(WX606), .B(WX537), .Z(II3390) ) ;
NAND2   gate12196  (.A(WX606), .B(II3390), .Z(II3391) ) ;
NAND2   gate12197  (.A(WX537), .B(II3390), .Z(II3392) ) ;
NAND2   gate12198  (.A(WX607), .B(WX539), .Z(II3403) ) ;
NAND2   gate12199  (.A(WX607), .B(II3403), .Z(II3404) ) ;
NAND2   gate12200  (.A(WX539), .B(II3403), .Z(II3405) ) ;
NAND2   gate12201  (.A(WX608), .B(WX541), .Z(II3416) ) ;
NAND2   gate12202  (.A(WX608), .B(II3416), .Z(II3417) ) ;
NAND2   gate12203  (.A(WX541), .B(II3416), .Z(II3418) ) ;
NAND2   gate12204  (.A(WX609), .B(WX543), .Z(II3429) ) ;
NAND2   gate12205  (.A(WX609), .B(II3429), .Z(II3430) ) ;
NAND2   gate12206  (.A(WX543), .B(II3429), .Z(II3431) ) ;
NAND2   gate12207  (.A(WX610), .B(WX545), .Z(II3442) ) ;
NAND2   gate12208  (.A(WX610), .B(II3442), .Z(II3443) ) ;
NAND2   gate12209  (.A(WX545), .B(II3442), .Z(II3444) ) ;
NAND2   gate12210  (.A(WX611), .B(WX547), .Z(II3455) ) ;
NAND2   gate12211  (.A(WX611), .B(II3455), .Z(II3456) ) ;
NAND2   gate12212  (.A(WX547), .B(II3455), .Z(II3457) ) ;
NAND2   gate12213  (.A(WX627), .B(CRC_OUT_9_31), .Z(II3470) ) ;
NAND2   gate12214  (.A(WX627), .B(II3470), .Z(II3471) ) ;
NAND2   gate12215  (.A(CRC_OUT_9_31), .B(II3470), .Z(II3472) ) ;
NAND2   gate12216  (.A(II3471), .B(II3472), .Z(II3469) ) ;
NAND2   gate12217  (.A(CRC_OUT_9_15), .B(II3469), .Z(II3477) ) ;
NAND2   gate12218  (.A(CRC_OUT_9_15), .B(II3477), .Z(II3478) ) ;
NAND2   gate12219  (.A(II3469), .B(II3477), .Z(II3479) ) ;
NAND2   gate12220  (.A(WX632), .B(CRC_OUT_9_31), .Z(II3485) ) ;
NAND2   gate12221  (.A(WX632), .B(II3485), .Z(II3486) ) ;
NAND2   gate12222  (.A(CRC_OUT_9_31), .B(II3485), .Z(II3487) ) ;
NAND2   gate12223  (.A(II3486), .B(II3487), .Z(II3484) ) ;
NAND2   gate12224  (.A(CRC_OUT_9_10), .B(II3484), .Z(II3492) ) ;
NAND2   gate12225  (.A(CRC_OUT_9_10), .B(II3492), .Z(II3493) ) ;
NAND2   gate12226  (.A(II3484), .B(II3492), .Z(II3494) ) ;
NAND2   gate12227  (.A(WX639), .B(CRC_OUT_9_31), .Z(II3500) ) ;
NAND2   gate12228  (.A(WX639), .B(II3500), .Z(II3501) ) ;
NAND2   gate12229  (.A(CRC_OUT_9_31), .B(II3500), .Z(II3502) ) ;
NAND2   gate12230  (.A(II3501), .B(II3502), .Z(II3499) ) ;
NAND2   gate12231  (.A(CRC_OUT_9_3), .B(II3499), .Z(II3507) ) ;
NAND2   gate12232  (.A(CRC_OUT_9_3), .B(II3507), .Z(II3508) ) ;
NAND2   gate12233  (.A(II3499), .B(II3507), .Z(II3509) ) ;
NAND2   gate12234  (.A(WX643), .B(CRC_OUT_9_31), .Z(II3514) ) ;
NAND2   gate12235  (.A(WX643), .B(II3514), .Z(II3515) ) ;
NAND2   gate12236  (.A(CRC_OUT_9_31), .B(II3514), .Z(II3516) ) ;
NAND2   gate12237  (.A(WX612), .B(CRC_OUT_9_30), .Z(II3521) ) ;
NAND2   gate12238  (.A(WX612), .B(II3521), .Z(II3522) ) ;
NAND2   gate12239  (.A(CRC_OUT_9_30), .B(II3521), .Z(II3523) ) ;
NAND2   gate12240  (.A(WX613), .B(CRC_OUT_9_29), .Z(II3528) ) ;
NAND2   gate12241  (.A(WX613), .B(II3528), .Z(II3529) ) ;
NAND2   gate12242  (.A(CRC_OUT_9_29), .B(II3528), .Z(II3530) ) ;
NAND2   gate12243  (.A(WX614), .B(CRC_OUT_9_28), .Z(II3535) ) ;
NAND2   gate12244  (.A(WX614), .B(II3535), .Z(II3536) ) ;
NAND2   gate12245  (.A(CRC_OUT_9_28), .B(II3535), .Z(II3537) ) ;
NAND2   gate12246  (.A(WX615), .B(CRC_OUT_9_27), .Z(II3542) ) ;
NAND2   gate12247  (.A(WX615), .B(II3542), .Z(II3543) ) ;
NAND2   gate12248  (.A(CRC_OUT_9_27), .B(II3542), .Z(II3544) ) ;
NAND2   gate12249  (.A(WX616), .B(CRC_OUT_9_26), .Z(II3549) ) ;
NAND2   gate12250  (.A(WX616), .B(II3549), .Z(II3550) ) ;
NAND2   gate12251  (.A(CRC_OUT_9_26), .B(II3549), .Z(II3551) ) ;
NAND2   gate12252  (.A(WX617), .B(CRC_OUT_9_25), .Z(II3556) ) ;
NAND2   gate12253  (.A(WX617), .B(II3556), .Z(II3557) ) ;
NAND2   gate12254  (.A(CRC_OUT_9_25), .B(II3556), .Z(II3558) ) ;
NAND2   gate12255  (.A(WX618), .B(CRC_OUT_9_24), .Z(II3563) ) ;
NAND2   gate12256  (.A(WX618), .B(II3563), .Z(II3564) ) ;
NAND2   gate12257  (.A(CRC_OUT_9_24), .B(II3563), .Z(II3565) ) ;
NAND2   gate12258  (.A(WX619), .B(CRC_OUT_9_23), .Z(II3570) ) ;
NAND2   gate12259  (.A(WX619), .B(II3570), .Z(II3571) ) ;
NAND2   gate12260  (.A(CRC_OUT_9_23), .B(II3570), .Z(II3572) ) ;
NAND2   gate12261  (.A(WX620), .B(CRC_OUT_9_22), .Z(II3577) ) ;
NAND2   gate12262  (.A(WX620), .B(II3577), .Z(II3578) ) ;
NAND2   gate12263  (.A(CRC_OUT_9_22), .B(II3577), .Z(II3579) ) ;
NAND2   gate12264  (.A(WX621), .B(CRC_OUT_9_21), .Z(II3584) ) ;
NAND2   gate12265  (.A(WX621), .B(II3584), .Z(II3585) ) ;
NAND2   gate12266  (.A(CRC_OUT_9_21), .B(II3584), .Z(II3586) ) ;
NAND2   gate12267  (.A(WX622), .B(CRC_OUT_9_20), .Z(II3591) ) ;
NAND2   gate12268  (.A(WX622), .B(II3591), .Z(II3592) ) ;
NAND2   gate12269  (.A(CRC_OUT_9_20), .B(II3591), .Z(II3593) ) ;
NAND2   gate12270  (.A(WX623), .B(CRC_OUT_9_19), .Z(II3598) ) ;
NAND2   gate12271  (.A(WX623), .B(II3598), .Z(II3599) ) ;
NAND2   gate12272  (.A(CRC_OUT_9_19), .B(II3598), .Z(II3600) ) ;
NAND2   gate12273  (.A(WX624), .B(CRC_OUT_9_18), .Z(II3605) ) ;
NAND2   gate12274  (.A(WX624), .B(II3605), .Z(II3606) ) ;
NAND2   gate12275  (.A(CRC_OUT_9_18), .B(II3605), .Z(II3607) ) ;
NAND2   gate12276  (.A(WX625), .B(CRC_OUT_9_17), .Z(II3612) ) ;
NAND2   gate12277  (.A(WX625), .B(II3612), .Z(II3613) ) ;
NAND2   gate12278  (.A(CRC_OUT_9_17), .B(II3612), .Z(II3614) ) ;
NAND2   gate12279  (.A(WX626), .B(CRC_OUT_9_16), .Z(II3619) ) ;
NAND2   gate12280  (.A(WX626), .B(II3619), .Z(II3620) ) ;
NAND2   gate12281  (.A(CRC_OUT_9_16), .B(II3619), .Z(II3621) ) ;
NAND2   gate12282  (.A(WX628), .B(CRC_OUT_9_14), .Z(II3626) ) ;
NAND2   gate12283  (.A(WX628), .B(II3626), .Z(II3627) ) ;
NAND2   gate12284  (.A(CRC_OUT_9_14), .B(II3626), .Z(II3628) ) ;
NAND2   gate12285  (.A(WX629), .B(CRC_OUT_9_13), .Z(II3633) ) ;
NAND2   gate12286  (.A(WX629), .B(II3633), .Z(II3634) ) ;
NAND2   gate12287  (.A(CRC_OUT_9_13), .B(II3633), .Z(II3635) ) ;
NAND2   gate12288  (.A(WX630), .B(CRC_OUT_9_12), .Z(II3640) ) ;
NAND2   gate12289  (.A(WX630), .B(II3640), .Z(II3641) ) ;
NAND2   gate12290  (.A(CRC_OUT_9_12), .B(II3640), .Z(II3642) ) ;
NAND2   gate12291  (.A(WX631), .B(CRC_OUT_9_11), .Z(II3647) ) ;
NAND2   gate12292  (.A(WX631), .B(II3647), .Z(II3648) ) ;
NAND2   gate12293  (.A(CRC_OUT_9_11), .B(II3647), .Z(II3649) ) ;
NAND2   gate12294  (.A(WX633), .B(CRC_OUT_9_9), .Z(II3654) ) ;
NAND2   gate12295  (.A(WX633), .B(II3654), .Z(II3655) ) ;
NAND2   gate12296  (.A(CRC_OUT_9_9), .B(II3654), .Z(II3656) ) ;
NAND2   gate12297  (.A(WX634), .B(CRC_OUT_9_8), .Z(II3661) ) ;
NAND2   gate12298  (.A(WX634), .B(II3661), .Z(II3662) ) ;
NAND2   gate12299  (.A(CRC_OUT_9_8), .B(II3661), .Z(II3663) ) ;
NAND2   gate12300  (.A(WX635), .B(CRC_OUT_9_7), .Z(II3668) ) ;
NAND2   gate12301  (.A(WX635), .B(II3668), .Z(II3669) ) ;
NAND2   gate12302  (.A(CRC_OUT_9_7), .B(II3668), .Z(II3670) ) ;
NAND2   gate12303  (.A(WX636), .B(CRC_OUT_9_6), .Z(II3675) ) ;
NAND2   gate12304  (.A(WX636), .B(II3675), .Z(II3676) ) ;
NAND2   gate12305  (.A(CRC_OUT_9_6), .B(II3675), .Z(II3677) ) ;
NAND2   gate12306  (.A(WX637), .B(CRC_OUT_9_5), .Z(II3682) ) ;
NAND2   gate12307  (.A(WX637), .B(II3682), .Z(II3683) ) ;
NAND2   gate12308  (.A(CRC_OUT_9_5), .B(II3682), .Z(II3684) ) ;
NAND2   gate12309  (.A(WX638), .B(CRC_OUT_9_4), .Z(II3689) ) ;
NAND2   gate12310  (.A(WX638), .B(II3689), .Z(II3690) ) ;
NAND2   gate12311  (.A(CRC_OUT_9_4), .B(II3689), .Z(II3691) ) ;
NAND2   gate12312  (.A(WX640), .B(CRC_OUT_9_2), .Z(II3696) ) ;
NAND2   gate12313  (.A(WX640), .B(II3696), .Z(II3697) ) ;
NAND2   gate12314  (.A(CRC_OUT_9_2), .B(II3696), .Z(II3698) ) ;
NAND2   gate12315  (.A(WX641), .B(CRC_OUT_9_1), .Z(II3703) ) ;
NAND2   gate12316  (.A(WX641), .B(II3703), .Z(II3704) ) ;
NAND2   gate12317  (.A(CRC_OUT_9_1), .B(II3703), .Z(II3705) ) ;
NAND2   gate12318  (.A(WX642), .B(CRC_OUT_9_0), .Z(II3710) ) ;
NAND2   gate12319  (.A(WX642), .B(II3710), .Z(II3711) ) ;
NAND2   gate12320  (.A(CRC_OUT_9_0), .B(II3710), .Z(II3712) ) ;
NAND2   gate12321  (.A(WX2294), .B(WX1938), .Z(II5993) ) ;
NAND2   gate12322  (.A(WX2294), .B(II5993), .Z(II5994) ) ;
NAND2   gate12323  (.A(WX1938), .B(II5993), .Z(II5995) ) ;
NAND2   gate12324  (.A(II5994), .B(II5995), .Z(II5992) ) ;
NAND2   gate12325  (.A(WX2002), .B(II5992), .Z(II6000) ) ;
NAND2   gate12326  (.A(WX2002), .B(II6000), .Z(II6001) ) ;
NAND2   gate12327  (.A(II5992), .B(II6000), .Z(II6002) ) ;
NAND2   gate12328  (.A(II6001), .B(II6002), .Z(II5991) ) ;
NAND2   gate12329  (.A(WX2066), .B(WX2130), .Z(II6008) ) ;
NAND2   gate12330  (.A(WX2066), .B(II6008), .Z(II6009) ) ;
NAND2   gate12331  (.A(WX2130), .B(II6008), .Z(II6010) ) ;
NAND2   gate12332  (.A(II6009), .B(II6010), .Z(II6007) ) ;
NAND2   gate12333  (.A(II5991), .B(II6007), .Z(II6015) ) ;
NAND2   gate12334  (.A(II5991), .B(II6015), .Z(II6016) ) ;
NAND2   gate12335  (.A(II6007), .B(II6015), .Z(II6017) ) ;
NAND2   gate12336  (.A(WX2294), .B(WX1940), .Z(II6024) ) ;
NAND2   gate12337  (.A(WX2294), .B(II6024), .Z(II6025) ) ;
NAND2   gate12338  (.A(WX1940), .B(II6024), .Z(II6026) ) ;
NAND2   gate12339  (.A(II6025), .B(II6026), .Z(II6023) ) ;
NAND2   gate12340  (.A(WX2004), .B(II6023), .Z(II6031) ) ;
NAND2   gate12341  (.A(WX2004), .B(II6031), .Z(II6032) ) ;
NAND2   gate12342  (.A(II6023), .B(II6031), .Z(II6033) ) ;
NAND2   gate12343  (.A(II6032), .B(II6033), .Z(II6022) ) ;
NAND2   gate12344  (.A(WX2068), .B(WX2132), .Z(II6039) ) ;
NAND2   gate12345  (.A(WX2068), .B(II6039), .Z(II6040) ) ;
NAND2   gate12346  (.A(WX2132), .B(II6039), .Z(II6041) ) ;
NAND2   gate12347  (.A(II6040), .B(II6041), .Z(II6038) ) ;
NAND2   gate12348  (.A(II6022), .B(II6038), .Z(II6046) ) ;
NAND2   gate12349  (.A(II6022), .B(II6046), .Z(II6047) ) ;
NAND2   gate12350  (.A(II6038), .B(II6046), .Z(II6048) ) ;
NAND2   gate12351  (.A(WX2294), .B(WX1942), .Z(II6055) ) ;
NAND2   gate12352  (.A(WX2294), .B(II6055), .Z(II6056) ) ;
NAND2   gate12353  (.A(WX1942), .B(II6055), .Z(II6057) ) ;
NAND2   gate12354  (.A(II6056), .B(II6057), .Z(II6054) ) ;
NAND2   gate12355  (.A(WX2006), .B(II6054), .Z(II6062) ) ;
NAND2   gate12356  (.A(WX2006), .B(II6062), .Z(II6063) ) ;
NAND2   gate12357  (.A(II6054), .B(II6062), .Z(II6064) ) ;
NAND2   gate12358  (.A(II6063), .B(II6064), .Z(II6053) ) ;
NAND2   gate12359  (.A(WX2070), .B(WX2134), .Z(II6070) ) ;
NAND2   gate12360  (.A(WX2070), .B(II6070), .Z(II6071) ) ;
NAND2   gate12361  (.A(WX2134), .B(II6070), .Z(II6072) ) ;
NAND2   gate12362  (.A(II6071), .B(II6072), .Z(II6069) ) ;
NAND2   gate12363  (.A(II6053), .B(II6069), .Z(II6077) ) ;
NAND2   gate12364  (.A(II6053), .B(II6077), .Z(II6078) ) ;
NAND2   gate12365  (.A(II6069), .B(II6077), .Z(II6079) ) ;
NAND2   gate12366  (.A(WX2294), .B(WX1944), .Z(II6086) ) ;
NAND2   gate12367  (.A(WX2294), .B(II6086), .Z(II6087) ) ;
NAND2   gate12368  (.A(WX1944), .B(II6086), .Z(II6088) ) ;
NAND2   gate12369  (.A(II6087), .B(II6088), .Z(II6085) ) ;
NAND2   gate12370  (.A(WX2008), .B(II6085), .Z(II6093) ) ;
NAND2   gate12371  (.A(WX2008), .B(II6093), .Z(II6094) ) ;
NAND2   gate12372  (.A(II6085), .B(II6093), .Z(II6095) ) ;
NAND2   gate12373  (.A(II6094), .B(II6095), .Z(II6084) ) ;
NAND2   gate12374  (.A(WX2072), .B(WX2136), .Z(II6101) ) ;
NAND2   gate12375  (.A(WX2072), .B(II6101), .Z(II6102) ) ;
NAND2   gate12376  (.A(WX2136), .B(II6101), .Z(II6103) ) ;
NAND2   gate12377  (.A(II6102), .B(II6103), .Z(II6100) ) ;
NAND2   gate12378  (.A(II6084), .B(II6100), .Z(II6108) ) ;
NAND2   gate12379  (.A(II6084), .B(II6108), .Z(II6109) ) ;
NAND2   gate12380  (.A(II6100), .B(II6108), .Z(II6110) ) ;
NAND2   gate12381  (.A(WX2294), .B(WX1946), .Z(II6117) ) ;
NAND2   gate12382  (.A(WX2294), .B(II6117), .Z(II6118) ) ;
NAND2   gate12383  (.A(WX1946), .B(II6117), .Z(II6119) ) ;
NAND2   gate12384  (.A(II6118), .B(II6119), .Z(II6116) ) ;
NAND2   gate12385  (.A(WX2010), .B(II6116), .Z(II6124) ) ;
NAND2   gate12386  (.A(WX2010), .B(II6124), .Z(II6125) ) ;
NAND2   gate12387  (.A(II6116), .B(II6124), .Z(II6126) ) ;
NAND2   gate12388  (.A(II6125), .B(II6126), .Z(II6115) ) ;
NAND2   gate12389  (.A(WX2074), .B(WX2138), .Z(II6132) ) ;
NAND2   gate12390  (.A(WX2074), .B(II6132), .Z(II6133) ) ;
NAND2   gate12391  (.A(WX2138), .B(II6132), .Z(II6134) ) ;
NAND2   gate12392  (.A(II6133), .B(II6134), .Z(II6131) ) ;
NAND2   gate12393  (.A(II6115), .B(II6131), .Z(II6139) ) ;
NAND2   gate12394  (.A(II6115), .B(II6139), .Z(II6140) ) ;
NAND2   gate12395  (.A(II6131), .B(II6139), .Z(II6141) ) ;
NAND2   gate12396  (.A(WX2294), .B(WX1948), .Z(II6148) ) ;
NAND2   gate12397  (.A(WX2294), .B(II6148), .Z(II6149) ) ;
NAND2   gate12398  (.A(WX1948), .B(II6148), .Z(II6150) ) ;
NAND2   gate12399  (.A(II6149), .B(II6150), .Z(II6147) ) ;
NAND2   gate12400  (.A(WX2012), .B(II6147), .Z(II6155) ) ;
NAND2   gate12401  (.A(WX2012), .B(II6155), .Z(II6156) ) ;
NAND2   gate12402  (.A(II6147), .B(II6155), .Z(II6157) ) ;
NAND2   gate12403  (.A(II6156), .B(II6157), .Z(II6146) ) ;
NAND2   gate12404  (.A(WX2076), .B(WX2140), .Z(II6163) ) ;
NAND2   gate12405  (.A(WX2076), .B(II6163), .Z(II6164) ) ;
NAND2   gate12406  (.A(WX2140), .B(II6163), .Z(II6165) ) ;
NAND2   gate12407  (.A(II6164), .B(II6165), .Z(II6162) ) ;
NAND2   gate12408  (.A(II6146), .B(II6162), .Z(II6170) ) ;
NAND2   gate12409  (.A(II6146), .B(II6170), .Z(II6171) ) ;
NAND2   gate12410  (.A(II6162), .B(II6170), .Z(II6172) ) ;
NAND2   gate12411  (.A(WX2294), .B(WX1950), .Z(II6179) ) ;
NAND2   gate12412  (.A(WX2294), .B(II6179), .Z(II6180) ) ;
NAND2   gate12413  (.A(WX1950), .B(II6179), .Z(II6181) ) ;
NAND2   gate12414  (.A(II6180), .B(II6181), .Z(II6178) ) ;
NAND2   gate12415  (.A(WX2014), .B(II6178), .Z(II6186) ) ;
NAND2   gate12416  (.A(WX2014), .B(II6186), .Z(II6187) ) ;
NAND2   gate12417  (.A(II6178), .B(II6186), .Z(II6188) ) ;
NAND2   gate12418  (.A(II6187), .B(II6188), .Z(II6177) ) ;
NAND2   gate12419  (.A(WX2078), .B(WX2142), .Z(II6194) ) ;
NAND2   gate12420  (.A(WX2078), .B(II6194), .Z(II6195) ) ;
NAND2   gate12421  (.A(WX2142), .B(II6194), .Z(II6196) ) ;
NAND2   gate12422  (.A(II6195), .B(II6196), .Z(II6193) ) ;
NAND2   gate12423  (.A(II6177), .B(II6193), .Z(II6201) ) ;
NAND2   gate12424  (.A(II6177), .B(II6201), .Z(II6202) ) ;
NAND2   gate12425  (.A(II6193), .B(II6201), .Z(II6203) ) ;
NAND2   gate12426  (.A(WX2294), .B(WX1952), .Z(II6210) ) ;
NAND2   gate12427  (.A(WX2294), .B(II6210), .Z(II6211) ) ;
NAND2   gate12428  (.A(WX1952), .B(II6210), .Z(II6212) ) ;
NAND2   gate12429  (.A(II6211), .B(II6212), .Z(II6209) ) ;
NAND2   gate12430  (.A(WX2016), .B(II6209), .Z(II6217) ) ;
NAND2   gate12431  (.A(WX2016), .B(II6217), .Z(II6218) ) ;
NAND2   gate12432  (.A(II6209), .B(II6217), .Z(II6219) ) ;
NAND2   gate12433  (.A(II6218), .B(II6219), .Z(II6208) ) ;
NAND2   gate12434  (.A(WX2080), .B(WX2144), .Z(II6225) ) ;
NAND2   gate12435  (.A(WX2080), .B(II6225), .Z(II6226) ) ;
NAND2   gate12436  (.A(WX2144), .B(II6225), .Z(II6227) ) ;
NAND2   gate12437  (.A(II6226), .B(II6227), .Z(II6224) ) ;
NAND2   gate12438  (.A(II6208), .B(II6224), .Z(II6232) ) ;
NAND2   gate12439  (.A(II6208), .B(II6232), .Z(II6233) ) ;
NAND2   gate12440  (.A(II6224), .B(II6232), .Z(II6234) ) ;
NAND2   gate12441  (.A(WX2294), .B(WX1954), .Z(II6241) ) ;
NAND2   gate12442  (.A(WX2294), .B(II6241), .Z(II6242) ) ;
NAND2   gate12443  (.A(WX1954), .B(II6241), .Z(II6243) ) ;
NAND2   gate12444  (.A(II6242), .B(II6243), .Z(II6240) ) ;
NAND2   gate12445  (.A(WX2018), .B(II6240), .Z(II6248) ) ;
NAND2   gate12446  (.A(WX2018), .B(II6248), .Z(II6249) ) ;
NAND2   gate12447  (.A(II6240), .B(II6248), .Z(II6250) ) ;
NAND2   gate12448  (.A(II6249), .B(II6250), .Z(II6239) ) ;
NAND2   gate12449  (.A(WX2082), .B(WX2146), .Z(II6256) ) ;
NAND2   gate12450  (.A(WX2082), .B(II6256), .Z(II6257) ) ;
NAND2   gate12451  (.A(WX2146), .B(II6256), .Z(II6258) ) ;
NAND2   gate12452  (.A(II6257), .B(II6258), .Z(II6255) ) ;
NAND2   gate12453  (.A(II6239), .B(II6255), .Z(II6263) ) ;
NAND2   gate12454  (.A(II6239), .B(II6263), .Z(II6264) ) ;
NAND2   gate12455  (.A(II6255), .B(II6263), .Z(II6265) ) ;
NAND2   gate12456  (.A(WX2294), .B(WX1956), .Z(II6272) ) ;
NAND2   gate12457  (.A(WX2294), .B(II6272), .Z(II6273) ) ;
NAND2   gate12458  (.A(WX1956), .B(II6272), .Z(II6274) ) ;
NAND2   gate12459  (.A(II6273), .B(II6274), .Z(II6271) ) ;
NAND2   gate12460  (.A(WX2020), .B(II6271), .Z(II6279) ) ;
NAND2   gate12461  (.A(WX2020), .B(II6279), .Z(II6280) ) ;
NAND2   gate12462  (.A(II6271), .B(II6279), .Z(II6281) ) ;
NAND2   gate12463  (.A(II6280), .B(II6281), .Z(II6270) ) ;
NAND2   gate12464  (.A(WX2084), .B(WX2148), .Z(II6287) ) ;
NAND2   gate12465  (.A(WX2084), .B(II6287), .Z(II6288) ) ;
NAND2   gate12466  (.A(WX2148), .B(II6287), .Z(II6289) ) ;
NAND2   gate12467  (.A(II6288), .B(II6289), .Z(II6286) ) ;
NAND2   gate12468  (.A(II6270), .B(II6286), .Z(II6294) ) ;
NAND2   gate12469  (.A(II6270), .B(II6294), .Z(II6295) ) ;
NAND2   gate12470  (.A(II6286), .B(II6294), .Z(II6296) ) ;
NAND2   gate12471  (.A(WX2294), .B(WX1958), .Z(II6303) ) ;
NAND2   gate12472  (.A(WX2294), .B(II6303), .Z(II6304) ) ;
NAND2   gate12473  (.A(WX1958), .B(II6303), .Z(II6305) ) ;
NAND2   gate12474  (.A(II6304), .B(II6305), .Z(II6302) ) ;
NAND2   gate12475  (.A(WX2022), .B(II6302), .Z(II6310) ) ;
NAND2   gate12476  (.A(WX2022), .B(II6310), .Z(II6311) ) ;
NAND2   gate12477  (.A(II6302), .B(II6310), .Z(II6312) ) ;
NAND2   gate12478  (.A(II6311), .B(II6312), .Z(II6301) ) ;
NAND2   gate12479  (.A(WX2086), .B(WX2150), .Z(II6318) ) ;
NAND2   gate12480  (.A(WX2086), .B(II6318), .Z(II6319) ) ;
NAND2   gate12481  (.A(WX2150), .B(II6318), .Z(II6320) ) ;
NAND2   gate12482  (.A(II6319), .B(II6320), .Z(II6317) ) ;
NAND2   gate12483  (.A(II6301), .B(II6317), .Z(II6325) ) ;
NAND2   gate12484  (.A(II6301), .B(II6325), .Z(II6326) ) ;
NAND2   gate12485  (.A(II6317), .B(II6325), .Z(II6327) ) ;
NAND2   gate12486  (.A(WX2294), .B(WX1960), .Z(II6334) ) ;
NAND2   gate12487  (.A(WX2294), .B(II6334), .Z(II6335) ) ;
NAND2   gate12488  (.A(WX1960), .B(II6334), .Z(II6336) ) ;
NAND2   gate12489  (.A(II6335), .B(II6336), .Z(II6333) ) ;
NAND2   gate12490  (.A(WX2024), .B(II6333), .Z(II6341) ) ;
NAND2   gate12491  (.A(WX2024), .B(II6341), .Z(II6342) ) ;
NAND2   gate12492  (.A(II6333), .B(II6341), .Z(II6343) ) ;
NAND2   gate12493  (.A(II6342), .B(II6343), .Z(II6332) ) ;
NAND2   gate12494  (.A(WX2088), .B(WX2152), .Z(II6349) ) ;
NAND2   gate12495  (.A(WX2088), .B(II6349), .Z(II6350) ) ;
NAND2   gate12496  (.A(WX2152), .B(II6349), .Z(II6351) ) ;
NAND2   gate12497  (.A(II6350), .B(II6351), .Z(II6348) ) ;
NAND2   gate12498  (.A(II6332), .B(II6348), .Z(II6356) ) ;
NAND2   gate12499  (.A(II6332), .B(II6356), .Z(II6357) ) ;
NAND2   gate12500  (.A(II6348), .B(II6356), .Z(II6358) ) ;
NAND2   gate12501  (.A(WX2294), .B(WX1962), .Z(II6365) ) ;
NAND2   gate12502  (.A(WX2294), .B(II6365), .Z(II6366) ) ;
NAND2   gate12503  (.A(WX1962), .B(II6365), .Z(II6367) ) ;
NAND2   gate12504  (.A(II6366), .B(II6367), .Z(II6364) ) ;
NAND2   gate12505  (.A(WX2026), .B(II6364), .Z(II6372) ) ;
NAND2   gate12506  (.A(WX2026), .B(II6372), .Z(II6373) ) ;
NAND2   gate12507  (.A(II6364), .B(II6372), .Z(II6374) ) ;
NAND2   gate12508  (.A(II6373), .B(II6374), .Z(II6363) ) ;
NAND2   gate12509  (.A(WX2090), .B(WX2154), .Z(II6380) ) ;
NAND2   gate12510  (.A(WX2090), .B(II6380), .Z(II6381) ) ;
NAND2   gate12511  (.A(WX2154), .B(II6380), .Z(II6382) ) ;
NAND2   gate12512  (.A(II6381), .B(II6382), .Z(II6379) ) ;
NAND2   gate12513  (.A(II6363), .B(II6379), .Z(II6387) ) ;
NAND2   gate12514  (.A(II6363), .B(II6387), .Z(II6388) ) ;
NAND2   gate12515  (.A(II6379), .B(II6387), .Z(II6389) ) ;
NAND2   gate12516  (.A(WX2294), .B(WX1964), .Z(II6396) ) ;
NAND2   gate12517  (.A(WX2294), .B(II6396), .Z(II6397) ) ;
NAND2   gate12518  (.A(WX1964), .B(II6396), .Z(II6398) ) ;
NAND2   gate12519  (.A(II6397), .B(II6398), .Z(II6395) ) ;
NAND2   gate12520  (.A(WX2028), .B(II6395), .Z(II6403) ) ;
NAND2   gate12521  (.A(WX2028), .B(II6403), .Z(II6404) ) ;
NAND2   gate12522  (.A(II6395), .B(II6403), .Z(II6405) ) ;
NAND2   gate12523  (.A(II6404), .B(II6405), .Z(II6394) ) ;
NAND2   gate12524  (.A(WX2092), .B(WX2156), .Z(II6411) ) ;
NAND2   gate12525  (.A(WX2092), .B(II6411), .Z(II6412) ) ;
NAND2   gate12526  (.A(WX2156), .B(II6411), .Z(II6413) ) ;
NAND2   gate12527  (.A(II6412), .B(II6413), .Z(II6410) ) ;
NAND2   gate12528  (.A(II6394), .B(II6410), .Z(II6418) ) ;
NAND2   gate12529  (.A(II6394), .B(II6418), .Z(II6419) ) ;
NAND2   gate12530  (.A(II6410), .B(II6418), .Z(II6420) ) ;
NAND2   gate12531  (.A(WX2294), .B(WX1966), .Z(II6427) ) ;
NAND2   gate12532  (.A(WX2294), .B(II6427), .Z(II6428) ) ;
NAND2   gate12533  (.A(WX1966), .B(II6427), .Z(II6429) ) ;
NAND2   gate12534  (.A(II6428), .B(II6429), .Z(II6426) ) ;
NAND2   gate12535  (.A(WX2030), .B(II6426), .Z(II6434) ) ;
NAND2   gate12536  (.A(WX2030), .B(II6434), .Z(II6435) ) ;
NAND2   gate12537  (.A(II6426), .B(II6434), .Z(II6436) ) ;
NAND2   gate12538  (.A(II6435), .B(II6436), .Z(II6425) ) ;
NAND2   gate12539  (.A(WX2094), .B(WX2158), .Z(II6442) ) ;
NAND2   gate12540  (.A(WX2094), .B(II6442), .Z(II6443) ) ;
NAND2   gate12541  (.A(WX2158), .B(II6442), .Z(II6444) ) ;
NAND2   gate12542  (.A(II6443), .B(II6444), .Z(II6441) ) ;
NAND2   gate12543  (.A(II6425), .B(II6441), .Z(II6449) ) ;
NAND2   gate12544  (.A(II6425), .B(II6449), .Z(II6450) ) ;
NAND2   gate12545  (.A(II6441), .B(II6449), .Z(II6451) ) ;
NAND2   gate12546  (.A(WX2294), .B(WX1968), .Z(II6458) ) ;
NAND2   gate12547  (.A(WX2294), .B(II6458), .Z(II6459) ) ;
NAND2   gate12548  (.A(WX1968), .B(II6458), .Z(II6460) ) ;
NAND2   gate12549  (.A(II6459), .B(II6460), .Z(II6457) ) ;
NAND2   gate12550  (.A(WX2032), .B(II6457), .Z(II6465) ) ;
NAND2   gate12551  (.A(WX2032), .B(II6465), .Z(II6466) ) ;
NAND2   gate12552  (.A(II6457), .B(II6465), .Z(II6467) ) ;
NAND2   gate12553  (.A(II6466), .B(II6467), .Z(II6456) ) ;
NAND2   gate12554  (.A(WX2096), .B(WX2160), .Z(II6473) ) ;
NAND2   gate12555  (.A(WX2096), .B(II6473), .Z(II6474) ) ;
NAND2   gate12556  (.A(WX2160), .B(II6473), .Z(II6475) ) ;
NAND2   gate12557  (.A(II6474), .B(II6475), .Z(II6472) ) ;
NAND2   gate12558  (.A(II6456), .B(II6472), .Z(II6480) ) ;
NAND2   gate12559  (.A(II6456), .B(II6480), .Z(II6481) ) ;
NAND2   gate12560  (.A(II6472), .B(II6480), .Z(II6482) ) ;
NAND2   gate12561  (.A(WX2295), .B(WX1970), .Z(II6489) ) ;
NAND2   gate12562  (.A(WX2295), .B(II6489), .Z(II6490) ) ;
NAND2   gate12563  (.A(WX1970), .B(II6489), .Z(II6491) ) ;
NAND2   gate12564  (.A(II6490), .B(II6491), .Z(II6488) ) ;
NAND2   gate12565  (.A(WX2034), .B(II6488), .Z(II6496) ) ;
NAND2   gate12566  (.A(WX2034), .B(II6496), .Z(II6497) ) ;
NAND2   gate12567  (.A(II6488), .B(II6496), .Z(II6498) ) ;
NAND2   gate12568  (.A(II6497), .B(II6498), .Z(II6487) ) ;
NAND2   gate12569  (.A(WX2098), .B(WX2162), .Z(II6504) ) ;
NAND2   gate12570  (.A(WX2098), .B(II6504), .Z(II6505) ) ;
NAND2   gate12571  (.A(WX2162), .B(II6504), .Z(II6506) ) ;
NAND2   gate12572  (.A(II6505), .B(II6506), .Z(II6503) ) ;
NAND2   gate12573  (.A(II6487), .B(II6503), .Z(II6511) ) ;
NAND2   gate12574  (.A(II6487), .B(II6511), .Z(II6512) ) ;
NAND2   gate12575  (.A(II6503), .B(II6511), .Z(II6513) ) ;
NAND2   gate12576  (.A(WX2295), .B(WX1972), .Z(II6520) ) ;
NAND2   gate12577  (.A(WX2295), .B(II6520), .Z(II6521) ) ;
NAND2   gate12578  (.A(WX1972), .B(II6520), .Z(II6522) ) ;
NAND2   gate12579  (.A(II6521), .B(II6522), .Z(II6519) ) ;
NAND2   gate12580  (.A(WX2036), .B(II6519), .Z(II6527) ) ;
NAND2   gate12581  (.A(WX2036), .B(II6527), .Z(II6528) ) ;
NAND2   gate12582  (.A(II6519), .B(II6527), .Z(II6529) ) ;
NAND2   gate12583  (.A(II6528), .B(II6529), .Z(II6518) ) ;
NAND2   gate12584  (.A(WX2100), .B(WX2164), .Z(II6535) ) ;
NAND2   gate12585  (.A(WX2100), .B(II6535), .Z(II6536) ) ;
NAND2   gate12586  (.A(WX2164), .B(II6535), .Z(II6537) ) ;
NAND2   gate12587  (.A(II6536), .B(II6537), .Z(II6534) ) ;
NAND2   gate12588  (.A(II6518), .B(II6534), .Z(II6542) ) ;
NAND2   gate12589  (.A(II6518), .B(II6542), .Z(II6543) ) ;
NAND2   gate12590  (.A(II6534), .B(II6542), .Z(II6544) ) ;
NAND2   gate12591  (.A(WX2295), .B(WX1974), .Z(II6551) ) ;
NAND2   gate12592  (.A(WX2295), .B(II6551), .Z(II6552) ) ;
NAND2   gate12593  (.A(WX1974), .B(II6551), .Z(II6553) ) ;
NAND2   gate12594  (.A(II6552), .B(II6553), .Z(II6550) ) ;
NAND2   gate12595  (.A(WX2038), .B(II6550), .Z(II6558) ) ;
NAND2   gate12596  (.A(WX2038), .B(II6558), .Z(II6559) ) ;
NAND2   gate12597  (.A(II6550), .B(II6558), .Z(II6560) ) ;
NAND2   gate12598  (.A(II6559), .B(II6560), .Z(II6549) ) ;
NAND2   gate12599  (.A(WX2102), .B(WX2166), .Z(II6566) ) ;
NAND2   gate12600  (.A(WX2102), .B(II6566), .Z(II6567) ) ;
NAND2   gate12601  (.A(WX2166), .B(II6566), .Z(II6568) ) ;
NAND2   gate12602  (.A(II6567), .B(II6568), .Z(II6565) ) ;
NAND2   gate12603  (.A(II6549), .B(II6565), .Z(II6573) ) ;
NAND2   gate12604  (.A(II6549), .B(II6573), .Z(II6574) ) ;
NAND2   gate12605  (.A(II6565), .B(II6573), .Z(II6575) ) ;
NAND2   gate12606  (.A(WX2295), .B(WX1976), .Z(II6582) ) ;
NAND2   gate12607  (.A(WX2295), .B(II6582), .Z(II6583) ) ;
NAND2   gate12608  (.A(WX1976), .B(II6582), .Z(II6584) ) ;
NAND2   gate12609  (.A(II6583), .B(II6584), .Z(II6581) ) ;
NAND2   gate12610  (.A(WX2040), .B(II6581), .Z(II6589) ) ;
NAND2   gate12611  (.A(WX2040), .B(II6589), .Z(II6590) ) ;
NAND2   gate12612  (.A(II6581), .B(II6589), .Z(II6591) ) ;
NAND2   gate12613  (.A(II6590), .B(II6591), .Z(II6580) ) ;
NAND2   gate12614  (.A(WX2104), .B(WX2168), .Z(II6597) ) ;
NAND2   gate12615  (.A(WX2104), .B(II6597), .Z(II6598) ) ;
NAND2   gate12616  (.A(WX2168), .B(II6597), .Z(II6599) ) ;
NAND2   gate12617  (.A(II6598), .B(II6599), .Z(II6596) ) ;
NAND2   gate12618  (.A(II6580), .B(II6596), .Z(II6604) ) ;
NAND2   gate12619  (.A(II6580), .B(II6604), .Z(II6605) ) ;
NAND2   gate12620  (.A(II6596), .B(II6604), .Z(II6606) ) ;
NAND2   gate12621  (.A(WX2295), .B(WX1978), .Z(II6613) ) ;
NAND2   gate12622  (.A(WX2295), .B(II6613), .Z(II6614) ) ;
NAND2   gate12623  (.A(WX1978), .B(II6613), .Z(II6615) ) ;
NAND2   gate12624  (.A(II6614), .B(II6615), .Z(II6612) ) ;
NAND2   gate12625  (.A(WX2042), .B(II6612), .Z(II6620) ) ;
NAND2   gate12626  (.A(WX2042), .B(II6620), .Z(II6621) ) ;
NAND2   gate12627  (.A(II6612), .B(II6620), .Z(II6622) ) ;
NAND2   gate12628  (.A(II6621), .B(II6622), .Z(II6611) ) ;
NAND2   gate12629  (.A(WX2106), .B(WX2170), .Z(II6628) ) ;
NAND2   gate12630  (.A(WX2106), .B(II6628), .Z(II6629) ) ;
NAND2   gate12631  (.A(WX2170), .B(II6628), .Z(II6630) ) ;
NAND2   gate12632  (.A(II6629), .B(II6630), .Z(II6627) ) ;
NAND2   gate12633  (.A(II6611), .B(II6627), .Z(II6635) ) ;
NAND2   gate12634  (.A(II6611), .B(II6635), .Z(II6636) ) ;
NAND2   gate12635  (.A(II6627), .B(II6635), .Z(II6637) ) ;
NAND2   gate12636  (.A(WX2295), .B(WX1980), .Z(II6644) ) ;
NAND2   gate12637  (.A(WX2295), .B(II6644), .Z(II6645) ) ;
NAND2   gate12638  (.A(WX1980), .B(II6644), .Z(II6646) ) ;
NAND2   gate12639  (.A(II6645), .B(II6646), .Z(II6643) ) ;
NAND2   gate12640  (.A(WX2044), .B(II6643), .Z(II6651) ) ;
NAND2   gate12641  (.A(WX2044), .B(II6651), .Z(II6652) ) ;
NAND2   gate12642  (.A(II6643), .B(II6651), .Z(II6653) ) ;
NAND2   gate12643  (.A(II6652), .B(II6653), .Z(II6642) ) ;
NAND2   gate12644  (.A(WX2108), .B(WX2172), .Z(II6659) ) ;
NAND2   gate12645  (.A(WX2108), .B(II6659), .Z(II6660) ) ;
NAND2   gate12646  (.A(WX2172), .B(II6659), .Z(II6661) ) ;
NAND2   gate12647  (.A(II6660), .B(II6661), .Z(II6658) ) ;
NAND2   gate12648  (.A(II6642), .B(II6658), .Z(II6666) ) ;
NAND2   gate12649  (.A(II6642), .B(II6666), .Z(II6667) ) ;
NAND2   gate12650  (.A(II6658), .B(II6666), .Z(II6668) ) ;
NAND2   gate12651  (.A(WX2295), .B(WX1982), .Z(II6675) ) ;
NAND2   gate12652  (.A(WX2295), .B(II6675), .Z(II6676) ) ;
NAND2   gate12653  (.A(WX1982), .B(II6675), .Z(II6677) ) ;
NAND2   gate12654  (.A(II6676), .B(II6677), .Z(II6674) ) ;
NAND2   gate12655  (.A(WX2046), .B(II6674), .Z(II6682) ) ;
NAND2   gate12656  (.A(WX2046), .B(II6682), .Z(II6683) ) ;
NAND2   gate12657  (.A(II6674), .B(II6682), .Z(II6684) ) ;
NAND2   gate12658  (.A(II6683), .B(II6684), .Z(II6673) ) ;
NAND2   gate12659  (.A(WX2110), .B(WX2174), .Z(II6690) ) ;
NAND2   gate12660  (.A(WX2110), .B(II6690), .Z(II6691) ) ;
NAND2   gate12661  (.A(WX2174), .B(II6690), .Z(II6692) ) ;
NAND2   gate12662  (.A(II6691), .B(II6692), .Z(II6689) ) ;
NAND2   gate12663  (.A(II6673), .B(II6689), .Z(II6697) ) ;
NAND2   gate12664  (.A(II6673), .B(II6697), .Z(II6698) ) ;
NAND2   gate12665  (.A(II6689), .B(II6697), .Z(II6699) ) ;
NAND2   gate12666  (.A(WX2295), .B(WX1984), .Z(II6706) ) ;
NAND2   gate12667  (.A(WX2295), .B(II6706), .Z(II6707) ) ;
NAND2   gate12668  (.A(WX1984), .B(II6706), .Z(II6708) ) ;
NAND2   gate12669  (.A(II6707), .B(II6708), .Z(II6705) ) ;
NAND2   gate12670  (.A(WX2048), .B(II6705), .Z(II6713) ) ;
NAND2   gate12671  (.A(WX2048), .B(II6713), .Z(II6714) ) ;
NAND2   gate12672  (.A(II6705), .B(II6713), .Z(II6715) ) ;
NAND2   gate12673  (.A(II6714), .B(II6715), .Z(II6704) ) ;
NAND2   gate12674  (.A(WX2112), .B(WX2176), .Z(II6721) ) ;
NAND2   gate12675  (.A(WX2112), .B(II6721), .Z(II6722) ) ;
NAND2   gate12676  (.A(WX2176), .B(II6721), .Z(II6723) ) ;
NAND2   gate12677  (.A(II6722), .B(II6723), .Z(II6720) ) ;
NAND2   gate12678  (.A(II6704), .B(II6720), .Z(II6728) ) ;
NAND2   gate12679  (.A(II6704), .B(II6728), .Z(II6729) ) ;
NAND2   gate12680  (.A(II6720), .B(II6728), .Z(II6730) ) ;
NAND2   gate12681  (.A(WX2295), .B(WX1986), .Z(II6737) ) ;
NAND2   gate12682  (.A(WX2295), .B(II6737), .Z(II6738) ) ;
NAND2   gate12683  (.A(WX1986), .B(II6737), .Z(II6739) ) ;
NAND2   gate12684  (.A(II6738), .B(II6739), .Z(II6736) ) ;
NAND2   gate12685  (.A(WX2050), .B(II6736), .Z(II6744) ) ;
NAND2   gate12686  (.A(WX2050), .B(II6744), .Z(II6745) ) ;
NAND2   gate12687  (.A(II6736), .B(II6744), .Z(II6746) ) ;
NAND2   gate12688  (.A(II6745), .B(II6746), .Z(II6735) ) ;
NAND2   gate12689  (.A(WX2114), .B(WX2178), .Z(II6752) ) ;
NAND2   gate12690  (.A(WX2114), .B(II6752), .Z(II6753) ) ;
NAND2   gate12691  (.A(WX2178), .B(II6752), .Z(II6754) ) ;
NAND2   gate12692  (.A(II6753), .B(II6754), .Z(II6751) ) ;
NAND2   gate12693  (.A(II6735), .B(II6751), .Z(II6759) ) ;
NAND2   gate12694  (.A(II6735), .B(II6759), .Z(II6760) ) ;
NAND2   gate12695  (.A(II6751), .B(II6759), .Z(II6761) ) ;
NAND2   gate12696  (.A(WX2295), .B(WX1988), .Z(II6768) ) ;
NAND2   gate12697  (.A(WX2295), .B(II6768), .Z(II6769) ) ;
NAND2   gate12698  (.A(WX1988), .B(II6768), .Z(II6770) ) ;
NAND2   gate12699  (.A(II6769), .B(II6770), .Z(II6767) ) ;
NAND2   gate12700  (.A(WX2052), .B(II6767), .Z(II6775) ) ;
NAND2   gate12701  (.A(WX2052), .B(II6775), .Z(II6776) ) ;
NAND2   gate12702  (.A(II6767), .B(II6775), .Z(II6777) ) ;
NAND2   gate12703  (.A(II6776), .B(II6777), .Z(II6766) ) ;
NAND2   gate12704  (.A(WX2116), .B(WX2180), .Z(II6783) ) ;
NAND2   gate12705  (.A(WX2116), .B(II6783), .Z(II6784) ) ;
NAND2   gate12706  (.A(WX2180), .B(II6783), .Z(II6785) ) ;
NAND2   gate12707  (.A(II6784), .B(II6785), .Z(II6782) ) ;
NAND2   gate12708  (.A(II6766), .B(II6782), .Z(II6790) ) ;
NAND2   gate12709  (.A(II6766), .B(II6790), .Z(II6791) ) ;
NAND2   gate12710  (.A(II6782), .B(II6790), .Z(II6792) ) ;
NAND2   gate12711  (.A(WX2295), .B(WX1990), .Z(II6799) ) ;
NAND2   gate12712  (.A(WX2295), .B(II6799), .Z(II6800) ) ;
NAND2   gate12713  (.A(WX1990), .B(II6799), .Z(II6801) ) ;
NAND2   gate12714  (.A(II6800), .B(II6801), .Z(II6798) ) ;
NAND2   gate12715  (.A(WX2054), .B(II6798), .Z(II6806) ) ;
NAND2   gate12716  (.A(WX2054), .B(II6806), .Z(II6807) ) ;
NAND2   gate12717  (.A(II6798), .B(II6806), .Z(II6808) ) ;
NAND2   gate12718  (.A(II6807), .B(II6808), .Z(II6797) ) ;
NAND2   gate12719  (.A(WX2118), .B(WX2182), .Z(II6814) ) ;
NAND2   gate12720  (.A(WX2118), .B(II6814), .Z(II6815) ) ;
NAND2   gate12721  (.A(WX2182), .B(II6814), .Z(II6816) ) ;
NAND2   gate12722  (.A(II6815), .B(II6816), .Z(II6813) ) ;
NAND2   gate12723  (.A(II6797), .B(II6813), .Z(II6821) ) ;
NAND2   gate12724  (.A(II6797), .B(II6821), .Z(II6822) ) ;
NAND2   gate12725  (.A(II6813), .B(II6821), .Z(II6823) ) ;
NAND2   gate12726  (.A(WX2295), .B(WX1992), .Z(II6830) ) ;
NAND2   gate12727  (.A(WX2295), .B(II6830), .Z(II6831) ) ;
NAND2   gate12728  (.A(WX1992), .B(II6830), .Z(II6832) ) ;
NAND2   gate12729  (.A(II6831), .B(II6832), .Z(II6829) ) ;
NAND2   gate12730  (.A(WX2056), .B(II6829), .Z(II6837) ) ;
NAND2   gate12731  (.A(WX2056), .B(II6837), .Z(II6838) ) ;
NAND2   gate12732  (.A(II6829), .B(II6837), .Z(II6839) ) ;
NAND2   gate12733  (.A(II6838), .B(II6839), .Z(II6828) ) ;
NAND2   gate12734  (.A(WX2120), .B(WX2184), .Z(II6845) ) ;
NAND2   gate12735  (.A(WX2120), .B(II6845), .Z(II6846) ) ;
NAND2   gate12736  (.A(WX2184), .B(II6845), .Z(II6847) ) ;
NAND2   gate12737  (.A(II6846), .B(II6847), .Z(II6844) ) ;
NAND2   gate12738  (.A(II6828), .B(II6844), .Z(II6852) ) ;
NAND2   gate12739  (.A(II6828), .B(II6852), .Z(II6853) ) ;
NAND2   gate12740  (.A(II6844), .B(II6852), .Z(II6854) ) ;
NAND2   gate12741  (.A(WX2295), .B(WX1994), .Z(II6861) ) ;
NAND2   gate12742  (.A(WX2295), .B(II6861), .Z(II6862) ) ;
NAND2   gate12743  (.A(WX1994), .B(II6861), .Z(II6863) ) ;
NAND2   gate12744  (.A(II6862), .B(II6863), .Z(II6860) ) ;
NAND2   gate12745  (.A(WX2058), .B(II6860), .Z(II6868) ) ;
NAND2   gate12746  (.A(WX2058), .B(II6868), .Z(II6869) ) ;
NAND2   gate12747  (.A(II6860), .B(II6868), .Z(II6870) ) ;
NAND2   gate12748  (.A(II6869), .B(II6870), .Z(II6859) ) ;
NAND2   gate12749  (.A(WX2122), .B(WX2186), .Z(II6876) ) ;
NAND2   gate12750  (.A(WX2122), .B(II6876), .Z(II6877) ) ;
NAND2   gate12751  (.A(WX2186), .B(II6876), .Z(II6878) ) ;
NAND2   gate12752  (.A(II6877), .B(II6878), .Z(II6875) ) ;
NAND2   gate12753  (.A(II6859), .B(II6875), .Z(II6883) ) ;
NAND2   gate12754  (.A(II6859), .B(II6883), .Z(II6884) ) ;
NAND2   gate12755  (.A(II6875), .B(II6883), .Z(II6885) ) ;
NAND2   gate12756  (.A(WX2295), .B(WX1996), .Z(II6892) ) ;
NAND2   gate12757  (.A(WX2295), .B(II6892), .Z(II6893) ) ;
NAND2   gate12758  (.A(WX1996), .B(II6892), .Z(II6894) ) ;
NAND2   gate12759  (.A(II6893), .B(II6894), .Z(II6891) ) ;
NAND2   gate12760  (.A(WX2060), .B(II6891), .Z(II6899) ) ;
NAND2   gate12761  (.A(WX2060), .B(II6899), .Z(II6900) ) ;
NAND2   gate12762  (.A(II6891), .B(II6899), .Z(II6901) ) ;
NAND2   gate12763  (.A(II6900), .B(II6901), .Z(II6890) ) ;
NAND2   gate12764  (.A(WX2124), .B(WX2188), .Z(II6907) ) ;
NAND2   gate12765  (.A(WX2124), .B(II6907), .Z(II6908) ) ;
NAND2   gate12766  (.A(WX2188), .B(II6907), .Z(II6909) ) ;
NAND2   gate12767  (.A(II6908), .B(II6909), .Z(II6906) ) ;
NAND2   gate12768  (.A(II6890), .B(II6906), .Z(II6914) ) ;
NAND2   gate12769  (.A(II6890), .B(II6914), .Z(II6915) ) ;
NAND2   gate12770  (.A(II6906), .B(II6914), .Z(II6916) ) ;
NAND2   gate12771  (.A(WX2295), .B(WX1998), .Z(II6923) ) ;
NAND2   gate12772  (.A(WX2295), .B(II6923), .Z(II6924) ) ;
NAND2   gate12773  (.A(WX1998), .B(II6923), .Z(II6925) ) ;
NAND2   gate12774  (.A(II6924), .B(II6925), .Z(II6922) ) ;
NAND2   gate12775  (.A(WX2062), .B(II6922), .Z(II6930) ) ;
NAND2   gate12776  (.A(WX2062), .B(II6930), .Z(II6931) ) ;
NAND2   gate12777  (.A(II6922), .B(II6930), .Z(II6932) ) ;
NAND2   gate12778  (.A(II6931), .B(II6932), .Z(II6921) ) ;
NAND2   gate12779  (.A(WX2126), .B(WX2190), .Z(II6938) ) ;
NAND2   gate12780  (.A(WX2126), .B(II6938), .Z(II6939) ) ;
NAND2   gate12781  (.A(WX2190), .B(II6938), .Z(II6940) ) ;
NAND2   gate12782  (.A(II6939), .B(II6940), .Z(II6937) ) ;
NAND2   gate12783  (.A(II6921), .B(II6937), .Z(II6945) ) ;
NAND2   gate12784  (.A(II6921), .B(II6945), .Z(II6946) ) ;
NAND2   gate12785  (.A(II6937), .B(II6945), .Z(II6947) ) ;
NAND2   gate12786  (.A(WX2295), .B(WX2000), .Z(II6954) ) ;
NAND2   gate12787  (.A(WX2295), .B(II6954), .Z(II6955) ) ;
NAND2   gate12788  (.A(WX2000), .B(II6954), .Z(II6956) ) ;
NAND2   gate12789  (.A(II6955), .B(II6956), .Z(II6953) ) ;
NAND2   gate12790  (.A(WX2064), .B(II6953), .Z(II6961) ) ;
NAND2   gate12791  (.A(WX2064), .B(II6961), .Z(II6962) ) ;
NAND2   gate12792  (.A(II6953), .B(II6961), .Z(II6963) ) ;
NAND2   gate12793  (.A(II6962), .B(II6963), .Z(II6952) ) ;
NAND2   gate12794  (.A(WX2128), .B(WX2192), .Z(II6969) ) ;
NAND2   gate12795  (.A(WX2128), .B(II6969), .Z(II6970) ) ;
NAND2   gate12796  (.A(WX2192), .B(II6969), .Z(II6971) ) ;
NAND2   gate12797  (.A(II6970), .B(II6971), .Z(II6968) ) ;
NAND2   gate12798  (.A(II6952), .B(II6968), .Z(II6976) ) ;
NAND2   gate12799  (.A(II6952), .B(II6976), .Z(II6977) ) ;
NAND2   gate12800  (.A(II6968), .B(II6976), .Z(II6978) ) ;
NAND2   gate12801  (.A(WX1873), .B(WX1778), .Z(II7057) ) ;
NAND2   gate12802  (.A(WX1873), .B(II7057), .Z(II7058) ) ;
NAND2   gate12803  (.A(WX1778), .B(II7057), .Z(II7059) ) ;
NAND2   gate12804  (.A(WX1874), .B(WX1780), .Z(II7070) ) ;
NAND2   gate12805  (.A(WX1874), .B(II7070), .Z(II7071) ) ;
NAND2   gate12806  (.A(WX1780), .B(II7070), .Z(II7072) ) ;
NAND2   gate12807  (.A(WX1875), .B(WX1782), .Z(II7083) ) ;
NAND2   gate12808  (.A(WX1875), .B(II7083), .Z(II7084) ) ;
NAND2   gate12809  (.A(WX1782), .B(II7083), .Z(II7085) ) ;
NAND2   gate12810  (.A(WX1876), .B(WX1784), .Z(II7096) ) ;
NAND2   gate12811  (.A(WX1876), .B(II7096), .Z(II7097) ) ;
NAND2   gate12812  (.A(WX1784), .B(II7096), .Z(II7098) ) ;
NAND2   gate12813  (.A(WX1877), .B(WX1786), .Z(II7109) ) ;
NAND2   gate12814  (.A(WX1877), .B(II7109), .Z(II7110) ) ;
NAND2   gate12815  (.A(WX1786), .B(II7109), .Z(II7111) ) ;
NAND2   gate12816  (.A(WX1878), .B(WX1788), .Z(II7122) ) ;
NAND2   gate12817  (.A(WX1878), .B(II7122), .Z(II7123) ) ;
NAND2   gate12818  (.A(WX1788), .B(II7122), .Z(II7124) ) ;
NAND2   gate12819  (.A(WX1879), .B(WX1790), .Z(II7135) ) ;
NAND2   gate12820  (.A(WX1879), .B(II7135), .Z(II7136) ) ;
NAND2   gate12821  (.A(WX1790), .B(II7135), .Z(II7137) ) ;
NAND2   gate12822  (.A(WX1880), .B(WX1792), .Z(II7148) ) ;
NAND2   gate12823  (.A(WX1880), .B(II7148), .Z(II7149) ) ;
NAND2   gate12824  (.A(WX1792), .B(II7148), .Z(II7150) ) ;
NAND2   gate12825  (.A(WX1881), .B(WX1794), .Z(II7161) ) ;
NAND2   gate12826  (.A(WX1881), .B(II7161), .Z(II7162) ) ;
NAND2   gate12827  (.A(WX1794), .B(II7161), .Z(II7163) ) ;
NAND2   gate12828  (.A(WX1882), .B(WX1796), .Z(II7174) ) ;
NAND2   gate12829  (.A(WX1882), .B(II7174), .Z(II7175) ) ;
NAND2   gate12830  (.A(WX1796), .B(II7174), .Z(II7176) ) ;
NAND2   gate12831  (.A(WX1883), .B(WX1798), .Z(II7187) ) ;
NAND2   gate12832  (.A(WX1883), .B(II7187), .Z(II7188) ) ;
NAND2   gate12833  (.A(WX1798), .B(II7187), .Z(II7189) ) ;
NAND2   gate12834  (.A(WX1884), .B(WX1800), .Z(II7200) ) ;
NAND2   gate12835  (.A(WX1884), .B(II7200), .Z(II7201) ) ;
NAND2   gate12836  (.A(WX1800), .B(II7200), .Z(II7202) ) ;
NAND2   gate12837  (.A(WX1885), .B(WX1802), .Z(II7213) ) ;
NAND2   gate12838  (.A(WX1885), .B(II7213), .Z(II7214) ) ;
NAND2   gate12839  (.A(WX1802), .B(II7213), .Z(II7215) ) ;
NAND2   gate12840  (.A(WX1886), .B(WX1804), .Z(II7226) ) ;
NAND2   gate12841  (.A(WX1886), .B(II7226), .Z(II7227) ) ;
NAND2   gate12842  (.A(WX1804), .B(II7226), .Z(II7228) ) ;
NAND2   gate12843  (.A(WX1887), .B(WX1806), .Z(II7239) ) ;
NAND2   gate12844  (.A(WX1887), .B(II7239), .Z(II7240) ) ;
NAND2   gate12845  (.A(WX1806), .B(II7239), .Z(II7241) ) ;
NAND2   gate12846  (.A(WX1888), .B(WX1808), .Z(II7252) ) ;
NAND2   gate12847  (.A(WX1888), .B(II7252), .Z(II7253) ) ;
NAND2   gate12848  (.A(WX1808), .B(II7252), .Z(II7254) ) ;
NAND2   gate12849  (.A(WX1889), .B(WX1810), .Z(II7265) ) ;
NAND2   gate12850  (.A(WX1889), .B(II7265), .Z(II7266) ) ;
NAND2   gate12851  (.A(WX1810), .B(II7265), .Z(II7267) ) ;
NAND2   gate12852  (.A(WX1890), .B(WX1812), .Z(II7278) ) ;
NAND2   gate12853  (.A(WX1890), .B(II7278), .Z(II7279) ) ;
NAND2   gate12854  (.A(WX1812), .B(II7278), .Z(II7280) ) ;
NAND2   gate12855  (.A(WX1891), .B(WX1814), .Z(II7291) ) ;
NAND2   gate12856  (.A(WX1891), .B(II7291), .Z(II7292) ) ;
NAND2   gate12857  (.A(WX1814), .B(II7291), .Z(II7293) ) ;
NAND2   gate12858  (.A(WX1892), .B(WX1816), .Z(II7304) ) ;
NAND2   gate12859  (.A(WX1892), .B(II7304), .Z(II7305) ) ;
NAND2   gate12860  (.A(WX1816), .B(II7304), .Z(II7306) ) ;
NAND2   gate12861  (.A(WX1893), .B(WX1818), .Z(II7317) ) ;
NAND2   gate12862  (.A(WX1893), .B(II7317), .Z(II7318) ) ;
NAND2   gate12863  (.A(WX1818), .B(II7317), .Z(II7319) ) ;
NAND2   gate12864  (.A(WX1894), .B(WX1820), .Z(II7330) ) ;
NAND2   gate12865  (.A(WX1894), .B(II7330), .Z(II7331) ) ;
NAND2   gate12866  (.A(WX1820), .B(II7330), .Z(II7332) ) ;
NAND2   gate12867  (.A(WX1895), .B(WX1822), .Z(II7343) ) ;
NAND2   gate12868  (.A(WX1895), .B(II7343), .Z(II7344) ) ;
NAND2   gate12869  (.A(WX1822), .B(II7343), .Z(II7345) ) ;
NAND2   gate12870  (.A(WX1896), .B(WX1824), .Z(II7356) ) ;
NAND2   gate12871  (.A(WX1896), .B(II7356), .Z(II7357) ) ;
NAND2   gate12872  (.A(WX1824), .B(II7356), .Z(II7358) ) ;
NAND2   gate12873  (.A(WX1897), .B(WX1826), .Z(II7369) ) ;
NAND2   gate12874  (.A(WX1897), .B(II7369), .Z(II7370) ) ;
NAND2   gate12875  (.A(WX1826), .B(II7369), .Z(II7371) ) ;
NAND2   gate12876  (.A(WX1898), .B(WX1828), .Z(II7382) ) ;
NAND2   gate12877  (.A(WX1898), .B(II7382), .Z(II7383) ) ;
NAND2   gate12878  (.A(WX1828), .B(II7382), .Z(II7384) ) ;
NAND2   gate12879  (.A(WX1899), .B(WX1830), .Z(II7395) ) ;
NAND2   gate12880  (.A(WX1899), .B(II7395), .Z(II7396) ) ;
NAND2   gate12881  (.A(WX1830), .B(II7395), .Z(II7397) ) ;
NAND2   gate12882  (.A(WX1900), .B(WX1832), .Z(II7408) ) ;
NAND2   gate12883  (.A(WX1900), .B(II7408), .Z(II7409) ) ;
NAND2   gate12884  (.A(WX1832), .B(II7408), .Z(II7410) ) ;
NAND2   gate12885  (.A(WX1901), .B(WX1834), .Z(II7421) ) ;
NAND2   gate12886  (.A(WX1901), .B(II7421), .Z(II7422) ) ;
NAND2   gate12887  (.A(WX1834), .B(II7421), .Z(II7423) ) ;
NAND2   gate12888  (.A(WX1902), .B(WX1836), .Z(II7434) ) ;
NAND2   gate12889  (.A(WX1902), .B(II7434), .Z(II7435) ) ;
NAND2   gate12890  (.A(WX1836), .B(II7434), .Z(II7436) ) ;
NAND2   gate12891  (.A(WX1903), .B(WX1838), .Z(II7447) ) ;
NAND2   gate12892  (.A(WX1903), .B(II7447), .Z(II7448) ) ;
NAND2   gate12893  (.A(WX1838), .B(II7447), .Z(II7449) ) ;
NAND2   gate12894  (.A(WX1904), .B(WX1840), .Z(II7460) ) ;
NAND2   gate12895  (.A(WX1904), .B(II7460), .Z(II7461) ) ;
NAND2   gate12896  (.A(WX1840), .B(II7460), .Z(II7462) ) ;
NAND2   gate12897  (.A(WX1920), .B(CRC_OUT_8_31), .Z(II7475) ) ;
NAND2   gate12898  (.A(WX1920), .B(II7475), .Z(II7476) ) ;
NAND2   gate12899  (.A(CRC_OUT_8_31), .B(II7475), .Z(II7477) ) ;
NAND2   gate12900  (.A(II7476), .B(II7477), .Z(II7474) ) ;
NAND2   gate12901  (.A(CRC_OUT_8_15), .B(II7474), .Z(II7482) ) ;
NAND2   gate12902  (.A(CRC_OUT_8_15), .B(II7482), .Z(II7483) ) ;
NAND2   gate12903  (.A(II7474), .B(II7482), .Z(II7484) ) ;
NAND2   gate12904  (.A(WX1925), .B(CRC_OUT_8_31), .Z(II7490) ) ;
NAND2   gate12905  (.A(WX1925), .B(II7490), .Z(II7491) ) ;
NAND2   gate12906  (.A(CRC_OUT_8_31), .B(II7490), .Z(II7492) ) ;
NAND2   gate12907  (.A(II7491), .B(II7492), .Z(II7489) ) ;
NAND2   gate12908  (.A(CRC_OUT_8_10), .B(II7489), .Z(II7497) ) ;
NAND2   gate12909  (.A(CRC_OUT_8_10), .B(II7497), .Z(II7498) ) ;
NAND2   gate12910  (.A(II7489), .B(II7497), .Z(II7499) ) ;
NAND2   gate12911  (.A(WX1932), .B(CRC_OUT_8_31), .Z(II7505) ) ;
NAND2   gate12912  (.A(WX1932), .B(II7505), .Z(II7506) ) ;
NAND2   gate12913  (.A(CRC_OUT_8_31), .B(II7505), .Z(II7507) ) ;
NAND2   gate12914  (.A(II7506), .B(II7507), .Z(II7504) ) ;
NAND2   gate12915  (.A(CRC_OUT_8_3), .B(II7504), .Z(II7512) ) ;
NAND2   gate12916  (.A(CRC_OUT_8_3), .B(II7512), .Z(II7513) ) ;
NAND2   gate12917  (.A(II7504), .B(II7512), .Z(II7514) ) ;
NAND2   gate12918  (.A(WX1936), .B(CRC_OUT_8_31), .Z(II7519) ) ;
NAND2   gate12919  (.A(WX1936), .B(II7519), .Z(II7520) ) ;
NAND2   gate12920  (.A(CRC_OUT_8_31), .B(II7519), .Z(II7521) ) ;
NAND2   gate12921  (.A(WX1905), .B(CRC_OUT_8_30), .Z(II7526) ) ;
NAND2   gate12922  (.A(WX1905), .B(II7526), .Z(II7527) ) ;
NAND2   gate12923  (.A(CRC_OUT_8_30), .B(II7526), .Z(II7528) ) ;
NAND2   gate12924  (.A(WX1906), .B(CRC_OUT_8_29), .Z(II7533) ) ;
NAND2   gate12925  (.A(WX1906), .B(II7533), .Z(II7534) ) ;
NAND2   gate12926  (.A(CRC_OUT_8_29), .B(II7533), .Z(II7535) ) ;
NAND2   gate12927  (.A(WX1907), .B(CRC_OUT_8_28), .Z(II7540) ) ;
NAND2   gate12928  (.A(WX1907), .B(II7540), .Z(II7541) ) ;
NAND2   gate12929  (.A(CRC_OUT_8_28), .B(II7540), .Z(II7542) ) ;
NAND2   gate12930  (.A(WX1908), .B(CRC_OUT_8_27), .Z(II7547) ) ;
NAND2   gate12931  (.A(WX1908), .B(II7547), .Z(II7548) ) ;
NAND2   gate12932  (.A(CRC_OUT_8_27), .B(II7547), .Z(II7549) ) ;
NAND2   gate12933  (.A(WX1909), .B(CRC_OUT_8_26), .Z(II7554) ) ;
NAND2   gate12934  (.A(WX1909), .B(II7554), .Z(II7555) ) ;
NAND2   gate12935  (.A(CRC_OUT_8_26), .B(II7554), .Z(II7556) ) ;
NAND2   gate12936  (.A(WX1910), .B(CRC_OUT_8_25), .Z(II7561) ) ;
NAND2   gate12937  (.A(WX1910), .B(II7561), .Z(II7562) ) ;
NAND2   gate12938  (.A(CRC_OUT_8_25), .B(II7561), .Z(II7563) ) ;
NAND2   gate12939  (.A(WX1911), .B(CRC_OUT_8_24), .Z(II7568) ) ;
NAND2   gate12940  (.A(WX1911), .B(II7568), .Z(II7569) ) ;
NAND2   gate12941  (.A(CRC_OUT_8_24), .B(II7568), .Z(II7570) ) ;
NAND2   gate12942  (.A(WX1912), .B(CRC_OUT_8_23), .Z(II7575) ) ;
NAND2   gate12943  (.A(WX1912), .B(II7575), .Z(II7576) ) ;
NAND2   gate12944  (.A(CRC_OUT_8_23), .B(II7575), .Z(II7577) ) ;
NAND2   gate12945  (.A(WX1913), .B(CRC_OUT_8_22), .Z(II7582) ) ;
NAND2   gate12946  (.A(WX1913), .B(II7582), .Z(II7583) ) ;
NAND2   gate12947  (.A(CRC_OUT_8_22), .B(II7582), .Z(II7584) ) ;
NAND2   gate12948  (.A(WX1914), .B(CRC_OUT_8_21), .Z(II7589) ) ;
NAND2   gate12949  (.A(WX1914), .B(II7589), .Z(II7590) ) ;
NAND2   gate12950  (.A(CRC_OUT_8_21), .B(II7589), .Z(II7591) ) ;
NAND2   gate12951  (.A(WX1915), .B(CRC_OUT_8_20), .Z(II7596) ) ;
NAND2   gate12952  (.A(WX1915), .B(II7596), .Z(II7597) ) ;
NAND2   gate12953  (.A(CRC_OUT_8_20), .B(II7596), .Z(II7598) ) ;
NAND2   gate12954  (.A(WX1916), .B(CRC_OUT_8_19), .Z(II7603) ) ;
NAND2   gate12955  (.A(WX1916), .B(II7603), .Z(II7604) ) ;
NAND2   gate12956  (.A(CRC_OUT_8_19), .B(II7603), .Z(II7605) ) ;
NAND2   gate12957  (.A(WX1917), .B(CRC_OUT_8_18), .Z(II7610) ) ;
NAND2   gate12958  (.A(WX1917), .B(II7610), .Z(II7611) ) ;
NAND2   gate12959  (.A(CRC_OUT_8_18), .B(II7610), .Z(II7612) ) ;
NAND2   gate12960  (.A(WX1918), .B(CRC_OUT_8_17), .Z(II7617) ) ;
NAND2   gate12961  (.A(WX1918), .B(II7617), .Z(II7618) ) ;
NAND2   gate12962  (.A(CRC_OUT_8_17), .B(II7617), .Z(II7619) ) ;
NAND2   gate12963  (.A(WX1919), .B(CRC_OUT_8_16), .Z(II7624) ) ;
NAND2   gate12964  (.A(WX1919), .B(II7624), .Z(II7625) ) ;
NAND2   gate12965  (.A(CRC_OUT_8_16), .B(II7624), .Z(II7626) ) ;
NAND2   gate12966  (.A(WX1921), .B(CRC_OUT_8_14), .Z(II7631) ) ;
NAND2   gate12967  (.A(WX1921), .B(II7631), .Z(II7632) ) ;
NAND2   gate12968  (.A(CRC_OUT_8_14), .B(II7631), .Z(II7633) ) ;
NAND2   gate12969  (.A(WX1922), .B(CRC_OUT_8_13), .Z(II7638) ) ;
NAND2   gate12970  (.A(WX1922), .B(II7638), .Z(II7639) ) ;
NAND2   gate12971  (.A(CRC_OUT_8_13), .B(II7638), .Z(II7640) ) ;
NAND2   gate12972  (.A(WX1923), .B(CRC_OUT_8_12), .Z(II7645) ) ;
NAND2   gate12973  (.A(WX1923), .B(II7645), .Z(II7646) ) ;
NAND2   gate12974  (.A(CRC_OUT_8_12), .B(II7645), .Z(II7647) ) ;
NAND2   gate12975  (.A(WX1924), .B(CRC_OUT_8_11), .Z(II7652) ) ;
NAND2   gate12976  (.A(WX1924), .B(II7652), .Z(II7653) ) ;
NAND2   gate12977  (.A(CRC_OUT_8_11), .B(II7652), .Z(II7654) ) ;
NAND2   gate12978  (.A(WX1926), .B(CRC_OUT_8_9), .Z(II7659) ) ;
NAND2   gate12979  (.A(WX1926), .B(II7659), .Z(II7660) ) ;
NAND2   gate12980  (.A(CRC_OUT_8_9), .B(II7659), .Z(II7661) ) ;
NAND2   gate12981  (.A(WX1927), .B(CRC_OUT_8_8), .Z(II7666) ) ;
NAND2   gate12982  (.A(WX1927), .B(II7666), .Z(II7667) ) ;
NAND2   gate12983  (.A(CRC_OUT_8_8), .B(II7666), .Z(II7668) ) ;
NAND2   gate12984  (.A(WX1928), .B(CRC_OUT_8_7), .Z(II7673) ) ;
NAND2   gate12985  (.A(WX1928), .B(II7673), .Z(II7674) ) ;
NAND2   gate12986  (.A(CRC_OUT_8_7), .B(II7673), .Z(II7675) ) ;
NAND2   gate12987  (.A(WX1929), .B(CRC_OUT_8_6), .Z(II7680) ) ;
NAND2   gate12988  (.A(WX1929), .B(II7680), .Z(II7681) ) ;
NAND2   gate12989  (.A(CRC_OUT_8_6), .B(II7680), .Z(II7682) ) ;
NAND2   gate12990  (.A(WX1930), .B(CRC_OUT_8_5), .Z(II7687) ) ;
NAND2   gate12991  (.A(WX1930), .B(II7687), .Z(II7688) ) ;
NAND2   gate12992  (.A(CRC_OUT_8_5), .B(II7687), .Z(II7689) ) ;
NAND2   gate12993  (.A(WX1931), .B(CRC_OUT_8_4), .Z(II7694) ) ;
NAND2   gate12994  (.A(WX1931), .B(II7694), .Z(II7695) ) ;
NAND2   gate12995  (.A(CRC_OUT_8_4), .B(II7694), .Z(II7696) ) ;
NAND2   gate12996  (.A(WX1933), .B(CRC_OUT_8_2), .Z(II7701) ) ;
NAND2   gate12997  (.A(WX1933), .B(II7701), .Z(II7702) ) ;
NAND2   gate12998  (.A(CRC_OUT_8_2), .B(II7701), .Z(II7703) ) ;
NAND2   gate12999  (.A(WX1934), .B(CRC_OUT_8_1), .Z(II7708) ) ;
NAND2   gate13000  (.A(WX1934), .B(II7708), .Z(II7709) ) ;
NAND2   gate13001  (.A(CRC_OUT_8_1), .B(II7708), .Z(II7710) ) ;
NAND2   gate13002  (.A(WX1935), .B(CRC_OUT_8_0), .Z(II7715) ) ;
NAND2   gate13003  (.A(WX1935), .B(II7715), .Z(II7716) ) ;
NAND2   gate13004  (.A(CRC_OUT_8_0), .B(II7715), .Z(II7717) ) ;
NAND2   gate13005  (.A(WX3587), .B(WX3231), .Z(II9998) ) ;
NAND2   gate13006  (.A(WX3587), .B(II9998), .Z(II9999) ) ;
NAND2   gate13007  (.A(WX3231), .B(II9998), .Z(II10000) ) ;
NAND2   gate13008  (.A(II9999), .B(II10000), .Z(II9997) ) ;
NAND2   gate13009  (.A(WX3295), .B(II9997), .Z(II10005) ) ;
NAND2   gate13010  (.A(WX3295), .B(II10005), .Z(II10006) ) ;
NAND2   gate13011  (.A(II9997), .B(II10005), .Z(II10007) ) ;
NAND2   gate13012  (.A(II10006), .B(II10007), .Z(II9996) ) ;
NAND2   gate13013  (.A(WX3359), .B(WX3423), .Z(II10013) ) ;
NAND2   gate13014  (.A(WX3359), .B(II10013), .Z(II10014) ) ;
NAND2   gate13015  (.A(WX3423), .B(II10013), .Z(II10015) ) ;
NAND2   gate13016  (.A(II10014), .B(II10015), .Z(II10012) ) ;
NAND2   gate13017  (.A(II9996), .B(II10012), .Z(II10020) ) ;
NAND2   gate13018  (.A(II9996), .B(II10020), .Z(II10021) ) ;
NAND2   gate13019  (.A(II10012), .B(II10020), .Z(II10022) ) ;
NAND2   gate13020  (.A(WX3587), .B(WX3233), .Z(II10029) ) ;
NAND2   gate13021  (.A(WX3587), .B(II10029), .Z(II10030) ) ;
NAND2   gate13022  (.A(WX3233), .B(II10029), .Z(II10031) ) ;
NAND2   gate13023  (.A(II10030), .B(II10031), .Z(II10028) ) ;
NAND2   gate13024  (.A(WX3297), .B(II10028), .Z(II10036) ) ;
NAND2   gate13025  (.A(WX3297), .B(II10036), .Z(II10037) ) ;
NAND2   gate13026  (.A(II10028), .B(II10036), .Z(II10038) ) ;
NAND2   gate13027  (.A(II10037), .B(II10038), .Z(II10027) ) ;
NAND2   gate13028  (.A(WX3361), .B(WX3425), .Z(II10044) ) ;
NAND2   gate13029  (.A(WX3361), .B(II10044), .Z(II10045) ) ;
NAND2   gate13030  (.A(WX3425), .B(II10044), .Z(II10046) ) ;
NAND2   gate13031  (.A(II10045), .B(II10046), .Z(II10043) ) ;
NAND2   gate13032  (.A(II10027), .B(II10043), .Z(II10051) ) ;
NAND2   gate13033  (.A(II10027), .B(II10051), .Z(II10052) ) ;
NAND2   gate13034  (.A(II10043), .B(II10051), .Z(II10053) ) ;
NAND2   gate13035  (.A(WX3587), .B(WX3235), .Z(II10060) ) ;
NAND2   gate13036  (.A(WX3587), .B(II10060), .Z(II10061) ) ;
NAND2   gate13037  (.A(WX3235), .B(II10060), .Z(II10062) ) ;
NAND2   gate13038  (.A(II10061), .B(II10062), .Z(II10059) ) ;
NAND2   gate13039  (.A(WX3299), .B(II10059), .Z(II10067) ) ;
NAND2   gate13040  (.A(WX3299), .B(II10067), .Z(II10068) ) ;
NAND2   gate13041  (.A(II10059), .B(II10067), .Z(II10069) ) ;
NAND2   gate13042  (.A(II10068), .B(II10069), .Z(II10058) ) ;
NAND2   gate13043  (.A(WX3363), .B(WX3427), .Z(II10075) ) ;
NAND2   gate13044  (.A(WX3363), .B(II10075), .Z(II10076) ) ;
NAND2   gate13045  (.A(WX3427), .B(II10075), .Z(II10077) ) ;
NAND2   gate13046  (.A(II10076), .B(II10077), .Z(II10074) ) ;
NAND2   gate13047  (.A(II10058), .B(II10074), .Z(II10082) ) ;
NAND2   gate13048  (.A(II10058), .B(II10082), .Z(II10083) ) ;
NAND2   gate13049  (.A(II10074), .B(II10082), .Z(II10084) ) ;
NAND2   gate13050  (.A(WX3587), .B(WX3237), .Z(II10091) ) ;
NAND2   gate13051  (.A(WX3587), .B(II10091), .Z(II10092) ) ;
NAND2   gate13052  (.A(WX3237), .B(II10091), .Z(II10093) ) ;
NAND2   gate13053  (.A(II10092), .B(II10093), .Z(II10090) ) ;
NAND2   gate13054  (.A(WX3301), .B(II10090), .Z(II10098) ) ;
NAND2   gate13055  (.A(WX3301), .B(II10098), .Z(II10099) ) ;
NAND2   gate13056  (.A(II10090), .B(II10098), .Z(II10100) ) ;
NAND2   gate13057  (.A(II10099), .B(II10100), .Z(II10089) ) ;
NAND2   gate13058  (.A(WX3365), .B(WX3429), .Z(II10106) ) ;
NAND2   gate13059  (.A(WX3365), .B(II10106), .Z(II10107) ) ;
NAND2   gate13060  (.A(WX3429), .B(II10106), .Z(II10108) ) ;
NAND2   gate13061  (.A(II10107), .B(II10108), .Z(II10105) ) ;
NAND2   gate13062  (.A(II10089), .B(II10105), .Z(II10113) ) ;
NAND2   gate13063  (.A(II10089), .B(II10113), .Z(II10114) ) ;
NAND2   gate13064  (.A(II10105), .B(II10113), .Z(II10115) ) ;
NAND2   gate13065  (.A(WX3587), .B(WX3239), .Z(II10122) ) ;
NAND2   gate13066  (.A(WX3587), .B(II10122), .Z(II10123) ) ;
NAND2   gate13067  (.A(WX3239), .B(II10122), .Z(II10124) ) ;
NAND2   gate13068  (.A(II10123), .B(II10124), .Z(II10121) ) ;
NAND2   gate13069  (.A(WX3303), .B(II10121), .Z(II10129) ) ;
NAND2   gate13070  (.A(WX3303), .B(II10129), .Z(II10130) ) ;
NAND2   gate13071  (.A(II10121), .B(II10129), .Z(II10131) ) ;
NAND2   gate13072  (.A(II10130), .B(II10131), .Z(II10120) ) ;
NAND2   gate13073  (.A(WX3367), .B(WX3431), .Z(II10137) ) ;
NAND2   gate13074  (.A(WX3367), .B(II10137), .Z(II10138) ) ;
NAND2   gate13075  (.A(WX3431), .B(II10137), .Z(II10139) ) ;
NAND2   gate13076  (.A(II10138), .B(II10139), .Z(II10136) ) ;
NAND2   gate13077  (.A(II10120), .B(II10136), .Z(II10144) ) ;
NAND2   gate13078  (.A(II10120), .B(II10144), .Z(II10145) ) ;
NAND2   gate13079  (.A(II10136), .B(II10144), .Z(II10146) ) ;
NAND2   gate13080  (.A(WX3587), .B(WX3241), .Z(II10153) ) ;
NAND2   gate13081  (.A(WX3587), .B(II10153), .Z(II10154) ) ;
NAND2   gate13082  (.A(WX3241), .B(II10153), .Z(II10155) ) ;
NAND2   gate13083  (.A(II10154), .B(II10155), .Z(II10152) ) ;
NAND2   gate13084  (.A(WX3305), .B(II10152), .Z(II10160) ) ;
NAND2   gate13085  (.A(WX3305), .B(II10160), .Z(II10161) ) ;
NAND2   gate13086  (.A(II10152), .B(II10160), .Z(II10162) ) ;
NAND2   gate13087  (.A(II10161), .B(II10162), .Z(II10151) ) ;
NAND2   gate13088  (.A(WX3369), .B(WX3433), .Z(II10168) ) ;
NAND2   gate13089  (.A(WX3369), .B(II10168), .Z(II10169) ) ;
NAND2   gate13090  (.A(WX3433), .B(II10168), .Z(II10170) ) ;
NAND2   gate13091  (.A(II10169), .B(II10170), .Z(II10167) ) ;
NAND2   gate13092  (.A(II10151), .B(II10167), .Z(II10175) ) ;
NAND2   gate13093  (.A(II10151), .B(II10175), .Z(II10176) ) ;
NAND2   gate13094  (.A(II10167), .B(II10175), .Z(II10177) ) ;
NAND2   gate13095  (.A(WX3587), .B(WX3243), .Z(II10184) ) ;
NAND2   gate13096  (.A(WX3587), .B(II10184), .Z(II10185) ) ;
NAND2   gate13097  (.A(WX3243), .B(II10184), .Z(II10186) ) ;
NAND2   gate13098  (.A(II10185), .B(II10186), .Z(II10183) ) ;
NAND2   gate13099  (.A(WX3307), .B(II10183), .Z(II10191) ) ;
NAND2   gate13100  (.A(WX3307), .B(II10191), .Z(II10192) ) ;
NAND2   gate13101  (.A(II10183), .B(II10191), .Z(II10193) ) ;
NAND2   gate13102  (.A(II10192), .B(II10193), .Z(II10182) ) ;
NAND2   gate13103  (.A(WX3371), .B(WX3435), .Z(II10199) ) ;
NAND2   gate13104  (.A(WX3371), .B(II10199), .Z(II10200) ) ;
NAND2   gate13105  (.A(WX3435), .B(II10199), .Z(II10201) ) ;
NAND2   gate13106  (.A(II10200), .B(II10201), .Z(II10198) ) ;
NAND2   gate13107  (.A(II10182), .B(II10198), .Z(II10206) ) ;
NAND2   gate13108  (.A(II10182), .B(II10206), .Z(II10207) ) ;
NAND2   gate13109  (.A(II10198), .B(II10206), .Z(II10208) ) ;
NAND2   gate13110  (.A(WX3587), .B(WX3245), .Z(II10215) ) ;
NAND2   gate13111  (.A(WX3587), .B(II10215), .Z(II10216) ) ;
NAND2   gate13112  (.A(WX3245), .B(II10215), .Z(II10217) ) ;
NAND2   gate13113  (.A(II10216), .B(II10217), .Z(II10214) ) ;
NAND2   gate13114  (.A(WX3309), .B(II10214), .Z(II10222) ) ;
NAND2   gate13115  (.A(WX3309), .B(II10222), .Z(II10223) ) ;
NAND2   gate13116  (.A(II10214), .B(II10222), .Z(II10224) ) ;
NAND2   gate13117  (.A(II10223), .B(II10224), .Z(II10213) ) ;
NAND2   gate13118  (.A(WX3373), .B(WX3437), .Z(II10230) ) ;
NAND2   gate13119  (.A(WX3373), .B(II10230), .Z(II10231) ) ;
NAND2   gate13120  (.A(WX3437), .B(II10230), .Z(II10232) ) ;
NAND2   gate13121  (.A(II10231), .B(II10232), .Z(II10229) ) ;
NAND2   gate13122  (.A(II10213), .B(II10229), .Z(II10237) ) ;
NAND2   gate13123  (.A(II10213), .B(II10237), .Z(II10238) ) ;
NAND2   gate13124  (.A(II10229), .B(II10237), .Z(II10239) ) ;
NAND2   gate13125  (.A(WX3587), .B(WX3247), .Z(II10246) ) ;
NAND2   gate13126  (.A(WX3587), .B(II10246), .Z(II10247) ) ;
NAND2   gate13127  (.A(WX3247), .B(II10246), .Z(II10248) ) ;
NAND2   gate13128  (.A(II10247), .B(II10248), .Z(II10245) ) ;
NAND2   gate13129  (.A(WX3311), .B(II10245), .Z(II10253) ) ;
NAND2   gate13130  (.A(WX3311), .B(II10253), .Z(II10254) ) ;
NAND2   gate13131  (.A(II10245), .B(II10253), .Z(II10255) ) ;
NAND2   gate13132  (.A(II10254), .B(II10255), .Z(II10244) ) ;
NAND2   gate13133  (.A(WX3375), .B(WX3439), .Z(II10261) ) ;
NAND2   gate13134  (.A(WX3375), .B(II10261), .Z(II10262) ) ;
NAND2   gate13135  (.A(WX3439), .B(II10261), .Z(II10263) ) ;
NAND2   gate13136  (.A(II10262), .B(II10263), .Z(II10260) ) ;
NAND2   gate13137  (.A(II10244), .B(II10260), .Z(II10268) ) ;
NAND2   gate13138  (.A(II10244), .B(II10268), .Z(II10269) ) ;
NAND2   gate13139  (.A(II10260), .B(II10268), .Z(II10270) ) ;
NAND2   gate13140  (.A(WX3587), .B(WX3249), .Z(II10277) ) ;
NAND2   gate13141  (.A(WX3587), .B(II10277), .Z(II10278) ) ;
NAND2   gate13142  (.A(WX3249), .B(II10277), .Z(II10279) ) ;
NAND2   gate13143  (.A(II10278), .B(II10279), .Z(II10276) ) ;
NAND2   gate13144  (.A(WX3313), .B(II10276), .Z(II10284) ) ;
NAND2   gate13145  (.A(WX3313), .B(II10284), .Z(II10285) ) ;
NAND2   gate13146  (.A(II10276), .B(II10284), .Z(II10286) ) ;
NAND2   gate13147  (.A(II10285), .B(II10286), .Z(II10275) ) ;
NAND2   gate13148  (.A(WX3377), .B(WX3441), .Z(II10292) ) ;
NAND2   gate13149  (.A(WX3377), .B(II10292), .Z(II10293) ) ;
NAND2   gate13150  (.A(WX3441), .B(II10292), .Z(II10294) ) ;
NAND2   gate13151  (.A(II10293), .B(II10294), .Z(II10291) ) ;
NAND2   gate13152  (.A(II10275), .B(II10291), .Z(II10299) ) ;
NAND2   gate13153  (.A(II10275), .B(II10299), .Z(II10300) ) ;
NAND2   gate13154  (.A(II10291), .B(II10299), .Z(II10301) ) ;
NAND2   gate13155  (.A(WX3587), .B(WX3251), .Z(II10308) ) ;
NAND2   gate13156  (.A(WX3587), .B(II10308), .Z(II10309) ) ;
NAND2   gate13157  (.A(WX3251), .B(II10308), .Z(II10310) ) ;
NAND2   gate13158  (.A(II10309), .B(II10310), .Z(II10307) ) ;
NAND2   gate13159  (.A(WX3315), .B(II10307), .Z(II10315) ) ;
NAND2   gate13160  (.A(WX3315), .B(II10315), .Z(II10316) ) ;
NAND2   gate13161  (.A(II10307), .B(II10315), .Z(II10317) ) ;
NAND2   gate13162  (.A(II10316), .B(II10317), .Z(II10306) ) ;
NAND2   gate13163  (.A(WX3379), .B(WX3443), .Z(II10323) ) ;
NAND2   gate13164  (.A(WX3379), .B(II10323), .Z(II10324) ) ;
NAND2   gate13165  (.A(WX3443), .B(II10323), .Z(II10325) ) ;
NAND2   gate13166  (.A(II10324), .B(II10325), .Z(II10322) ) ;
NAND2   gate13167  (.A(II10306), .B(II10322), .Z(II10330) ) ;
NAND2   gate13168  (.A(II10306), .B(II10330), .Z(II10331) ) ;
NAND2   gate13169  (.A(II10322), .B(II10330), .Z(II10332) ) ;
NAND2   gate13170  (.A(WX3587), .B(WX3253), .Z(II10339) ) ;
NAND2   gate13171  (.A(WX3587), .B(II10339), .Z(II10340) ) ;
NAND2   gate13172  (.A(WX3253), .B(II10339), .Z(II10341) ) ;
NAND2   gate13173  (.A(II10340), .B(II10341), .Z(II10338) ) ;
NAND2   gate13174  (.A(WX3317), .B(II10338), .Z(II10346) ) ;
NAND2   gate13175  (.A(WX3317), .B(II10346), .Z(II10347) ) ;
NAND2   gate13176  (.A(II10338), .B(II10346), .Z(II10348) ) ;
NAND2   gate13177  (.A(II10347), .B(II10348), .Z(II10337) ) ;
NAND2   gate13178  (.A(WX3381), .B(WX3445), .Z(II10354) ) ;
NAND2   gate13179  (.A(WX3381), .B(II10354), .Z(II10355) ) ;
NAND2   gate13180  (.A(WX3445), .B(II10354), .Z(II10356) ) ;
NAND2   gate13181  (.A(II10355), .B(II10356), .Z(II10353) ) ;
NAND2   gate13182  (.A(II10337), .B(II10353), .Z(II10361) ) ;
NAND2   gate13183  (.A(II10337), .B(II10361), .Z(II10362) ) ;
NAND2   gate13184  (.A(II10353), .B(II10361), .Z(II10363) ) ;
NAND2   gate13185  (.A(WX3587), .B(WX3255), .Z(II10370) ) ;
NAND2   gate13186  (.A(WX3587), .B(II10370), .Z(II10371) ) ;
NAND2   gate13187  (.A(WX3255), .B(II10370), .Z(II10372) ) ;
NAND2   gate13188  (.A(II10371), .B(II10372), .Z(II10369) ) ;
NAND2   gate13189  (.A(WX3319), .B(II10369), .Z(II10377) ) ;
NAND2   gate13190  (.A(WX3319), .B(II10377), .Z(II10378) ) ;
NAND2   gate13191  (.A(II10369), .B(II10377), .Z(II10379) ) ;
NAND2   gate13192  (.A(II10378), .B(II10379), .Z(II10368) ) ;
NAND2   gate13193  (.A(WX3383), .B(WX3447), .Z(II10385) ) ;
NAND2   gate13194  (.A(WX3383), .B(II10385), .Z(II10386) ) ;
NAND2   gate13195  (.A(WX3447), .B(II10385), .Z(II10387) ) ;
NAND2   gate13196  (.A(II10386), .B(II10387), .Z(II10384) ) ;
NAND2   gate13197  (.A(II10368), .B(II10384), .Z(II10392) ) ;
NAND2   gate13198  (.A(II10368), .B(II10392), .Z(II10393) ) ;
NAND2   gate13199  (.A(II10384), .B(II10392), .Z(II10394) ) ;
NAND2   gate13200  (.A(WX3587), .B(WX3257), .Z(II10401) ) ;
NAND2   gate13201  (.A(WX3587), .B(II10401), .Z(II10402) ) ;
NAND2   gate13202  (.A(WX3257), .B(II10401), .Z(II10403) ) ;
NAND2   gate13203  (.A(II10402), .B(II10403), .Z(II10400) ) ;
NAND2   gate13204  (.A(WX3321), .B(II10400), .Z(II10408) ) ;
NAND2   gate13205  (.A(WX3321), .B(II10408), .Z(II10409) ) ;
NAND2   gate13206  (.A(II10400), .B(II10408), .Z(II10410) ) ;
NAND2   gate13207  (.A(II10409), .B(II10410), .Z(II10399) ) ;
NAND2   gate13208  (.A(WX3385), .B(WX3449), .Z(II10416) ) ;
NAND2   gate13209  (.A(WX3385), .B(II10416), .Z(II10417) ) ;
NAND2   gate13210  (.A(WX3449), .B(II10416), .Z(II10418) ) ;
NAND2   gate13211  (.A(II10417), .B(II10418), .Z(II10415) ) ;
NAND2   gate13212  (.A(II10399), .B(II10415), .Z(II10423) ) ;
NAND2   gate13213  (.A(II10399), .B(II10423), .Z(II10424) ) ;
NAND2   gate13214  (.A(II10415), .B(II10423), .Z(II10425) ) ;
NAND2   gate13215  (.A(WX3587), .B(WX3259), .Z(II10432) ) ;
NAND2   gate13216  (.A(WX3587), .B(II10432), .Z(II10433) ) ;
NAND2   gate13217  (.A(WX3259), .B(II10432), .Z(II10434) ) ;
NAND2   gate13218  (.A(II10433), .B(II10434), .Z(II10431) ) ;
NAND2   gate13219  (.A(WX3323), .B(II10431), .Z(II10439) ) ;
NAND2   gate13220  (.A(WX3323), .B(II10439), .Z(II10440) ) ;
NAND2   gate13221  (.A(II10431), .B(II10439), .Z(II10441) ) ;
NAND2   gate13222  (.A(II10440), .B(II10441), .Z(II10430) ) ;
NAND2   gate13223  (.A(WX3387), .B(WX3451), .Z(II10447) ) ;
NAND2   gate13224  (.A(WX3387), .B(II10447), .Z(II10448) ) ;
NAND2   gate13225  (.A(WX3451), .B(II10447), .Z(II10449) ) ;
NAND2   gate13226  (.A(II10448), .B(II10449), .Z(II10446) ) ;
NAND2   gate13227  (.A(II10430), .B(II10446), .Z(II10454) ) ;
NAND2   gate13228  (.A(II10430), .B(II10454), .Z(II10455) ) ;
NAND2   gate13229  (.A(II10446), .B(II10454), .Z(II10456) ) ;
NAND2   gate13230  (.A(WX3587), .B(WX3261), .Z(II10463) ) ;
NAND2   gate13231  (.A(WX3587), .B(II10463), .Z(II10464) ) ;
NAND2   gate13232  (.A(WX3261), .B(II10463), .Z(II10465) ) ;
NAND2   gate13233  (.A(II10464), .B(II10465), .Z(II10462) ) ;
NAND2   gate13234  (.A(WX3325), .B(II10462), .Z(II10470) ) ;
NAND2   gate13235  (.A(WX3325), .B(II10470), .Z(II10471) ) ;
NAND2   gate13236  (.A(II10462), .B(II10470), .Z(II10472) ) ;
NAND2   gate13237  (.A(II10471), .B(II10472), .Z(II10461) ) ;
NAND2   gate13238  (.A(WX3389), .B(WX3453), .Z(II10478) ) ;
NAND2   gate13239  (.A(WX3389), .B(II10478), .Z(II10479) ) ;
NAND2   gate13240  (.A(WX3453), .B(II10478), .Z(II10480) ) ;
NAND2   gate13241  (.A(II10479), .B(II10480), .Z(II10477) ) ;
NAND2   gate13242  (.A(II10461), .B(II10477), .Z(II10485) ) ;
NAND2   gate13243  (.A(II10461), .B(II10485), .Z(II10486) ) ;
NAND2   gate13244  (.A(II10477), .B(II10485), .Z(II10487) ) ;
NAND2   gate13245  (.A(WX3588), .B(WX3263), .Z(II10494) ) ;
NAND2   gate13246  (.A(WX3588), .B(II10494), .Z(II10495) ) ;
NAND2   gate13247  (.A(WX3263), .B(II10494), .Z(II10496) ) ;
NAND2   gate13248  (.A(II10495), .B(II10496), .Z(II10493) ) ;
NAND2   gate13249  (.A(WX3327), .B(II10493), .Z(II10501) ) ;
NAND2   gate13250  (.A(WX3327), .B(II10501), .Z(II10502) ) ;
NAND2   gate13251  (.A(II10493), .B(II10501), .Z(II10503) ) ;
NAND2   gate13252  (.A(II10502), .B(II10503), .Z(II10492) ) ;
NAND2   gate13253  (.A(WX3391), .B(WX3455), .Z(II10509) ) ;
NAND2   gate13254  (.A(WX3391), .B(II10509), .Z(II10510) ) ;
NAND2   gate13255  (.A(WX3455), .B(II10509), .Z(II10511) ) ;
NAND2   gate13256  (.A(II10510), .B(II10511), .Z(II10508) ) ;
NAND2   gate13257  (.A(II10492), .B(II10508), .Z(II10516) ) ;
NAND2   gate13258  (.A(II10492), .B(II10516), .Z(II10517) ) ;
NAND2   gate13259  (.A(II10508), .B(II10516), .Z(II10518) ) ;
NAND2   gate13260  (.A(WX3588), .B(WX3265), .Z(II10525) ) ;
NAND2   gate13261  (.A(WX3588), .B(II10525), .Z(II10526) ) ;
NAND2   gate13262  (.A(WX3265), .B(II10525), .Z(II10527) ) ;
NAND2   gate13263  (.A(II10526), .B(II10527), .Z(II10524) ) ;
NAND2   gate13264  (.A(WX3329), .B(II10524), .Z(II10532) ) ;
NAND2   gate13265  (.A(WX3329), .B(II10532), .Z(II10533) ) ;
NAND2   gate13266  (.A(II10524), .B(II10532), .Z(II10534) ) ;
NAND2   gate13267  (.A(II10533), .B(II10534), .Z(II10523) ) ;
NAND2   gate13268  (.A(WX3393), .B(WX3457), .Z(II10540) ) ;
NAND2   gate13269  (.A(WX3393), .B(II10540), .Z(II10541) ) ;
NAND2   gate13270  (.A(WX3457), .B(II10540), .Z(II10542) ) ;
NAND2   gate13271  (.A(II10541), .B(II10542), .Z(II10539) ) ;
NAND2   gate13272  (.A(II10523), .B(II10539), .Z(II10547) ) ;
NAND2   gate13273  (.A(II10523), .B(II10547), .Z(II10548) ) ;
NAND2   gate13274  (.A(II10539), .B(II10547), .Z(II10549) ) ;
NAND2   gate13275  (.A(WX3588), .B(WX3267), .Z(II10556) ) ;
NAND2   gate13276  (.A(WX3588), .B(II10556), .Z(II10557) ) ;
NAND2   gate13277  (.A(WX3267), .B(II10556), .Z(II10558) ) ;
NAND2   gate13278  (.A(II10557), .B(II10558), .Z(II10555) ) ;
NAND2   gate13279  (.A(WX3331), .B(II10555), .Z(II10563) ) ;
NAND2   gate13280  (.A(WX3331), .B(II10563), .Z(II10564) ) ;
NAND2   gate13281  (.A(II10555), .B(II10563), .Z(II10565) ) ;
NAND2   gate13282  (.A(II10564), .B(II10565), .Z(II10554) ) ;
NAND2   gate13283  (.A(WX3395), .B(WX3459), .Z(II10571) ) ;
NAND2   gate13284  (.A(WX3395), .B(II10571), .Z(II10572) ) ;
NAND2   gate13285  (.A(WX3459), .B(II10571), .Z(II10573) ) ;
NAND2   gate13286  (.A(II10572), .B(II10573), .Z(II10570) ) ;
NAND2   gate13287  (.A(II10554), .B(II10570), .Z(II10578) ) ;
NAND2   gate13288  (.A(II10554), .B(II10578), .Z(II10579) ) ;
NAND2   gate13289  (.A(II10570), .B(II10578), .Z(II10580) ) ;
NAND2   gate13290  (.A(WX3588), .B(WX3269), .Z(II10587) ) ;
NAND2   gate13291  (.A(WX3588), .B(II10587), .Z(II10588) ) ;
NAND2   gate13292  (.A(WX3269), .B(II10587), .Z(II10589) ) ;
NAND2   gate13293  (.A(II10588), .B(II10589), .Z(II10586) ) ;
NAND2   gate13294  (.A(WX3333), .B(II10586), .Z(II10594) ) ;
NAND2   gate13295  (.A(WX3333), .B(II10594), .Z(II10595) ) ;
NAND2   gate13296  (.A(II10586), .B(II10594), .Z(II10596) ) ;
NAND2   gate13297  (.A(II10595), .B(II10596), .Z(II10585) ) ;
NAND2   gate13298  (.A(WX3397), .B(WX3461), .Z(II10602) ) ;
NAND2   gate13299  (.A(WX3397), .B(II10602), .Z(II10603) ) ;
NAND2   gate13300  (.A(WX3461), .B(II10602), .Z(II10604) ) ;
NAND2   gate13301  (.A(II10603), .B(II10604), .Z(II10601) ) ;
NAND2   gate13302  (.A(II10585), .B(II10601), .Z(II10609) ) ;
NAND2   gate13303  (.A(II10585), .B(II10609), .Z(II10610) ) ;
NAND2   gate13304  (.A(II10601), .B(II10609), .Z(II10611) ) ;
NAND2   gate13305  (.A(WX3588), .B(WX3271), .Z(II10618) ) ;
NAND2   gate13306  (.A(WX3588), .B(II10618), .Z(II10619) ) ;
NAND2   gate13307  (.A(WX3271), .B(II10618), .Z(II10620) ) ;
NAND2   gate13308  (.A(II10619), .B(II10620), .Z(II10617) ) ;
NAND2   gate13309  (.A(WX3335), .B(II10617), .Z(II10625) ) ;
NAND2   gate13310  (.A(WX3335), .B(II10625), .Z(II10626) ) ;
NAND2   gate13311  (.A(II10617), .B(II10625), .Z(II10627) ) ;
NAND2   gate13312  (.A(II10626), .B(II10627), .Z(II10616) ) ;
NAND2   gate13313  (.A(WX3399), .B(WX3463), .Z(II10633) ) ;
NAND2   gate13314  (.A(WX3399), .B(II10633), .Z(II10634) ) ;
NAND2   gate13315  (.A(WX3463), .B(II10633), .Z(II10635) ) ;
NAND2   gate13316  (.A(II10634), .B(II10635), .Z(II10632) ) ;
NAND2   gate13317  (.A(II10616), .B(II10632), .Z(II10640) ) ;
NAND2   gate13318  (.A(II10616), .B(II10640), .Z(II10641) ) ;
NAND2   gate13319  (.A(II10632), .B(II10640), .Z(II10642) ) ;
NAND2   gate13320  (.A(WX3588), .B(WX3273), .Z(II10649) ) ;
NAND2   gate13321  (.A(WX3588), .B(II10649), .Z(II10650) ) ;
NAND2   gate13322  (.A(WX3273), .B(II10649), .Z(II10651) ) ;
NAND2   gate13323  (.A(II10650), .B(II10651), .Z(II10648) ) ;
NAND2   gate13324  (.A(WX3337), .B(II10648), .Z(II10656) ) ;
NAND2   gate13325  (.A(WX3337), .B(II10656), .Z(II10657) ) ;
NAND2   gate13326  (.A(II10648), .B(II10656), .Z(II10658) ) ;
NAND2   gate13327  (.A(II10657), .B(II10658), .Z(II10647) ) ;
NAND2   gate13328  (.A(WX3401), .B(WX3465), .Z(II10664) ) ;
NAND2   gate13329  (.A(WX3401), .B(II10664), .Z(II10665) ) ;
NAND2   gate13330  (.A(WX3465), .B(II10664), .Z(II10666) ) ;
NAND2   gate13331  (.A(II10665), .B(II10666), .Z(II10663) ) ;
NAND2   gate13332  (.A(II10647), .B(II10663), .Z(II10671) ) ;
NAND2   gate13333  (.A(II10647), .B(II10671), .Z(II10672) ) ;
NAND2   gate13334  (.A(II10663), .B(II10671), .Z(II10673) ) ;
NAND2   gate13335  (.A(WX3588), .B(WX3275), .Z(II10680) ) ;
NAND2   gate13336  (.A(WX3588), .B(II10680), .Z(II10681) ) ;
NAND2   gate13337  (.A(WX3275), .B(II10680), .Z(II10682) ) ;
NAND2   gate13338  (.A(II10681), .B(II10682), .Z(II10679) ) ;
NAND2   gate13339  (.A(WX3339), .B(II10679), .Z(II10687) ) ;
NAND2   gate13340  (.A(WX3339), .B(II10687), .Z(II10688) ) ;
NAND2   gate13341  (.A(II10679), .B(II10687), .Z(II10689) ) ;
NAND2   gate13342  (.A(II10688), .B(II10689), .Z(II10678) ) ;
NAND2   gate13343  (.A(WX3403), .B(WX3467), .Z(II10695) ) ;
NAND2   gate13344  (.A(WX3403), .B(II10695), .Z(II10696) ) ;
NAND2   gate13345  (.A(WX3467), .B(II10695), .Z(II10697) ) ;
NAND2   gate13346  (.A(II10696), .B(II10697), .Z(II10694) ) ;
NAND2   gate13347  (.A(II10678), .B(II10694), .Z(II10702) ) ;
NAND2   gate13348  (.A(II10678), .B(II10702), .Z(II10703) ) ;
NAND2   gate13349  (.A(II10694), .B(II10702), .Z(II10704) ) ;
NAND2   gate13350  (.A(WX3588), .B(WX3277), .Z(II10711) ) ;
NAND2   gate13351  (.A(WX3588), .B(II10711), .Z(II10712) ) ;
NAND2   gate13352  (.A(WX3277), .B(II10711), .Z(II10713) ) ;
NAND2   gate13353  (.A(II10712), .B(II10713), .Z(II10710) ) ;
NAND2   gate13354  (.A(WX3341), .B(II10710), .Z(II10718) ) ;
NAND2   gate13355  (.A(WX3341), .B(II10718), .Z(II10719) ) ;
NAND2   gate13356  (.A(II10710), .B(II10718), .Z(II10720) ) ;
NAND2   gate13357  (.A(II10719), .B(II10720), .Z(II10709) ) ;
NAND2   gate13358  (.A(WX3405), .B(WX3469), .Z(II10726) ) ;
NAND2   gate13359  (.A(WX3405), .B(II10726), .Z(II10727) ) ;
NAND2   gate13360  (.A(WX3469), .B(II10726), .Z(II10728) ) ;
NAND2   gate13361  (.A(II10727), .B(II10728), .Z(II10725) ) ;
NAND2   gate13362  (.A(II10709), .B(II10725), .Z(II10733) ) ;
NAND2   gate13363  (.A(II10709), .B(II10733), .Z(II10734) ) ;
NAND2   gate13364  (.A(II10725), .B(II10733), .Z(II10735) ) ;
NAND2   gate13365  (.A(WX3588), .B(WX3279), .Z(II10742) ) ;
NAND2   gate13366  (.A(WX3588), .B(II10742), .Z(II10743) ) ;
NAND2   gate13367  (.A(WX3279), .B(II10742), .Z(II10744) ) ;
NAND2   gate13368  (.A(II10743), .B(II10744), .Z(II10741) ) ;
NAND2   gate13369  (.A(WX3343), .B(II10741), .Z(II10749) ) ;
NAND2   gate13370  (.A(WX3343), .B(II10749), .Z(II10750) ) ;
NAND2   gate13371  (.A(II10741), .B(II10749), .Z(II10751) ) ;
NAND2   gate13372  (.A(II10750), .B(II10751), .Z(II10740) ) ;
NAND2   gate13373  (.A(WX3407), .B(WX3471), .Z(II10757) ) ;
NAND2   gate13374  (.A(WX3407), .B(II10757), .Z(II10758) ) ;
NAND2   gate13375  (.A(WX3471), .B(II10757), .Z(II10759) ) ;
NAND2   gate13376  (.A(II10758), .B(II10759), .Z(II10756) ) ;
NAND2   gate13377  (.A(II10740), .B(II10756), .Z(II10764) ) ;
NAND2   gate13378  (.A(II10740), .B(II10764), .Z(II10765) ) ;
NAND2   gate13379  (.A(II10756), .B(II10764), .Z(II10766) ) ;
NAND2   gate13380  (.A(WX3588), .B(WX3281), .Z(II10773) ) ;
NAND2   gate13381  (.A(WX3588), .B(II10773), .Z(II10774) ) ;
NAND2   gate13382  (.A(WX3281), .B(II10773), .Z(II10775) ) ;
NAND2   gate13383  (.A(II10774), .B(II10775), .Z(II10772) ) ;
NAND2   gate13384  (.A(WX3345), .B(II10772), .Z(II10780) ) ;
NAND2   gate13385  (.A(WX3345), .B(II10780), .Z(II10781) ) ;
NAND2   gate13386  (.A(II10772), .B(II10780), .Z(II10782) ) ;
NAND2   gate13387  (.A(II10781), .B(II10782), .Z(II10771) ) ;
NAND2   gate13388  (.A(WX3409), .B(WX3473), .Z(II10788) ) ;
NAND2   gate13389  (.A(WX3409), .B(II10788), .Z(II10789) ) ;
NAND2   gate13390  (.A(WX3473), .B(II10788), .Z(II10790) ) ;
NAND2   gate13391  (.A(II10789), .B(II10790), .Z(II10787) ) ;
NAND2   gate13392  (.A(II10771), .B(II10787), .Z(II10795) ) ;
NAND2   gate13393  (.A(II10771), .B(II10795), .Z(II10796) ) ;
NAND2   gate13394  (.A(II10787), .B(II10795), .Z(II10797) ) ;
NAND2   gate13395  (.A(WX3588), .B(WX3283), .Z(II10804) ) ;
NAND2   gate13396  (.A(WX3588), .B(II10804), .Z(II10805) ) ;
NAND2   gate13397  (.A(WX3283), .B(II10804), .Z(II10806) ) ;
NAND2   gate13398  (.A(II10805), .B(II10806), .Z(II10803) ) ;
NAND2   gate13399  (.A(WX3347), .B(II10803), .Z(II10811) ) ;
NAND2   gate13400  (.A(WX3347), .B(II10811), .Z(II10812) ) ;
NAND2   gate13401  (.A(II10803), .B(II10811), .Z(II10813) ) ;
NAND2   gate13402  (.A(II10812), .B(II10813), .Z(II10802) ) ;
NAND2   gate13403  (.A(WX3411), .B(WX3475), .Z(II10819) ) ;
NAND2   gate13404  (.A(WX3411), .B(II10819), .Z(II10820) ) ;
NAND2   gate13405  (.A(WX3475), .B(II10819), .Z(II10821) ) ;
NAND2   gate13406  (.A(II10820), .B(II10821), .Z(II10818) ) ;
NAND2   gate13407  (.A(II10802), .B(II10818), .Z(II10826) ) ;
NAND2   gate13408  (.A(II10802), .B(II10826), .Z(II10827) ) ;
NAND2   gate13409  (.A(II10818), .B(II10826), .Z(II10828) ) ;
NAND2   gate13410  (.A(WX3588), .B(WX3285), .Z(II10835) ) ;
NAND2   gate13411  (.A(WX3588), .B(II10835), .Z(II10836) ) ;
NAND2   gate13412  (.A(WX3285), .B(II10835), .Z(II10837) ) ;
NAND2   gate13413  (.A(II10836), .B(II10837), .Z(II10834) ) ;
NAND2   gate13414  (.A(WX3349), .B(II10834), .Z(II10842) ) ;
NAND2   gate13415  (.A(WX3349), .B(II10842), .Z(II10843) ) ;
NAND2   gate13416  (.A(II10834), .B(II10842), .Z(II10844) ) ;
NAND2   gate13417  (.A(II10843), .B(II10844), .Z(II10833) ) ;
NAND2   gate13418  (.A(WX3413), .B(WX3477), .Z(II10850) ) ;
NAND2   gate13419  (.A(WX3413), .B(II10850), .Z(II10851) ) ;
NAND2   gate13420  (.A(WX3477), .B(II10850), .Z(II10852) ) ;
NAND2   gate13421  (.A(II10851), .B(II10852), .Z(II10849) ) ;
NAND2   gate13422  (.A(II10833), .B(II10849), .Z(II10857) ) ;
NAND2   gate13423  (.A(II10833), .B(II10857), .Z(II10858) ) ;
NAND2   gate13424  (.A(II10849), .B(II10857), .Z(II10859) ) ;
NAND2   gate13425  (.A(WX3588), .B(WX3287), .Z(II10866) ) ;
NAND2   gate13426  (.A(WX3588), .B(II10866), .Z(II10867) ) ;
NAND2   gate13427  (.A(WX3287), .B(II10866), .Z(II10868) ) ;
NAND2   gate13428  (.A(II10867), .B(II10868), .Z(II10865) ) ;
NAND2   gate13429  (.A(WX3351), .B(II10865), .Z(II10873) ) ;
NAND2   gate13430  (.A(WX3351), .B(II10873), .Z(II10874) ) ;
NAND2   gate13431  (.A(II10865), .B(II10873), .Z(II10875) ) ;
NAND2   gate13432  (.A(II10874), .B(II10875), .Z(II10864) ) ;
NAND2   gate13433  (.A(WX3415), .B(WX3479), .Z(II10881) ) ;
NAND2   gate13434  (.A(WX3415), .B(II10881), .Z(II10882) ) ;
NAND2   gate13435  (.A(WX3479), .B(II10881), .Z(II10883) ) ;
NAND2   gate13436  (.A(II10882), .B(II10883), .Z(II10880) ) ;
NAND2   gate13437  (.A(II10864), .B(II10880), .Z(II10888) ) ;
NAND2   gate13438  (.A(II10864), .B(II10888), .Z(II10889) ) ;
NAND2   gate13439  (.A(II10880), .B(II10888), .Z(II10890) ) ;
NAND2   gate13440  (.A(WX3588), .B(WX3289), .Z(II10897) ) ;
NAND2   gate13441  (.A(WX3588), .B(II10897), .Z(II10898) ) ;
NAND2   gate13442  (.A(WX3289), .B(II10897), .Z(II10899) ) ;
NAND2   gate13443  (.A(II10898), .B(II10899), .Z(II10896) ) ;
NAND2   gate13444  (.A(WX3353), .B(II10896), .Z(II10904) ) ;
NAND2   gate13445  (.A(WX3353), .B(II10904), .Z(II10905) ) ;
NAND2   gate13446  (.A(II10896), .B(II10904), .Z(II10906) ) ;
NAND2   gate13447  (.A(II10905), .B(II10906), .Z(II10895) ) ;
NAND2   gate13448  (.A(WX3417), .B(WX3481), .Z(II10912) ) ;
NAND2   gate13449  (.A(WX3417), .B(II10912), .Z(II10913) ) ;
NAND2   gate13450  (.A(WX3481), .B(II10912), .Z(II10914) ) ;
NAND2   gate13451  (.A(II10913), .B(II10914), .Z(II10911) ) ;
NAND2   gate13452  (.A(II10895), .B(II10911), .Z(II10919) ) ;
NAND2   gate13453  (.A(II10895), .B(II10919), .Z(II10920) ) ;
NAND2   gate13454  (.A(II10911), .B(II10919), .Z(II10921) ) ;
NAND2   gate13455  (.A(WX3588), .B(WX3291), .Z(II10928) ) ;
NAND2   gate13456  (.A(WX3588), .B(II10928), .Z(II10929) ) ;
NAND2   gate13457  (.A(WX3291), .B(II10928), .Z(II10930) ) ;
NAND2   gate13458  (.A(II10929), .B(II10930), .Z(II10927) ) ;
NAND2   gate13459  (.A(WX3355), .B(II10927), .Z(II10935) ) ;
NAND2   gate13460  (.A(WX3355), .B(II10935), .Z(II10936) ) ;
NAND2   gate13461  (.A(II10927), .B(II10935), .Z(II10937) ) ;
NAND2   gate13462  (.A(II10936), .B(II10937), .Z(II10926) ) ;
NAND2   gate13463  (.A(WX3419), .B(WX3483), .Z(II10943) ) ;
NAND2   gate13464  (.A(WX3419), .B(II10943), .Z(II10944) ) ;
NAND2   gate13465  (.A(WX3483), .B(II10943), .Z(II10945) ) ;
NAND2   gate13466  (.A(II10944), .B(II10945), .Z(II10942) ) ;
NAND2   gate13467  (.A(II10926), .B(II10942), .Z(II10950) ) ;
NAND2   gate13468  (.A(II10926), .B(II10950), .Z(II10951) ) ;
NAND2   gate13469  (.A(II10942), .B(II10950), .Z(II10952) ) ;
NAND2   gate13470  (.A(WX3588), .B(WX3293), .Z(II10959) ) ;
NAND2   gate13471  (.A(WX3588), .B(II10959), .Z(II10960) ) ;
NAND2   gate13472  (.A(WX3293), .B(II10959), .Z(II10961) ) ;
NAND2   gate13473  (.A(II10960), .B(II10961), .Z(II10958) ) ;
NAND2   gate13474  (.A(WX3357), .B(II10958), .Z(II10966) ) ;
NAND2   gate13475  (.A(WX3357), .B(II10966), .Z(II10967) ) ;
NAND2   gate13476  (.A(II10958), .B(II10966), .Z(II10968) ) ;
NAND2   gate13477  (.A(II10967), .B(II10968), .Z(II10957) ) ;
NAND2   gate13478  (.A(WX3421), .B(WX3485), .Z(II10974) ) ;
NAND2   gate13479  (.A(WX3421), .B(II10974), .Z(II10975) ) ;
NAND2   gate13480  (.A(WX3485), .B(II10974), .Z(II10976) ) ;
NAND2   gate13481  (.A(II10975), .B(II10976), .Z(II10973) ) ;
NAND2   gate13482  (.A(II10957), .B(II10973), .Z(II10981) ) ;
NAND2   gate13483  (.A(II10957), .B(II10981), .Z(II10982) ) ;
NAND2   gate13484  (.A(II10973), .B(II10981), .Z(II10983) ) ;
NAND2   gate13485  (.A(WX3166), .B(WX3071), .Z(II11062) ) ;
NAND2   gate13486  (.A(WX3166), .B(II11062), .Z(II11063) ) ;
NAND2   gate13487  (.A(WX3071), .B(II11062), .Z(II11064) ) ;
NAND2   gate13488  (.A(WX3167), .B(WX3073), .Z(II11075) ) ;
NAND2   gate13489  (.A(WX3167), .B(II11075), .Z(II11076) ) ;
NAND2   gate13490  (.A(WX3073), .B(II11075), .Z(II11077) ) ;
NAND2   gate13491  (.A(WX3168), .B(WX3075), .Z(II11088) ) ;
NAND2   gate13492  (.A(WX3168), .B(II11088), .Z(II11089) ) ;
NAND2   gate13493  (.A(WX3075), .B(II11088), .Z(II11090) ) ;
NAND2   gate13494  (.A(WX3169), .B(WX3077), .Z(II11101) ) ;
NAND2   gate13495  (.A(WX3169), .B(II11101), .Z(II11102) ) ;
NAND2   gate13496  (.A(WX3077), .B(II11101), .Z(II11103) ) ;
NAND2   gate13497  (.A(WX3170), .B(WX3079), .Z(II11114) ) ;
NAND2   gate13498  (.A(WX3170), .B(II11114), .Z(II11115) ) ;
NAND2   gate13499  (.A(WX3079), .B(II11114), .Z(II11116) ) ;
NAND2   gate13500  (.A(WX3171), .B(WX3081), .Z(II11127) ) ;
NAND2   gate13501  (.A(WX3171), .B(II11127), .Z(II11128) ) ;
NAND2   gate13502  (.A(WX3081), .B(II11127), .Z(II11129) ) ;
NAND2   gate13503  (.A(WX3172), .B(WX3083), .Z(II11140) ) ;
NAND2   gate13504  (.A(WX3172), .B(II11140), .Z(II11141) ) ;
NAND2   gate13505  (.A(WX3083), .B(II11140), .Z(II11142) ) ;
NAND2   gate13506  (.A(WX3173), .B(WX3085), .Z(II11153) ) ;
NAND2   gate13507  (.A(WX3173), .B(II11153), .Z(II11154) ) ;
NAND2   gate13508  (.A(WX3085), .B(II11153), .Z(II11155) ) ;
NAND2   gate13509  (.A(WX3174), .B(WX3087), .Z(II11166) ) ;
NAND2   gate13510  (.A(WX3174), .B(II11166), .Z(II11167) ) ;
NAND2   gate13511  (.A(WX3087), .B(II11166), .Z(II11168) ) ;
NAND2   gate13512  (.A(WX3175), .B(WX3089), .Z(II11179) ) ;
NAND2   gate13513  (.A(WX3175), .B(II11179), .Z(II11180) ) ;
NAND2   gate13514  (.A(WX3089), .B(II11179), .Z(II11181) ) ;
NAND2   gate13515  (.A(WX3176), .B(WX3091), .Z(II11192) ) ;
NAND2   gate13516  (.A(WX3176), .B(II11192), .Z(II11193) ) ;
NAND2   gate13517  (.A(WX3091), .B(II11192), .Z(II11194) ) ;
NAND2   gate13518  (.A(WX3177), .B(WX3093), .Z(II11205) ) ;
NAND2   gate13519  (.A(WX3177), .B(II11205), .Z(II11206) ) ;
NAND2   gate13520  (.A(WX3093), .B(II11205), .Z(II11207) ) ;
NAND2   gate13521  (.A(WX3178), .B(WX3095), .Z(II11218) ) ;
NAND2   gate13522  (.A(WX3178), .B(II11218), .Z(II11219) ) ;
NAND2   gate13523  (.A(WX3095), .B(II11218), .Z(II11220) ) ;
NAND2   gate13524  (.A(WX3179), .B(WX3097), .Z(II11231) ) ;
NAND2   gate13525  (.A(WX3179), .B(II11231), .Z(II11232) ) ;
NAND2   gate13526  (.A(WX3097), .B(II11231), .Z(II11233) ) ;
NAND2   gate13527  (.A(WX3180), .B(WX3099), .Z(II11244) ) ;
NAND2   gate13528  (.A(WX3180), .B(II11244), .Z(II11245) ) ;
NAND2   gate13529  (.A(WX3099), .B(II11244), .Z(II11246) ) ;
NAND2   gate13530  (.A(WX3181), .B(WX3101), .Z(II11257) ) ;
NAND2   gate13531  (.A(WX3181), .B(II11257), .Z(II11258) ) ;
NAND2   gate13532  (.A(WX3101), .B(II11257), .Z(II11259) ) ;
NAND2   gate13533  (.A(WX3182), .B(WX3103), .Z(II11270) ) ;
NAND2   gate13534  (.A(WX3182), .B(II11270), .Z(II11271) ) ;
NAND2   gate13535  (.A(WX3103), .B(II11270), .Z(II11272) ) ;
NAND2   gate13536  (.A(WX3183), .B(WX3105), .Z(II11283) ) ;
NAND2   gate13537  (.A(WX3183), .B(II11283), .Z(II11284) ) ;
NAND2   gate13538  (.A(WX3105), .B(II11283), .Z(II11285) ) ;
NAND2   gate13539  (.A(WX3184), .B(WX3107), .Z(II11296) ) ;
NAND2   gate13540  (.A(WX3184), .B(II11296), .Z(II11297) ) ;
NAND2   gate13541  (.A(WX3107), .B(II11296), .Z(II11298) ) ;
NAND2   gate13542  (.A(WX3185), .B(WX3109), .Z(II11309) ) ;
NAND2   gate13543  (.A(WX3185), .B(II11309), .Z(II11310) ) ;
NAND2   gate13544  (.A(WX3109), .B(II11309), .Z(II11311) ) ;
NAND2   gate13545  (.A(WX3186), .B(WX3111), .Z(II11322) ) ;
NAND2   gate13546  (.A(WX3186), .B(II11322), .Z(II11323) ) ;
NAND2   gate13547  (.A(WX3111), .B(II11322), .Z(II11324) ) ;
NAND2   gate13548  (.A(WX3187), .B(WX3113), .Z(II11335) ) ;
NAND2   gate13549  (.A(WX3187), .B(II11335), .Z(II11336) ) ;
NAND2   gate13550  (.A(WX3113), .B(II11335), .Z(II11337) ) ;
NAND2   gate13551  (.A(WX3188), .B(WX3115), .Z(II11348) ) ;
NAND2   gate13552  (.A(WX3188), .B(II11348), .Z(II11349) ) ;
NAND2   gate13553  (.A(WX3115), .B(II11348), .Z(II11350) ) ;
NAND2   gate13554  (.A(WX3189), .B(WX3117), .Z(II11361) ) ;
NAND2   gate13555  (.A(WX3189), .B(II11361), .Z(II11362) ) ;
NAND2   gate13556  (.A(WX3117), .B(II11361), .Z(II11363) ) ;
NAND2   gate13557  (.A(WX3190), .B(WX3119), .Z(II11374) ) ;
NAND2   gate13558  (.A(WX3190), .B(II11374), .Z(II11375) ) ;
NAND2   gate13559  (.A(WX3119), .B(II11374), .Z(II11376) ) ;
NAND2   gate13560  (.A(WX3191), .B(WX3121), .Z(II11387) ) ;
NAND2   gate13561  (.A(WX3191), .B(II11387), .Z(II11388) ) ;
NAND2   gate13562  (.A(WX3121), .B(II11387), .Z(II11389) ) ;
NAND2   gate13563  (.A(WX3192), .B(WX3123), .Z(II11400) ) ;
NAND2   gate13564  (.A(WX3192), .B(II11400), .Z(II11401) ) ;
NAND2   gate13565  (.A(WX3123), .B(II11400), .Z(II11402) ) ;
NAND2   gate13566  (.A(WX3193), .B(WX3125), .Z(II11413) ) ;
NAND2   gate13567  (.A(WX3193), .B(II11413), .Z(II11414) ) ;
NAND2   gate13568  (.A(WX3125), .B(II11413), .Z(II11415) ) ;
NAND2   gate13569  (.A(WX3194), .B(WX3127), .Z(II11426) ) ;
NAND2   gate13570  (.A(WX3194), .B(II11426), .Z(II11427) ) ;
NAND2   gate13571  (.A(WX3127), .B(II11426), .Z(II11428) ) ;
NAND2   gate13572  (.A(WX3195), .B(WX3129), .Z(II11439) ) ;
NAND2   gate13573  (.A(WX3195), .B(II11439), .Z(II11440) ) ;
NAND2   gate13574  (.A(WX3129), .B(II11439), .Z(II11441) ) ;
NAND2   gate13575  (.A(WX3196), .B(WX3131), .Z(II11452) ) ;
NAND2   gate13576  (.A(WX3196), .B(II11452), .Z(II11453) ) ;
NAND2   gate13577  (.A(WX3131), .B(II11452), .Z(II11454) ) ;
NAND2   gate13578  (.A(WX3197), .B(WX3133), .Z(II11465) ) ;
NAND2   gate13579  (.A(WX3197), .B(II11465), .Z(II11466) ) ;
NAND2   gate13580  (.A(WX3133), .B(II11465), .Z(II11467) ) ;
NAND2   gate13581  (.A(WX3213), .B(CRC_OUT_7_31), .Z(II11480) ) ;
NAND2   gate13582  (.A(WX3213), .B(II11480), .Z(II11481) ) ;
NAND2   gate13583  (.A(CRC_OUT_7_31), .B(II11480), .Z(II11482) ) ;
NAND2   gate13584  (.A(II11481), .B(II11482), .Z(II11479) ) ;
NAND2   gate13585  (.A(CRC_OUT_7_15), .B(II11479), .Z(II11487) ) ;
NAND2   gate13586  (.A(CRC_OUT_7_15), .B(II11487), .Z(II11488) ) ;
NAND2   gate13587  (.A(II11479), .B(II11487), .Z(II11489) ) ;
NAND2   gate13588  (.A(WX3218), .B(CRC_OUT_7_31), .Z(II11495) ) ;
NAND2   gate13589  (.A(WX3218), .B(II11495), .Z(II11496) ) ;
NAND2   gate13590  (.A(CRC_OUT_7_31), .B(II11495), .Z(II11497) ) ;
NAND2   gate13591  (.A(II11496), .B(II11497), .Z(II11494) ) ;
NAND2   gate13592  (.A(CRC_OUT_7_10), .B(II11494), .Z(II11502) ) ;
NAND2   gate13593  (.A(CRC_OUT_7_10), .B(II11502), .Z(II11503) ) ;
NAND2   gate13594  (.A(II11494), .B(II11502), .Z(II11504) ) ;
NAND2   gate13595  (.A(WX3225), .B(CRC_OUT_7_31), .Z(II11510) ) ;
NAND2   gate13596  (.A(WX3225), .B(II11510), .Z(II11511) ) ;
NAND2   gate13597  (.A(CRC_OUT_7_31), .B(II11510), .Z(II11512) ) ;
NAND2   gate13598  (.A(II11511), .B(II11512), .Z(II11509) ) ;
NAND2   gate13599  (.A(CRC_OUT_7_3), .B(II11509), .Z(II11517) ) ;
NAND2   gate13600  (.A(CRC_OUT_7_3), .B(II11517), .Z(II11518) ) ;
NAND2   gate13601  (.A(II11509), .B(II11517), .Z(II11519) ) ;
NAND2   gate13602  (.A(WX3229), .B(CRC_OUT_7_31), .Z(II11524) ) ;
NAND2   gate13603  (.A(WX3229), .B(II11524), .Z(II11525) ) ;
NAND2   gate13604  (.A(CRC_OUT_7_31), .B(II11524), .Z(II11526) ) ;
NAND2   gate13605  (.A(WX3198), .B(CRC_OUT_7_30), .Z(II11531) ) ;
NAND2   gate13606  (.A(WX3198), .B(II11531), .Z(II11532) ) ;
NAND2   gate13607  (.A(CRC_OUT_7_30), .B(II11531), .Z(II11533) ) ;
NAND2   gate13608  (.A(WX3199), .B(CRC_OUT_7_29), .Z(II11538) ) ;
NAND2   gate13609  (.A(WX3199), .B(II11538), .Z(II11539) ) ;
NAND2   gate13610  (.A(CRC_OUT_7_29), .B(II11538), .Z(II11540) ) ;
NAND2   gate13611  (.A(WX3200), .B(CRC_OUT_7_28), .Z(II11545) ) ;
NAND2   gate13612  (.A(WX3200), .B(II11545), .Z(II11546) ) ;
NAND2   gate13613  (.A(CRC_OUT_7_28), .B(II11545), .Z(II11547) ) ;
NAND2   gate13614  (.A(WX3201), .B(CRC_OUT_7_27), .Z(II11552) ) ;
NAND2   gate13615  (.A(WX3201), .B(II11552), .Z(II11553) ) ;
NAND2   gate13616  (.A(CRC_OUT_7_27), .B(II11552), .Z(II11554) ) ;
NAND2   gate13617  (.A(WX3202), .B(CRC_OUT_7_26), .Z(II11559) ) ;
NAND2   gate13618  (.A(WX3202), .B(II11559), .Z(II11560) ) ;
NAND2   gate13619  (.A(CRC_OUT_7_26), .B(II11559), .Z(II11561) ) ;
NAND2   gate13620  (.A(WX3203), .B(CRC_OUT_7_25), .Z(II11566) ) ;
NAND2   gate13621  (.A(WX3203), .B(II11566), .Z(II11567) ) ;
NAND2   gate13622  (.A(CRC_OUT_7_25), .B(II11566), .Z(II11568) ) ;
NAND2   gate13623  (.A(WX3204), .B(CRC_OUT_7_24), .Z(II11573) ) ;
NAND2   gate13624  (.A(WX3204), .B(II11573), .Z(II11574) ) ;
NAND2   gate13625  (.A(CRC_OUT_7_24), .B(II11573), .Z(II11575) ) ;
NAND2   gate13626  (.A(WX3205), .B(CRC_OUT_7_23), .Z(II11580) ) ;
NAND2   gate13627  (.A(WX3205), .B(II11580), .Z(II11581) ) ;
NAND2   gate13628  (.A(CRC_OUT_7_23), .B(II11580), .Z(II11582) ) ;
NAND2   gate13629  (.A(WX3206), .B(CRC_OUT_7_22), .Z(II11587) ) ;
NAND2   gate13630  (.A(WX3206), .B(II11587), .Z(II11588) ) ;
NAND2   gate13631  (.A(CRC_OUT_7_22), .B(II11587), .Z(II11589) ) ;
NAND2   gate13632  (.A(WX3207), .B(CRC_OUT_7_21), .Z(II11594) ) ;
NAND2   gate13633  (.A(WX3207), .B(II11594), .Z(II11595) ) ;
NAND2   gate13634  (.A(CRC_OUT_7_21), .B(II11594), .Z(II11596) ) ;
NAND2   gate13635  (.A(WX3208), .B(CRC_OUT_7_20), .Z(II11601) ) ;
NAND2   gate13636  (.A(WX3208), .B(II11601), .Z(II11602) ) ;
NAND2   gate13637  (.A(CRC_OUT_7_20), .B(II11601), .Z(II11603) ) ;
NAND2   gate13638  (.A(WX3209), .B(CRC_OUT_7_19), .Z(II11608) ) ;
NAND2   gate13639  (.A(WX3209), .B(II11608), .Z(II11609) ) ;
NAND2   gate13640  (.A(CRC_OUT_7_19), .B(II11608), .Z(II11610) ) ;
NAND2   gate13641  (.A(WX3210), .B(CRC_OUT_7_18), .Z(II11615) ) ;
NAND2   gate13642  (.A(WX3210), .B(II11615), .Z(II11616) ) ;
NAND2   gate13643  (.A(CRC_OUT_7_18), .B(II11615), .Z(II11617) ) ;
NAND2   gate13644  (.A(WX3211), .B(CRC_OUT_7_17), .Z(II11622) ) ;
NAND2   gate13645  (.A(WX3211), .B(II11622), .Z(II11623) ) ;
NAND2   gate13646  (.A(CRC_OUT_7_17), .B(II11622), .Z(II11624) ) ;
NAND2   gate13647  (.A(WX3212), .B(CRC_OUT_7_16), .Z(II11629) ) ;
NAND2   gate13648  (.A(WX3212), .B(II11629), .Z(II11630) ) ;
NAND2   gate13649  (.A(CRC_OUT_7_16), .B(II11629), .Z(II11631) ) ;
NAND2   gate13650  (.A(WX3214), .B(CRC_OUT_7_14), .Z(II11636) ) ;
NAND2   gate13651  (.A(WX3214), .B(II11636), .Z(II11637) ) ;
NAND2   gate13652  (.A(CRC_OUT_7_14), .B(II11636), .Z(II11638) ) ;
NAND2   gate13653  (.A(WX3215), .B(CRC_OUT_7_13), .Z(II11643) ) ;
NAND2   gate13654  (.A(WX3215), .B(II11643), .Z(II11644) ) ;
NAND2   gate13655  (.A(CRC_OUT_7_13), .B(II11643), .Z(II11645) ) ;
NAND2   gate13656  (.A(WX3216), .B(CRC_OUT_7_12), .Z(II11650) ) ;
NAND2   gate13657  (.A(WX3216), .B(II11650), .Z(II11651) ) ;
NAND2   gate13658  (.A(CRC_OUT_7_12), .B(II11650), .Z(II11652) ) ;
NAND2   gate13659  (.A(WX3217), .B(CRC_OUT_7_11), .Z(II11657) ) ;
NAND2   gate13660  (.A(WX3217), .B(II11657), .Z(II11658) ) ;
NAND2   gate13661  (.A(CRC_OUT_7_11), .B(II11657), .Z(II11659) ) ;
NAND2   gate13662  (.A(WX3219), .B(CRC_OUT_7_9), .Z(II11664) ) ;
NAND2   gate13663  (.A(WX3219), .B(II11664), .Z(II11665) ) ;
NAND2   gate13664  (.A(CRC_OUT_7_9), .B(II11664), .Z(II11666) ) ;
NAND2   gate13665  (.A(WX3220), .B(CRC_OUT_7_8), .Z(II11671) ) ;
NAND2   gate13666  (.A(WX3220), .B(II11671), .Z(II11672) ) ;
NAND2   gate13667  (.A(CRC_OUT_7_8), .B(II11671), .Z(II11673) ) ;
NAND2   gate13668  (.A(WX3221), .B(CRC_OUT_7_7), .Z(II11678) ) ;
NAND2   gate13669  (.A(WX3221), .B(II11678), .Z(II11679) ) ;
NAND2   gate13670  (.A(CRC_OUT_7_7), .B(II11678), .Z(II11680) ) ;
NAND2   gate13671  (.A(WX3222), .B(CRC_OUT_7_6), .Z(II11685) ) ;
NAND2   gate13672  (.A(WX3222), .B(II11685), .Z(II11686) ) ;
NAND2   gate13673  (.A(CRC_OUT_7_6), .B(II11685), .Z(II11687) ) ;
NAND2   gate13674  (.A(WX3223), .B(CRC_OUT_7_5), .Z(II11692) ) ;
NAND2   gate13675  (.A(WX3223), .B(II11692), .Z(II11693) ) ;
NAND2   gate13676  (.A(CRC_OUT_7_5), .B(II11692), .Z(II11694) ) ;
NAND2   gate13677  (.A(WX3224), .B(CRC_OUT_7_4), .Z(II11699) ) ;
NAND2   gate13678  (.A(WX3224), .B(II11699), .Z(II11700) ) ;
NAND2   gate13679  (.A(CRC_OUT_7_4), .B(II11699), .Z(II11701) ) ;
NAND2   gate13680  (.A(WX3226), .B(CRC_OUT_7_2), .Z(II11706) ) ;
NAND2   gate13681  (.A(WX3226), .B(II11706), .Z(II11707) ) ;
NAND2   gate13682  (.A(CRC_OUT_7_2), .B(II11706), .Z(II11708) ) ;
NAND2   gate13683  (.A(WX3227), .B(CRC_OUT_7_1), .Z(II11713) ) ;
NAND2   gate13684  (.A(WX3227), .B(II11713), .Z(II11714) ) ;
NAND2   gate13685  (.A(CRC_OUT_7_1), .B(II11713), .Z(II11715) ) ;
NAND2   gate13686  (.A(WX3228), .B(CRC_OUT_7_0), .Z(II11720) ) ;
NAND2   gate13687  (.A(WX3228), .B(II11720), .Z(II11721) ) ;
NAND2   gate13688  (.A(CRC_OUT_7_0), .B(II11720), .Z(II11722) ) ;
NAND2   gate13689  (.A(WX4880), .B(WX4524), .Z(II14003) ) ;
NAND2   gate13690  (.A(WX4880), .B(II14003), .Z(II14004) ) ;
NAND2   gate13691  (.A(WX4524), .B(II14003), .Z(II14005) ) ;
NAND2   gate13692  (.A(II14004), .B(II14005), .Z(II14002) ) ;
NAND2   gate13693  (.A(WX4588), .B(II14002), .Z(II14010) ) ;
NAND2   gate13694  (.A(WX4588), .B(II14010), .Z(II14011) ) ;
NAND2   gate13695  (.A(II14002), .B(II14010), .Z(II14012) ) ;
NAND2   gate13696  (.A(II14011), .B(II14012), .Z(II14001) ) ;
NAND2   gate13697  (.A(WX4652), .B(WX4716), .Z(II14018) ) ;
NAND2   gate13698  (.A(WX4652), .B(II14018), .Z(II14019) ) ;
NAND2   gate13699  (.A(WX4716), .B(II14018), .Z(II14020) ) ;
NAND2   gate13700  (.A(II14019), .B(II14020), .Z(II14017) ) ;
NAND2   gate13701  (.A(II14001), .B(II14017), .Z(II14025) ) ;
NAND2   gate13702  (.A(II14001), .B(II14025), .Z(II14026) ) ;
NAND2   gate13703  (.A(II14017), .B(II14025), .Z(II14027) ) ;
NAND2   gate13704  (.A(WX4880), .B(WX4526), .Z(II14034) ) ;
NAND2   gate13705  (.A(WX4880), .B(II14034), .Z(II14035) ) ;
NAND2   gate13706  (.A(WX4526), .B(II14034), .Z(II14036) ) ;
NAND2   gate13707  (.A(II14035), .B(II14036), .Z(II14033) ) ;
NAND2   gate13708  (.A(WX4590), .B(II14033), .Z(II14041) ) ;
NAND2   gate13709  (.A(WX4590), .B(II14041), .Z(II14042) ) ;
NAND2   gate13710  (.A(II14033), .B(II14041), .Z(II14043) ) ;
NAND2   gate13711  (.A(II14042), .B(II14043), .Z(II14032) ) ;
NAND2   gate13712  (.A(WX4654), .B(WX4718), .Z(II14049) ) ;
NAND2   gate13713  (.A(WX4654), .B(II14049), .Z(II14050) ) ;
NAND2   gate13714  (.A(WX4718), .B(II14049), .Z(II14051) ) ;
NAND2   gate13715  (.A(II14050), .B(II14051), .Z(II14048) ) ;
NAND2   gate13716  (.A(II14032), .B(II14048), .Z(II14056) ) ;
NAND2   gate13717  (.A(II14032), .B(II14056), .Z(II14057) ) ;
NAND2   gate13718  (.A(II14048), .B(II14056), .Z(II14058) ) ;
NAND2   gate13719  (.A(WX4880), .B(WX4528), .Z(II14065) ) ;
NAND2   gate13720  (.A(WX4880), .B(II14065), .Z(II14066) ) ;
NAND2   gate13721  (.A(WX4528), .B(II14065), .Z(II14067) ) ;
NAND2   gate13722  (.A(II14066), .B(II14067), .Z(II14064) ) ;
NAND2   gate13723  (.A(WX4592), .B(II14064), .Z(II14072) ) ;
NAND2   gate13724  (.A(WX4592), .B(II14072), .Z(II14073) ) ;
NAND2   gate13725  (.A(II14064), .B(II14072), .Z(II14074) ) ;
NAND2   gate13726  (.A(II14073), .B(II14074), .Z(II14063) ) ;
NAND2   gate13727  (.A(WX4656), .B(WX4720), .Z(II14080) ) ;
NAND2   gate13728  (.A(WX4656), .B(II14080), .Z(II14081) ) ;
NAND2   gate13729  (.A(WX4720), .B(II14080), .Z(II14082) ) ;
NAND2   gate13730  (.A(II14081), .B(II14082), .Z(II14079) ) ;
NAND2   gate13731  (.A(II14063), .B(II14079), .Z(II14087) ) ;
NAND2   gate13732  (.A(II14063), .B(II14087), .Z(II14088) ) ;
NAND2   gate13733  (.A(II14079), .B(II14087), .Z(II14089) ) ;
NAND2   gate13734  (.A(WX4880), .B(WX4530), .Z(II14096) ) ;
NAND2   gate13735  (.A(WX4880), .B(II14096), .Z(II14097) ) ;
NAND2   gate13736  (.A(WX4530), .B(II14096), .Z(II14098) ) ;
NAND2   gate13737  (.A(II14097), .B(II14098), .Z(II14095) ) ;
NAND2   gate13738  (.A(WX4594), .B(II14095), .Z(II14103) ) ;
NAND2   gate13739  (.A(WX4594), .B(II14103), .Z(II14104) ) ;
NAND2   gate13740  (.A(II14095), .B(II14103), .Z(II14105) ) ;
NAND2   gate13741  (.A(II14104), .B(II14105), .Z(II14094) ) ;
NAND2   gate13742  (.A(WX4658), .B(WX4722), .Z(II14111) ) ;
NAND2   gate13743  (.A(WX4658), .B(II14111), .Z(II14112) ) ;
NAND2   gate13744  (.A(WX4722), .B(II14111), .Z(II14113) ) ;
NAND2   gate13745  (.A(II14112), .B(II14113), .Z(II14110) ) ;
NAND2   gate13746  (.A(II14094), .B(II14110), .Z(II14118) ) ;
NAND2   gate13747  (.A(II14094), .B(II14118), .Z(II14119) ) ;
NAND2   gate13748  (.A(II14110), .B(II14118), .Z(II14120) ) ;
NAND2   gate13749  (.A(WX4880), .B(WX4532), .Z(II14127) ) ;
NAND2   gate13750  (.A(WX4880), .B(II14127), .Z(II14128) ) ;
NAND2   gate13751  (.A(WX4532), .B(II14127), .Z(II14129) ) ;
NAND2   gate13752  (.A(II14128), .B(II14129), .Z(II14126) ) ;
NAND2   gate13753  (.A(WX4596), .B(II14126), .Z(II14134) ) ;
NAND2   gate13754  (.A(WX4596), .B(II14134), .Z(II14135) ) ;
NAND2   gate13755  (.A(II14126), .B(II14134), .Z(II14136) ) ;
NAND2   gate13756  (.A(II14135), .B(II14136), .Z(II14125) ) ;
NAND2   gate13757  (.A(WX4660), .B(WX4724), .Z(II14142) ) ;
NAND2   gate13758  (.A(WX4660), .B(II14142), .Z(II14143) ) ;
NAND2   gate13759  (.A(WX4724), .B(II14142), .Z(II14144) ) ;
NAND2   gate13760  (.A(II14143), .B(II14144), .Z(II14141) ) ;
NAND2   gate13761  (.A(II14125), .B(II14141), .Z(II14149) ) ;
NAND2   gate13762  (.A(II14125), .B(II14149), .Z(II14150) ) ;
NAND2   gate13763  (.A(II14141), .B(II14149), .Z(II14151) ) ;
NAND2   gate13764  (.A(WX4880), .B(WX4534), .Z(II14158) ) ;
NAND2   gate13765  (.A(WX4880), .B(II14158), .Z(II14159) ) ;
NAND2   gate13766  (.A(WX4534), .B(II14158), .Z(II14160) ) ;
NAND2   gate13767  (.A(II14159), .B(II14160), .Z(II14157) ) ;
NAND2   gate13768  (.A(WX4598), .B(II14157), .Z(II14165) ) ;
NAND2   gate13769  (.A(WX4598), .B(II14165), .Z(II14166) ) ;
NAND2   gate13770  (.A(II14157), .B(II14165), .Z(II14167) ) ;
NAND2   gate13771  (.A(II14166), .B(II14167), .Z(II14156) ) ;
NAND2   gate13772  (.A(WX4662), .B(WX4726), .Z(II14173) ) ;
NAND2   gate13773  (.A(WX4662), .B(II14173), .Z(II14174) ) ;
NAND2   gate13774  (.A(WX4726), .B(II14173), .Z(II14175) ) ;
NAND2   gate13775  (.A(II14174), .B(II14175), .Z(II14172) ) ;
NAND2   gate13776  (.A(II14156), .B(II14172), .Z(II14180) ) ;
NAND2   gate13777  (.A(II14156), .B(II14180), .Z(II14181) ) ;
NAND2   gate13778  (.A(II14172), .B(II14180), .Z(II14182) ) ;
NAND2   gate13779  (.A(WX4880), .B(WX4536), .Z(II14189) ) ;
NAND2   gate13780  (.A(WX4880), .B(II14189), .Z(II14190) ) ;
NAND2   gate13781  (.A(WX4536), .B(II14189), .Z(II14191) ) ;
NAND2   gate13782  (.A(II14190), .B(II14191), .Z(II14188) ) ;
NAND2   gate13783  (.A(WX4600), .B(II14188), .Z(II14196) ) ;
NAND2   gate13784  (.A(WX4600), .B(II14196), .Z(II14197) ) ;
NAND2   gate13785  (.A(II14188), .B(II14196), .Z(II14198) ) ;
NAND2   gate13786  (.A(II14197), .B(II14198), .Z(II14187) ) ;
NAND2   gate13787  (.A(WX4664), .B(WX4728), .Z(II14204) ) ;
NAND2   gate13788  (.A(WX4664), .B(II14204), .Z(II14205) ) ;
NAND2   gate13789  (.A(WX4728), .B(II14204), .Z(II14206) ) ;
NAND2   gate13790  (.A(II14205), .B(II14206), .Z(II14203) ) ;
NAND2   gate13791  (.A(II14187), .B(II14203), .Z(II14211) ) ;
NAND2   gate13792  (.A(II14187), .B(II14211), .Z(II14212) ) ;
NAND2   gate13793  (.A(II14203), .B(II14211), .Z(II14213) ) ;
NAND2   gate13794  (.A(WX4880), .B(WX4538), .Z(II14220) ) ;
NAND2   gate13795  (.A(WX4880), .B(II14220), .Z(II14221) ) ;
NAND2   gate13796  (.A(WX4538), .B(II14220), .Z(II14222) ) ;
NAND2   gate13797  (.A(II14221), .B(II14222), .Z(II14219) ) ;
NAND2   gate13798  (.A(WX4602), .B(II14219), .Z(II14227) ) ;
NAND2   gate13799  (.A(WX4602), .B(II14227), .Z(II14228) ) ;
NAND2   gate13800  (.A(II14219), .B(II14227), .Z(II14229) ) ;
NAND2   gate13801  (.A(II14228), .B(II14229), .Z(II14218) ) ;
NAND2   gate13802  (.A(WX4666), .B(WX4730), .Z(II14235) ) ;
NAND2   gate13803  (.A(WX4666), .B(II14235), .Z(II14236) ) ;
NAND2   gate13804  (.A(WX4730), .B(II14235), .Z(II14237) ) ;
NAND2   gate13805  (.A(II14236), .B(II14237), .Z(II14234) ) ;
NAND2   gate13806  (.A(II14218), .B(II14234), .Z(II14242) ) ;
NAND2   gate13807  (.A(II14218), .B(II14242), .Z(II14243) ) ;
NAND2   gate13808  (.A(II14234), .B(II14242), .Z(II14244) ) ;
NAND2   gate13809  (.A(WX4880), .B(WX4540), .Z(II14251) ) ;
NAND2   gate13810  (.A(WX4880), .B(II14251), .Z(II14252) ) ;
NAND2   gate13811  (.A(WX4540), .B(II14251), .Z(II14253) ) ;
NAND2   gate13812  (.A(II14252), .B(II14253), .Z(II14250) ) ;
NAND2   gate13813  (.A(WX4604), .B(II14250), .Z(II14258) ) ;
NAND2   gate13814  (.A(WX4604), .B(II14258), .Z(II14259) ) ;
NAND2   gate13815  (.A(II14250), .B(II14258), .Z(II14260) ) ;
NAND2   gate13816  (.A(II14259), .B(II14260), .Z(II14249) ) ;
NAND2   gate13817  (.A(WX4668), .B(WX4732), .Z(II14266) ) ;
NAND2   gate13818  (.A(WX4668), .B(II14266), .Z(II14267) ) ;
NAND2   gate13819  (.A(WX4732), .B(II14266), .Z(II14268) ) ;
NAND2   gate13820  (.A(II14267), .B(II14268), .Z(II14265) ) ;
NAND2   gate13821  (.A(II14249), .B(II14265), .Z(II14273) ) ;
NAND2   gate13822  (.A(II14249), .B(II14273), .Z(II14274) ) ;
NAND2   gate13823  (.A(II14265), .B(II14273), .Z(II14275) ) ;
NAND2   gate13824  (.A(WX4880), .B(WX4542), .Z(II14282) ) ;
NAND2   gate13825  (.A(WX4880), .B(II14282), .Z(II14283) ) ;
NAND2   gate13826  (.A(WX4542), .B(II14282), .Z(II14284) ) ;
NAND2   gate13827  (.A(II14283), .B(II14284), .Z(II14281) ) ;
NAND2   gate13828  (.A(WX4606), .B(II14281), .Z(II14289) ) ;
NAND2   gate13829  (.A(WX4606), .B(II14289), .Z(II14290) ) ;
NAND2   gate13830  (.A(II14281), .B(II14289), .Z(II14291) ) ;
NAND2   gate13831  (.A(II14290), .B(II14291), .Z(II14280) ) ;
NAND2   gate13832  (.A(WX4670), .B(WX4734), .Z(II14297) ) ;
NAND2   gate13833  (.A(WX4670), .B(II14297), .Z(II14298) ) ;
NAND2   gate13834  (.A(WX4734), .B(II14297), .Z(II14299) ) ;
NAND2   gate13835  (.A(II14298), .B(II14299), .Z(II14296) ) ;
NAND2   gate13836  (.A(II14280), .B(II14296), .Z(II14304) ) ;
NAND2   gate13837  (.A(II14280), .B(II14304), .Z(II14305) ) ;
NAND2   gate13838  (.A(II14296), .B(II14304), .Z(II14306) ) ;
NAND2   gate13839  (.A(WX4880), .B(WX4544), .Z(II14313) ) ;
NAND2   gate13840  (.A(WX4880), .B(II14313), .Z(II14314) ) ;
NAND2   gate13841  (.A(WX4544), .B(II14313), .Z(II14315) ) ;
NAND2   gate13842  (.A(II14314), .B(II14315), .Z(II14312) ) ;
NAND2   gate13843  (.A(WX4608), .B(II14312), .Z(II14320) ) ;
NAND2   gate13844  (.A(WX4608), .B(II14320), .Z(II14321) ) ;
NAND2   gate13845  (.A(II14312), .B(II14320), .Z(II14322) ) ;
NAND2   gate13846  (.A(II14321), .B(II14322), .Z(II14311) ) ;
NAND2   gate13847  (.A(WX4672), .B(WX4736), .Z(II14328) ) ;
NAND2   gate13848  (.A(WX4672), .B(II14328), .Z(II14329) ) ;
NAND2   gate13849  (.A(WX4736), .B(II14328), .Z(II14330) ) ;
NAND2   gate13850  (.A(II14329), .B(II14330), .Z(II14327) ) ;
NAND2   gate13851  (.A(II14311), .B(II14327), .Z(II14335) ) ;
NAND2   gate13852  (.A(II14311), .B(II14335), .Z(II14336) ) ;
NAND2   gate13853  (.A(II14327), .B(II14335), .Z(II14337) ) ;
NAND2   gate13854  (.A(WX4880), .B(WX4546), .Z(II14344) ) ;
NAND2   gate13855  (.A(WX4880), .B(II14344), .Z(II14345) ) ;
NAND2   gate13856  (.A(WX4546), .B(II14344), .Z(II14346) ) ;
NAND2   gate13857  (.A(II14345), .B(II14346), .Z(II14343) ) ;
NAND2   gate13858  (.A(WX4610), .B(II14343), .Z(II14351) ) ;
NAND2   gate13859  (.A(WX4610), .B(II14351), .Z(II14352) ) ;
NAND2   gate13860  (.A(II14343), .B(II14351), .Z(II14353) ) ;
NAND2   gate13861  (.A(II14352), .B(II14353), .Z(II14342) ) ;
NAND2   gate13862  (.A(WX4674), .B(WX4738), .Z(II14359) ) ;
NAND2   gate13863  (.A(WX4674), .B(II14359), .Z(II14360) ) ;
NAND2   gate13864  (.A(WX4738), .B(II14359), .Z(II14361) ) ;
NAND2   gate13865  (.A(II14360), .B(II14361), .Z(II14358) ) ;
NAND2   gate13866  (.A(II14342), .B(II14358), .Z(II14366) ) ;
NAND2   gate13867  (.A(II14342), .B(II14366), .Z(II14367) ) ;
NAND2   gate13868  (.A(II14358), .B(II14366), .Z(II14368) ) ;
NAND2   gate13869  (.A(WX4880), .B(WX4548), .Z(II14375) ) ;
NAND2   gate13870  (.A(WX4880), .B(II14375), .Z(II14376) ) ;
NAND2   gate13871  (.A(WX4548), .B(II14375), .Z(II14377) ) ;
NAND2   gate13872  (.A(II14376), .B(II14377), .Z(II14374) ) ;
NAND2   gate13873  (.A(WX4612), .B(II14374), .Z(II14382) ) ;
NAND2   gate13874  (.A(WX4612), .B(II14382), .Z(II14383) ) ;
NAND2   gate13875  (.A(II14374), .B(II14382), .Z(II14384) ) ;
NAND2   gate13876  (.A(II14383), .B(II14384), .Z(II14373) ) ;
NAND2   gate13877  (.A(WX4676), .B(WX4740), .Z(II14390) ) ;
NAND2   gate13878  (.A(WX4676), .B(II14390), .Z(II14391) ) ;
NAND2   gate13879  (.A(WX4740), .B(II14390), .Z(II14392) ) ;
NAND2   gate13880  (.A(II14391), .B(II14392), .Z(II14389) ) ;
NAND2   gate13881  (.A(II14373), .B(II14389), .Z(II14397) ) ;
NAND2   gate13882  (.A(II14373), .B(II14397), .Z(II14398) ) ;
NAND2   gate13883  (.A(II14389), .B(II14397), .Z(II14399) ) ;
NAND2   gate13884  (.A(WX4880), .B(WX4550), .Z(II14406) ) ;
NAND2   gate13885  (.A(WX4880), .B(II14406), .Z(II14407) ) ;
NAND2   gate13886  (.A(WX4550), .B(II14406), .Z(II14408) ) ;
NAND2   gate13887  (.A(II14407), .B(II14408), .Z(II14405) ) ;
NAND2   gate13888  (.A(WX4614), .B(II14405), .Z(II14413) ) ;
NAND2   gate13889  (.A(WX4614), .B(II14413), .Z(II14414) ) ;
NAND2   gate13890  (.A(II14405), .B(II14413), .Z(II14415) ) ;
NAND2   gate13891  (.A(II14414), .B(II14415), .Z(II14404) ) ;
NAND2   gate13892  (.A(WX4678), .B(WX4742), .Z(II14421) ) ;
NAND2   gate13893  (.A(WX4678), .B(II14421), .Z(II14422) ) ;
NAND2   gate13894  (.A(WX4742), .B(II14421), .Z(II14423) ) ;
NAND2   gate13895  (.A(II14422), .B(II14423), .Z(II14420) ) ;
NAND2   gate13896  (.A(II14404), .B(II14420), .Z(II14428) ) ;
NAND2   gate13897  (.A(II14404), .B(II14428), .Z(II14429) ) ;
NAND2   gate13898  (.A(II14420), .B(II14428), .Z(II14430) ) ;
NAND2   gate13899  (.A(WX4880), .B(WX4552), .Z(II14437) ) ;
NAND2   gate13900  (.A(WX4880), .B(II14437), .Z(II14438) ) ;
NAND2   gate13901  (.A(WX4552), .B(II14437), .Z(II14439) ) ;
NAND2   gate13902  (.A(II14438), .B(II14439), .Z(II14436) ) ;
NAND2   gate13903  (.A(WX4616), .B(II14436), .Z(II14444) ) ;
NAND2   gate13904  (.A(WX4616), .B(II14444), .Z(II14445) ) ;
NAND2   gate13905  (.A(II14436), .B(II14444), .Z(II14446) ) ;
NAND2   gate13906  (.A(II14445), .B(II14446), .Z(II14435) ) ;
NAND2   gate13907  (.A(WX4680), .B(WX4744), .Z(II14452) ) ;
NAND2   gate13908  (.A(WX4680), .B(II14452), .Z(II14453) ) ;
NAND2   gate13909  (.A(WX4744), .B(II14452), .Z(II14454) ) ;
NAND2   gate13910  (.A(II14453), .B(II14454), .Z(II14451) ) ;
NAND2   gate13911  (.A(II14435), .B(II14451), .Z(II14459) ) ;
NAND2   gate13912  (.A(II14435), .B(II14459), .Z(II14460) ) ;
NAND2   gate13913  (.A(II14451), .B(II14459), .Z(II14461) ) ;
NAND2   gate13914  (.A(WX4880), .B(WX4554), .Z(II14468) ) ;
NAND2   gate13915  (.A(WX4880), .B(II14468), .Z(II14469) ) ;
NAND2   gate13916  (.A(WX4554), .B(II14468), .Z(II14470) ) ;
NAND2   gate13917  (.A(II14469), .B(II14470), .Z(II14467) ) ;
NAND2   gate13918  (.A(WX4618), .B(II14467), .Z(II14475) ) ;
NAND2   gate13919  (.A(WX4618), .B(II14475), .Z(II14476) ) ;
NAND2   gate13920  (.A(II14467), .B(II14475), .Z(II14477) ) ;
NAND2   gate13921  (.A(II14476), .B(II14477), .Z(II14466) ) ;
NAND2   gate13922  (.A(WX4682), .B(WX4746), .Z(II14483) ) ;
NAND2   gate13923  (.A(WX4682), .B(II14483), .Z(II14484) ) ;
NAND2   gate13924  (.A(WX4746), .B(II14483), .Z(II14485) ) ;
NAND2   gate13925  (.A(II14484), .B(II14485), .Z(II14482) ) ;
NAND2   gate13926  (.A(II14466), .B(II14482), .Z(II14490) ) ;
NAND2   gate13927  (.A(II14466), .B(II14490), .Z(II14491) ) ;
NAND2   gate13928  (.A(II14482), .B(II14490), .Z(II14492) ) ;
NAND2   gate13929  (.A(WX4881), .B(WX4556), .Z(II14499) ) ;
NAND2   gate13930  (.A(WX4881), .B(II14499), .Z(II14500) ) ;
NAND2   gate13931  (.A(WX4556), .B(II14499), .Z(II14501) ) ;
NAND2   gate13932  (.A(II14500), .B(II14501), .Z(II14498) ) ;
NAND2   gate13933  (.A(WX4620), .B(II14498), .Z(II14506) ) ;
NAND2   gate13934  (.A(WX4620), .B(II14506), .Z(II14507) ) ;
NAND2   gate13935  (.A(II14498), .B(II14506), .Z(II14508) ) ;
NAND2   gate13936  (.A(II14507), .B(II14508), .Z(II14497) ) ;
NAND2   gate13937  (.A(WX4684), .B(WX4748), .Z(II14514) ) ;
NAND2   gate13938  (.A(WX4684), .B(II14514), .Z(II14515) ) ;
NAND2   gate13939  (.A(WX4748), .B(II14514), .Z(II14516) ) ;
NAND2   gate13940  (.A(II14515), .B(II14516), .Z(II14513) ) ;
NAND2   gate13941  (.A(II14497), .B(II14513), .Z(II14521) ) ;
NAND2   gate13942  (.A(II14497), .B(II14521), .Z(II14522) ) ;
NAND2   gate13943  (.A(II14513), .B(II14521), .Z(II14523) ) ;
NAND2   gate13944  (.A(WX4881), .B(WX4558), .Z(II14530) ) ;
NAND2   gate13945  (.A(WX4881), .B(II14530), .Z(II14531) ) ;
NAND2   gate13946  (.A(WX4558), .B(II14530), .Z(II14532) ) ;
NAND2   gate13947  (.A(II14531), .B(II14532), .Z(II14529) ) ;
NAND2   gate13948  (.A(WX4622), .B(II14529), .Z(II14537) ) ;
NAND2   gate13949  (.A(WX4622), .B(II14537), .Z(II14538) ) ;
NAND2   gate13950  (.A(II14529), .B(II14537), .Z(II14539) ) ;
NAND2   gate13951  (.A(II14538), .B(II14539), .Z(II14528) ) ;
NAND2   gate13952  (.A(WX4686), .B(WX4750), .Z(II14545) ) ;
NAND2   gate13953  (.A(WX4686), .B(II14545), .Z(II14546) ) ;
NAND2   gate13954  (.A(WX4750), .B(II14545), .Z(II14547) ) ;
NAND2   gate13955  (.A(II14546), .B(II14547), .Z(II14544) ) ;
NAND2   gate13956  (.A(II14528), .B(II14544), .Z(II14552) ) ;
NAND2   gate13957  (.A(II14528), .B(II14552), .Z(II14553) ) ;
NAND2   gate13958  (.A(II14544), .B(II14552), .Z(II14554) ) ;
NAND2   gate13959  (.A(WX4881), .B(WX4560), .Z(II14561) ) ;
NAND2   gate13960  (.A(WX4881), .B(II14561), .Z(II14562) ) ;
NAND2   gate13961  (.A(WX4560), .B(II14561), .Z(II14563) ) ;
NAND2   gate13962  (.A(II14562), .B(II14563), .Z(II14560) ) ;
NAND2   gate13963  (.A(WX4624), .B(II14560), .Z(II14568) ) ;
NAND2   gate13964  (.A(WX4624), .B(II14568), .Z(II14569) ) ;
NAND2   gate13965  (.A(II14560), .B(II14568), .Z(II14570) ) ;
NAND2   gate13966  (.A(II14569), .B(II14570), .Z(II14559) ) ;
NAND2   gate13967  (.A(WX4688), .B(WX4752), .Z(II14576) ) ;
NAND2   gate13968  (.A(WX4688), .B(II14576), .Z(II14577) ) ;
NAND2   gate13969  (.A(WX4752), .B(II14576), .Z(II14578) ) ;
NAND2   gate13970  (.A(II14577), .B(II14578), .Z(II14575) ) ;
NAND2   gate13971  (.A(II14559), .B(II14575), .Z(II14583) ) ;
NAND2   gate13972  (.A(II14559), .B(II14583), .Z(II14584) ) ;
NAND2   gate13973  (.A(II14575), .B(II14583), .Z(II14585) ) ;
NAND2   gate13974  (.A(WX4881), .B(WX4562), .Z(II14592) ) ;
NAND2   gate13975  (.A(WX4881), .B(II14592), .Z(II14593) ) ;
NAND2   gate13976  (.A(WX4562), .B(II14592), .Z(II14594) ) ;
NAND2   gate13977  (.A(II14593), .B(II14594), .Z(II14591) ) ;
NAND2   gate13978  (.A(WX4626), .B(II14591), .Z(II14599) ) ;
NAND2   gate13979  (.A(WX4626), .B(II14599), .Z(II14600) ) ;
NAND2   gate13980  (.A(II14591), .B(II14599), .Z(II14601) ) ;
NAND2   gate13981  (.A(II14600), .B(II14601), .Z(II14590) ) ;
NAND2   gate13982  (.A(WX4690), .B(WX4754), .Z(II14607) ) ;
NAND2   gate13983  (.A(WX4690), .B(II14607), .Z(II14608) ) ;
NAND2   gate13984  (.A(WX4754), .B(II14607), .Z(II14609) ) ;
NAND2   gate13985  (.A(II14608), .B(II14609), .Z(II14606) ) ;
NAND2   gate13986  (.A(II14590), .B(II14606), .Z(II14614) ) ;
NAND2   gate13987  (.A(II14590), .B(II14614), .Z(II14615) ) ;
NAND2   gate13988  (.A(II14606), .B(II14614), .Z(II14616) ) ;
NAND2   gate13989  (.A(WX4881), .B(WX4564), .Z(II14623) ) ;
NAND2   gate13990  (.A(WX4881), .B(II14623), .Z(II14624) ) ;
NAND2   gate13991  (.A(WX4564), .B(II14623), .Z(II14625) ) ;
NAND2   gate13992  (.A(II14624), .B(II14625), .Z(II14622) ) ;
NAND2   gate13993  (.A(WX4628), .B(II14622), .Z(II14630) ) ;
NAND2   gate13994  (.A(WX4628), .B(II14630), .Z(II14631) ) ;
NAND2   gate13995  (.A(II14622), .B(II14630), .Z(II14632) ) ;
NAND2   gate13996  (.A(II14631), .B(II14632), .Z(II14621) ) ;
NAND2   gate13997  (.A(WX4692), .B(WX4756), .Z(II14638) ) ;
NAND2   gate13998  (.A(WX4692), .B(II14638), .Z(II14639) ) ;
NAND2   gate13999  (.A(WX4756), .B(II14638), .Z(II14640) ) ;
NAND2   gate14000  (.A(II14639), .B(II14640), .Z(II14637) ) ;
NAND2   gate14001  (.A(II14621), .B(II14637), .Z(II14645) ) ;
NAND2   gate14002  (.A(II14621), .B(II14645), .Z(II14646) ) ;
NAND2   gate14003  (.A(II14637), .B(II14645), .Z(II14647) ) ;
NAND2   gate14004  (.A(WX4881), .B(WX4566), .Z(II14654) ) ;
NAND2   gate14005  (.A(WX4881), .B(II14654), .Z(II14655) ) ;
NAND2   gate14006  (.A(WX4566), .B(II14654), .Z(II14656) ) ;
NAND2   gate14007  (.A(II14655), .B(II14656), .Z(II14653) ) ;
NAND2   gate14008  (.A(WX4630), .B(II14653), .Z(II14661) ) ;
NAND2   gate14009  (.A(WX4630), .B(II14661), .Z(II14662) ) ;
NAND2   gate14010  (.A(II14653), .B(II14661), .Z(II14663) ) ;
NAND2   gate14011  (.A(II14662), .B(II14663), .Z(II14652) ) ;
NAND2   gate14012  (.A(WX4694), .B(WX4758), .Z(II14669) ) ;
NAND2   gate14013  (.A(WX4694), .B(II14669), .Z(II14670) ) ;
NAND2   gate14014  (.A(WX4758), .B(II14669), .Z(II14671) ) ;
NAND2   gate14015  (.A(II14670), .B(II14671), .Z(II14668) ) ;
NAND2   gate14016  (.A(II14652), .B(II14668), .Z(II14676) ) ;
NAND2   gate14017  (.A(II14652), .B(II14676), .Z(II14677) ) ;
NAND2   gate14018  (.A(II14668), .B(II14676), .Z(II14678) ) ;
NAND2   gate14019  (.A(WX4881), .B(WX4568), .Z(II14685) ) ;
NAND2   gate14020  (.A(WX4881), .B(II14685), .Z(II14686) ) ;
NAND2   gate14021  (.A(WX4568), .B(II14685), .Z(II14687) ) ;
NAND2   gate14022  (.A(II14686), .B(II14687), .Z(II14684) ) ;
NAND2   gate14023  (.A(WX4632), .B(II14684), .Z(II14692) ) ;
NAND2   gate14024  (.A(WX4632), .B(II14692), .Z(II14693) ) ;
NAND2   gate14025  (.A(II14684), .B(II14692), .Z(II14694) ) ;
NAND2   gate14026  (.A(II14693), .B(II14694), .Z(II14683) ) ;
NAND2   gate14027  (.A(WX4696), .B(WX4760), .Z(II14700) ) ;
NAND2   gate14028  (.A(WX4696), .B(II14700), .Z(II14701) ) ;
NAND2   gate14029  (.A(WX4760), .B(II14700), .Z(II14702) ) ;
NAND2   gate14030  (.A(II14701), .B(II14702), .Z(II14699) ) ;
NAND2   gate14031  (.A(II14683), .B(II14699), .Z(II14707) ) ;
NAND2   gate14032  (.A(II14683), .B(II14707), .Z(II14708) ) ;
NAND2   gate14033  (.A(II14699), .B(II14707), .Z(II14709) ) ;
NAND2   gate14034  (.A(WX4881), .B(WX4570), .Z(II14716) ) ;
NAND2   gate14035  (.A(WX4881), .B(II14716), .Z(II14717) ) ;
NAND2   gate14036  (.A(WX4570), .B(II14716), .Z(II14718) ) ;
NAND2   gate14037  (.A(II14717), .B(II14718), .Z(II14715) ) ;
NAND2   gate14038  (.A(WX4634), .B(II14715), .Z(II14723) ) ;
NAND2   gate14039  (.A(WX4634), .B(II14723), .Z(II14724) ) ;
NAND2   gate14040  (.A(II14715), .B(II14723), .Z(II14725) ) ;
NAND2   gate14041  (.A(II14724), .B(II14725), .Z(II14714) ) ;
NAND2   gate14042  (.A(WX4698), .B(WX4762), .Z(II14731) ) ;
NAND2   gate14043  (.A(WX4698), .B(II14731), .Z(II14732) ) ;
NAND2   gate14044  (.A(WX4762), .B(II14731), .Z(II14733) ) ;
NAND2   gate14045  (.A(II14732), .B(II14733), .Z(II14730) ) ;
NAND2   gate14046  (.A(II14714), .B(II14730), .Z(II14738) ) ;
NAND2   gate14047  (.A(II14714), .B(II14738), .Z(II14739) ) ;
NAND2   gate14048  (.A(II14730), .B(II14738), .Z(II14740) ) ;
NAND2   gate14049  (.A(WX4881), .B(WX4572), .Z(II14747) ) ;
NAND2   gate14050  (.A(WX4881), .B(II14747), .Z(II14748) ) ;
NAND2   gate14051  (.A(WX4572), .B(II14747), .Z(II14749) ) ;
NAND2   gate14052  (.A(II14748), .B(II14749), .Z(II14746) ) ;
NAND2   gate14053  (.A(WX4636), .B(II14746), .Z(II14754) ) ;
NAND2   gate14054  (.A(WX4636), .B(II14754), .Z(II14755) ) ;
NAND2   gate14055  (.A(II14746), .B(II14754), .Z(II14756) ) ;
NAND2   gate14056  (.A(II14755), .B(II14756), .Z(II14745) ) ;
NAND2   gate14057  (.A(WX4700), .B(WX4764), .Z(II14762) ) ;
NAND2   gate14058  (.A(WX4700), .B(II14762), .Z(II14763) ) ;
NAND2   gate14059  (.A(WX4764), .B(II14762), .Z(II14764) ) ;
NAND2   gate14060  (.A(II14763), .B(II14764), .Z(II14761) ) ;
NAND2   gate14061  (.A(II14745), .B(II14761), .Z(II14769) ) ;
NAND2   gate14062  (.A(II14745), .B(II14769), .Z(II14770) ) ;
NAND2   gate14063  (.A(II14761), .B(II14769), .Z(II14771) ) ;
NAND2   gate14064  (.A(WX4881), .B(WX4574), .Z(II14778) ) ;
NAND2   gate14065  (.A(WX4881), .B(II14778), .Z(II14779) ) ;
NAND2   gate14066  (.A(WX4574), .B(II14778), .Z(II14780) ) ;
NAND2   gate14067  (.A(II14779), .B(II14780), .Z(II14777) ) ;
NAND2   gate14068  (.A(WX4638), .B(II14777), .Z(II14785) ) ;
NAND2   gate14069  (.A(WX4638), .B(II14785), .Z(II14786) ) ;
NAND2   gate14070  (.A(II14777), .B(II14785), .Z(II14787) ) ;
NAND2   gate14071  (.A(II14786), .B(II14787), .Z(II14776) ) ;
NAND2   gate14072  (.A(WX4702), .B(WX4766), .Z(II14793) ) ;
NAND2   gate14073  (.A(WX4702), .B(II14793), .Z(II14794) ) ;
NAND2   gate14074  (.A(WX4766), .B(II14793), .Z(II14795) ) ;
NAND2   gate14075  (.A(II14794), .B(II14795), .Z(II14792) ) ;
NAND2   gate14076  (.A(II14776), .B(II14792), .Z(II14800) ) ;
NAND2   gate14077  (.A(II14776), .B(II14800), .Z(II14801) ) ;
NAND2   gate14078  (.A(II14792), .B(II14800), .Z(II14802) ) ;
NAND2   gate14079  (.A(WX4881), .B(WX4576), .Z(II14809) ) ;
NAND2   gate14080  (.A(WX4881), .B(II14809), .Z(II14810) ) ;
NAND2   gate14081  (.A(WX4576), .B(II14809), .Z(II14811) ) ;
NAND2   gate14082  (.A(II14810), .B(II14811), .Z(II14808) ) ;
NAND2   gate14083  (.A(WX4640), .B(II14808), .Z(II14816) ) ;
NAND2   gate14084  (.A(WX4640), .B(II14816), .Z(II14817) ) ;
NAND2   gate14085  (.A(II14808), .B(II14816), .Z(II14818) ) ;
NAND2   gate14086  (.A(II14817), .B(II14818), .Z(II14807) ) ;
NAND2   gate14087  (.A(WX4704), .B(WX4768), .Z(II14824) ) ;
NAND2   gate14088  (.A(WX4704), .B(II14824), .Z(II14825) ) ;
NAND2   gate14089  (.A(WX4768), .B(II14824), .Z(II14826) ) ;
NAND2   gate14090  (.A(II14825), .B(II14826), .Z(II14823) ) ;
NAND2   gate14091  (.A(II14807), .B(II14823), .Z(II14831) ) ;
NAND2   gate14092  (.A(II14807), .B(II14831), .Z(II14832) ) ;
NAND2   gate14093  (.A(II14823), .B(II14831), .Z(II14833) ) ;
NAND2   gate14094  (.A(WX4881), .B(WX4578), .Z(II14840) ) ;
NAND2   gate14095  (.A(WX4881), .B(II14840), .Z(II14841) ) ;
NAND2   gate14096  (.A(WX4578), .B(II14840), .Z(II14842) ) ;
NAND2   gate14097  (.A(II14841), .B(II14842), .Z(II14839) ) ;
NAND2   gate14098  (.A(WX4642), .B(II14839), .Z(II14847) ) ;
NAND2   gate14099  (.A(WX4642), .B(II14847), .Z(II14848) ) ;
NAND2   gate14100  (.A(II14839), .B(II14847), .Z(II14849) ) ;
NAND2   gate14101  (.A(II14848), .B(II14849), .Z(II14838) ) ;
NAND2   gate14102  (.A(WX4706), .B(WX4770), .Z(II14855) ) ;
NAND2   gate14103  (.A(WX4706), .B(II14855), .Z(II14856) ) ;
NAND2   gate14104  (.A(WX4770), .B(II14855), .Z(II14857) ) ;
NAND2   gate14105  (.A(II14856), .B(II14857), .Z(II14854) ) ;
NAND2   gate14106  (.A(II14838), .B(II14854), .Z(II14862) ) ;
NAND2   gate14107  (.A(II14838), .B(II14862), .Z(II14863) ) ;
NAND2   gate14108  (.A(II14854), .B(II14862), .Z(II14864) ) ;
NAND2   gate14109  (.A(WX4881), .B(WX4580), .Z(II14871) ) ;
NAND2   gate14110  (.A(WX4881), .B(II14871), .Z(II14872) ) ;
NAND2   gate14111  (.A(WX4580), .B(II14871), .Z(II14873) ) ;
NAND2   gate14112  (.A(II14872), .B(II14873), .Z(II14870) ) ;
NAND2   gate14113  (.A(WX4644), .B(II14870), .Z(II14878) ) ;
NAND2   gate14114  (.A(WX4644), .B(II14878), .Z(II14879) ) ;
NAND2   gate14115  (.A(II14870), .B(II14878), .Z(II14880) ) ;
NAND2   gate14116  (.A(II14879), .B(II14880), .Z(II14869) ) ;
NAND2   gate14117  (.A(WX4708), .B(WX4772), .Z(II14886) ) ;
NAND2   gate14118  (.A(WX4708), .B(II14886), .Z(II14887) ) ;
NAND2   gate14119  (.A(WX4772), .B(II14886), .Z(II14888) ) ;
NAND2   gate14120  (.A(II14887), .B(II14888), .Z(II14885) ) ;
NAND2   gate14121  (.A(II14869), .B(II14885), .Z(II14893) ) ;
NAND2   gate14122  (.A(II14869), .B(II14893), .Z(II14894) ) ;
NAND2   gate14123  (.A(II14885), .B(II14893), .Z(II14895) ) ;
NAND2   gate14124  (.A(WX4881), .B(WX4582), .Z(II14902) ) ;
NAND2   gate14125  (.A(WX4881), .B(II14902), .Z(II14903) ) ;
NAND2   gate14126  (.A(WX4582), .B(II14902), .Z(II14904) ) ;
NAND2   gate14127  (.A(II14903), .B(II14904), .Z(II14901) ) ;
NAND2   gate14128  (.A(WX4646), .B(II14901), .Z(II14909) ) ;
NAND2   gate14129  (.A(WX4646), .B(II14909), .Z(II14910) ) ;
NAND2   gate14130  (.A(II14901), .B(II14909), .Z(II14911) ) ;
NAND2   gate14131  (.A(II14910), .B(II14911), .Z(II14900) ) ;
NAND2   gate14132  (.A(WX4710), .B(WX4774), .Z(II14917) ) ;
NAND2   gate14133  (.A(WX4710), .B(II14917), .Z(II14918) ) ;
NAND2   gate14134  (.A(WX4774), .B(II14917), .Z(II14919) ) ;
NAND2   gate14135  (.A(II14918), .B(II14919), .Z(II14916) ) ;
NAND2   gate14136  (.A(II14900), .B(II14916), .Z(II14924) ) ;
NAND2   gate14137  (.A(II14900), .B(II14924), .Z(II14925) ) ;
NAND2   gate14138  (.A(II14916), .B(II14924), .Z(II14926) ) ;
NAND2   gate14139  (.A(WX4881), .B(WX4584), .Z(II14933) ) ;
NAND2   gate14140  (.A(WX4881), .B(II14933), .Z(II14934) ) ;
NAND2   gate14141  (.A(WX4584), .B(II14933), .Z(II14935) ) ;
NAND2   gate14142  (.A(II14934), .B(II14935), .Z(II14932) ) ;
NAND2   gate14143  (.A(WX4648), .B(II14932), .Z(II14940) ) ;
NAND2   gate14144  (.A(WX4648), .B(II14940), .Z(II14941) ) ;
NAND2   gate14145  (.A(II14932), .B(II14940), .Z(II14942) ) ;
NAND2   gate14146  (.A(II14941), .B(II14942), .Z(II14931) ) ;
NAND2   gate14147  (.A(WX4712), .B(WX4776), .Z(II14948) ) ;
NAND2   gate14148  (.A(WX4712), .B(II14948), .Z(II14949) ) ;
NAND2   gate14149  (.A(WX4776), .B(II14948), .Z(II14950) ) ;
NAND2   gate14150  (.A(II14949), .B(II14950), .Z(II14947) ) ;
NAND2   gate14151  (.A(II14931), .B(II14947), .Z(II14955) ) ;
NAND2   gate14152  (.A(II14931), .B(II14955), .Z(II14956) ) ;
NAND2   gate14153  (.A(II14947), .B(II14955), .Z(II14957) ) ;
NAND2   gate14154  (.A(WX4881), .B(WX4586), .Z(II14964) ) ;
NAND2   gate14155  (.A(WX4881), .B(II14964), .Z(II14965) ) ;
NAND2   gate14156  (.A(WX4586), .B(II14964), .Z(II14966) ) ;
NAND2   gate14157  (.A(II14965), .B(II14966), .Z(II14963) ) ;
NAND2   gate14158  (.A(WX4650), .B(II14963), .Z(II14971) ) ;
NAND2   gate14159  (.A(WX4650), .B(II14971), .Z(II14972) ) ;
NAND2   gate14160  (.A(II14963), .B(II14971), .Z(II14973) ) ;
NAND2   gate14161  (.A(II14972), .B(II14973), .Z(II14962) ) ;
NAND2   gate14162  (.A(WX4714), .B(WX4778), .Z(II14979) ) ;
NAND2   gate14163  (.A(WX4714), .B(II14979), .Z(II14980) ) ;
NAND2   gate14164  (.A(WX4778), .B(II14979), .Z(II14981) ) ;
NAND2   gate14165  (.A(II14980), .B(II14981), .Z(II14978) ) ;
NAND2   gate14166  (.A(II14962), .B(II14978), .Z(II14986) ) ;
NAND2   gate14167  (.A(II14962), .B(II14986), .Z(II14987) ) ;
NAND2   gate14168  (.A(II14978), .B(II14986), .Z(II14988) ) ;
NAND2   gate14169  (.A(WX4459), .B(WX4364), .Z(II15067) ) ;
NAND2   gate14170  (.A(WX4459), .B(II15067), .Z(II15068) ) ;
NAND2   gate14171  (.A(WX4364), .B(II15067), .Z(II15069) ) ;
NAND2   gate14172  (.A(WX4460), .B(WX4366), .Z(II15080) ) ;
NAND2   gate14173  (.A(WX4460), .B(II15080), .Z(II15081) ) ;
NAND2   gate14174  (.A(WX4366), .B(II15080), .Z(II15082) ) ;
NAND2   gate14175  (.A(WX4461), .B(WX4368), .Z(II15093) ) ;
NAND2   gate14176  (.A(WX4461), .B(II15093), .Z(II15094) ) ;
NAND2   gate14177  (.A(WX4368), .B(II15093), .Z(II15095) ) ;
NAND2   gate14178  (.A(WX4462), .B(WX4370), .Z(II15106) ) ;
NAND2   gate14179  (.A(WX4462), .B(II15106), .Z(II15107) ) ;
NAND2   gate14180  (.A(WX4370), .B(II15106), .Z(II15108) ) ;
NAND2   gate14181  (.A(WX4463), .B(WX4372), .Z(II15119) ) ;
NAND2   gate14182  (.A(WX4463), .B(II15119), .Z(II15120) ) ;
NAND2   gate14183  (.A(WX4372), .B(II15119), .Z(II15121) ) ;
NAND2   gate14184  (.A(WX4464), .B(WX4374), .Z(II15132) ) ;
NAND2   gate14185  (.A(WX4464), .B(II15132), .Z(II15133) ) ;
NAND2   gate14186  (.A(WX4374), .B(II15132), .Z(II15134) ) ;
NAND2   gate14187  (.A(WX4465), .B(WX4376), .Z(II15145) ) ;
NAND2   gate14188  (.A(WX4465), .B(II15145), .Z(II15146) ) ;
NAND2   gate14189  (.A(WX4376), .B(II15145), .Z(II15147) ) ;
NAND2   gate14190  (.A(WX4466), .B(WX4378), .Z(II15158) ) ;
NAND2   gate14191  (.A(WX4466), .B(II15158), .Z(II15159) ) ;
NAND2   gate14192  (.A(WX4378), .B(II15158), .Z(II15160) ) ;
NAND2   gate14193  (.A(WX4467), .B(WX4380), .Z(II15171) ) ;
NAND2   gate14194  (.A(WX4467), .B(II15171), .Z(II15172) ) ;
NAND2   gate14195  (.A(WX4380), .B(II15171), .Z(II15173) ) ;
NAND2   gate14196  (.A(WX4468), .B(WX4382), .Z(II15184) ) ;
NAND2   gate14197  (.A(WX4468), .B(II15184), .Z(II15185) ) ;
NAND2   gate14198  (.A(WX4382), .B(II15184), .Z(II15186) ) ;
NAND2   gate14199  (.A(WX4469), .B(WX4384), .Z(II15197) ) ;
NAND2   gate14200  (.A(WX4469), .B(II15197), .Z(II15198) ) ;
NAND2   gate14201  (.A(WX4384), .B(II15197), .Z(II15199) ) ;
NAND2   gate14202  (.A(WX4470), .B(WX4386), .Z(II15210) ) ;
NAND2   gate14203  (.A(WX4470), .B(II15210), .Z(II15211) ) ;
NAND2   gate14204  (.A(WX4386), .B(II15210), .Z(II15212) ) ;
NAND2   gate14205  (.A(WX4471), .B(WX4388), .Z(II15223) ) ;
NAND2   gate14206  (.A(WX4471), .B(II15223), .Z(II15224) ) ;
NAND2   gate14207  (.A(WX4388), .B(II15223), .Z(II15225) ) ;
NAND2   gate14208  (.A(WX4472), .B(WX4390), .Z(II15236) ) ;
NAND2   gate14209  (.A(WX4472), .B(II15236), .Z(II15237) ) ;
NAND2   gate14210  (.A(WX4390), .B(II15236), .Z(II15238) ) ;
NAND2   gate14211  (.A(WX4473), .B(WX4392), .Z(II15249) ) ;
NAND2   gate14212  (.A(WX4473), .B(II15249), .Z(II15250) ) ;
NAND2   gate14213  (.A(WX4392), .B(II15249), .Z(II15251) ) ;
NAND2   gate14214  (.A(WX4474), .B(WX4394), .Z(II15262) ) ;
NAND2   gate14215  (.A(WX4474), .B(II15262), .Z(II15263) ) ;
NAND2   gate14216  (.A(WX4394), .B(II15262), .Z(II15264) ) ;
NAND2   gate14217  (.A(WX4475), .B(WX4396), .Z(II15275) ) ;
NAND2   gate14218  (.A(WX4475), .B(II15275), .Z(II15276) ) ;
NAND2   gate14219  (.A(WX4396), .B(II15275), .Z(II15277) ) ;
NAND2   gate14220  (.A(WX4476), .B(WX4398), .Z(II15288) ) ;
NAND2   gate14221  (.A(WX4476), .B(II15288), .Z(II15289) ) ;
NAND2   gate14222  (.A(WX4398), .B(II15288), .Z(II15290) ) ;
NAND2   gate14223  (.A(WX4477), .B(WX4400), .Z(II15301) ) ;
NAND2   gate14224  (.A(WX4477), .B(II15301), .Z(II15302) ) ;
NAND2   gate14225  (.A(WX4400), .B(II15301), .Z(II15303) ) ;
NAND2   gate14226  (.A(WX4478), .B(WX4402), .Z(II15314) ) ;
NAND2   gate14227  (.A(WX4478), .B(II15314), .Z(II15315) ) ;
NAND2   gate14228  (.A(WX4402), .B(II15314), .Z(II15316) ) ;
NAND2   gate14229  (.A(WX4479), .B(WX4404), .Z(II15327) ) ;
NAND2   gate14230  (.A(WX4479), .B(II15327), .Z(II15328) ) ;
NAND2   gate14231  (.A(WX4404), .B(II15327), .Z(II15329) ) ;
NAND2   gate14232  (.A(WX4480), .B(WX4406), .Z(II15340) ) ;
NAND2   gate14233  (.A(WX4480), .B(II15340), .Z(II15341) ) ;
NAND2   gate14234  (.A(WX4406), .B(II15340), .Z(II15342) ) ;
NAND2   gate14235  (.A(WX4481), .B(WX4408), .Z(II15353) ) ;
NAND2   gate14236  (.A(WX4481), .B(II15353), .Z(II15354) ) ;
NAND2   gate14237  (.A(WX4408), .B(II15353), .Z(II15355) ) ;
NAND2   gate14238  (.A(WX4482), .B(WX4410), .Z(II15366) ) ;
NAND2   gate14239  (.A(WX4482), .B(II15366), .Z(II15367) ) ;
NAND2   gate14240  (.A(WX4410), .B(II15366), .Z(II15368) ) ;
NAND2   gate14241  (.A(WX4483), .B(WX4412), .Z(II15379) ) ;
NAND2   gate14242  (.A(WX4483), .B(II15379), .Z(II15380) ) ;
NAND2   gate14243  (.A(WX4412), .B(II15379), .Z(II15381) ) ;
NAND2   gate14244  (.A(WX4484), .B(WX4414), .Z(II15392) ) ;
NAND2   gate14245  (.A(WX4484), .B(II15392), .Z(II15393) ) ;
NAND2   gate14246  (.A(WX4414), .B(II15392), .Z(II15394) ) ;
NAND2   gate14247  (.A(WX4485), .B(WX4416), .Z(II15405) ) ;
NAND2   gate14248  (.A(WX4485), .B(II15405), .Z(II15406) ) ;
NAND2   gate14249  (.A(WX4416), .B(II15405), .Z(II15407) ) ;
NAND2   gate14250  (.A(WX4486), .B(WX4418), .Z(II15418) ) ;
NAND2   gate14251  (.A(WX4486), .B(II15418), .Z(II15419) ) ;
NAND2   gate14252  (.A(WX4418), .B(II15418), .Z(II15420) ) ;
NAND2   gate14253  (.A(WX4487), .B(WX4420), .Z(II15431) ) ;
NAND2   gate14254  (.A(WX4487), .B(II15431), .Z(II15432) ) ;
NAND2   gate14255  (.A(WX4420), .B(II15431), .Z(II15433) ) ;
NAND2   gate14256  (.A(WX4488), .B(WX4422), .Z(II15444) ) ;
NAND2   gate14257  (.A(WX4488), .B(II15444), .Z(II15445) ) ;
NAND2   gate14258  (.A(WX4422), .B(II15444), .Z(II15446) ) ;
NAND2   gate14259  (.A(WX4489), .B(WX4424), .Z(II15457) ) ;
NAND2   gate14260  (.A(WX4489), .B(II15457), .Z(II15458) ) ;
NAND2   gate14261  (.A(WX4424), .B(II15457), .Z(II15459) ) ;
NAND2   gate14262  (.A(WX4490), .B(WX4426), .Z(II15470) ) ;
NAND2   gate14263  (.A(WX4490), .B(II15470), .Z(II15471) ) ;
NAND2   gate14264  (.A(WX4426), .B(II15470), .Z(II15472) ) ;
NAND2   gate14265  (.A(WX4506), .B(CRC_OUT_6_31), .Z(II15485) ) ;
NAND2   gate14266  (.A(WX4506), .B(II15485), .Z(II15486) ) ;
NAND2   gate14267  (.A(CRC_OUT_6_31), .B(II15485), .Z(II15487) ) ;
NAND2   gate14268  (.A(II15486), .B(II15487), .Z(II15484) ) ;
NAND2   gate14269  (.A(CRC_OUT_6_15), .B(II15484), .Z(II15492) ) ;
NAND2   gate14270  (.A(CRC_OUT_6_15), .B(II15492), .Z(II15493) ) ;
NAND2   gate14271  (.A(II15484), .B(II15492), .Z(II15494) ) ;
NAND2   gate14272  (.A(WX4511), .B(CRC_OUT_6_31), .Z(II15500) ) ;
NAND2   gate14273  (.A(WX4511), .B(II15500), .Z(II15501) ) ;
NAND2   gate14274  (.A(CRC_OUT_6_31), .B(II15500), .Z(II15502) ) ;
NAND2   gate14275  (.A(II15501), .B(II15502), .Z(II15499) ) ;
NAND2   gate14276  (.A(CRC_OUT_6_10), .B(II15499), .Z(II15507) ) ;
NAND2   gate14277  (.A(CRC_OUT_6_10), .B(II15507), .Z(II15508) ) ;
NAND2   gate14278  (.A(II15499), .B(II15507), .Z(II15509) ) ;
NAND2   gate14279  (.A(WX4518), .B(CRC_OUT_6_31), .Z(II15515) ) ;
NAND2   gate14280  (.A(WX4518), .B(II15515), .Z(II15516) ) ;
NAND2   gate14281  (.A(CRC_OUT_6_31), .B(II15515), .Z(II15517) ) ;
NAND2   gate14282  (.A(II15516), .B(II15517), .Z(II15514) ) ;
NAND2   gate14283  (.A(CRC_OUT_6_3), .B(II15514), .Z(II15522) ) ;
NAND2   gate14284  (.A(CRC_OUT_6_3), .B(II15522), .Z(II15523) ) ;
NAND2   gate14285  (.A(II15514), .B(II15522), .Z(II15524) ) ;
NAND2   gate14286  (.A(WX4522), .B(CRC_OUT_6_31), .Z(II15529) ) ;
NAND2   gate14287  (.A(WX4522), .B(II15529), .Z(II15530) ) ;
NAND2   gate14288  (.A(CRC_OUT_6_31), .B(II15529), .Z(II15531) ) ;
NAND2   gate14289  (.A(WX4491), .B(CRC_OUT_6_30), .Z(II15536) ) ;
NAND2   gate14290  (.A(WX4491), .B(II15536), .Z(II15537) ) ;
NAND2   gate14291  (.A(CRC_OUT_6_30), .B(II15536), .Z(II15538) ) ;
NAND2   gate14292  (.A(WX4492), .B(CRC_OUT_6_29), .Z(II15543) ) ;
NAND2   gate14293  (.A(WX4492), .B(II15543), .Z(II15544) ) ;
NAND2   gate14294  (.A(CRC_OUT_6_29), .B(II15543), .Z(II15545) ) ;
NAND2   gate14295  (.A(WX4493), .B(CRC_OUT_6_28), .Z(II15550) ) ;
NAND2   gate14296  (.A(WX4493), .B(II15550), .Z(II15551) ) ;
NAND2   gate14297  (.A(CRC_OUT_6_28), .B(II15550), .Z(II15552) ) ;
NAND2   gate14298  (.A(WX4494), .B(CRC_OUT_6_27), .Z(II15557) ) ;
NAND2   gate14299  (.A(WX4494), .B(II15557), .Z(II15558) ) ;
NAND2   gate14300  (.A(CRC_OUT_6_27), .B(II15557), .Z(II15559) ) ;
NAND2   gate14301  (.A(WX4495), .B(CRC_OUT_6_26), .Z(II15564) ) ;
NAND2   gate14302  (.A(WX4495), .B(II15564), .Z(II15565) ) ;
NAND2   gate14303  (.A(CRC_OUT_6_26), .B(II15564), .Z(II15566) ) ;
NAND2   gate14304  (.A(WX4496), .B(CRC_OUT_6_25), .Z(II15571) ) ;
NAND2   gate14305  (.A(WX4496), .B(II15571), .Z(II15572) ) ;
NAND2   gate14306  (.A(CRC_OUT_6_25), .B(II15571), .Z(II15573) ) ;
NAND2   gate14307  (.A(WX4497), .B(CRC_OUT_6_24), .Z(II15578) ) ;
NAND2   gate14308  (.A(WX4497), .B(II15578), .Z(II15579) ) ;
NAND2   gate14309  (.A(CRC_OUT_6_24), .B(II15578), .Z(II15580) ) ;
NAND2   gate14310  (.A(WX4498), .B(CRC_OUT_6_23), .Z(II15585) ) ;
NAND2   gate14311  (.A(WX4498), .B(II15585), .Z(II15586) ) ;
NAND2   gate14312  (.A(CRC_OUT_6_23), .B(II15585), .Z(II15587) ) ;
NAND2   gate14313  (.A(WX4499), .B(CRC_OUT_6_22), .Z(II15592) ) ;
NAND2   gate14314  (.A(WX4499), .B(II15592), .Z(II15593) ) ;
NAND2   gate14315  (.A(CRC_OUT_6_22), .B(II15592), .Z(II15594) ) ;
NAND2   gate14316  (.A(WX4500), .B(CRC_OUT_6_21), .Z(II15599) ) ;
NAND2   gate14317  (.A(WX4500), .B(II15599), .Z(II15600) ) ;
NAND2   gate14318  (.A(CRC_OUT_6_21), .B(II15599), .Z(II15601) ) ;
NAND2   gate14319  (.A(WX4501), .B(CRC_OUT_6_20), .Z(II15606) ) ;
NAND2   gate14320  (.A(WX4501), .B(II15606), .Z(II15607) ) ;
NAND2   gate14321  (.A(CRC_OUT_6_20), .B(II15606), .Z(II15608) ) ;
NAND2   gate14322  (.A(WX4502), .B(CRC_OUT_6_19), .Z(II15613) ) ;
NAND2   gate14323  (.A(WX4502), .B(II15613), .Z(II15614) ) ;
NAND2   gate14324  (.A(CRC_OUT_6_19), .B(II15613), .Z(II15615) ) ;
NAND2   gate14325  (.A(WX4503), .B(CRC_OUT_6_18), .Z(II15620) ) ;
NAND2   gate14326  (.A(WX4503), .B(II15620), .Z(II15621) ) ;
NAND2   gate14327  (.A(CRC_OUT_6_18), .B(II15620), .Z(II15622) ) ;
NAND2   gate14328  (.A(WX4504), .B(CRC_OUT_6_17), .Z(II15627) ) ;
NAND2   gate14329  (.A(WX4504), .B(II15627), .Z(II15628) ) ;
NAND2   gate14330  (.A(CRC_OUT_6_17), .B(II15627), .Z(II15629) ) ;
NAND2   gate14331  (.A(WX4505), .B(CRC_OUT_6_16), .Z(II15634) ) ;
NAND2   gate14332  (.A(WX4505), .B(II15634), .Z(II15635) ) ;
NAND2   gate14333  (.A(CRC_OUT_6_16), .B(II15634), .Z(II15636) ) ;
NAND2   gate14334  (.A(WX4507), .B(CRC_OUT_6_14), .Z(II15641) ) ;
NAND2   gate14335  (.A(WX4507), .B(II15641), .Z(II15642) ) ;
NAND2   gate14336  (.A(CRC_OUT_6_14), .B(II15641), .Z(II15643) ) ;
NAND2   gate14337  (.A(WX4508), .B(CRC_OUT_6_13), .Z(II15648) ) ;
NAND2   gate14338  (.A(WX4508), .B(II15648), .Z(II15649) ) ;
NAND2   gate14339  (.A(CRC_OUT_6_13), .B(II15648), .Z(II15650) ) ;
NAND2   gate14340  (.A(WX4509), .B(CRC_OUT_6_12), .Z(II15655) ) ;
NAND2   gate14341  (.A(WX4509), .B(II15655), .Z(II15656) ) ;
NAND2   gate14342  (.A(CRC_OUT_6_12), .B(II15655), .Z(II15657) ) ;
NAND2   gate14343  (.A(WX4510), .B(CRC_OUT_6_11), .Z(II15662) ) ;
NAND2   gate14344  (.A(WX4510), .B(II15662), .Z(II15663) ) ;
NAND2   gate14345  (.A(CRC_OUT_6_11), .B(II15662), .Z(II15664) ) ;
NAND2   gate14346  (.A(WX4512), .B(CRC_OUT_6_9), .Z(II15669) ) ;
NAND2   gate14347  (.A(WX4512), .B(II15669), .Z(II15670) ) ;
NAND2   gate14348  (.A(CRC_OUT_6_9), .B(II15669), .Z(II15671) ) ;
NAND2   gate14349  (.A(WX4513), .B(CRC_OUT_6_8), .Z(II15676) ) ;
NAND2   gate14350  (.A(WX4513), .B(II15676), .Z(II15677) ) ;
NAND2   gate14351  (.A(CRC_OUT_6_8), .B(II15676), .Z(II15678) ) ;
NAND2   gate14352  (.A(WX4514), .B(CRC_OUT_6_7), .Z(II15683) ) ;
NAND2   gate14353  (.A(WX4514), .B(II15683), .Z(II15684) ) ;
NAND2   gate14354  (.A(CRC_OUT_6_7), .B(II15683), .Z(II15685) ) ;
NAND2   gate14355  (.A(WX4515), .B(CRC_OUT_6_6), .Z(II15690) ) ;
NAND2   gate14356  (.A(WX4515), .B(II15690), .Z(II15691) ) ;
NAND2   gate14357  (.A(CRC_OUT_6_6), .B(II15690), .Z(II15692) ) ;
NAND2   gate14358  (.A(WX4516), .B(CRC_OUT_6_5), .Z(II15697) ) ;
NAND2   gate14359  (.A(WX4516), .B(II15697), .Z(II15698) ) ;
NAND2   gate14360  (.A(CRC_OUT_6_5), .B(II15697), .Z(II15699) ) ;
NAND2   gate14361  (.A(WX4517), .B(CRC_OUT_6_4), .Z(II15704) ) ;
NAND2   gate14362  (.A(WX4517), .B(II15704), .Z(II15705) ) ;
NAND2   gate14363  (.A(CRC_OUT_6_4), .B(II15704), .Z(II15706) ) ;
NAND2   gate14364  (.A(WX4519), .B(CRC_OUT_6_2), .Z(II15711) ) ;
NAND2   gate14365  (.A(WX4519), .B(II15711), .Z(II15712) ) ;
NAND2   gate14366  (.A(CRC_OUT_6_2), .B(II15711), .Z(II15713) ) ;
NAND2   gate14367  (.A(WX4520), .B(CRC_OUT_6_1), .Z(II15718) ) ;
NAND2   gate14368  (.A(WX4520), .B(II15718), .Z(II15719) ) ;
NAND2   gate14369  (.A(CRC_OUT_6_1), .B(II15718), .Z(II15720) ) ;
NAND2   gate14370  (.A(WX4521), .B(CRC_OUT_6_0), .Z(II15725) ) ;
NAND2   gate14371  (.A(WX4521), .B(II15725), .Z(II15726) ) ;
NAND2   gate14372  (.A(CRC_OUT_6_0), .B(II15725), .Z(II15727) ) ;
NAND2   gate14373  (.A(WX6173), .B(WX5817), .Z(II18008) ) ;
NAND2   gate14374  (.A(WX6173), .B(II18008), .Z(II18009) ) ;
NAND2   gate14375  (.A(WX5817), .B(II18008), .Z(II18010) ) ;
NAND2   gate14376  (.A(II18009), .B(II18010), .Z(II18007) ) ;
NAND2   gate14377  (.A(WX5881), .B(II18007), .Z(II18015) ) ;
NAND2   gate14378  (.A(WX5881), .B(II18015), .Z(II18016) ) ;
NAND2   gate14379  (.A(II18007), .B(II18015), .Z(II18017) ) ;
NAND2   gate14380  (.A(II18016), .B(II18017), .Z(II18006) ) ;
NAND2   gate14381  (.A(WX5945), .B(WX6009), .Z(II18023) ) ;
NAND2   gate14382  (.A(WX5945), .B(II18023), .Z(II18024) ) ;
NAND2   gate14383  (.A(WX6009), .B(II18023), .Z(II18025) ) ;
NAND2   gate14384  (.A(II18024), .B(II18025), .Z(II18022) ) ;
NAND2   gate14385  (.A(II18006), .B(II18022), .Z(II18030) ) ;
NAND2   gate14386  (.A(II18006), .B(II18030), .Z(II18031) ) ;
NAND2   gate14387  (.A(II18022), .B(II18030), .Z(II18032) ) ;
NAND2   gate14388  (.A(WX6173), .B(WX5819), .Z(II18039) ) ;
NAND2   gate14389  (.A(WX6173), .B(II18039), .Z(II18040) ) ;
NAND2   gate14390  (.A(WX5819), .B(II18039), .Z(II18041) ) ;
NAND2   gate14391  (.A(II18040), .B(II18041), .Z(II18038) ) ;
NAND2   gate14392  (.A(WX5883), .B(II18038), .Z(II18046) ) ;
NAND2   gate14393  (.A(WX5883), .B(II18046), .Z(II18047) ) ;
NAND2   gate14394  (.A(II18038), .B(II18046), .Z(II18048) ) ;
NAND2   gate14395  (.A(II18047), .B(II18048), .Z(II18037) ) ;
NAND2   gate14396  (.A(WX5947), .B(WX6011), .Z(II18054) ) ;
NAND2   gate14397  (.A(WX5947), .B(II18054), .Z(II18055) ) ;
NAND2   gate14398  (.A(WX6011), .B(II18054), .Z(II18056) ) ;
NAND2   gate14399  (.A(II18055), .B(II18056), .Z(II18053) ) ;
NAND2   gate14400  (.A(II18037), .B(II18053), .Z(II18061) ) ;
NAND2   gate14401  (.A(II18037), .B(II18061), .Z(II18062) ) ;
NAND2   gate14402  (.A(II18053), .B(II18061), .Z(II18063) ) ;
NAND2   gate14403  (.A(WX6173), .B(WX5821), .Z(II18070) ) ;
NAND2   gate14404  (.A(WX6173), .B(II18070), .Z(II18071) ) ;
NAND2   gate14405  (.A(WX5821), .B(II18070), .Z(II18072) ) ;
NAND2   gate14406  (.A(II18071), .B(II18072), .Z(II18069) ) ;
NAND2   gate14407  (.A(WX5885), .B(II18069), .Z(II18077) ) ;
NAND2   gate14408  (.A(WX5885), .B(II18077), .Z(II18078) ) ;
NAND2   gate14409  (.A(II18069), .B(II18077), .Z(II18079) ) ;
NAND2   gate14410  (.A(II18078), .B(II18079), .Z(II18068) ) ;
NAND2   gate14411  (.A(WX5949), .B(WX6013), .Z(II18085) ) ;
NAND2   gate14412  (.A(WX5949), .B(II18085), .Z(II18086) ) ;
NAND2   gate14413  (.A(WX6013), .B(II18085), .Z(II18087) ) ;
NAND2   gate14414  (.A(II18086), .B(II18087), .Z(II18084) ) ;
NAND2   gate14415  (.A(II18068), .B(II18084), .Z(II18092) ) ;
NAND2   gate14416  (.A(II18068), .B(II18092), .Z(II18093) ) ;
NAND2   gate14417  (.A(II18084), .B(II18092), .Z(II18094) ) ;
NAND2   gate14418  (.A(WX6173), .B(WX5823), .Z(II18101) ) ;
NAND2   gate14419  (.A(WX6173), .B(II18101), .Z(II18102) ) ;
NAND2   gate14420  (.A(WX5823), .B(II18101), .Z(II18103) ) ;
NAND2   gate14421  (.A(II18102), .B(II18103), .Z(II18100) ) ;
NAND2   gate14422  (.A(WX5887), .B(II18100), .Z(II18108) ) ;
NAND2   gate14423  (.A(WX5887), .B(II18108), .Z(II18109) ) ;
NAND2   gate14424  (.A(II18100), .B(II18108), .Z(II18110) ) ;
NAND2   gate14425  (.A(II18109), .B(II18110), .Z(II18099) ) ;
NAND2   gate14426  (.A(WX5951), .B(WX6015), .Z(II18116) ) ;
NAND2   gate14427  (.A(WX5951), .B(II18116), .Z(II18117) ) ;
NAND2   gate14428  (.A(WX6015), .B(II18116), .Z(II18118) ) ;
NAND2   gate14429  (.A(II18117), .B(II18118), .Z(II18115) ) ;
NAND2   gate14430  (.A(II18099), .B(II18115), .Z(II18123) ) ;
NAND2   gate14431  (.A(II18099), .B(II18123), .Z(II18124) ) ;
NAND2   gate14432  (.A(II18115), .B(II18123), .Z(II18125) ) ;
NAND2   gate14433  (.A(WX6173), .B(WX5825), .Z(II18132) ) ;
NAND2   gate14434  (.A(WX6173), .B(II18132), .Z(II18133) ) ;
NAND2   gate14435  (.A(WX5825), .B(II18132), .Z(II18134) ) ;
NAND2   gate14436  (.A(II18133), .B(II18134), .Z(II18131) ) ;
NAND2   gate14437  (.A(WX5889), .B(II18131), .Z(II18139) ) ;
NAND2   gate14438  (.A(WX5889), .B(II18139), .Z(II18140) ) ;
NAND2   gate14439  (.A(II18131), .B(II18139), .Z(II18141) ) ;
NAND2   gate14440  (.A(II18140), .B(II18141), .Z(II18130) ) ;
NAND2   gate14441  (.A(WX5953), .B(WX6017), .Z(II18147) ) ;
NAND2   gate14442  (.A(WX5953), .B(II18147), .Z(II18148) ) ;
NAND2   gate14443  (.A(WX6017), .B(II18147), .Z(II18149) ) ;
NAND2   gate14444  (.A(II18148), .B(II18149), .Z(II18146) ) ;
NAND2   gate14445  (.A(II18130), .B(II18146), .Z(II18154) ) ;
NAND2   gate14446  (.A(II18130), .B(II18154), .Z(II18155) ) ;
NAND2   gate14447  (.A(II18146), .B(II18154), .Z(II18156) ) ;
NAND2   gate14448  (.A(WX6173), .B(WX5827), .Z(II18163) ) ;
NAND2   gate14449  (.A(WX6173), .B(II18163), .Z(II18164) ) ;
NAND2   gate14450  (.A(WX5827), .B(II18163), .Z(II18165) ) ;
NAND2   gate14451  (.A(II18164), .B(II18165), .Z(II18162) ) ;
NAND2   gate14452  (.A(WX5891), .B(II18162), .Z(II18170) ) ;
NAND2   gate14453  (.A(WX5891), .B(II18170), .Z(II18171) ) ;
NAND2   gate14454  (.A(II18162), .B(II18170), .Z(II18172) ) ;
NAND2   gate14455  (.A(II18171), .B(II18172), .Z(II18161) ) ;
NAND2   gate14456  (.A(WX5955), .B(WX6019), .Z(II18178) ) ;
NAND2   gate14457  (.A(WX5955), .B(II18178), .Z(II18179) ) ;
NAND2   gate14458  (.A(WX6019), .B(II18178), .Z(II18180) ) ;
NAND2   gate14459  (.A(II18179), .B(II18180), .Z(II18177) ) ;
NAND2   gate14460  (.A(II18161), .B(II18177), .Z(II18185) ) ;
NAND2   gate14461  (.A(II18161), .B(II18185), .Z(II18186) ) ;
NAND2   gate14462  (.A(II18177), .B(II18185), .Z(II18187) ) ;
NAND2   gate14463  (.A(WX6173), .B(WX5829), .Z(II18194) ) ;
NAND2   gate14464  (.A(WX6173), .B(II18194), .Z(II18195) ) ;
NAND2   gate14465  (.A(WX5829), .B(II18194), .Z(II18196) ) ;
NAND2   gate14466  (.A(II18195), .B(II18196), .Z(II18193) ) ;
NAND2   gate14467  (.A(WX5893), .B(II18193), .Z(II18201) ) ;
NAND2   gate14468  (.A(WX5893), .B(II18201), .Z(II18202) ) ;
NAND2   gate14469  (.A(II18193), .B(II18201), .Z(II18203) ) ;
NAND2   gate14470  (.A(II18202), .B(II18203), .Z(II18192) ) ;
NAND2   gate14471  (.A(WX5957), .B(WX6021), .Z(II18209) ) ;
NAND2   gate14472  (.A(WX5957), .B(II18209), .Z(II18210) ) ;
NAND2   gate14473  (.A(WX6021), .B(II18209), .Z(II18211) ) ;
NAND2   gate14474  (.A(II18210), .B(II18211), .Z(II18208) ) ;
NAND2   gate14475  (.A(II18192), .B(II18208), .Z(II18216) ) ;
NAND2   gate14476  (.A(II18192), .B(II18216), .Z(II18217) ) ;
NAND2   gate14477  (.A(II18208), .B(II18216), .Z(II18218) ) ;
NAND2   gate14478  (.A(WX6173), .B(WX5831), .Z(II18225) ) ;
NAND2   gate14479  (.A(WX6173), .B(II18225), .Z(II18226) ) ;
NAND2   gate14480  (.A(WX5831), .B(II18225), .Z(II18227) ) ;
NAND2   gate14481  (.A(II18226), .B(II18227), .Z(II18224) ) ;
NAND2   gate14482  (.A(WX5895), .B(II18224), .Z(II18232) ) ;
NAND2   gate14483  (.A(WX5895), .B(II18232), .Z(II18233) ) ;
NAND2   gate14484  (.A(II18224), .B(II18232), .Z(II18234) ) ;
NAND2   gate14485  (.A(II18233), .B(II18234), .Z(II18223) ) ;
NAND2   gate14486  (.A(WX5959), .B(WX6023), .Z(II18240) ) ;
NAND2   gate14487  (.A(WX5959), .B(II18240), .Z(II18241) ) ;
NAND2   gate14488  (.A(WX6023), .B(II18240), .Z(II18242) ) ;
NAND2   gate14489  (.A(II18241), .B(II18242), .Z(II18239) ) ;
NAND2   gate14490  (.A(II18223), .B(II18239), .Z(II18247) ) ;
NAND2   gate14491  (.A(II18223), .B(II18247), .Z(II18248) ) ;
NAND2   gate14492  (.A(II18239), .B(II18247), .Z(II18249) ) ;
NAND2   gate14493  (.A(WX6173), .B(WX5833), .Z(II18256) ) ;
NAND2   gate14494  (.A(WX6173), .B(II18256), .Z(II18257) ) ;
NAND2   gate14495  (.A(WX5833), .B(II18256), .Z(II18258) ) ;
NAND2   gate14496  (.A(II18257), .B(II18258), .Z(II18255) ) ;
NAND2   gate14497  (.A(WX5897), .B(II18255), .Z(II18263) ) ;
NAND2   gate14498  (.A(WX5897), .B(II18263), .Z(II18264) ) ;
NAND2   gate14499  (.A(II18255), .B(II18263), .Z(II18265) ) ;
NAND2   gate14500  (.A(II18264), .B(II18265), .Z(II18254) ) ;
NAND2   gate14501  (.A(WX5961), .B(WX6025), .Z(II18271) ) ;
NAND2   gate14502  (.A(WX5961), .B(II18271), .Z(II18272) ) ;
NAND2   gate14503  (.A(WX6025), .B(II18271), .Z(II18273) ) ;
NAND2   gate14504  (.A(II18272), .B(II18273), .Z(II18270) ) ;
NAND2   gate14505  (.A(II18254), .B(II18270), .Z(II18278) ) ;
NAND2   gate14506  (.A(II18254), .B(II18278), .Z(II18279) ) ;
NAND2   gate14507  (.A(II18270), .B(II18278), .Z(II18280) ) ;
NAND2   gate14508  (.A(WX6173), .B(WX5835), .Z(II18287) ) ;
NAND2   gate14509  (.A(WX6173), .B(II18287), .Z(II18288) ) ;
NAND2   gate14510  (.A(WX5835), .B(II18287), .Z(II18289) ) ;
NAND2   gate14511  (.A(II18288), .B(II18289), .Z(II18286) ) ;
NAND2   gate14512  (.A(WX5899), .B(II18286), .Z(II18294) ) ;
NAND2   gate14513  (.A(WX5899), .B(II18294), .Z(II18295) ) ;
NAND2   gate14514  (.A(II18286), .B(II18294), .Z(II18296) ) ;
NAND2   gate14515  (.A(II18295), .B(II18296), .Z(II18285) ) ;
NAND2   gate14516  (.A(WX5963), .B(WX6027), .Z(II18302) ) ;
NAND2   gate14517  (.A(WX5963), .B(II18302), .Z(II18303) ) ;
NAND2   gate14518  (.A(WX6027), .B(II18302), .Z(II18304) ) ;
NAND2   gate14519  (.A(II18303), .B(II18304), .Z(II18301) ) ;
NAND2   gate14520  (.A(II18285), .B(II18301), .Z(II18309) ) ;
NAND2   gate14521  (.A(II18285), .B(II18309), .Z(II18310) ) ;
NAND2   gate14522  (.A(II18301), .B(II18309), .Z(II18311) ) ;
NAND2   gate14523  (.A(WX6173), .B(WX5837), .Z(II18318) ) ;
NAND2   gate14524  (.A(WX6173), .B(II18318), .Z(II18319) ) ;
NAND2   gate14525  (.A(WX5837), .B(II18318), .Z(II18320) ) ;
NAND2   gate14526  (.A(II18319), .B(II18320), .Z(II18317) ) ;
NAND2   gate14527  (.A(WX5901), .B(II18317), .Z(II18325) ) ;
NAND2   gate14528  (.A(WX5901), .B(II18325), .Z(II18326) ) ;
NAND2   gate14529  (.A(II18317), .B(II18325), .Z(II18327) ) ;
NAND2   gate14530  (.A(II18326), .B(II18327), .Z(II18316) ) ;
NAND2   gate14531  (.A(WX5965), .B(WX6029), .Z(II18333) ) ;
NAND2   gate14532  (.A(WX5965), .B(II18333), .Z(II18334) ) ;
NAND2   gate14533  (.A(WX6029), .B(II18333), .Z(II18335) ) ;
NAND2   gate14534  (.A(II18334), .B(II18335), .Z(II18332) ) ;
NAND2   gate14535  (.A(II18316), .B(II18332), .Z(II18340) ) ;
NAND2   gate14536  (.A(II18316), .B(II18340), .Z(II18341) ) ;
NAND2   gate14537  (.A(II18332), .B(II18340), .Z(II18342) ) ;
NAND2   gate14538  (.A(WX6173), .B(WX5839), .Z(II18349) ) ;
NAND2   gate14539  (.A(WX6173), .B(II18349), .Z(II18350) ) ;
NAND2   gate14540  (.A(WX5839), .B(II18349), .Z(II18351) ) ;
NAND2   gate14541  (.A(II18350), .B(II18351), .Z(II18348) ) ;
NAND2   gate14542  (.A(WX5903), .B(II18348), .Z(II18356) ) ;
NAND2   gate14543  (.A(WX5903), .B(II18356), .Z(II18357) ) ;
NAND2   gate14544  (.A(II18348), .B(II18356), .Z(II18358) ) ;
NAND2   gate14545  (.A(II18357), .B(II18358), .Z(II18347) ) ;
NAND2   gate14546  (.A(WX5967), .B(WX6031), .Z(II18364) ) ;
NAND2   gate14547  (.A(WX5967), .B(II18364), .Z(II18365) ) ;
NAND2   gate14548  (.A(WX6031), .B(II18364), .Z(II18366) ) ;
NAND2   gate14549  (.A(II18365), .B(II18366), .Z(II18363) ) ;
NAND2   gate14550  (.A(II18347), .B(II18363), .Z(II18371) ) ;
NAND2   gate14551  (.A(II18347), .B(II18371), .Z(II18372) ) ;
NAND2   gate14552  (.A(II18363), .B(II18371), .Z(II18373) ) ;
NAND2   gate14553  (.A(WX6173), .B(WX5841), .Z(II18380) ) ;
NAND2   gate14554  (.A(WX6173), .B(II18380), .Z(II18381) ) ;
NAND2   gate14555  (.A(WX5841), .B(II18380), .Z(II18382) ) ;
NAND2   gate14556  (.A(II18381), .B(II18382), .Z(II18379) ) ;
NAND2   gate14557  (.A(WX5905), .B(II18379), .Z(II18387) ) ;
NAND2   gate14558  (.A(WX5905), .B(II18387), .Z(II18388) ) ;
NAND2   gate14559  (.A(II18379), .B(II18387), .Z(II18389) ) ;
NAND2   gate14560  (.A(II18388), .B(II18389), .Z(II18378) ) ;
NAND2   gate14561  (.A(WX5969), .B(WX6033), .Z(II18395) ) ;
NAND2   gate14562  (.A(WX5969), .B(II18395), .Z(II18396) ) ;
NAND2   gate14563  (.A(WX6033), .B(II18395), .Z(II18397) ) ;
NAND2   gate14564  (.A(II18396), .B(II18397), .Z(II18394) ) ;
NAND2   gate14565  (.A(II18378), .B(II18394), .Z(II18402) ) ;
NAND2   gate14566  (.A(II18378), .B(II18402), .Z(II18403) ) ;
NAND2   gate14567  (.A(II18394), .B(II18402), .Z(II18404) ) ;
NAND2   gate14568  (.A(WX6173), .B(WX5843), .Z(II18411) ) ;
NAND2   gate14569  (.A(WX6173), .B(II18411), .Z(II18412) ) ;
NAND2   gate14570  (.A(WX5843), .B(II18411), .Z(II18413) ) ;
NAND2   gate14571  (.A(II18412), .B(II18413), .Z(II18410) ) ;
NAND2   gate14572  (.A(WX5907), .B(II18410), .Z(II18418) ) ;
NAND2   gate14573  (.A(WX5907), .B(II18418), .Z(II18419) ) ;
NAND2   gate14574  (.A(II18410), .B(II18418), .Z(II18420) ) ;
NAND2   gate14575  (.A(II18419), .B(II18420), .Z(II18409) ) ;
NAND2   gate14576  (.A(WX5971), .B(WX6035), .Z(II18426) ) ;
NAND2   gate14577  (.A(WX5971), .B(II18426), .Z(II18427) ) ;
NAND2   gate14578  (.A(WX6035), .B(II18426), .Z(II18428) ) ;
NAND2   gate14579  (.A(II18427), .B(II18428), .Z(II18425) ) ;
NAND2   gate14580  (.A(II18409), .B(II18425), .Z(II18433) ) ;
NAND2   gate14581  (.A(II18409), .B(II18433), .Z(II18434) ) ;
NAND2   gate14582  (.A(II18425), .B(II18433), .Z(II18435) ) ;
NAND2   gate14583  (.A(WX6173), .B(WX5845), .Z(II18442) ) ;
NAND2   gate14584  (.A(WX6173), .B(II18442), .Z(II18443) ) ;
NAND2   gate14585  (.A(WX5845), .B(II18442), .Z(II18444) ) ;
NAND2   gate14586  (.A(II18443), .B(II18444), .Z(II18441) ) ;
NAND2   gate14587  (.A(WX5909), .B(II18441), .Z(II18449) ) ;
NAND2   gate14588  (.A(WX5909), .B(II18449), .Z(II18450) ) ;
NAND2   gate14589  (.A(II18441), .B(II18449), .Z(II18451) ) ;
NAND2   gate14590  (.A(II18450), .B(II18451), .Z(II18440) ) ;
NAND2   gate14591  (.A(WX5973), .B(WX6037), .Z(II18457) ) ;
NAND2   gate14592  (.A(WX5973), .B(II18457), .Z(II18458) ) ;
NAND2   gate14593  (.A(WX6037), .B(II18457), .Z(II18459) ) ;
NAND2   gate14594  (.A(II18458), .B(II18459), .Z(II18456) ) ;
NAND2   gate14595  (.A(II18440), .B(II18456), .Z(II18464) ) ;
NAND2   gate14596  (.A(II18440), .B(II18464), .Z(II18465) ) ;
NAND2   gate14597  (.A(II18456), .B(II18464), .Z(II18466) ) ;
NAND2   gate14598  (.A(WX6173), .B(WX5847), .Z(II18473) ) ;
NAND2   gate14599  (.A(WX6173), .B(II18473), .Z(II18474) ) ;
NAND2   gate14600  (.A(WX5847), .B(II18473), .Z(II18475) ) ;
NAND2   gate14601  (.A(II18474), .B(II18475), .Z(II18472) ) ;
NAND2   gate14602  (.A(WX5911), .B(II18472), .Z(II18480) ) ;
NAND2   gate14603  (.A(WX5911), .B(II18480), .Z(II18481) ) ;
NAND2   gate14604  (.A(II18472), .B(II18480), .Z(II18482) ) ;
NAND2   gate14605  (.A(II18481), .B(II18482), .Z(II18471) ) ;
NAND2   gate14606  (.A(WX5975), .B(WX6039), .Z(II18488) ) ;
NAND2   gate14607  (.A(WX5975), .B(II18488), .Z(II18489) ) ;
NAND2   gate14608  (.A(WX6039), .B(II18488), .Z(II18490) ) ;
NAND2   gate14609  (.A(II18489), .B(II18490), .Z(II18487) ) ;
NAND2   gate14610  (.A(II18471), .B(II18487), .Z(II18495) ) ;
NAND2   gate14611  (.A(II18471), .B(II18495), .Z(II18496) ) ;
NAND2   gate14612  (.A(II18487), .B(II18495), .Z(II18497) ) ;
NAND2   gate14613  (.A(WX6174), .B(WX5849), .Z(II18504) ) ;
NAND2   gate14614  (.A(WX6174), .B(II18504), .Z(II18505) ) ;
NAND2   gate14615  (.A(WX5849), .B(II18504), .Z(II18506) ) ;
NAND2   gate14616  (.A(II18505), .B(II18506), .Z(II18503) ) ;
NAND2   gate14617  (.A(WX5913), .B(II18503), .Z(II18511) ) ;
NAND2   gate14618  (.A(WX5913), .B(II18511), .Z(II18512) ) ;
NAND2   gate14619  (.A(II18503), .B(II18511), .Z(II18513) ) ;
NAND2   gate14620  (.A(II18512), .B(II18513), .Z(II18502) ) ;
NAND2   gate14621  (.A(WX5977), .B(WX6041), .Z(II18519) ) ;
NAND2   gate14622  (.A(WX5977), .B(II18519), .Z(II18520) ) ;
NAND2   gate14623  (.A(WX6041), .B(II18519), .Z(II18521) ) ;
NAND2   gate14624  (.A(II18520), .B(II18521), .Z(II18518) ) ;
NAND2   gate14625  (.A(II18502), .B(II18518), .Z(II18526) ) ;
NAND2   gate14626  (.A(II18502), .B(II18526), .Z(II18527) ) ;
NAND2   gate14627  (.A(II18518), .B(II18526), .Z(II18528) ) ;
NAND2   gate14628  (.A(WX6174), .B(WX5851), .Z(II18535) ) ;
NAND2   gate14629  (.A(WX6174), .B(II18535), .Z(II18536) ) ;
NAND2   gate14630  (.A(WX5851), .B(II18535), .Z(II18537) ) ;
NAND2   gate14631  (.A(II18536), .B(II18537), .Z(II18534) ) ;
NAND2   gate14632  (.A(WX5915), .B(II18534), .Z(II18542) ) ;
NAND2   gate14633  (.A(WX5915), .B(II18542), .Z(II18543) ) ;
NAND2   gate14634  (.A(II18534), .B(II18542), .Z(II18544) ) ;
NAND2   gate14635  (.A(II18543), .B(II18544), .Z(II18533) ) ;
NAND2   gate14636  (.A(WX5979), .B(WX6043), .Z(II18550) ) ;
NAND2   gate14637  (.A(WX5979), .B(II18550), .Z(II18551) ) ;
NAND2   gate14638  (.A(WX6043), .B(II18550), .Z(II18552) ) ;
NAND2   gate14639  (.A(II18551), .B(II18552), .Z(II18549) ) ;
NAND2   gate14640  (.A(II18533), .B(II18549), .Z(II18557) ) ;
NAND2   gate14641  (.A(II18533), .B(II18557), .Z(II18558) ) ;
NAND2   gate14642  (.A(II18549), .B(II18557), .Z(II18559) ) ;
NAND2   gate14643  (.A(WX6174), .B(WX5853), .Z(II18566) ) ;
NAND2   gate14644  (.A(WX6174), .B(II18566), .Z(II18567) ) ;
NAND2   gate14645  (.A(WX5853), .B(II18566), .Z(II18568) ) ;
NAND2   gate14646  (.A(II18567), .B(II18568), .Z(II18565) ) ;
NAND2   gate14647  (.A(WX5917), .B(II18565), .Z(II18573) ) ;
NAND2   gate14648  (.A(WX5917), .B(II18573), .Z(II18574) ) ;
NAND2   gate14649  (.A(II18565), .B(II18573), .Z(II18575) ) ;
NAND2   gate14650  (.A(II18574), .B(II18575), .Z(II18564) ) ;
NAND2   gate14651  (.A(WX5981), .B(WX6045), .Z(II18581) ) ;
NAND2   gate14652  (.A(WX5981), .B(II18581), .Z(II18582) ) ;
NAND2   gate14653  (.A(WX6045), .B(II18581), .Z(II18583) ) ;
NAND2   gate14654  (.A(II18582), .B(II18583), .Z(II18580) ) ;
NAND2   gate14655  (.A(II18564), .B(II18580), .Z(II18588) ) ;
NAND2   gate14656  (.A(II18564), .B(II18588), .Z(II18589) ) ;
NAND2   gate14657  (.A(II18580), .B(II18588), .Z(II18590) ) ;
NAND2   gate14658  (.A(WX6174), .B(WX5855), .Z(II18597) ) ;
NAND2   gate14659  (.A(WX6174), .B(II18597), .Z(II18598) ) ;
NAND2   gate14660  (.A(WX5855), .B(II18597), .Z(II18599) ) ;
NAND2   gate14661  (.A(II18598), .B(II18599), .Z(II18596) ) ;
NAND2   gate14662  (.A(WX5919), .B(II18596), .Z(II18604) ) ;
NAND2   gate14663  (.A(WX5919), .B(II18604), .Z(II18605) ) ;
NAND2   gate14664  (.A(II18596), .B(II18604), .Z(II18606) ) ;
NAND2   gate14665  (.A(II18605), .B(II18606), .Z(II18595) ) ;
NAND2   gate14666  (.A(WX5983), .B(WX6047), .Z(II18612) ) ;
NAND2   gate14667  (.A(WX5983), .B(II18612), .Z(II18613) ) ;
NAND2   gate14668  (.A(WX6047), .B(II18612), .Z(II18614) ) ;
NAND2   gate14669  (.A(II18613), .B(II18614), .Z(II18611) ) ;
NAND2   gate14670  (.A(II18595), .B(II18611), .Z(II18619) ) ;
NAND2   gate14671  (.A(II18595), .B(II18619), .Z(II18620) ) ;
NAND2   gate14672  (.A(II18611), .B(II18619), .Z(II18621) ) ;
NAND2   gate14673  (.A(WX6174), .B(WX5857), .Z(II18628) ) ;
NAND2   gate14674  (.A(WX6174), .B(II18628), .Z(II18629) ) ;
NAND2   gate14675  (.A(WX5857), .B(II18628), .Z(II18630) ) ;
NAND2   gate14676  (.A(II18629), .B(II18630), .Z(II18627) ) ;
NAND2   gate14677  (.A(WX5921), .B(II18627), .Z(II18635) ) ;
NAND2   gate14678  (.A(WX5921), .B(II18635), .Z(II18636) ) ;
NAND2   gate14679  (.A(II18627), .B(II18635), .Z(II18637) ) ;
NAND2   gate14680  (.A(II18636), .B(II18637), .Z(II18626) ) ;
NAND2   gate14681  (.A(WX5985), .B(WX6049), .Z(II18643) ) ;
NAND2   gate14682  (.A(WX5985), .B(II18643), .Z(II18644) ) ;
NAND2   gate14683  (.A(WX6049), .B(II18643), .Z(II18645) ) ;
NAND2   gate14684  (.A(II18644), .B(II18645), .Z(II18642) ) ;
NAND2   gate14685  (.A(II18626), .B(II18642), .Z(II18650) ) ;
NAND2   gate14686  (.A(II18626), .B(II18650), .Z(II18651) ) ;
NAND2   gate14687  (.A(II18642), .B(II18650), .Z(II18652) ) ;
NAND2   gate14688  (.A(WX6174), .B(WX5859), .Z(II18659) ) ;
NAND2   gate14689  (.A(WX6174), .B(II18659), .Z(II18660) ) ;
NAND2   gate14690  (.A(WX5859), .B(II18659), .Z(II18661) ) ;
NAND2   gate14691  (.A(II18660), .B(II18661), .Z(II18658) ) ;
NAND2   gate14692  (.A(WX5923), .B(II18658), .Z(II18666) ) ;
NAND2   gate14693  (.A(WX5923), .B(II18666), .Z(II18667) ) ;
NAND2   gate14694  (.A(II18658), .B(II18666), .Z(II18668) ) ;
NAND2   gate14695  (.A(II18667), .B(II18668), .Z(II18657) ) ;
NAND2   gate14696  (.A(WX5987), .B(WX6051), .Z(II18674) ) ;
NAND2   gate14697  (.A(WX5987), .B(II18674), .Z(II18675) ) ;
NAND2   gate14698  (.A(WX6051), .B(II18674), .Z(II18676) ) ;
NAND2   gate14699  (.A(II18675), .B(II18676), .Z(II18673) ) ;
NAND2   gate14700  (.A(II18657), .B(II18673), .Z(II18681) ) ;
NAND2   gate14701  (.A(II18657), .B(II18681), .Z(II18682) ) ;
NAND2   gate14702  (.A(II18673), .B(II18681), .Z(II18683) ) ;
NAND2   gate14703  (.A(WX6174), .B(WX5861), .Z(II18690) ) ;
NAND2   gate14704  (.A(WX6174), .B(II18690), .Z(II18691) ) ;
NAND2   gate14705  (.A(WX5861), .B(II18690), .Z(II18692) ) ;
NAND2   gate14706  (.A(II18691), .B(II18692), .Z(II18689) ) ;
NAND2   gate14707  (.A(WX5925), .B(II18689), .Z(II18697) ) ;
NAND2   gate14708  (.A(WX5925), .B(II18697), .Z(II18698) ) ;
NAND2   gate14709  (.A(II18689), .B(II18697), .Z(II18699) ) ;
NAND2   gate14710  (.A(II18698), .B(II18699), .Z(II18688) ) ;
NAND2   gate14711  (.A(WX5989), .B(WX6053), .Z(II18705) ) ;
NAND2   gate14712  (.A(WX5989), .B(II18705), .Z(II18706) ) ;
NAND2   gate14713  (.A(WX6053), .B(II18705), .Z(II18707) ) ;
NAND2   gate14714  (.A(II18706), .B(II18707), .Z(II18704) ) ;
NAND2   gate14715  (.A(II18688), .B(II18704), .Z(II18712) ) ;
NAND2   gate14716  (.A(II18688), .B(II18712), .Z(II18713) ) ;
NAND2   gate14717  (.A(II18704), .B(II18712), .Z(II18714) ) ;
NAND2   gate14718  (.A(WX6174), .B(WX5863), .Z(II18721) ) ;
NAND2   gate14719  (.A(WX6174), .B(II18721), .Z(II18722) ) ;
NAND2   gate14720  (.A(WX5863), .B(II18721), .Z(II18723) ) ;
NAND2   gate14721  (.A(II18722), .B(II18723), .Z(II18720) ) ;
NAND2   gate14722  (.A(WX5927), .B(II18720), .Z(II18728) ) ;
NAND2   gate14723  (.A(WX5927), .B(II18728), .Z(II18729) ) ;
NAND2   gate14724  (.A(II18720), .B(II18728), .Z(II18730) ) ;
NAND2   gate14725  (.A(II18729), .B(II18730), .Z(II18719) ) ;
NAND2   gate14726  (.A(WX5991), .B(WX6055), .Z(II18736) ) ;
NAND2   gate14727  (.A(WX5991), .B(II18736), .Z(II18737) ) ;
NAND2   gate14728  (.A(WX6055), .B(II18736), .Z(II18738) ) ;
NAND2   gate14729  (.A(II18737), .B(II18738), .Z(II18735) ) ;
NAND2   gate14730  (.A(II18719), .B(II18735), .Z(II18743) ) ;
NAND2   gate14731  (.A(II18719), .B(II18743), .Z(II18744) ) ;
NAND2   gate14732  (.A(II18735), .B(II18743), .Z(II18745) ) ;
NAND2   gate14733  (.A(WX6174), .B(WX5865), .Z(II18752) ) ;
NAND2   gate14734  (.A(WX6174), .B(II18752), .Z(II18753) ) ;
NAND2   gate14735  (.A(WX5865), .B(II18752), .Z(II18754) ) ;
NAND2   gate14736  (.A(II18753), .B(II18754), .Z(II18751) ) ;
NAND2   gate14737  (.A(WX5929), .B(II18751), .Z(II18759) ) ;
NAND2   gate14738  (.A(WX5929), .B(II18759), .Z(II18760) ) ;
NAND2   gate14739  (.A(II18751), .B(II18759), .Z(II18761) ) ;
NAND2   gate14740  (.A(II18760), .B(II18761), .Z(II18750) ) ;
NAND2   gate14741  (.A(WX5993), .B(WX6057), .Z(II18767) ) ;
NAND2   gate14742  (.A(WX5993), .B(II18767), .Z(II18768) ) ;
NAND2   gate14743  (.A(WX6057), .B(II18767), .Z(II18769) ) ;
NAND2   gate14744  (.A(II18768), .B(II18769), .Z(II18766) ) ;
NAND2   gate14745  (.A(II18750), .B(II18766), .Z(II18774) ) ;
NAND2   gate14746  (.A(II18750), .B(II18774), .Z(II18775) ) ;
NAND2   gate14747  (.A(II18766), .B(II18774), .Z(II18776) ) ;
NAND2   gate14748  (.A(WX6174), .B(WX5867), .Z(II18783) ) ;
NAND2   gate14749  (.A(WX6174), .B(II18783), .Z(II18784) ) ;
NAND2   gate14750  (.A(WX5867), .B(II18783), .Z(II18785) ) ;
NAND2   gate14751  (.A(II18784), .B(II18785), .Z(II18782) ) ;
NAND2   gate14752  (.A(WX5931), .B(II18782), .Z(II18790) ) ;
NAND2   gate14753  (.A(WX5931), .B(II18790), .Z(II18791) ) ;
NAND2   gate14754  (.A(II18782), .B(II18790), .Z(II18792) ) ;
NAND2   gate14755  (.A(II18791), .B(II18792), .Z(II18781) ) ;
NAND2   gate14756  (.A(WX5995), .B(WX6059), .Z(II18798) ) ;
NAND2   gate14757  (.A(WX5995), .B(II18798), .Z(II18799) ) ;
NAND2   gate14758  (.A(WX6059), .B(II18798), .Z(II18800) ) ;
NAND2   gate14759  (.A(II18799), .B(II18800), .Z(II18797) ) ;
NAND2   gate14760  (.A(II18781), .B(II18797), .Z(II18805) ) ;
NAND2   gate14761  (.A(II18781), .B(II18805), .Z(II18806) ) ;
NAND2   gate14762  (.A(II18797), .B(II18805), .Z(II18807) ) ;
NAND2   gate14763  (.A(WX6174), .B(WX5869), .Z(II18814) ) ;
NAND2   gate14764  (.A(WX6174), .B(II18814), .Z(II18815) ) ;
NAND2   gate14765  (.A(WX5869), .B(II18814), .Z(II18816) ) ;
NAND2   gate14766  (.A(II18815), .B(II18816), .Z(II18813) ) ;
NAND2   gate14767  (.A(WX5933), .B(II18813), .Z(II18821) ) ;
NAND2   gate14768  (.A(WX5933), .B(II18821), .Z(II18822) ) ;
NAND2   gate14769  (.A(II18813), .B(II18821), .Z(II18823) ) ;
NAND2   gate14770  (.A(II18822), .B(II18823), .Z(II18812) ) ;
NAND2   gate14771  (.A(WX5997), .B(WX6061), .Z(II18829) ) ;
NAND2   gate14772  (.A(WX5997), .B(II18829), .Z(II18830) ) ;
NAND2   gate14773  (.A(WX6061), .B(II18829), .Z(II18831) ) ;
NAND2   gate14774  (.A(II18830), .B(II18831), .Z(II18828) ) ;
NAND2   gate14775  (.A(II18812), .B(II18828), .Z(II18836) ) ;
NAND2   gate14776  (.A(II18812), .B(II18836), .Z(II18837) ) ;
NAND2   gate14777  (.A(II18828), .B(II18836), .Z(II18838) ) ;
NAND2   gate14778  (.A(WX6174), .B(WX5871), .Z(II18845) ) ;
NAND2   gate14779  (.A(WX6174), .B(II18845), .Z(II18846) ) ;
NAND2   gate14780  (.A(WX5871), .B(II18845), .Z(II18847) ) ;
NAND2   gate14781  (.A(II18846), .B(II18847), .Z(II18844) ) ;
NAND2   gate14782  (.A(WX5935), .B(II18844), .Z(II18852) ) ;
NAND2   gate14783  (.A(WX5935), .B(II18852), .Z(II18853) ) ;
NAND2   gate14784  (.A(II18844), .B(II18852), .Z(II18854) ) ;
NAND2   gate14785  (.A(II18853), .B(II18854), .Z(II18843) ) ;
NAND2   gate14786  (.A(WX5999), .B(WX6063), .Z(II18860) ) ;
NAND2   gate14787  (.A(WX5999), .B(II18860), .Z(II18861) ) ;
NAND2   gate14788  (.A(WX6063), .B(II18860), .Z(II18862) ) ;
NAND2   gate14789  (.A(II18861), .B(II18862), .Z(II18859) ) ;
NAND2   gate14790  (.A(II18843), .B(II18859), .Z(II18867) ) ;
NAND2   gate14791  (.A(II18843), .B(II18867), .Z(II18868) ) ;
NAND2   gate14792  (.A(II18859), .B(II18867), .Z(II18869) ) ;
NAND2   gate14793  (.A(WX6174), .B(WX5873), .Z(II18876) ) ;
NAND2   gate14794  (.A(WX6174), .B(II18876), .Z(II18877) ) ;
NAND2   gate14795  (.A(WX5873), .B(II18876), .Z(II18878) ) ;
NAND2   gate14796  (.A(II18877), .B(II18878), .Z(II18875) ) ;
NAND2   gate14797  (.A(WX5937), .B(II18875), .Z(II18883) ) ;
NAND2   gate14798  (.A(WX5937), .B(II18883), .Z(II18884) ) ;
NAND2   gate14799  (.A(II18875), .B(II18883), .Z(II18885) ) ;
NAND2   gate14800  (.A(II18884), .B(II18885), .Z(II18874) ) ;
NAND2   gate14801  (.A(WX6001), .B(WX6065), .Z(II18891) ) ;
NAND2   gate14802  (.A(WX6001), .B(II18891), .Z(II18892) ) ;
NAND2   gate14803  (.A(WX6065), .B(II18891), .Z(II18893) ) ;
NAND2   gate14804  (.A(II18892), .B(II18893), .Z(II18890) ) ;
NAND2   gate14805  (.A(II18874), .B(II18890), .Z(II18898) ) ;
NAND2   gate14806  (.A(II18874), .B(II18898), .Z(II18899) ) ;
NAND2   gate14807  (.A(II18890), .B(II18898), .Z(II18900) ) ;
NAND2   gate14808  (.A(WX6174), .B(WX5875), .Z(II18907) ) ;
NAND2   gate14809  (.A(WX6174), .B(II18907), .Z(II18908) ) ;
NAND2   gate14810  (.A(WX5875), .B(II18907), .Z(II18909) ) ;
NAND2   gate14811  (.A(II18908), .B(II18909), .Z(II18906) ) ;
NAND2   gate14812  (.A(WX5939), .B(II18906), .Z(II18914) ) ;
NAND2   gate14813  (.A(WX5939), .B(II18914), .Z(II18915) ) ;
NAND2   gate14814  (.A(II18906), .B(II18914), .Z(II18916) ) ;
NAND2   gate14815  (.A(II18915), .B(II18916), .Z(II18905) ) ;
NAND2   gate14816  (.A(WX6003), .B(WX6067), .Z(II18922) ) ;
NAND2   gate14817  (.A(WX6003), .B(II18922), .Z(II18923) ) ;
NAND2   gate14818  (.A(WX6067), .B(II18922), .Z(II18924) ) ;
NAND2   gate14819  (.A(II18923), .B(II18924), .Z(II18921) ) ;
NAND2   gate14820  (.A(II18905), .B(II18921), .Z(II18929) ) ;
NAND2   gate14821  (.A(II18905), .B(II18929), .Z(II18930) ) ;
NAND2   gate14822  (.A(II18921), .B(II18929), .Z(II18931) ) ;
NAND2   gate14823  (.A(WX6174), .B(WX5877), .Z(II18938) ) ;
NAND2   gate14824  (.A(WX6174), .B(II18938), .Z(II18939) ) ;
NAND2   gate14825  (.A(WX5877), .B(II18938), .Z(II18940) ) ;
NAND2   gate14826  (.A(II18939), .B(II18940), .Z(II18937) ) ;
NAND2   gate14827  (.A(WX5941), .B(II18937), .Z(II18945) ) ;
NAND2   gate14828  (.A(WX5941), .B(II18945), .Z(II18946) ) ;
NAND2   gate14829  (.A(II18937), .B(II18945), .Z(II18947) ) ;
NAND2   gate14830  (.A(II18946), .B(II18947), .Z(II18936) ) ;
NAND2   gate14831  (.A(WX6005), .B(WX6069), .Z(II18953) ) ;
NAND2   gate14832  (.A(WX6005), .B(II18953), .Z(II18954) ) ;
NAND2   gate14833  (.A(WX6069), .B(II18953), .Z(II18955) ) ;
NAND2   gate14834  (.A(II18954), .B(II18955), .Z(II18952) ) ;
NAND2   gate14835  (.A(II18936), .B(II18952), .Z(II18960) ) ;
NAND2   gate14836  (.A(II18936), .B(II18960), .Z(II18961) ) ;
NAND2   gate14837  (.A(II18952), .B(II18960), .Z(II18962) ) ;
NAND2   gate14838  (.A(WX6174), .B(WX5879), .Z(II18969) ) ;
NAND2   gate14839  (.A(WX6174), .B(II18969), .Z(II18970) ) ;
NAND2   gate14840  (.A(WX5879), .B(II18969), .Z(II18971) ) ;
NAND2   gate14841  (.A(II18970), .B(II18971), .Z(II18968) ) ;
NAND2   gate14842  (.A(WX5943), .B(II18968), .Z(II18976) ) ;
NAND2   gate14843  (.A(WX5943), .B(II18976), .Z(II18977) ) ;
NAND2   gate14844  (.A(II18968), .B(II18976), .Z(II18978) ) ;
NAND2   gate14845  (.A(II18977), .B(II18978), .Z(II18967) ) ;
NAND2   gate14846  (.A(WX6007), .B(WX6071), .Z(II18984) ) ;
NAND2   gate14847  (.A(WX6007), .B(II18984), .Z(II18985) ) ;
NAND2   gate14848  (.A(WX6071), .B(II18984), .Z(II18986) ) ;
NAND2   gate14849  (.A(II18985), .B(II18986), .Z(II18983) ) ;
NAND2   gate14850  (.A(II18967), .B(II18983), .Z(II18991) ) ;
NAND2   gate14851  (.A(II18967), .B(II18991), .Z(II18992) ) ;
NAND2   gate14852  (.A(II18983), .B(II18991), .Z(II18993) ) ;
NAND2   gate14853  (.A(WX5752), .B(WX5657), .Z(II19072) ) ;
NAND2   gate14854  (.A(WX5752), .B(II19072), .Z(II19073) ) ;
NAND2   gate14855  (.A(WX5657), .B(II19072), .Z(II19074) ) ;
NAND2   gate14856  (.A(WX5753), .B(WX5659), .Z(II19085) ) ;
NAND2   gate14857  (.A(WX5753), .B(II19085), .Z(II19086) ) ;
NAND2   gate14858  (.A(WX5659), .B(II19085), .Z(II19087) ) ;
NAND2   gate14859  (.A(WX5754), .B(WX5661), .Z(II19098) ) ;
NAND2   gate14860  (.A(WX5754), .B(II19098), .Z(II19099) ) ;
NAND2   gate14861  (.A(WX5661), .B(II19098), .Z(II19100) ) ;
NAND2   gate14862  (.A(WX5755), .B(WX5663), .Z(II19111) ) ;
NAND2   gate14863  (.A(WX5755), .B(II19111), .Z(II19112) ) ;
NAND2   gate14864  (.A(WX5663), .B(II19111), .Z(II19113) ) ;
NAND2   gate14865  (.A(WX5756), .B(WX5665), .Z(II19124) ) ;
NAND2   gate14866  (.A(WX5756), .B(II19124), .Z(II19125) ) ;
NAND2   gate14867  (.A(WX5665), .B(II19124), .Z(II19126) ) ;
NAND2   gate14868  (.A(WX5757), .B(WX5667), .Z(II19137) ) ;
NAND2   gate14869  (.A(WX5757), .B(II19137), .Z(II19138) ) ;
NAND2   gate14870  (.A(WX5667), .B(II19137), .Z(II19139) ) ;
NAND2   gate14871  (.A(WX5758), .B(WX5669), .Z(II19150) ) ;
NAND2   gate14872  (.A(WX5758), .B(II19150), .Z(II19151) ) ;
NAND2   gate14873  (.A(WX5669), .B(II19150), .Z(II19152) ) ;
NAND2   gate14874  (.A(WX5759), .B(WX5671), .Z(II19163) ) ;
NAND2   gate14875  (.A(WX5759), .B(II19163), .Z(II19164) ) ;
NAND2   gate14876  (.A(WX5671), .B(II19163), .Z(II19165) ) ;
NAND2   gate14877  (.A(WX5760), .B(WX5673), .Z(II19176) ) ;
NAND2   gate14878  (.A(WX5760), .B(II19176), .Z(II19177) ) ;
NAND2   gate14879  (.A(WX5673), .B(II19176), .Z(II19178) ) ;
NAND2   gate14880  (.A(WX5761), .B(WX5675), .Z(II19189) ) ;
NAND2   gate14881  (.A(WX5761), .B(II19189), .Z(II19190) ) ;
NAND2   gate14882  (.A(WX5675), .B(II19189), .Z(II19191) ) ;
NAND2   gate14883  (.A(WX5762), .B(WX5677), .Z(II19202) ) ;
NAND2   gate14884  (.A(WX5762), .B(II19202), .Z(II19203) ) ;
NAND2   gate14885  (.A(WX5677), .B(II19202), .Z(II19204) ) ;
NAND2   gate14886  (.A(WX5763), .B(WX5679), .Z(II19215) ) ;
NAND2   gate14887  (.A(WX5763), .B(II19215), .Z(II19216) ) ;
NAND2   gate14888  (.A(WX5679), .B(II19215), .Z(II19217) ) ;
NAND2   gate14889  (.A(WX5764), .B(WX5681), .Z(II19228) ) ;
NAND2   gate14890  (.A(WX5764), .B(II19228), .Z(II19229) ) ;
NAND2   gate14891  (.A(WX5681), .B(II19228), .Z(II19230) ) ;
NAND2   gate14892  (.A(WX5765), .B(WX5683), .Z(II19241) ) ;
NAND2   gate14893  (.A(WX5765), .B(II19241), .Z(II19242) ) ;
NAND2   gate14894  (.A(WX5683), .B(II19241), .Z(II19243) ) ;
NAND2   gate14895  (.A(WX5766), .B(WX5685), .Z(II19254) ) ;
NAND2   gate14896  (.A(WX5766), .B(II19254), .Z(II19255) ) ;
NAND2   gate14897  (.A(WX5685), .B(II19254), .Z(II19256) ) ;
NAND2   gate14898  (.A(WX5767), .B(WX5687), .Z(II19267) ) ;
NAND2   gate14899  (.A(WX5767), .B(II19267), .Z(II19268) ) ;
NAND2   gate14900  (.A(WX5687), .B(II19267), .Z(II19269) ) ;
NAND2   gate14901  (.A(WX5768), .B(WX5689), .Z(II19280) ) ;
NAND2   gate14902  (.A(WX5768), .B(II19280), .Z(II19281) ) ;
NAND2   gate14903  (.A(WX5689), .B(II19280), .Z(II19282) ) ;
NAND2   gate14904  (.A(WX5769), .B(WX5691), .Z(II19293) ) ;
NAND2   gate14905  (.A(WX5769), .B(II19293), .Z(II19294) ) ;
NAND2   gate14906  (.A(WX5691), .B(II19293), .Z(II19295) ) ;
NAND2   gate14907  (.A(WX5770), .B(WX5693), .Z(II19306) ) ;
NAND2   gate14908  (.A(WX5770), .B(II19306), .Z(II19307) ) ;
NAND2   gate14909  (.A(WX5693), .B(II19306), .Z(II19308) ) ;
NAND2   gate14910  (.A(WX5771), .B(WX5695), .Z(II19319) ) ;
NAND2   gate14911  (.A(WX5771), .B(II19319), .Z(II19320) ) ;
NAND2   gate14912  (.A(WX5695), .B(II19319), .Z(II19321) ) ;
NAND2   gate14913  (.A(WX5772), .B(WX5697), .Z(II19332) ) ;
NAND2   gate14914  (.A(WX5772), .B(II19332), .Z(II19333) ) ;
NAND2   gate14915  (.A(WX5697), .B(II19332), .Z(II19334) ) ;
NAND2   gate14916  (.A(WX5773), .B(WX5699), .Z(II19345) ) ;
NAND2   gate14917  (.A(WX5773), .B(II19345), .Z(II19346) ) ;
NAND2   gate14918  (.A(WX5699), .B(II19345), .Z(II19347) ) ;
NAND2   gate14919  (.A(WX5774), .B(WX5701), .Z(II19358) ) ;
NAND2   gate14920  (.A(WX5774), .B(II19358), .Z(II19359) ) ;
NAND2   gate14921  (.A(WX5701), .B(II19358), .Z(II19360) ) ;
NAND2   gate14922  (.A(WX5775), .B(WX5703), .Z(II19371) ) ;
NAND2   gate14923  (.A(WX5775), .B(II19371), .Z(II19372) ) ;
NAND2   gate14924  (.A(WX5703), .B(II19371), .Z(II19373) ) ;
NAND2   gate14925  (.A(WX5776), .B(WX5705), .Z(II19384) ) ;
NAND2   gate14926  (.A(WX5776), .B(II19384), .Z(II19385) ) ;
NAND2   gate14927  (.A(WX5705), .B(II19384), .Z(II19386) ) ;
NAND2   gate14928  (.A(WX5777), .B(WX5707), .Z(II19397) ) ;
NAND2   gate14929  (.A(WX5777), .B(II19397), .Z(II19398) ) ;
NAND2   gate14930  (.A(WX5707), .B(II19397), .Z(II19399) ) ;
NAND2   gate14931  (.A(WX5778), .B(WX5709), .Z(II19410) ) ;
NAND2   gate14932  (.A(WX5778), .B(II19410), .Z(II19411) ) ;
NAND2   gate14933  (.A(WX5709), .B(II19410), .Z(II19412) ) ;
NAND2   gate14934  (.A(WX5779), .B(WX5711), .Z(II19423) ) ;
NAND2   gate14935  (.A(WX5779), .B(II19423), .Z(II19424) ) ;
NAND2   gate14936  (.A(WX5711), .B(II19423), .Z(II19425) ) ;
NAND2   gate14937  (.A(WX5780), .B(WX5713), .Z(II19436) ) ;
NAND2   gate14938  (.A(WX5780), .B(II19436), .Z(II19437) ) ;
NAND2   gate14939  (.A(WX5713), .B(II19436), .Z(II19438) ) ;
NAND2   gate14940  (.A(WX5781), .B(WX5715), .Z(II19449) ) ;
NAND2   gate14941  (.A(WX5781), .B(II19449), .Z(II19450) ) ;
NAND2   gate14942  (.A(WX5715), .B(II19449), .Z(II19451) ) ;
NAND2   gate14943  (.A(WX5782), .B(WX5717), .Z(II19462) ) ;
NAND2   gate14944  (.A(WX5782), .B(II19462), .Z(II19463) ) ;
NAND2   gate14945  (.A(WX5717), .B(II19462), .Z(II19464) ) ;
NAND2   gate14946  (.A(WX5783), .B(WX5719), .Z(II19475) ) ;
NAND2   gate14947  (.A(WX5783), .B(II19475), .Z(II19476) ) ;
NAND2   gate14948  (.A(WX5719), .B(II19475), .Z(II19477) ) ;
NAND2   gate14949  (.A(WX5799), .B(CRC_OUT_5_31), .Z(II19490) ) ;
NAND2   gate14950  (.A(WX5799), .B(II19490), .Z(II19491) ) ;
NAND2   gate14951  (.A(CRC_OUT_5_31), .B(II19490), .Z(II19492) ) ;
NAND2   gate14952  (.A(II19491), .B(II19492), .Z(II19489) ) ;
NAND2   gate14953  (.A(CRC_OUT_5_15), .B(II19489), .Z(II19497) ) ;
NAND2   gate14954  (.A(CRC_OUT_5_15), .B(II19497), .Z(II19498) ) ;
NAND2   gate14955  (.A(II19489), .B(II19497), .Z(II19499) ) ;
NAND2   gate14956  (.A(WX5804), .B(CRC_OUT_5_31), .Z(II19505) ) ;
NAND2   gate14957  (.A(WX5804), .B(II19505), .Z(II19506) ) ;
NAND2   gate14958  (.A(CRC_OUT_5_31), .B(II19505), .Z(II19507) ) ;
NAND2   gate14959  (.A(II19506), .B(II19507), .Z(II19504) ) ;
NAND2   gate14960  (.A(CRC_OUT_5_10), .B(II19504), .Z(II19512) ) ;
NAND2   gate14961  (.A(CRC_OUT_5_10), .B(II19512), .Z(II19513) ) ;
NAND2   gate14962  (.A(II19504), .B(II19512), .Z(II19514) ) ;
NAND2   gate14963  (.A(WX5811), .B(CRC_OUT_5_31), .Z(II19520) ) ;
NAND2   gate14964  (.A(WX5811), .B(II19520), .Z(II19521) ) ;
NAND2   gate14965  (.A(CRC_OUT_5_31), .B(II19520), .Z(II19522) ) ;
NAND2   gate14966  (.A(II19521), .B(II19522), .Z(II19519) ) ;
NAND2   gate14967  (.A(CRC_OUT_5_3), .B(II19519), .Z(II19527) ) ;
NAND2   gate14968  (.A(CRC_OUT_5_3), .B(II19527), .Z(II19528) ) ;
NAND2   gate14969  (.A(II19519), .B(II19527), .Z(II19529) ) ;
NAND2   gate14970  (.A(WX5815), .B(CRC_OUT_5_31), .Z(II19534) ) ;
NAND2   gate14971  (.A(WX5815), .B(II19534), .Z(II19535) ) ;
NAND2   gate14972  (.A(CRC_OUT_5_31), .B(II19534), .Z(II19536) ) ;
NAND2   gate14973  (.A(WX5784), .B(CRC_OUT_5_30), .Z(II19541) ) ;
NAND2   gate14974  (.A(WX5784), .B(II19541), .Z(II19542) ) ;
NAND2   gate14975  (.A(CRC_OUT_5_30), .B(II19541), .Z(II19543) ) ;
NAND2   gate14976  (.A(WX5785), .B(CRC_OUT_5_29), .Z(II19548) ) ;
NAND2   gate14977  (.A(WX5785), .B(II19548), .Z(II19549) ) ;
NAND2   gate14978  (.A(CRC_OUT_5_29), .B(II19548), .Z(II19550) ) ;
NAND2   gate14979  (.A(WX5786), .B(CRC_OUT_5_28), .Z(II19555) ) ;
NAND2   gate14980  (.A(WX5786), .B(II19555), .Z(II19556) ) ;
NAND2   gate14981  (.A(CRC_OUT_5_28), .B(II19555), .Z(II19557) ) ;
NAND2   gate14982  (.A(WX5787), .B(CRC_OUT_5_27), .Z(II19562) ) ;
NAND2   gate14983  (.A(WX5787), .B(II19562), .Z(II19563) ) ;
NAND2   gate14984  (.A(CRC_OUT_5_27), .B(II19562), .Z(II19564) ) ;
NAND2   gate14985  (.A(WX5788), .B(CRC_OUT_5_26), .Z(II19569) ) ;
NAND2   gate14986  (.A(WX5788), .B(II19569), .Z(II19570) ) ;
NAND2   gate14987  (.A(CRC_OUT_5_26), .B(II19569), .Z(II19571) ) ;
NAND2   gate14988  (.A(WX5789), .B(CRC_OUT_5_25), .Z(II19576) ) ;
NAND2   gate14989  (.A(WX5789), .B(II19576), .Z(II19577) ) ;
NAND2   gate14990  (.A(CRC_OUT_5_25), .B(II19576), .Z(II19578) ) ;
NAND2   gate14991  (.A(WX5790), .B(CRC_OUT_5_24), .Z(II19583) ) ;
NAND2   gate14992  (.A(WX5790), .B(II19583), .Z(II19584) ) ;
NAND2   gate14993  (.A(CRC_OUT_5_24), .B(II19583), .Z(II19585) ) ;
NAND2   gate14994  (.A(WX5791), .B(CRC_OUT_5_23), .Z(II19590) ) ;
NAND2   gate14995  (.A(WX5791), .B(II19590), .Z(II19591) ) ;
NAND2   gate14996  (.A(CRC_OUT_5_23), .B(II19590), .Z(II19592) ) ;
NAND2   gate14997  (.A(WX5792), .B(CRC_OUT_5_22), .Z(II19597) ) ;
NAND2   gate14998  (.A(WX5792), .B(II19597), .Z(II19598) ) ;
NAND2   gate14999  (.A(CRC_OUT_5_22), .B(II19597), .Z(II19599) ) ;
NAND2   gate15000  (.A(WX5793), .B(CRC_OUT_5_21), .Z(II19604) ) ;
NAND2   gate15001  (.A(WX5793), .B(II19604), .Z(II19605) ) ;
NAND2   gate15002  (.A(CRC_OUT_5_21), .B(II19604), .Z(II19606) ) ;
NAND2   gate15003  (.A(WX5794), .B(CRC_OUT_5_20), .Z(II19611) ) ;
NAND2   gate15004  (.A(WX5794), .B(II19611), .Z(II19612) ) ;
NAND2   gate15005  (.A(CRC_OUT_5_20), .B(II19611), .Z(II19613) ) ;
NAND2   gate15006  (.A(WX5795), .B(CRC_OUT_5_19), .Z(II19618) ) ;
NAND2   gate15007  (.A(WX5795), .B(II19618), .Z(II19619) ) ;
NAND2   gate15008  (.A(CRC_OUT_5_19), .B(II19618), .Z(II19620) ) ;
NAND2   gate15009  (.A(WX5796), .B(CRC_OUT_5_18), .Z(II19625) ) ;
NAND2   gate15010  (.A(WX5796), .B(II19625), .Z(II19626) ) ;
NAND2   gate15011  (.A(CRC_OUT_5_18), .B(II19625), .Z(II19627) ) ;
NAND2   gate15012  (.A(WX5797), .B(CRC_OUT_5_17), .Z(II19632) ) ;
NAND2   gate15013  (.A(WX5797), .B(II19632), .Z(II19633) ) ;
NAND2   gate15014  (.A(CRC_OUT_5_17), .B(II19632), .Z(II19634) ) ;
NAND2   gate15015  (.A(WX5798), .B(CRC_OUT_5_16), .Z(II19639) ) ;
NAND2   gate15016  (.A(WX5798), .B(II19639), .Z(II19640) ) ;
NAND2   gate15017  (.A(CRC_OUT_5_16), .B(II19639), .Z(II19641) ) ;
NAND2   gate15018  (.A(WX5800), .B(CRC_OUT_5_14), .Z(II19646) ) ;
NAND2   gate15019  (.A(WX5800), .B(II19646), .Z(II19647) ) ;
NAND2   gate15020  (.A(CRC_OUT_5_14), .B(II19646), .Z(II19648) ) ;
NAND2   gate15021  (.A(WX5801), .B(CRC_OUT_5_13), .Z(II19653) ) ;
NAND2   gate15022  (.A(WX5801), .B(II19653), .Z(II19654) ) ;
NAND2   gate15023  (.A(CRC_OUT_5_13), .B(II19653), .Z(II19655) ) ;
NAND2   gate15024  (.A(WX5802), .B(CRC_OUT_5_12), .Z(II19660) ) ;
NAND2   gate15025  (.A(WX5802), .B(II19660), .Z(II19661) ) ;
NAND2   gate15026  (.A(CRC_OUT_5_12), .B(II19660), .Z(II19662) ) ;
NAND2   gate15027  (.A(WX5803), .B(CRC_OUT_5_11), .Z(II19667) ) ;
NAND2   gate15028  (.A(WX5803), .B(II19667), .Z(II19668) ) ;
NAND2   gate15029  (.A(CRC_OUT_5_11), .B(II19667), .Z(II19669) ) ;
NAND2   gate15030  (.A(WX5805), .B(CRC_OUT_5_9), .Z(II19674) ) ;
NAND2   gate15031  (.A(WX5805), .B(II19674), .Z(II19675) ) ;
NAND2   gate15032  (.A(CRC_OUT_5_9), .B(II19674), .Z(II19676) ) ;
NAND2   gate15033  (.A(WX5806), .B(CRC_OUT_5_8), .Z(II19681) ) ;
NAND2   gate15034  (.A(WX5806), .B(II19681), .Z(II19682) ) ;
NAND2   gate15035  (.A(CRC_OUT_5_8), .B(II19681), .Z(II19683) ) ;
NAND2   gate15036  (.A(WX5807), .B(CRC_OUT_5_7), .Z(II19688) ) ;
NAND2   gate15037  (.A(WX5807), .B(II19688), .Z(II19689) ) ;
NAND2   gate15038  (.A(CRC_OUT_5_7), .B(II19688), .Z(II19690) ) ;
NAND2   gate15039  (.A(WX5808), .B(CRC_OUT_5_6), .Z(II19695) ) ;
NAND2   gate15040  (.A(WX5808), .B(II19695), .Z(II19696) ) ;
NAND2   gate15041  (.A(CRC_OUT_5_6), .B(II19695), .Z(II19697) ) ;
NAND2   gate15042  (.A(WX5809), .B(CRC_OUT_5_5), .Z(II19702) ) ;
NAND2   gate15043  (.A(WX5809), .B(II19702), .Z(II19703) ) ;
NAND2   gate15044  (.A(CRC_OUT_5_5), .B(II19702), .Z(II19704) ) ;
NAND2   gate15045  (.A(WX5810), .B(CRC_OUT_5_4), .Z(II19709) ) ;
NAND2   gate15046  (.A(WX5810), .B(II19709), .Z(II19710) ) ;
NAND2   gate15047  (.A(CRC_OUT_5_4), .B(II19709), .Z(II19711) ) ;
NAND2   gate15048  (.A(WX5812), .B(CRC_OUT_5_2), .Z(II19716) ) ;
NAND2   gate15049  (.A(WX5812), .B(II19716), .Z(II19717) ) ;
NAND2   gate15050  (.A(CRC_OUT_5_2), .B(II19716), .Z(II19718) ) ;
NAND2   gate15051  (.A(WX5813), .B(CRC_OUT_5_1), .Z(II19723) ) ;
NAND2   gate15052  (.A(WX5813), .B(II19723), .Z(II19724) ) ;
NAND2   gate15053  (.A(CRC_OUT_5_1), .B(II19723), .Z(II19725) ) ;
NAND2   gate15054  (.A(WX5814), .B(CRC_OUT_5_0), .Z(II19730) ) ;
NAND2   gate15055  (.A(WX5814), .B(II19730), .Z(II19731) ) ;
NAND2   gate15056  (.A(CRC_OUT_5_0), .B(II19730), .Z(II19732) ) ;
NAND2   gate15057  (.A(WX7466), .B(WX7110), .Z(II22013) ) ;
NAND2   gate15058  (.A(WX7466), .B(II22013), .Z(II22014) ) ;
NAND2   gate15059  (.A(WX7110), .B(II22013), .Z(II22015) ) ;
NAND2   gate15060  (.A(II22014), .B(II22015), .Z(II22012) ) ;
NAND2   gate15061  (.A(WX7174), .B(II22012), .Z(II22020) ) ;
NAND2   gate15062  (.A(WX7174), .B(II22020), .Z(II22021) ) ;
NAND2   gate15063  (.A(II22012), .B(II22020), .Z(II22022) ) ;
NAND2   gate15064  (.A(II22021), .B(II22022), .Z(II22011) ) ;
NAND2   gate15065  (.A(WX7238), .B(WX7302), .Z(II22028) ) ;
NAND2   gate15066  (.A(WX7238), .B(II22028), .Z(II22029) ) ;
NAND2   gate15067  (.A(WX7302), .B(II22028), .Z(II22030) ) ;
NAND2   gate15068  (.A(II22029), .B(II22030), .Z(II22027) ) ;
NAND2   gate15069  (.A(II22011), .B(II22027), .Z(II22035) ) ;
NAND2   gate15070  (.A(II22011), .B(II22035), .Z(II22036) ) ;
NAND2   gate15071  (.A(II22027), .B(II22035), .Z(II22037) ) ;
NAND2   gate15072  (.A(WX7466), .B(WX7112), .Z(II22044) ) ;
NAND2   gate15073  (.A(WX7466), .B(II22044), .Z(II22045) ) ;
NAND2   gate15074  (.A(WX7112), .B(II22044), .Z(II22046) ) ;
NAND2   gate15075  (.A(II22045), .B(II22046), .Z(II22043) ) ;
NAND2   gate15076  (.A(WX7176), .B(II22043), .Z(II22051) ) ;
NAND2   gate15077  (.A(WX7176), .B(II22051), .Z(II22052) ) ;
NAND2   gate15078  (.A(II22043), .B(II22051), .Z(II22053) ) ;
NAND2   gate15079  (.A(II22052), .B(II22053), .Z(II22042) ) ;
NAND2   gate15080  (.A(WX7240), .B(WX7304), .Z(II22059) ) ;
NAND2   gate15081  (.A(WX7240), .B(II22059), .Z(II22060) ) ;
NAND2   gate15082  (.A(WX7304), .B(II22059), .Z(II22061) ) ;
NAND2   gate15083  (.A(II22060), .B(II22061), .Z(II22058) ) ;
NAND2   gate15084  (.A(II22042), .B(II22058), .Z(II22066) ) ;
NAND2   gate15085  (.A(II22042), .B(II22066), .Z(II22067) ) ;
NAND2   gate15086  (.A(II22058), .B(II22066), .Z(II22068) ) ;
NAND2   gate15087  (.A(WX7466), .B(WX7114), .Z(II22075) ) ;
NAND2   gate15088  (.A(WX7466), .B(II22075), .Z(II22076) ) ;
NAND2   gate15089  (.A(WX7114), .B(II22075), .Z(II22077) ) ;
NAND2   gate15090  (.A(II22076), .B(II22077), .Z(II22074) ) ;
NAND2   gate15091  (.A(WX7178), .B(II22074), .Z(II22082) ) ;
NAND2   gate15092  (.A(WX7178), .B(II22082), .Z(II22083) ) ;
NAND2   gate15093  (.A(II22074), .B(II22082), .Z(II22084) ) ;
NAND2   gate15094  (.A(II22083), .B(II22084), .Z(II22073) ) ;
NAND2   gate15095  (.A(WX7242), .B(WX7306), .Z(II22090) ) ;
NAND2   gate15096  (.A(WX7242), .B(II22090), .Z(II22091) ) ;
NAND2   gate15097  (.A(WX7306), .B(II22090), .Z(II22092) ) ;
NAND2   gate15098  (.A(II22091), .B(II22092), .Z(II22089) ) ;
NAND2   gate15099  (.A(II22073), .B(II22089), .Z(II22097) ) ;
NAND2   gate15100  (.A(II22073), .B(II22097), .Z(II22098) ) ;
NAND2   gate15101  (.A(II22089), .B(II22097), .Z(II22099) ) ;
NAND2   gate15102  (.A(WX7466), .B(WX7116), .Z(II22106) ) ;
NAND2   gate15103  (.A(WX7466), .B(II22106), .Z(II22107) ) ;
NAND2   gate15104  (.A(WX7116), .B(II22106), .Z(II22108) ) ;
NAND2   gate15105  (.A(II22107), .B(II22108), .Z(II22105) ) ;
NAND2   gate15106  (.A(WX7180), .B(II22105), .Z(II22113) ) ;
NAND2   gate15107  (.A(WX7180), .B(II22113), .Z(II22114) ) ;
NAND2   gate15108  (.A(II22105), .B(II22113), .Z(II22115) ) ;
NAND2   gate15109  (.A(II22114), .B(II22115), .Z(II22104) ) ;
NAND2   gate15110  (.A(WX7244), .B(WX7308), .Z(II22121) ) ;
NAND2   gate15111  (.A(WX7244), .B(II22121), .Z(II22122) ) ;
NAND2   gate15112  (.A(WX7308), .B(II22121), .Z(II22123) ) ;
NAND2   gate15113  (.A(II22122), .B(II22123), .Z(II22120) ) ;
NAND2   gate15114  (.A(II22104), .B(II22120), .Z(II22128) ) ;
NAND2   gate15115  (.A(II22104), .B(II22128), .Z(II22129) ) ;
NAND2   gate15116  (.A(II22120), .B(II22128), .Z(II22130) ) ;
NAND2   gate15117  (.A(WX7466), .B(WX7118), .Z(II22137) ) ;
NAND2   gate15118  (.A(WX7466), .B(II22137), .Z(II22138) ) ;
NAND2   gate15119  (.A(WX7118), .B(II22137), .Z(II22139) ) ;
NAND2   gate15120  (.A(II22138), .B(II22139), .Z(II22136) ) ;
NAND2   gate15121  (.A(WX7182), .B(II22136), .Z(II22144) ) ;
NAND2   gate15122  (.A(WX7182), .B(II22144), .Z(II22145) ) ;
NAND2   gate15123  (.A(II22136), .B(II22144), .Z(II22146) ) ;
NAND2   gate15124  (.A(II22145), .B(II22146), .Z(II22135) ) ;
NAND2   gate15125  (.A(WX7246), .B(WX7310), .Z(II22152) ) ;
NAND2   gate15126  (.A(WX7246), .B(II22152), .Z(II22153) ) ;
NAND2   gate15127  (.A(WX7310), .B(II22152), .Z(II22154) ) ;
NAND2   gate15128  (.A(II22153), .B(II22154), .Z(II22151) ) ;
NAND2   gate15129  (.A(II22135), .B(II22151), .Z(II22159) ) ;
NAND2   gate15130  (.A(II22135), .B(II22159), .Z(II22160) ) ;
NAND2   gate15131  (.A(II22151), .B(II22159), .Z(II22161) ) ;
NAND2   gate15132  (.A(WX7466), .B(WX7120), .Z(II22168) ) ;
NAND2   gate15133  (.A(WX7466), .B(II22168), .Z(II22169) ) ;
NAND2   gate15134  (.A(WX7120), .B(II22168), .Z(II22170) ) ;
NAND2   gate15135  (.A(II22169), .B(II22170), .Z(II22167) ) ;
NAND2   gate15136  (.A(WX7184), .B(II22167), .Z(II22175) ) ;
NAND2   gate15137  (.A(WX7184), .B(II22175), .Z(II22176) ) ;
NAND2   gate15138  (.A(II22167), .B(II22175), .Z(II22177) ) ;
NAND2   gate15139  (.A(II22176), .B(II22177), .Z(II22166) ) ;
NAND2   gate15140  (.A(WX7248), .B(WX7312), .Z(II22183) ) ;
NAND2   gate15141  (.A(WX7248), .B(II22183), .Z(II22184) ) ;
NAND2   gate15142  (.A(WX7312), .B(II22183), .Z(II22185) ) ;
NAND2   gate15143  (.A(II22184), .B(II22185), .Z(II22182) ) ;
NAND2   gate15144  (.A(II22166), .B(II22182), .Z(II22190) ) ;
NAND2   gate15145  (.A(II22166), .B(II22190), .Z(II22191) ) ;
NAND2   gate15146  (.A(II22182), .B(II22190), .Z(II22192) ) ;
NAND2   gate15147  (.A(WX7466), .B(WX7122), .Z(II22199) ) ;
NAND2   gate15148  (.A(WX7466), .B(II22199), .Z(II22200) ) ;
NAND2   gate15149  (.A(WX7122), .B(II22199), .Z(II22201) ) ;
NAND2   gate15150  (.A(II22200), .B(II22201), .Z(II22198) ) ;
NAND2   gate15151  (.A(WX7186), .B(II22198), .Z(II22206) ) ;
NAND2   gate15152  (.A(WX7186), .B(II22206), .Z(II22207) ) ;
NAND2   gate15153  (.A(II22198), .B(II22206), .Z(II22208) ) ;
NAND2   gate15154  (.A(II22207), .B(II22208), .Z(II22197) ) ;
NAND2   gate15155  (.A(WX7250), .B(WX7314), .Z(II22214) ) ;
NAND2   gate15156  (.A(WX7250), .B(II22214), .Z(II22215) ) ;
NAND2   gate15157  (.A(WX7314), .B(II22214), .Z(II22216) ) ;
NAND2   gate15158  (.A(II22215), .B(II22216), .Z(II22213) ) ;
NAND2   gate15159  (.A(II22197), .B(II22213), .Z(II22221) ) ;
NAND2   gate15160  (.A(II22197), .B(II22221), .Z(II22222) ) ;
NAND2   gate15161  (.A(II22213), .B(II22221), .Z(II22223) ) ;
NAND2   gate15162  (.A(WX7466), .B(WX7124), .Z(II22230) ) ;
NAND2   gate15163  (.A(WX7466), .B(II22230), .Z(II22231) ) ;
NAND2   gate15164  (.A(WX7124), .B(II22230), .Z(II22232) ) ;
NAND2   gate15165  (.A(II22231), .B(II22232), .Z(II22229) ) ;
NAND2   gate15166  (.A(WX7188), .B(II22229), .Z(II22237) ) ;
NAND2   gate15167  (.A(WX7188), .B(II22237), .Z(II22238) ) ;
NAND2   gate15168  (.A(II22229), .B(II22237), .Z(II22239) ) ;
NAND2   gate15169  (.A(II22238), .B(II22239), .Z(II22228) ) ;
NAND2   gate15170  (.A(WX7252), .B(WX7316), .Z(II22245) ) ;
NAND2   gate15171  (.A(WX7252), .B(II22245), .Z(II22246) ) ;
NAND2   gate15172  (.A(WX7316), .B(II22245), .Z(II22247) ) ;
NAND2   gate15173  (.A(II22246), .B(II22247), .Z(II22244) ) ;
NAND2   gate15174  (.A(II22228), .B(II22244), .Z(II22252) ) ;
NAND2   gate15175  (.A(II22228), .B(II22252), .Z(II22253) ) ;
NAND2   gate15176  (.A(II22244), .B(II22252), .Z(II22254) ) ;
NAND2   gate15177  (.A(WX7466), .B(WX7126), .Z(II22261) ) ;
NAND2   gate15178  (.A(WX7466), .B(II22261), .Z(II22262) ) ;
NAND2   gate15179  (.A(WX7126), .B(II22261), .Z(II22263) ) ;
NAND2   gate15180  (.A(II22262), .B(II22263), .Z(II22260) ) ;
NAND2   gate15181  (.A(WX7190), .B(II22260), .Z(II22268) ) ;
NAND2   gate15182  (.A(WX7190), .B(II22268), .Z(II22269) ) ;
NAND2   gate15183  (.A(II22260), .B(II22268), .Z(II22270) ) ;
NAND2   gate15184  (.A(II22269), .B(II22270), .Z(II22259) ) ;
NAND2   gate15185  (.A(WX7254), .B(WX7318), .Z(II22276) ) ;
NAND2   gate15186  (.A(WX7254), .B(II22276), .Z(II22277) ) ;
NAND2   gate15187  (.A(WX7318), .B(II22276), .Z(II22278) ) ;
NAND2   gate15188  (.A(II22277), .B(II22278), .Z(II22275) ) ;
NAND2   gate15189  (.A(II22259), .B(II22275), .Z(II22283) ) ;
NAND2   gate15190  (.A(II22259), .B(II22283), .Z(II22284) ) ;
NAND2   gate15191  (.A(II22275), .B(II22283), .Z(II22285) ) ;
NAND2   gate15192  (.A(WX7466), .B(WX7128), .Z(II22292) ) ;
NAND2   gate15193  (.A(WX7466), .B(II22292), .Z(II22293) ) ;
NAND2   gate15194  (.A(WX7128), .B(II22292), .Z(II22294) ) ;
NAND2   gate15195  (.A(II22293), .B(II22294), .Z(II22291) ) ;
NAND2   gate15196  (.A(WX7192), .B(II22291), .Z(II22299) ) ;
NAND2   gate15197  (.A(WX7192), .B(II22299), .Z(II22300) ) ;
NAND2   gate15198  (.A(II22291), .B(II22299), .Z(II22301) ) ;
NAND2   gate15199  (.A(II22300), .B(II22301), .Z(II22290) ) ;
NAND2   gate15200  (.A(WX7256), .B(WX7320), .Z(II22307) ) ;
NAND2   gate15201  (.A(WX7256), .B(II22307), .Z(II22308) ) ;
NAND2   gate15202  (.A(WX7320), .B(II22307), .Z(II22309) ) ;
NAND2   gate15203  (.A(II22308), .B(II22309), .Z(II22306) ) ;
NAND2   gate15204  (.A(II22290), .B(II22306), .Z(II22314) ) ;
NAND2   gate15205  (.A(II22290), .B(II22314), .Z(II22315) ) ;
NAND2   gate15206  (.A(II22306), .B(II22314), .Z(II22316) ) ;
NAND2   gate15207  (.A(WX7466), .B(WX7130), .Z(II22323) ) ;
NAND2   gate15208  (.A(WX7466), .B(II22323), .Z(II22324) ) ;
NAND2   gate15209  (.A(WX7130), .B(II22323), .Z(II22325) ) ;
NAND2   gate15210  (.A(II22324), .B(II22325), .Z(II22322) ) ;
NAND2   gate15211  (.A(WX7194), .B(II22322), .Z(II22330) ) ;
NAND2   gate15212  (.A(WX7194), .B(II22330), .Z(II22331) ) ;
NAND2   gate15213  (.A(II22322), .B(II22330), .Z(II22332) ) ;
NAND2   gate15214  (.A(II22331), .B(II22332), .Z(II22321) ) ;
NAND2   gate15215  (.A(WX7258), .B(WX7322), .Z(II22338) ) ;
NAND2   gate15216  (.A(WX7258), .B(II22338), .Z(II22339) ) ;
NAND2   gate15217  (.A(WX7322), .B(II22338), .Z(II22340) ) ;
NAND2   gate15218  (.A(II22339), .B(II22340), .Z(II22337) ) ;
NAND2   gate15219  (.A(II22321), .B(II22337), .Z(II22345) ) ;
NAND2   gate15220  (.A(II22321), .B(II22345), .Z(II22346) ) ;
NAND2   gate15221  (.A(II22337), .B(II22345), .Z(II22347) ) ;
NAND2   gate15222  (.A(WX7466), .B(WX7132), .Z(II22354) ) ;
NAND2   gate15223  (.A(WX7466), .B(II22354), .Z(II22355) ) ;
NAND2   gate15224  (.A(WX7132), .B(II22354), .Z(II22356) ) ;
NAND2   gate15225  (.A(II22355), .B(II22356), .Z(II22353) ) ;
NAND2   gate15226  (.A(WX7196), .B(II22353), .Z(II22361) ) ;
NAND2   gate15227  (.A(WX7196), .B(II22361), .Z(II22362) ) ;
NAND2   gate15228  (.A(II22353), .B(II22361), .Z(II22363) ) ;
NAND2   gate15229  (.A(II22362), .B(II22363), .Z(II22352) ) ;
NAND2   gate15230  (.A(WX7260), .B(WX7324), .Z(II22369) ) ;
NAND2   gate15231  (.A(WX7260), .B(II22369), .Z(II22370) ) ;
NAND2   gate15232  (.A(WX7324), .B(II22369), .Z(II22371) ) ;
NAND2   gate15233  (.A(II22370), .B(II22371), .Z(II22368) ) ;
NAND2   gate15234  (.A(II22352), .B(II22368), .Z(II22376) ) ;
NAND2   gate15235  (.A(II22352), .B(II22376), .Z(II22377) ) ;
NAND2   gate15236  (.A(II22368), .B(II22376), .Z(II22378) ) ;
NAND2   gate15237  (.A(WX7466), .B(WX7134), .Z(II22385) ) ;
NAND2   gate15238  (.A(WX7466), .B(II22385), .Z(II22386) ) ;
NAND2   gate15239  (.A(WX7134), .B(II22385), .Z(II22387) ) ;
NAND2   gate15240  (.A(II22386), .B(II22387), .Z(II22384) ) ;
NAND2   gate15241  (.A(WX7198), .B(II22384), .Z(II22392) ) ;
NAND2   gate15242  (.A(WX7198), .B(II22392), .Z(II22393) ) ;
NAND2   gate15243  (.A(II22384), .B(II22392), .Z(II22394) ) ;
NAND2   gate15244  (.A(II22393), .B(II22394), .Z(II22383) ) ;
NAND2   gate15245  (.A(WX7262), .B(WX7326), .Z(II22400) ) ;
NAND2   gate15246  (.A(WX7262), .B(II22400), .Z(II22401) ) ;
NAND2   gate15247  (.A(WX7326), .B(II22400), .Z(II22402) ) ;
NAND2   gate15248  (.A(II22401), .B(II22402), .Z(II22399) ) ;
NAND2   gate15249  (.A(II22383), .B(II22399), .Z(II22407) ) ;
NAND2   gate15250  (.A(II22383), .B(II22407), .Z(II22408) ) ;
NAND2   gate15251  (.A(II22399), .B(II22407), .Z(II22409) ) ;
NAND2   gate15252  (.A(WX7466), .B(WX7136), .Z(II22416) ) ;
NAND2   gate15253  (.A(WX7466), .B(II22416), .Z(II22417) ) ;
NAND2   gate15254  (.A(WX7136), .B(II22416), .Z(II22418) ) ;
NAND2   gate15255  (.A(II22417), .B(II22418), .Z(II22415) ) ;
NAND2   gate15256  (.A(WX7200), .B(II22415), .Z(II22423) ) ;
NAND2   gate15257  (.A(WX7200), .B(II22423), .Z(II22424) ) ;
NAND2   gate15258  (.A(II22415), .B(II22423), .Z(II22425) ) ;
NAND2   gate15259  (.A(II22424), .B(II22425), .Z(II22414) ) ;
NAND2   gate15260  (.A(WX7264), .B(WX7328), .Z(II22431) ) ;
NAND2   gate15261  (.A(WX7264), .B(II22431), .Z(II22432) ) ;
NAND2   gate15262  (.A(WX7328), .B(II22431), .Z(II22433) ) ;
NAND2   gate15263  (.A(II22432), .B(II22433), .Z(II22430) ) ;
NAND2   gate15264  (.A(II22414), .B(II22430), .Z(II22438) ) ;
NAND2   gate15265  (.A(II22414), .B(II22438), .Z(II22439) ) ;
NAND2   gate15266  (.A(II22430), .B(II22438), .Z(II22440) ) ;
NAND2   gate15267  (.A(WX7466), .B(WX7138), .Z(II22447) ) ;
NAND2   gate15268  (.A(WX7466), .B(II22447), .Z(II22448) ) ;
NAND2   gate15269  (.A(WX7138), .B(II22447), .Z(II22449) ) ;
NAND2   gate15270  (.A(II22448), .B(II22449), .Z(II22446) ) ;
NAND2   gate15271  (.A(WX7202), .B(II22446), .Z(II22454) ) ;
NAND2   gate15272  (.A(WX7202), .B(II22454), .Z(II22455) ) ;
NAND2   gate15273  (.A(II22446), .B(II22454), .Z(II22456) ) ;
NAND2   gate15274  (.A(II22455), .B(II22456), .Z(II22445) ) ;
NAND2   gate15275  (.A(WX7266), .B(WX7330), .Z(II22462) ) ;
NAND2   gate15276  (.A(WX7266), .B(II22462), .Z(II22463) ) ;
NAND2   gate15277  (.A(WX7330), .B(II22462), .Z(II22464) ) ;
NAND2   gate15278  (.A(II22463), .B(II22464), .Z(II22461) ) ;
NAND2   gate15279  (.A(II22445), .B(II22461), .Z(II22469) ) ;
NAND2   gate15280  (.A(II22445), .B(II22469), .Z(II22470) ) ;
NAND2   gate15281  (.A(II22461), .B(II22469), .Z(II22471) ) ;
NAND2   gate15282  (.A(WX7466), .B(WX7140), .Z(II22478) ) ;
NAND2   gate15283  (.A(WX7466), .B(II22478), .Z(II22479) ) ;
NAND2   gate15284  (.A(WX7140), .B(II22478), .Z(II22480) ) ;
NAND2   gate15285  (.A(II22479), .B(II22480), .Z(II22477) ) ;
NAND2   gate15286  (.A(WX7204), .B(II22477), .Z(II22485) ) ;
NAND2   gate15287  (.A(WX7204), .B(II22485), .Z(II22486) ) ;
NAND2   gate15288  (.A(II22477), .B(II22485), .Z(II22487) ) ;
NAND2   gate15289  (.A(II22486), .B(II22487), .Z(II22476) ) ;
NAND2   gate15290  (.A(WX7268), .B(WX7332), .Z(II22493) ) ;
NAND2   gate15291  (.A(WX7268), .B(II22493), .Z(II22494) ) ;
NAND2   gate15292  (.A(WX7332), .B(II22493), .Z(II22495) ) ;
NAND2   gate15293  (.A(II22494), .B(II22495), .Z(II22492) ) ;
NAND2   gate15294  (.A(II22476), .B(II22492), .Z(II22500) ) ;
NAND2   gate15295  (.A(II22476), .B(II22500), .Z(II22501) ) ;
NAND2   gate15296  (.A(II22492), .B(II22500), .Z(II22502) ) ;
NAND2   gate15297  (.A(WX7467), .B(WX7142), .Z(II22509) ) ;
NAND2   gate15298  (.A(WX7467), .B(II22509), .Z(II22510) ) ;
NAND2   gate15299  (.A(WX7142), .B(II22509), .Z(II22511) ) ;
NAND2   gate15300  (.A(II22510), .B(II22511), .Z(II22508) ) ;
NAND2   gate15301  (.A(WX7206), .B(II22508), .Z(II22516) ) ;
NAND2   gate15302  (.A(WX7206), .B(II22516), .Z(II22517) ) ;
NAND2   gate15303  (.A(II22508), .B(II22516), .Z(II22518) ) ;
NAND2   gate15304  (.A(II22517), .B(II22518), .Z(II22507) ) ;
NAND2   gate15305  (.A(WX7270), .B(WX7334), .Z(II22524) ) ;
NAND2   gate15306  (.A(WX7270), .B(II22524), .Z(II22525) ) ;
NAND2   gate15307  (.A(WX7334), .B(II22524), .Z(II22526) ) ;
NAND2   gate15308  (.A(II22525), .B(II22526), .Z(II22523) ) ;
NAND2   gate15309  (.A(II22507), .B(II22523), .Z(II22531) ) ;
NAND2   gate15310  (.A(II22507), .B(II22531), .Z(II22532) ) ;
NAND2   gate15311  (.A(II22523), .B(II22531), .Z(II22533) ) ;
NAND2   gate15312  (.A(WX7467), .B(WX7144), .Z(II22540) ) ;
NAND2   gate15313  (.A(WX7467), .B(II22540), .Z(II22541) ) ;
NAND2   gate15314  (.A(WX7144), .B(II22540), .Z(II22542) ) ;
NAND2   gate15315  (.A(II22541), .B(II22542), .Z(II22539) ) ;
NAND2   gate15316  (.A(WX7208), .B(II22539), .Z(II22547) ) ;
NAND2   gate15317  (.A(WX7208), .B(II22547), .Z(II22548) ) ;
NAND2   gate15318  (.A(II22539), .B(II22547), .Z(II22549) ) ;
NAND2   gate15319  (.A(II22548), .B(II22549), .Z(II22538) ) ;
NAND2   gate15320  (.A(WX7272), .B(WX7336), .Z(II22555) ) ;
NAND2   gate15321  (.A(WX7272), .B(II22555), .Z(II22556) ) ;
NAND2   gate15322  (.A(WX7336), .B(II22555), .Z(II22557) ) ;
NAND2   gate15323  (.A(II22556), .B(II22557), .Z(II22554) ) ;
NAND2   gate15324  (.A(II22538), .B(II22554), .Z(II22562) ) ;
NAND2   gate15325  (.A(II22538), .B(II22562), .Z(II22563) ) ;
NAND2   gate15326  (.A(II22554), .B(II22562), .Z(II22564) ) ;
NAND2   gate15327  (.A(WX7467), .B(WX7146), .Z(II22571) ) ;
NAND2   gate15328  (.A(WX7467), .B(II22571), .Z(II22572) ) ;
NAND2   gate15329  (.A(WX7146), .B(II22571), .Z(II22573) ) ;
NAND2   gate15330  (.A(II22572), .B(II22573), .Z(II22570) ) ;
NAND2   gate15331  (.A(WX7210), .B(II22570), .Z(II22578) ) ;
NAND2   gate15332  (.A(WX7210), .B(II22578), .Z(II22579) ) ;
NAND2   gate15333  (.A(II22570), .B(II22578), .Z(II22580) ) ;
NAND2   gate15334  (.A(II22579), .B(II22580), .Z(II22569) ) ;
NAND2   gate15335  (.A(WX7274), .B(WX7338), .Z(II22586) ) ;
NAND2   gate15336  (.A(WX7274), .B(II22586), .Z(II22587) ) ;
NAND2   gate15337  (.A(WX7338), .B(II22586), .Z(II22588) ) ;
NAND2   gate15338  (.A(II22587), .B(II22588), .Z(II22585) ) ;
NAND2   gate15339  (.A(II22569), .B(II22585), .Z(II22593) ) ;
NAND2   gate15340  (.A(II22569), .B(II22593), .Z(II22594) ) ;
NAND2   gate15341  (.A(II22585), .B(II22593), .Z(II22595) ) ;
NAND2   gate15342  (.A(WX7467), .B(WX7148), .Z(II22602) ) ;
NAND2   gate15343  (.A(WX7467), .B(II22602), .Z(II22603) ) ;
NAND2   gate15344  (.A(WX7148), .B(II22602), .Z(II22604) ) ;
NAND2   gate15345  (.A(II22603), .B(II22604), .Z(II22601) ) ;
NAND2   gate15346  (.A(WX7212), .B(II22601), .Z(II22609) ) ;
NAND2   gate15347  (.A(WX7212), .B(II22609), .Z(II22610) ) ;
NAND2   gate15348  (.A(II22601), .B(II22609), .Z(II22611) ) ;
NAND2   gate15349  (.A(II22610), .B(II22611), .Z(II22600) ) ;
NAND2   gate15350  (.A(WX7276), .B(WX7340), .Z(II22617) ) ;
NAND2   gate15351  (.A(WX7276), .B(II22617), .Z(II22618) ) ;
NAND2   gate15352  (.A(WX7340), .B(II22617), .Z(II22619) ) ;
NAND2   gate15353  (.A(II22618), .B(II22619), .Z(II22616) ) ;
NAND2   gate15354  (.A(II22600), .B(II22616), .Z(II22624) ) ;
NAND2   gate15355  (.A(II22600), .B(II22624), .Z(II22625) ) ;
NAND2   gate15356  (.A(II22616), .B(II22624), .Z(II22626) ) ;
NAND2   gate15357  (.A(WX7467), .B(WX7150), .Z(II22633) ) ;
NAND2   gate15358  (.A(WX7467), .B(II22633), .Z(II22634) ) ;
NAND2   gate15359  (.A(WX7150), .B(II22633), .Z(II22635) ) ;
NAND2   gate15360  (.A(II22634), .B(II22635), .Z(II22632) ) ;
NAND2   gate15361  (.A(WX7214), .B(II22632), .Z(II22640) ) ;
NAND2   gate15362  (.A(WX7214), .B(II22640), .Z(II22641) ) ;
NAND2   gate15363  (.A(II22632), .B(II22640), .Z(II22642) ) ;
NAND2   gate15364  (.A(II22641), .B(II22642), .Z(II22631) ) ;
NAND2   gate15365  (.A(WX7278), .B(WX7342), .Z(II22648) ) ;
NAND2   gate15366  (.A(WX7278), .B(II22648), .Z(II22649) ) ;
NAND2   gate15367  (.A(WX7342), .B(II22648), .Z(II22650) ) ;
NAND2   gate15368  (.A(II22649), .B(II22650), .Z(II22647) ) ;
NAND2   gate15369  (.A(II22631), .B(II22647), .Z(II22655) ) ;
NAND2   gate15370  (.A(II22631), .B(II22655), .Z(II22656) ) ;
NAND2   gate15371  (.A(II22647), .B(II22655), .Z(II22657) ) ;
NAND2   gate15372  (.A(WX7467), .B(WX7152), .Z(II22664) ) ;
NAND2   gate15373  (.A(WX7467), .B(II22664), .Z(II22665) ) ;
NAND2   gate15374  (.A(WX7152), .B(II22664), .Z(II22666) ) ;
NAND2   gate15375  (.A(II22665), .B(II22666), .Z(II22663) ) ;
NAND2   gate15376  (.A(WX7216), .B(II22663), .Z(II22671) ) ;
NAND2   gate15377  (.A(WX7216), .B(II22671), .Z(II22672) ) ;
NAND2   gate15378  (.A(II22663), .B(II22671), .Z(II22673) ) ;
NAND2   gate15379  (.A(II22672), .B(II22673), .Z(II22662) ) ;
NAND2   gate15380  (.A(WX7280), .B(WX7344), .Z(II22679) ) ;
NAND2   gate15381  (.A(WX7280), .B(II22679), .Z(II22680) ) ;
NAND2   gate15382  (.A(WX7344), .B(II22679), .Z(II22681) ) ;
NAND2   gate15383  (.A(II22680), .B(II22681), .Z(II22678) ) ;
NAND2   gate15384  (.A(II22662), .B(II22678), .Z(II22686) ) ;
NAND2   gate15385  (.A(II22662), .B(II22686), .Z(II22687) ) ;
NAND2   gate15386  (.A(II22678), .B(II22686), .Z(II22688) ) ;
NAND2   gate15387  (.A(WX7467), .B(WX7154), .Z(II22695) ) ;
NAND2   gate15388  (.A(WX7467), .B(II22695), .Z(II22696) ) ;
NAND2   gate15389  (.A(WX7154), .B(II22695), .Z(II22697) ) ;
NAND2   gate15390  (.A(II22696), .B(II22697), .Z(II22694) ) ;
NAND2   gate15391  (.A(WX7218), .B(II22694), .Z(II22702) ) ;
NAND2   gate15392  (.A(WX7218), .B(II22702), .Z(II22703) ) ;
NAND2   gate15393  (.A(II22694), .B(II22702), .Z(II22704) ) ;
NAND2   gate15394  (.A(II22703), .B(II22704), .Z(II22693) ) ;
NAND2   gate15395  (.A(WX7282), .B(WX7346), .Z(II22710) ) ;
NAND2   gate15396  (.A(WX7282), .B(II22710), .Z(II22711) ) ;
NAND2   gate15397  (.A(WX7346), .B(II22710), .Z(II22712) ) ;
NAND2   gate15398  (.A(II22711), .B(II22712), .Z(II22709) ) ;
NAND2   gate15399  (.A(II22693), .B(II22709), .Z(II22717) ) ;
NAND2   gate15400  (.A(II22693), .B(II22717), .Z(II22718) ) ;
NAND2   gate15401  (.A(II22709), .B(II22717), .Z(II22719) ) ;
NAND2   gate15402  (.A(WX7467), .B(WX7156), .Z(II22726) ) ;
NAND2   gate15403  (.A(WX7467), .B(II22726), .Z(II22727) ) ;
NAND2   gate15404  (.A(WX7156), .B(II22726), .Z(II22728) ) ;
NAND2   gate15405  (.A(II22727), .B(II22728), .Z(II22725) ) ;
NAND2   gate15406  (.A(WX7220), .B(II22725), .Z(II22733) ) ;
NAND2   gate15407  (.A(WX7220), .B(II22733), .Z(II22734) ) ;
NAND2   gate15408  (.A(II22725), .B(II22733), .Z(II22735) ) ;
NAND2   gate15409  (.A(II22734), .B(II22735), .Z(II22724) ) ;
NAND2   gate15410  (.A(WX7284), .B(WX7348), .Z(II22741) ) ;
NAND2   gate15411  (.A(WX7284), .B(II22741), .Z(II22742) ) ;
NAND2   gate15412  (.A(WX7348), .B(II22741), .Z(II22743) ) ;
NAND2   gate15413  (.A(II22742), .B(II22743), .Z(II22740) ) ;
NAND2   gate15414  (.A(II22724), .B(II22740), .Z(II22748) ) ;
NAND2   gate15415  (.A(II22724), .B(II22748), .Z(II22749) ) ;
NAND2   gate15416  (.A(II22740), .B(II22748), .Z(II22750) ) ;
NAND2   gate15417  (.A(WX7467), .B(WX7158), .Z(II22757) ) ;
NAND2   gate15418  (.A(WX7467), .B(II22757), .Z(II22758) ) ;
NAND2   gate15419  (.A(WX7158), .B(II22757), .Z(II22759) ) ;
NAND2   gate15420  (.A(II22758), .B(II22759), .Z(II22756) ) ;
NAND2   gate15421  (.A(WX7222), .B(II22756), .Z(II22764) ) ;
NAND2   gate15422  (.A(WX7222), .B(II22764), .Z(II22765) ) ;
NAND2   gate15423  (.A(II22756), .B(II22764), .Z(II22766) ) ;
NAND2   gate15424  (.A(II22765), .B(II22766), .Z(II22755) ) ;
NAND2   gate15425  (.A(WX7286), .B(WX7350), .Z(II22772) ) ;
NAND2   gate15426  (.A(WX7286), .B(II22772), .Z(II22773) ) ;
NAND2   gate15427  (.A(WX7350), .B(II22772), .Z(II22774) ) ;
NAND2   gate15428  (.A(II22773), .B(II22774), .Z(II22771) ) ;
NAND2   gate15429  (.A(II22755), .B(II22771), .Z(II22779) ) ;
NAND2   gate15430  (.A(II22755), .B(II22779), .Z(II22780) ) ;
NAND2   gate15431  (.A(II22771), .B(II22779), .Z(II22781) ) ;
NAND2   gate15432  (.A(WX7467), .B(WX7160), .Z(II22788) ) ;
NAND2   gate15433  (.A(WX7467), .B(II22788), .Z(II22789) ) ;
NAND2   gate15434  (.A(WX7160), .B(II22788), .Z(II22790) ) ;
NAND2   gate15435  (.A(II22789), .B(II22790), .Z(II22787) ) ;
NAND2   gate15436  (.A(WX7224), .B(II22787), .Z(II22795) ) ;
NAND2   gate15437  (.A(WX7224), .B(II22795), .Z(II22796) ) ;
NAND2   gate15438  (.A(II22787), .B(II22795), .Z(II22797) ) ;
NAND2   gate15439  (.A(II22796), .B(II22797), .Z(II22786) ) ;
NAND2   gate15440  (.A(WX7288), .B(WX7352), .Z(II22803) ) ;
NAND2   gate15441  (.A(WX7288), .B(II22803), .Z(II22804) ) ;
NAND2   gate15442  (.A(WX7352), .B(II22803), .Z(II22805) ) ;
NAND2   gate15443  (.A(II22804), .B(II22805), .Z(II22802) ) ;
NAND2   gate15444  (.A(II22786), .B(II22802), .Z(II22810) ) ;
NAND2   gate15445  (.A(II22786), .B(II22810), .Z(II22811) ) ;
NAND2   gate15446  (.A(II22802), .B(II22810), .Z(II22812) ) ;
NAND2   gate15447  (.A(WX7467), .B(WX7162), .Z(II22819) ) ;
NAND2   gate15448  (.A(WX7467), .B(II22819), .Z(II22820) ) ;
NAND2   gate15449  (.A(WX7162), .B(II22819), .Z(II22821) ) ;
NAND2   gate15450  (.A(II22820), .B(II22821), .Z(II22818) ) ;
NAND2   gate15451  (.A(WX7226), .B(II22818), .Z(II22826) ) ;
NAND2   gate15452  (.A(WX7226), .B(II22826), .Z(II22827) ) ;
NAND2   gate15453  (.A(II22818), .B(II22826), .Z(II22828) ) ;
NAND2   gate15454  (.A(II22827), .B(II22828), .Z(II22817) ) ;
NAND2   gate15455  (.A(WX7290), .B(WX7354), .Z(II22834) ) ;
NAND2   gate15456  (.A(WX7290), .B(II22834), .Z(II22835) ) ;
NAND2   gate15457  (.A(WX7354), .B(II22834), .Z(II22836) ) ;
NAND2   gate15458  (.A(II22835), .B(II22836), .Z(II22833) ) ;
NAND2   gate15459  (.A(II22817), .B(II22833), .Z(II22841) ) ;
NAND2   gate15460  (.A(II22817), .B(II22841), .Z(II22842) ) ;
NAND2   gate15461  (.A(II22833), .B(II22841), .Z(II22843) ) ;
NAND2   gate15462  (.A(WX7467), .B(WX7164), .Z(II22850) ) ;
NAND2   gate15463  (.A(WX7467), .B(II22850), .Z(II22851) ) ;
NAND2   gate15464  (.A(WX7164), .B(II22850), .Z(II22852) ) ;
NAND2   gate15465  (.A(II22851), .B(II22852), .Z(II22849) ) ;
NAND2   gate15466  (.A(WX7228), .B(II22849), .Z(II22857) ) ;
NAND2   gate15467  (.A(WX7228), .B(II22857), .Z(II22858) ) ;
NAND2   gate15468  (.A(II22849), .B(II22857), .Z(II22859) ) ;
NAND2   gate15469  (.A(II22858), .B(II22859), .Z(II22848) ) ;
NAND2   gate15470  (.A(WX7292), .B(WX7356), .Z(II22865) ) ;
NAND2   gate15471  (.A(WX7292), .B(II22865), .Z(II22866) ) ;
NAND2   gate15472  (.A(WX7356), .B(II22865), .Z(II22867) ) ;
NAND2   gate15473  (.A(II22866), .B(II22867), .Z(II22864) ) ;
NAND2   gate15474  (.A(II22848), .B(II22864), .Z(II22872) ) ;
NAND2   gate15475  (.A(II22848), .B(II22872), .Z(II22873) ) ;
NAND2   gate15476  (.A(II22864), .B(II22872), .Z(II22874) ) ;
NAND2   gate15477  (.A(WX7467), .B(WX7166), .Z(II22881) ) ;
NAND2   gate15478  (.A(WX7467), .B(II22881), .Z(II22882) ) ;
NAND2   gate15479  (.A(WX7166), .B(II22881), .Z(II22883) ) ;
NAND2   gate15480  (.A(II22882), .B(II22883), .Z(II22880) ) ;
NAND2   gate15481  (.A(WX7230), .B(II22880), .Z(II22888) ) ;
NAND2   gate15482  (.A(WX7230), .B(II22888), .Z(II22889) ) ;
NAND2   gate15483  (.A(II22880), .B(II22888), .Z(II22890) ) ;
NAND2   gate15484  (.A(II22889), .B(II22890), .Z(II22879) ) ;
NAND2   gate15485  (.A(WX7294), .B(WX7358), .Z(II22896) ) ;
NAND2   gate15486  (.A(WX7294), .B(II22896), .Z(II22897) ) ;
NAND2   gate15487  (.A(WX7358), .B(II22896), .Z(II22898) ) ;
NAND2   gate15488  (.A(II22897), .B(II22898), .Z(II22895) ) ;
NAND2   gate15489  (.A(II22879), .B(II22895), .Z(II22903) ) ;
NAND2   gate15490  (.A(II22879), .B(II22903), .Z(II22904) ) ;
NAND2   gate15491  (.A(II22895), .B(II22903), .Z(II22905) ) ;
NAND2   gate15492  (.A(WX7467), .B(WX7168), .Z(II22912) ) ;
NAND2   gate15493  (.A(WX7467), .B(II22912), .Z(II22913) ) ;
NAND2   gate15494  (.A(WX7168), .B(II22912), .Z(II22914) ) ;
NAND2   gate15495  (.A(II22913), .B(II22914), .Z(II22911) ) ;
NAND2   gate15496  (.A(WX7232), .B(II22911), .Z(II22919) ) ;
NAND2   gate15497  (.A(WX7232), .B(II22919), .Z(II22920) ) ;
NAND2   gate15498  (.A(II22911), .B(II22919), .Z(II22921) ) ;
NAND2   gate15499  (.A(II22920), .B(II22921), .Z(II22910) ) ;
NAND2   gate15500  (.A(WX7296), .B(WX7360), .Z(II22927) ) ;
NAND2   gate15501  (.A(WX7296), .B(II22927), .Z(II22928) ) ;
NAND2   gate15502  (.A(WX7360), .B(II22927), .Z(II22929) ) ;
NAND2   gate15503  (.A(II22928), .B(II22929), .Z(II22926) ) ;
NAND2   gate15504  (.A(II22910), .B(II22926), .Z(II22934) ) ;
NAND2   gate15505  (.A(II22910), .B(II22934), .Z(II22935) ) ;
NAND2   gate15506  (.A(II22926), .B(II22934), .Z(II22936) ) ;
NAND2   gate15507  (.A(WX7467), .B(WX7170), .Z(II22943) ) ;
NAND2   gate15508  (.A(WX7467), .B(II22943), .Z(II22944) ) ;
NAND2   gate15509  (.A(WX7170), .B(II22943), .Z(II22945) ) ;
NAND2   gate15510  (.A(II22944), .B(II22945), .Z(II22942) ) ;
NAND2   gate15511  (.A(WX7234), .B(II22942), .Z(II22950) ) ;
NAND2   gate15512  (.A(WX7234), .B(II22950), .Z(II22951) ) ;
NAND2   gate15513  (.A(II22942), .B(II22950), .Z(II22952) ) ;
NAND2   gate15514  (.A(II22951), .B(II22952), .Z(II22941) ) ;
NAND2   gate15515  (.A(WX7298), .B(WX7362), .Z(II22958) ) ;
NAND2   gate15516  (.A(WX7298), .B(II22958), .Z(II22959) ) ;
NAND2   gate15517  (.A(WX7362), .B(II22958), .Z(II22960) ) ;
NAND2   gate15518  (.A(II22959), .B(II22960), .Z(II22957) ) ;
NAND2   gate15519  (.A(II22941), .B(II22957), .Z(II22965) ) ;
NAND2   gate15520  (.A(II22941), .B(II22965), .Z(II22966) ) ;
NAND2   gate15521  (.A(II22957), .B(II22965), .Z(II22967) ) ;
NAND2   gate15522  (.A(WX7467), .B(WX7172), .Z(II22974) ) ;
NAND2   gate15523  (.A(WX7467), .B(II22974), .Z(II22975) ) ;
NAND2   gate15524  (.A(WX7172), .B(II22974), .Z(II22976) ) ;
NAND2   gate15525  (.A(II22975), .B(II22976), .Z(II22973) ) ;
NAND2   gate15526  (.A(WX7236), .B(II22973), .Z(II22981) ) ;
NAND2   gate15527  (.A(WX7236), .B(II22981), .Z(II22982) ) ;
NAND2   gate15528  (.A(II22973), .B(II22981), .Z(II22983) ) ;
NAND2   gate15529  (.A(II22982), .B(II22983), .Z(II22972) ) ;
NAND2   gate15530  (.A(WX7300), .B(WX7364), .Z(II22989) ) ;
NAND2   gate15531  (.A(WX7300), .B(II22989), .Z(II22990) ) ;
NAND2   gate15532  (.A(WX7364), .B(II22989), .Z(II22991) ) ;
NAND2   gate15533  (.A(II22990), .B(II22991), .Z(II22988) ) ;
NAND2   gate15534  (.A(II22972), .B(II22988), .Z(II22996) ) ;
NAND2   gate15535  (.A(II22972), .B(II22996), .Z(II22997) ) ;
NAND2   gate15536  (.A(II22988), .B(II22996), .Z(II22998) ) ;
NAND2   gate15537  (.A(WX7045), .B(WX6950), .Z(II23077) ) ;
NAND2   gate15538  (.A(WX7045), .B(II23077), .Z(II23078) ) ;
NAND2   gate15539  (.A(WX6950), .B(II23077), .Z(II23079) ) ;
NAND2   gate15540  (.A(WX7046), .B(WX6952), .Z(II23090) ) ;
NAND2   gate15541  (.A(WX7046), .B(II23090), .Z(II23091) ) ;
NAND2   gate15542  (.A(WX6952), .B(II23090), .Z(II23092) ) ;
NAND2   gate15543  (.A(WX7047), .B(WX6954), .Z(II23103) ) ;
NAND2   gate15544  (.A(WX7047), .B(II23103), .Z(II23104) ) ;
NAND2   gate15545  (.A(WX6954), .B(II23103), .Z(II23105) ) ;
NAND2   gate15546  (.A(WX7048), .B(WX6956), .Z(II23116) ) ;
NAND2   gate15547  (.A(WX7048), .B(II23116), .Z(II23117) ) ;
NAND2   gate15548  (.A(WX6956), .B(II23116), .Z(II23118) ) ;
NAND2   gate15549  (.A(WX7049), .B(WX6958), .Z(II23129) ) ;
NAND2   gate15550  (.A(WX7049), .B(II23129), .Z(II23130) ) ;
NAND2   gate15551  (.A(WX6958), .B(II23129), .Z(II23131) ) ;
NAND2   gate15552  (.A(WX7050), .B(WX6960), .Z(II23142) ) ;
NAND2   gate15553  (.A(WX7050), .B(II23142), .Z(II23143) ) ;
NAND2   gate15554  (.A(WX6960), .B(II23142), .Z(II23144) ) ;
NAND2   gate15555  (.A(WX7051), .B(WX6962), .Z(II23155) ) ;
NAND2   gate15556  (.A(WX7051), .B(II23155), .Z(II23156) ) ;
NAND2   gate15557  (.A(WX6962), .B(II23155), .Z(II23157) ) ;
NAND2   gate15558  (.A(WX7052), .B(WX6964), .Z(II23168) ) ;
NAND2   gate15559  (.A(WX7052), .B(II23168), .Z(II23169) ) ;
NAND2   gate15560  (.A(WX6964), .B(II23168), .Z(II23170) ) ;
NAND2   gate15561  (.A(WX7053), .B(WX6966), .Z(II23181) ) ;
NAND2   gate15562  (.A(WX7053), .B(II23181), .Z(II23182) ) ;
NAND2   gate15563  (.A(WX6966), .B(II23181), .Z(II23183) ) ;
NAND2   gate15564  (.A(WX7054), .B(WX6968), .Z(II23194) ) ;
NAND2   gate15565  (.A(WX7054), .B(II23194), .Z(II23195) ) ;
NAND2   gate15566  (.A(WX6968), .B(II23194), .Z(II23196) ) ;
NAND2   gate15567  (.A(WX7055), .B(WX6970), .Z(II23207) ) ;
NAND2   gate15568  (.A(WX7055), .B(II23207), .Z(II23208) ) ;
NAND2   gate15569  (.A(WX6970), .B(II23207), .Z(II23209) ) ;
NAND2   gate15570  (.A(WX7056), .B(WX6972), .Z(II23220) ) ;
NAND2   gate15571  (.A(WX7056), .B(II23220), .Z(II23221) ) ;
NAND2   gate15572  (.A(WX6972), .B(II23220), .Z(II23222) ) ;
NAND2   gate15573  (.A(WX7057), .B(WX6974), .Z(II23233) ) ;
NAND2   gate15574  (.A(WX7057), .B(II23233), .Z(II23234) ) ;
NAND2   gate15575  (.A(WX6974), .B(II23233), .Z(II23235) ) ;
NAND2   gate15576  (.A(WX7058), .B(WX6976), .Z(II23246) ) ;
NAND2   gate15577  (.A(WX7058), .B(II23246), .Z(II23247) ) ;
NAND2   gate15578  (.A(WX6976), .B(II23246), .Z(II23248) ) ;
NAND2   gate15579  (.A(WX7059), .B(WX6978), .Z(II23259) ) ;
NAND2   gate15580  (.A(WX7059), .B(II23259), .Z(II23260) ) ;
NAND2   gate15581  (.A(WX6978), .B(II23259), .Z(II23261) ) ;
NAND2   gate15582  (.A(WX7060), .B(WX6980), .Z(II23272) ) ;
NAND2   gate15583  (.A(WX7060), .B(II23272), .Z(II23273) ) ;
NAND2   gate15584  (.A(WX6980), .B(II23272), .Z(II23274) ) ;
NAND2   gate15585  (.A(WX7061), .B(WX6982), .Z(II23285) ) ;
NAND2   gate15586  (.A(WX7061), .B(II23285), .Z(II23286) ) ;
NAND2   gate15587  (.A(WX6982), .B(II23285), .Z(II23287) ) ;
NAND2   gate15588  (.A(WX7062), .B(WX6984), .Z(II23298) ) ;
NAND2   gate15589  (.A(WX7062), .B(II23298), .Z(II23299) ) ;
NAND2   gate15590  (.A(WX6984), .B(II23298), .Z(II23300) ) ;
NAND2   gate15591  (.A(WX7063), .B(WX6986), .Z(II23311) ) ;
NAND2   gate15592  (.A(WX7063), .B(II23311), .Z(II23312) ) ;
NAND2   gate15593  (.A(WX6986), .B(II23311), .Z(II23313) ) ;
NAND2   gate15594  (.A(WX7064), .B(WX6988), .Z(II23324) ) ;
NAND2   gate15595  (.A(WX7064), .B(II23324), .Z(II23325) ) ;
NAND2   gate15596  (.A(WX6988), .B(II23324), .Z(II23326) ) ;
NAND2   gate15597  (.A(WX7065), .B(WX6990), .Z(II23337) ) ;
NAND2   gate15598  (.A(WX7065), .B(II23337), .Z(II23338) ) ;
NAND2   gate15599  (.A(WX6990), .B(II23337), .Z(II23339) ) ;
NAND2   gate15600  (.A(WX7066), .B(WX6992), .Z(II23350) ) ;
NAND2   gate15601  (.A(WX7066), .B(II23350), .Z(II23351) ) ;
NAND2   gate15602  (.A(WX6992), .B(II23350), .Z(II23352) ) ;
NAND2   gate15603  (.A(WX7067), .B(WX6994), .Z(II23363) ) ;
NAND2   gate15604  (.A(WX7067), .B(II23363), .Z(II23364) ) ;
NAND2   gate15605  (.A(WX6994), .B(II23363), .Z(II23365) ) ;
NAND2   gate15606  (.A(WX7068), .B(WX6996), .Z(II23376) ) ;
NAND2   gate15607  (.A(WX7068), .B(II23376), .Z(II23377) ) ;
NAND2   gate15608  (.A(WX6996), .B(II23376), .Z(II23378) ) ;
NAND2   gate15609  (.A(WX7069), .B(WX6998), .Z(II23389) ) ;
NAND2   gate15610  (.A(WX7069), .B(II23389), .Z(II23390) ) ;
NAND2   gate15611  (.A(WX6998), .B(II23389), .Z(II23391) ) ;
NAND2   gate15612  (.A(WX7070), .B(WX7000), .Z(II23402) ) ;
NAND2   gate15613  (.A(WX7070), .B(II23402), .Z(II23403) ) ;
NAND2   gate15614  (.A(WX7000), .B(II23402), .Z(II23404) ) ;
NAND2   gate15615  (.A(WX7071), .B(WX7002), .Z(II23415) ) ;
NAND2   gate15616  (.A(WX7071), .B(II23415), .Z(II23416) ) ;
NAND2   gate15617  (.A(WX7002), .B(II23415), .Z(II23417) ) ;
NAND2   gate15618  (.A(WX7072), .B(WX7004), .Z(II23428) ) ;
NAND2   gate15619  (.A(WX7072), .B(II23428), .Z(II23429) ) ;
NAND2   gate15620  (.A(WX7004), .B(II23428), .Z(II23430) ) ;
NAND2   gate15621  (.A(WX7073), .B(WX7006), .Z(II23441) ) ;
NAND2   gate15622  (.A(WX7073), .B(II23441), .Z(II23442) ) ;
NAND2   gate15623  (.A(WX7006), .B(II23441), .Z(II23443) ) ;
NAND2   gate15624  (.A(WX7074), .B(WX7008), .Z(II23454) ) ;
NAND2   gate15625  (.A(WX7074), .B(II23454), .Z(II23455) ) ;
NAND2   gate15626  (.A(WX7008), .B(II23454), .Z(II23456) ) ;
NAND2   gate15627  (.A(WX7075), .B(WX7010), .Z(II23467) ) ;
NAND2   gate15628  (.A(WX7075), .B(II23467), .Z(II23468) ) ;
NAND2   gate15629  (.A(WX7010), .B(II23467), .Z(II23469) ) ;
NAND2   gate15630  (.A(WX7076), .B(WX7012), .Z(II23480) ) ;
NAND2   gate15631  (.A(WX7076), .B(II23480), .Z(II23481) ) ;
NAND2   gate15632  (.A(WX7012), .B(II23480), .Z(II23482) ) ;
NAND2   gate15633  (.A(WX7092), .B(CRC_OUT_4_31), .Z(II23495) ) ;
NAND2   gate15634  (.A(WX7092), .B(II23495), .Z(II23496) ) ;
NAND2   gate15635  (.A(CRC_OUT_4_31), .B(II23495), .Z(II23497) ) ;
NAND2   gate15636  (.A(II23496), .B(II23497), .Z(II23494) ) ;
NAND2   gate15637  (.A(CRC_OUT_4_15), .B(II23494), .Z(II23502) ) ;
NAND2   gate15638  (.A(CRC_OUT_4_15), .B(II23502), .Z(II23503) ) ;
NAND2   gate15639  (.A(II23494), .B(II23502), .Z(II23504) ) ;
NAND2   gate15640  (.A(WX7097), .B(CRC_OUT_4_31), .Z(II23510) ) ;
NAND2   gate15641  (.A(WX7097), .B(II23510), .Z(II23511) ) ;
NAND2   gate15642  (.A(CRC_OUT_4_31), .B(II23510), .Z(II23512) ) ;
NAND2   gate15643  (.A(II23511), .B(II23512), .Z(II23509) ) ;
NAND2   gate15644  (.A(CRC_OUT_4_10), .B(II23509), .Z(II23517) ) ;
NAND2   gate15645  (.A(CRC_OUT_4_10), .B(II23517), .Z(II23518) ) ;
NAND2   gate15646  (.A(II23509), .B(II23517), .Z(II23519) ) ;
NAND2   gate15647  (.A(WX7104), .B(CRC_OUT_4_31), .Z(II23525) ) ;
NAND2   gate15648  (.A(WX7104), .B(II23525), .Z(II23526) ) ;
NAND2   gate15649  (.A(CRC_OUT_4_31), .B(II23525), .Z(II23527) ) ;
NAND2   gate15650  (.A(II23526), .B(II23527), .Z(II23524) ) ;
NAND2   gate15651  (.A(CRC_OUT_4_3), .B(II23524), .Z(II23532) ) ;
NAND2   gate15652  (.A(CRC_OUT_4_3), .B(II23532), .Z(II23533) ) ;
NAND2   gate15653  (.A(II23524), .B(II23532), .Z(II23534) ) ;
NAND2   gate15654  (.A(WX7108), .B(CRC_OUT_4_31), .Z(II23539) ) ;
NAND2   gate15655  (.A(WX7108), .B(II23539), .Z(II23540) ) ;
NAND2   gate15656  (.A(CRC_OUT_4_31), .B(II23539), .Z(II23541) ) ;
NAND2   gate15657  (.A(WX7077), .B(CRC_OUT_4_30), .Z(II23546) ) ;
NAND2   gate15658  (.A(WX7077), .B(II23546), .Z(II23547) ) ;
NAND2   gate15659  (.A(CRC_OUT_4_30), .B(II23546), .Z(II23548) ) ;
NAND2   gate15660  (.A(WX7078), .B(CRC_OUT_4_29), .Z(II23553) ) ;
NAND2   gate15661  (.A(WX7078), .B(II23553), .Z(II23554) ) ;
NAND2   gate15662  (.A(CRC_OUT_4_29), .B(II23553), .Z(II23555) ) ;
NAND2   gate15663  (.A(WX7079), .B(CRC_OUT_4_28), .Z(II23560) ) ;
NAND2   gate15664  (.A(WX7079), .B(II23560), .Z(II23561) ) ;
NAND2   gate15665  (.A(CRC_OUT_4_28), .B(II23560), .Z(II23562) ) ;
NAND2   gate15666  (.A(WX7080), .B(CRC_OUT_4_27), .Z(II23567) ) ;
NAND2   gate15667  (.A(WX7080), .B(II23567), .Z(II23568) ) ;
NAND2   gate15668  (.A(CRC_OUT_4_27), .B(II23567), .Z(II23569) ) ;
NAND2   gate15669  (.A(WX7081), .B(CRC_OUT_4_26), .Z(II23574) ) ;
NAND2   gate15670  (.A(WX7081), .B(II23574), .Z(II23575) ) ;
NAND2   gate15671  (.A(CRC_OUT_4_26), .B(II23574), .Z(II23576) ) ;
NAND2   gate15672  (.A(WX7082), .B(CRC_OUT_4_25), .Z(II23581) ) ;
NAND2   gate15673  (.A(WX7082), .B(II23581), .Z(II23582) ) ;
NAND2   gate15674  (.A(CRC_OUT_4_25), .B(II23581), .Z(II23583) ) ;
NAND2   gate15675  (.A(WX7083), .B(CRC_OUT_4_24), .Z(II23588) ) ;
NAND2   gate15676  (.A(WX7083), .B(II23588), .Z(II23589) ) ;
NAND2   gate15677  (.A(CRC_OUT_4_24), .B(II23588), .Z(II23590) ) ;
NAND2   gate15678  (.A(WX7084), .B(CRC_OUT_4_23), .Z(II23595) ) ;
NAND2   gate15679  (.A(WX7084), .B(II23595), .Z(II23596) ) ;
NAND2   gate15680  (.A(CRC_OUT_4_23), .B(II23595), .Z(II23597) ) ;
NAND2   gate15681  (.A(WX7085), .B(CRC_OUT_4_22), .Z(II23602) ) ;
NAND2   gate15682  (.A(WX7085), .B(II23602), .Z(II23603) ) ;
NAND2   gate15683  (.A(CRC_OUT_4_22), .B(II23602), .Z(II23604) ) ;
NAND2   gate15684  (.A(WX7086), .B(CRC_OUT_4_21), .Z(II23609) ) ;
NAND2   gate15685  (.A(WX7086), .B(II23609), .Z(II23610) ) ;
NAND2   gate15686  (.A(CRC_OUT_4_21), .B(II23609), .Z(II23611) ) ;
NAND2   gate15687  (.A(WX7087), .B(CRC_OUT_4_20), .Z(II23616) ) ;
NAND2   gate15688  (.A(WX7087), .B(II23616), .Z(II23617) ) ;
NAND2   gate15689  (.A(CRC_OUT_4_20), .B(II23616), .Z(II23618) ) ;
NAND2   gate15690  (.A(WX7088), .B(CRC_OUT_4_19), .Z(II23623) ) ;
NAND2   gate15691  (.A(WX7088), .B(II23623), .Z(II23624) ) ;
NAND2   gate15692  (.A(CRC_OUT_4_19), .B(II23623), .Z(II23625) ) ;
NAND2   gate15693  (.A(WX7089), .B(CRC_OUT_4_18), .Z(II23630) ) ;
NAND2   gate15694  (.A(WX7089), .B(II23630), .Z(II23631) ) ;
NAND2   gate15695  (.A(CRC_OUT_4_18), .B(II23630), .Z(II23632) ) ;
NAND2   gate15696  (.A(WX7090), .B(CRC_OUT_4_17), .Z(II23637) ) ;
NAND2   gate15697  (.A(WX7090), .B(II23637), .Z(II23638) ) ;
NAND2   gate15698  (.A(CRC_OUT_4_17), .B(II23637), .Z(II23639) ) ;
NAND2   gate15699  (.A(WX7091), .B(CRC_OUT_4_16), .Z(II23644) ) ;
NAND2   gate15700  (.A(WX7091), .B(II23644), .Z(II23645) ) ;
NAND2   gate15701  (.A(CRC_OUT_4_16), .B(II23644), .Z(II23646) ) ;
NAND2   gate15702  (.A(WX7093), .B(CRC_OUT_4_14), .Z(II23651) ) ;
NAND2   gate15703  (.A(WX7093), .B(II23651), .Z(II23652) ) ;
NAND2   gate15704  (.A(CRC_OUT_4_14), .B(II23651), .Z(II23653) ) ;
NAND2   gate15705  (.A(WX7094), .B(CRC_OUT_4_13), .Z(II23658) ) ;
NAND2   gate15706  (.A(WX7094), .B(II23658), .Z(II23659) ) ;
NAND2   gate15707  (.A(CRC_OUT_4_13), .B(II23658), .Z(II23660) ) ;
NAND2   gate15708  (.A(WX7095), .B(CRC_OUT_4_12), .Z(II23665) ) ;
NAND2   gate15709  (.A(WX7095), .B(II23665), .Z(II23666) ) ;
NAND2   gate15710  (.A(CRC_OUT_4_12), .B(II23665), .Z(II23667) ) ;
NAND2   gate15711  (.A(WX7096), .B(CRC_OUT_4_11), .Z(II23672) ) ;
NAND2   gate15712  (.A(WX7096), .B(II23672), .Z(II23673) ) ;
NAND2   gate15713  (.A(CRC_OUT_4_11), .B(II23672), .Z(II23674) ) ;
NAND2   gate15714  (.A(WX7098), .B(CRC_OUT_4_9), .Z(II23679) ) ;
NAND2   gate15715  (.A(WX7098), .B(II23679), .Z(II23680) ) ;
NAND2   gate15716  (.A(CRC_OUT_4_9), .B(II23679), .Z(II23681) ) ;
NAND2   gate15717  (.A(WX7099), .B(CRC_OUT_4_8), .Z(II23686) ) ;
NAND2   gate15718  (.A(WX7099), .B(II23686), .Z(II23687) ) ;
NAND2   gate15719  (.A(CRC_OUT_4_8), .B(II23686), .Z(II23688) ) ;
NAND2   gate15720  (.A(WX7100), .B(CRC_OUT_4_7), .Z(II23693) ) ;
NAND2   gate15721  (.A(WX7100), .B(II23693), .Z(II23694) ) ;
NAND2   gate15722  (.A(CRC_OUT_4_7), .B(II23693), .Z(II23695) ) ;
NAND2   gate15723  (.A(WX7101), .B(CRC_OUT_4_6), .Z(II23700) ) ;
NAND2   gate15724  (.A(WX7101), .B(II23700), .Z(II23701) ) ;
NAND2   gate15725  (.A(CRC_OUT_4_6), .B(II23700), .Z(II23702) ) ;
NAND2   gate15726  (.A(WX7102), .B(CRC_OUT_4_5), .Z(II23707) ) ;
NAND2   gate15727  (.A(WX7102), .B(II23707), .Z(II23708) ) ;
NAND2   gate15728  (.A(CRC_OUT_4_5), .B(II23707), .Z(II23709) ) ;
NAND2   gate15729  (.A(WX7103), .B(CRC_OUT_4_4), .Z(II23714) ) ;
NAND2   gate15730  (.A(WX7103), .B(II23714), .Z(II23715) ) ;
NAND2   gate15731  (.A(CRC_OUT_4_4), .B(II23714), .Z(II23716) ) ;
NAND2   gate15732  (.A(WX7105), .B(CRC_OUT_4_2), .Z(II23721) ) ;
NAND2   gate15733  (.A(WX7105), .B(II23721), .Z(II23722) ) ;
NAND2   gate15734  (.A(CRC_OUT_4_2), .B(II23721), .Z(II23723) ) ;
NAND2   gate15735  (.A(WX7106), .B(CRC_OUT_4_1), .Z(II23728) ) ;
NAND2   gate15736  (.A(WX7106), .B(II23728), .Z(II23729) ) ;
NAND2   gate15737  (.A(CRC_OUT_4_1), .B(II23728), .Z(II23730) ) ;
NAND2   gate15738  (.A(WX7107), .B(CRC_OUT_4_0), .Z(II23735) ) ;
NAND2   gate15739  (.A(WX7107), .B(II23735), .Z(II23736) ) ;
NAND2   gate15740  (.A(CRC_OUT_4_0), .B(II23735), .Z(II23737) ) ;
NAND2   gate15741  (.A(WX8759), .B(WX8403), .Z(II26018) ) ;
NAND2   gate15742  (.A(WX8759), .B(II26018), .Z(II26019) ) ;
NAND2   gate15743  (.A(WX8403), .B(II26018), .Z(II26020) ) ;
NAND2   gate15744  (.A(II26019), .B(II26020), .Z(II26017) ) ;
NAND2   gate15745  (.A(WX8467), .B(II26017), .Z(II26025) ) ;
NAND2   gate15746  (.A(WX8467), .B(II26025), .Z(II26026) ) ;
NAND2   gate15747  (.A(II26017), .B(II26025), .Z(II26027) ) ;
NAND2   gate15748  (.A(II26026), .B(II26027), .Z(II26016) ) ;
NAND2   gate15749  (.A(WX8531), .B(WX8595), .Z(II26033) ) ;
NAND2   gate15750  (.A(WX8531), .B(II26033), .Z(II26034) ) ;
NAND2   gate15751  (.A(WX8595), .B(II26033), .Z(II26035) ) ;
NAND2   gate15752  (.A(II26034), .B(II26035), .Z(II26032) ) ;
NAND2   gate15753  (.A(II26016), .B(II26032), .Z(II26040) ) ;
NAND2   gate15754  (.A(II26016), .B(II26040), .Z(II26041) ) ;
NAND2   gate15755  (.A(II26032), .B(II26040), .Z(II26042) ) ;
NAND2   gate15756  (.A(WX8759), .B(WX8405), .Z(II26049) ) ;
NAND2   gate15757  (.A(WX8759), .B(II26049), .Z(II26050) ) ;
NAND2   gate15758  (.A(WX8405), .B(II26049), .Z(II26051) ) ;
NAND2   gate15759  (.A(II26050), .B(II26051), .Z(II26048) ) ;
NAND2   gate15760  (.A(WX8469), .B(II26048), .Z(II26056) ) ;
NAND2   gate15761  (.A(WX8469), .B(II26056), .Z(II26057) ) ;
NAND2   gate15762  (.A(II26048), .B(II26056), .Z(II26058) ) ;
NAND2   gate15763  (.A(II26057), .B(II26058), .Z(II26047) ) ;
NAND2   gate15764  (.A(WX8533), .B(WX8597), .Z(II26064) ) ;
NAND2   gate15765  (.A(WX8533), .B(II26064), .Z(II26065) ) ;
NAND2   gate15766  (.A(WX8597), .B(II26064), .Z(II26066) ) ;
NAND2   gate15767  (.A(II26065), .B(II26066), .Z(II26063) ) ;
NAND2   gate15768  (.A(II26047), .B(II26063), .Z(II26071) ) ;
NAND2   gate15769  (.A(II26047), .B(II26071), .Z(II26072) ) ;
NAND2   gate15770  (.A(II26063), .B(II26071), .Z(II26073) ) ;
NAND2   gate15771  (.A(WX8759), .B(WX8407), .Z(II26080) ) ;
NAND2   gate15772  (.A(WX8759), .B(II26080), .Z(II26081) ) ;
NAND2   gate15773  (.A(WX8407), .B(II26080), .Z(II26082) ) ;
NAND2   gate15774  (.A(II26081), .B(II26082), .Z(II26079) ) ;
NAND2   gate15775  (.A(WX8471), .B(II26079), .Z(II26087) ) ;
NAND2   gate15776  (.A(WX8471), .B(II26087), .Z(II26088) ) ;
NAND2   gate15777  (.A(II26079), .B(II26087), .Z(II26089) ) ;
NAND2   gate15778  (.A(II26088), .B(II26089), .Z(II26078) ) ;
NAND2   gate15779  (.A(WX8535), .B(WX8599), .Z(II26095) ) ;
NAND2   gate15780  (.A(WX8535), .B(II26095), .Z(II26096) ) ;
NAND2   gate15781  (.A(WX8599), .B(II26095), .Z(II26097) ) ;
NAND2   gate15782  (.A(II26096), .B(II26097), .Z(II26094) ) ;
NAND2   gate15783  (.A(II26078), .B(II26094), .Z(II26102) ) ;
NAND2   gate15784  (.A(II26078), .B(II26102), .Z(II26103) ) ;
NAND2   gate15785  (.A(II26094), .B(II26102), .Z(II26104) ) ;
NAND2   gate15786  (.A(WX8759), .B(WX8409), .Z(II26111) ) ;
NAND2   gate15787  (.A(WX8759), .B(II26111), .Z(II26112) ) ;
NAND2   gate15788  (.A(WX8409), .B(II26111), .Z(II26113) ) ;
NAND2   gate15789  (.A(II26112), .B(II26113), .Z(II26110) ) ;
NAND2   gate15790  (.A(WX8473), .B(II26110), .Z(II26118) ) ;
NAND2   gate15791  (.A(WX8473), .B(II26118), .Z(II26119) ) ;
NAND2   gate15792  (.A(II26110), .B(II26118), .Z(II26120) ) ;
NAND2   gate15793  (.A(II26119), .B(II26120), .Z(II26109) ) ;
NAND2   gate15794  (.A(WX8537), .B(WX8601), .Z(II26126) ) ;
NAND2   gate15795  (.A(WX8537), .B(II26126), .Z(II26127) ) ;
NAND2   gate15796  (.A(WX8601), .B(II26126), .Z(II26128) ) ;
NAND2   gate15797  (.A(II26127), .B(II26128), .Z(II26125) ) ;
NAND2   gate15798  (.A(II26109), .B(II26125), .Z(II26133) ) ;
NAND2   gate15799  (.A(II26109), .B(II26133), .Z(II26134) ) ;
NAND2   gate15800  (.A(II26125), .B(II26133), .Z(II26135) ) ;
NAND2   gate15801  (.A(WX8759), .B(WX8411), .Z(II26142) ) ;
NAND2   gate15802  (.A(WX8759), .B(II26142), .Z(II26143) ) ;
NAND2   gate15803  (.A(WX8411), .B(II26142), .Z(II26144) ) ;
NAND2   gate15804  (.A(II26143), .B(II26144), .Z(II26141) ) ;
NAND2   gate15805  (.A(WX8475), .B(II26141), .Z(II26149) ) ;
NAND2   gate15806  (.A(WX8475), .B(II26149), .Z(II26150) ) ;
NAND2   gate15807  (.A(II26141), .B(II26149), .Z(II26151) ) ;
NAND2   gate15808  (.A(II26150), .B(II26151), .Z(II26140) ) ;
NAND2   gate15809  (.A(WX8539), .B(WX8603), .Z(II26157) ) ;
NAND2   gate15810  (.A(WX8539), .B(II26157), .Z(II26158) ) ;
NAND2   gate15811  (.A(WX8603), .B(II26157), .Z(II26159) ) ;
NAND2   gate15812  (.A(II26158), .B(II26159), .Z(II26156) ) ;
NAND2   gate15813  (.A(II26140), .B(II26156), .Z(II26164) ) ;
NAND2   gate15814  (.A(II26140), .B(II26164), .Z(II26165) ) ;
NAND2   gate15815  (.A(II26156), .B(II26164), .Z(II26166) ) ;
NAND2   gate15816  (.A(WX8759), .B(WX8413), .Z(II26173) ) ;
NAND2   gate15817  (.A(WX8759), .B(II26173), .Z(II26174) ) ;
NAND2   gate15818  (.A(WX8413), .B(II26173), .Z(II26175) ) ;
NAND2   gate15819  (.A(II26174), .B(II26175), .Z(II26172) ) ;
NAND2   gate15820  (.A(WX8477), .B(II26172), .Z(II26180) ) ;
NAND2   gate15821  (.A(WX8477), .B(II26180), .Z(II26181) ) ;
NAND2   gate15822  (.A(II26172), .B(II26180), .Z(II26182) ) ;
NAND2   gate15823  (.A(II26181), .B(II26182), .Z(II26171) ) ;
NAND2   gate15824  (.A(WX8541), .B(WX8605), .Z(II26188) ) ;
NAND2   gate15825  (.A(WX8541), .B(II26188), .Z(II26189) ) ;
NAND2   gate15826  (.A(WX8605), .B(II26188), .Z(II26190) ) ;
NAND2   gate15827  (.A(II26189), .B(II26190), .Z(II26187) ) ;
NAND2   gate15828  (.A(II26171), .B(II26187), .Z(II26195) ) ;
NAND2   gate15829  (.A(II26171), .B(II26195), .Z(II26196) ) ;
NAND2   gate15830  (.A(II26187), .B(II26195), .Z(II26197) ) ;
NAND2   gate15831  (.A(WX8759), .B(WX8415), .Z(II26204) ) ;
NAND2   gate15832  (.A(WX8759), .B(II26204), .Z(II26205) ) ;
NAND2   gate15833  (.A(WX8415), .B(II26204), .Z(II26206) ) ;
NAND2   gate15834  (.A(II26205), .B(II26206), .Z(II26203) ) ;
NAND2   gate15835  (.A(WX8479), .B(II26203), .Z(II26211) ) ;
NAND2   gate15836  (.A(WX8479), .B(II26211), .Z(II26212) ) ;
NAND2   gate15837  (.A(II26203), .B(II26211), .Z(II26213) ) ;
NAND2   gate15838  (.A(II26212), .B(II26213), .Z(II26202) ) ;
NAND2   gate15839  (.A(WX8543), .B(WX8607), .Z(II26219) ) ;
NAND2   gate15840  (.A(WX8543), .B(II26219), .Z(II26220) ) ;
NAND2   gate15841  (.A(WX8607), .B(II26219), .Z(II26221) ) ;
NAND2   gate15842  (.A(II26220), .B(II26221), .Z(II26218) ) ;
NAND2   gate15843  (.A(II26202), .B(II26218), .Z(II26226) ) ;
NAND2   gate15844  (.A(II26202), .B(II26226), .Z(II26227) ) ;
NAND2   gate15845  (.A(II26218), .B(II26226), .Z(II26228) ) ;
NAND2   gate15846  (.A(WX8759), .B(WX8417), .Z(II26235) ) ;
NAND2   gate15847  (.A(WX8759), .B(II26235), .Z(II26236) ) ;
NAND2   gate15848  (.A(WX8417), .B(II26235), .Z(II26237) ) ;
NAND2   gate15849  (.A(II26236), .B(II26237), .Z(II26234) ) ;
NAND2   gate15850  (.A(WX8481), .B(II26234), .Z(II26242) ) ;
NAND2   gate15851  (.A(WX8481), .B(II26242), .Z(II26243) ) ;
NAND2   gate15852  (.A(II26234), .B(II26242), .Z(II26244) ) ;
NAND2   gate15853  (.A(II26243), .B(II26244), .Z(II26233) ) ;
NAND2   gate15854  (.A(WX8545), .B(WX8609), .Z(II26250) ) ;
NAND2   gate15855  (.A(WX8545), .B(II26250), .Z(II26251) ) ;
NAND2   gate15856  (.A(WX8609), .B(II26250), .Z(II26252) ) ;
NAND2   gate15857  (.A(II26251), .B(II26252), .Z(II26249) ) ;
NAND2   gate15858  (.A(II26233), .B(II26249), .Z(II26257) ) ;
NAND2   gate15859  (.A(II26233), .B(II26257), .Z(II26258) ) ;
NAND2   gate15860  (.A(II26249), .B(II26257), .Z(II26259) ) ;
NAND2   gate15861  (.A(WX8759), .B(WX8419), .Z(II26266) ) ;
NAND2   gate15862  (.A(WX8759), .B(II26266), .Z(II26267) ) ;
NAND2   gate15863  (.A(WX8419), .B(II26266), .Z(II26268) ) ;
NAND2   gate15864  (.A(II26267), .B(II26268), .Z(II26265) ) ;
NAND2   gate15865  (.A(WX8483), .B(II26265), .Z(II26273) ) ;
NAND2   gate15866  (.A(WX8483), .B(II26273), .Z(II26274) ) ;
NAND2   gate15867  (.A(II26265), .B(II26273), .Z(II26275) ) ;
NAND2   gate15868  (.A(II26274), .B(II26275), .Z(II26264) ) ;
NAND2   gate15869  (.A(WX8547), .B(WX8611), .Z(II26281) ) ;
NAND2   gate15870  (.A(WX8547), .B(II26281), .Z(II26282) ) ;
NAND2   gate15871  (.A(WX8611), .B(II26281), .Z(II26283) ) ;
NAND2   gate15872  (.A(II26282), .B(II26283), .Z(II26280) ) ;
NAND2   gate15873  (.A(II26264), .B(II26280), .Z(II26288) ) ;
NAND2   gate15874  (.A(II26264), .B(II26288), .Z(II26289) ) ;
NAND2   gate15875  (.A(II26280), .B(II26288), .Z(II26290) ) ;
NAND2   gate15876  (.A(WX8759), .B(WX8421), .Z(II26297) ) ;
NAND2   gate15877  (.A(WX8759), .B(II26297), .Z(II26298) ) ;
NAND2   gate15878  (.A(WX8421), .B(II26297), .Z(II26299) ) ;
NAND2   gate15879  (.A(II26298), .B(II26299), .Z(II26296) ) ;
NAND2   gate15880  (.A(WX8485), .B(II26296), .Z(II26304) ) ;
NAND2   gate15881  (.A(WX8485), .B(II26304), .Z(II26305) ) ;
NAND2   gate15882  (.A(II26296), .B(II26304), .Z(II26306) ) ;
NAND2   gate15883  (.A(II26305), .B(II26306), .Z(II26295) ) ;
NAND2   gate15884  (.A(WX8549), .B(WX8613), .Z(II26312) ) ;
NAND2   gate15885  (.A(WX8549), .B(II26312), .Z(II26313) ) ;
NAND2   gate15886  (.A(WX8613), .B(II26312), .Z(II26314) ) ;
NAND2   gate15887  (.A(II26313), .B(II26314), .Z(II26311) ) ;
NAND2   gate15888  (.A(II26295), .B(II26311), .Z(II26319) ) ;
NAND2   gate15889  (.A(II26295), .B(II26319), .Z(II26320) ) ;
NAND2   gate15890  (.A(II26311), .B(II26319), .Z(II26321) ) ;
NAND2   gate15891  (.A(WX8759), .B(WX8423), .Z(II26328) ) ;
NAND2   gate15892  (.A(WX8759), .B(II26328), .Z(II26329) ) ;
NAND2   gate15893  (.A(WX8423), .B(II26328), .Z(II26330) ) ;
NAND2   gate15894  (.A(II26329), .B(II26330), .Z(II26327) ) ;
NAND2   gate15895  (.A(WX8487), .B(II26327), .Z(II26335) ) ;
NAND2   gate15896  (.A(WX8487), .B(II26335), .Z(II26336) ) ;
NAND2   gate15897  (.A(II26327), .B(II26335), .Z(II26337) ) ;
NAND2   gate15898  (.A(II26336), .B(II26337), .Z(II26326) ) ;
NAND2   gate15899  (.A(WX8551), .B(WX8615), .Z(II26343) ) ;
NAND2   gate15900  (.A(WX8551), .B(II26343), .Z(II26344) ) ;
NAND2   gate15901  (.A(WX8615), .B(II26343), .Z(II26345) ) ;
NAND2   gate15902  (.A(II26344), .B(II26345), .Z(II26342) ) ;
NAND2   gate15903  (.A(II26326), .B(II26342), .Z(II26350) ) ;
NAND2   gate15904  (.A(II26326), .B(II26350), .Z(II26351) ) ;
NAND2   gate15905  (.A(II26342), .B(II26350), .Z(II26352) ) ;
NAND2   gate15906  (.A(WX8759), .B(WX8425), .Z(II26359) ) ;
NAND2   gate15907  (.A(WX8759), .B(II26359), .Z(II26360) ) ;
NAND2   gate15908  (.A(WX8425), .B(II26359), .Z(II26361) ) ;
NAND2   gate15909  (.A(II26360), .B(II26361), .Z(II26358) ) ;
NAND2   gate15910  (.A(WX8489), .B(II26358), .Z(II26366) ) ;
NAND2   gate15911  (.A(WX8489), .B(II26366), .Z(II26367) ) ;
NAND2   gate15912  (.A(II26358), .B(II26366), .Z(II26368) ) ;
NAND2   gate15913  (.A(II26367), .B(II26368), .Z(II26357) ) ;
NAND2   gate15914  (.A(WX8553), .B(WX8617), .Z(II26374) ) ;
NAND2   gate15915  (.A(WX8553), .B(II26374), .Z(II26375) ) ;
NAND2   gate15916  (.A(WX8617), .B(II26374), .Z(II26376) ) ;
NAND2   gate15917  (.A(II26375), .B(II26376), .Z(II26373) ) ;
NAND2   gate15918  (.A(II26357), .B(II26373), .Z(II26381) ) ;
NAND2   gate15919  (.A(II26357), .B(II26381), .Z(II26382) ) ;
NAND2   gate15920  (.A(II26373), .B(II26381), .Z(II26383) ) ;
NAND2   gate15921  (.A(WX8759), .B(WX8427), .Z(II26390) ) ;
NAND2   gate15922  (.A(WX8759), .B(II26390), .Z(II26391) ) ;
NAND2   gate15923  (.A(WX8427), .B(II26390), .Z(II26392) ) ;
NAND2   gate15924  (.A(II26391), .B(II26392), .Z(II26389) ) ;
NAND2   gate15925  (.A(WX8491), .B(II26389), .Z(II26397) ) ;
NAND2   gate15926  (.A(WX8491), .B(II26397), .Z(II26398) ) ;
NAND2   gate15927  (.A(II26389), .B(II26397), .Z(II26399) ) ;
NAND2   gate15928  (.A(II26398), .B(II26399), .Z(II26388) ) ;
NAND2   gate15929  (.A(WX8555), .B(WX8619), .Z(II26405) ) ;
NAND2   gate15930  (.A(WX8555), .B(II26405), .Z(II26406) ) ;
NAND2   gate15931  (.A(WX8619), .B(II26405), .Z(II26407) ) ;
NAND2   gate15932  (.A(II26406), .B(II26407), .Z(II26404) ) ;
NAND2   gate15933  (.A(II26388), .B(II26404), .Z(II26412) ) ;
NAND2   gate15934  (.A(II26388), .B(II26412), .Z(II26413) ) ;
NAND2   gate15935  (.A(II26404), .B(II26412), .Z(II26414) ) ;
NAND2   gate15936  (.A(WX8759), .B(WX8429), .Z(II26421) ) ;
NAND2   gate15937  (.A(WX8759), .B(II26421), .Z(II26422) ) ;
NAND2   gate15938  (.A(WX8429), .B(II26421), .Z(II26423) ) ;
NAND2   gate15939  (.A(II26422), .B(II26423), .Z(II26420) ) ;
NAND2   gate15940  (.A(WX8493), .B(II26420), .Z(II26428) ) ;
NAND2   gate15941  (.A(WX8493), .B(II26428), .Z(II26429) ) ;
NAND2   gate15942  (.A(II26420), .B(II26428), .Z(II26430) ) ;
NAND2   gate15943  (.A(II26429), .B(II26430), .Z(II26419) ) ;
NAND2   gate15944  (.A(WX8557), .B(WX8621), .Z(II26436) ) ;
NAND2   gate15945  (.A(WX8557), .B(II26436), .Z(II26437) ) ;
NAND2   gate15946  (.A(WX8621), .B(II26436), .Z(II26438) ) ;
NAND2   gate15947  (.A(II26437), .B(II26438), .Z(II26435) ) ;
NAND2   gate15948  (.A(II26419), .B(II26435), .Z(II26443) ) ;
NAND2   gate15949  (.A(II26419), .B(II26443), .Z(II26444) ) ;
NAND2   gate15950  (.A(II26435), .B(II26443), .Z(II26445) ) ;
NAND2   gate15951  (.A(WX8759), .B(WX8431), .Z(II26452) ) ;
NAND2   gate15952  (.A(WX8759), .B(II26452), .Z(II26453) ) ;
NAND2   gate15953  (.A(WX8431), .B(II26452), .Z(II26454) ) ;
NAND2   gate15954  (.A(II26453), .B(II26454), .Z(II26451) ) ;
NAND2   gate15955  (.A(WX8495), .B(II26451), .Z(II26459) ) ;
NAND2   gate15956  (.A(WX8495), .B(II26459), .Z(II26460) ) ;
NAND2   gate15957  (.A(II26451), .B(II26459), .Z(II26461) ) ;
NAND2   gate15958  (.A(II26460), .B(II26461), .Z(II26450) ) ;
NAND2   gate15959  (.A(WX8559), .B(WX8623), .Z(II26467) ) ;
NAND2   gate15960  (.A(WX8559), .B(II26467), .Z(II26468) ) ;
NAND2   gate15961  (.A(WX8623), .B(II26467), .Z(II26469) ) ;
NAND2   gate15962  (.A(II26468), .B(II26469), .Z(II26466) ) ;
NAND2   gate15963  (.A(II26450), .B(II26466), .Z(II26474) ) ;
NAND2   gate15964  (.A(II26450), .B(II26474), .Z(II26475) ) ;
NAND2   gate15965  (.A(II26466), .B(II26474), .Z(II26476) ) ;
NAND2   gate15966  (.A(WX8759), .B(WX8433), .Z(II26483) ) ;
NAND2   gate15967  (.A(WX8759), .B(II26483), .Z(II26484) ) ;
NAND2   gate15968  (.A(WX8433), .B(II26483), .Z(II26485) ) ;
NAND2   gate15969  (.A(II26484), .B(II26485), .Z(II26482) ) ;
NAND2   gate15970  (.A(WX8497), .B(II26482), .Z(II26490) ) ;
NAND2   gate15971  (.A(WX8497), .B(II26490), .Z(II26491) ) ;
NAND2   gate15972  (.A(II26482), .B(II26490), .Z(II26492) ) ;
NAND2   gate15973  (.A(II26491), .B(II26492), .Z(II26481) ) ;
NAND2   gate15974  (.A(WX8561), .B(WX8625), .Z(II26498) ) ;
NAND2   gate15975  (.A(WX8561), .B(II26498), .Z(II26499) ) ;
NAND2   gate15976  (.A(WX8625), .B(II26498), .Z(II26500) ) ;
NAND2   gate15977  (.A(II26499), .B(II26500), .Z(II26497) ) ;
NAND2   gate15978  (.A(II26481), .B(II26497), .Z(II26505) ) ;
NAND2   gate15979  (.A(II26481), .B(II26505), .Z(II26506) ) ;
NAND2   gate15980  (.A(II26497), .B(II26505), .Z(II26507) ) ;
NAND2   gate15981  (.A(WX8760), .B(WX8435), .Z(II26514) ) ;
NAND2   gate15982  (.A(WX8760), .B(II26514), .Z(II26515) ) ;
NAND2   gate15983  (.A(WX8435), .B(II26514), .Z(II26516) ) ;
NAND2   gate15984  (.A(II26515), .B(II26516), .Z(II26513) ) ;
NAND2   gate15985  (.A(WX8499), .B(II26513), .Z(II26521) ) ;
NAND2   gate15986  (.A(WX8499), .B(II26521), .Z(II26522) ) ;
NAND2   gate15987  (.A(II26513), .B(II26521), .Z(II26523) ) ;
NAND2   gate15988  (.A(II26522), .B(II26523), .Z(II26512) ) ;
NAND2   gate15989  (.A(WX8563), .B(WX8627), .Z(II26529) ) ;
NAND2   gate15990  (.A(WX8563), .B(II26529), .Z(II26530) ) ;
NAND2   gate15991  (.A(WX8627), .B(II26529), .Z(II26531) ) ;
NAND2   gate15992  (.A(II26530), .B(II26531), .Z(II26528) ) ;
NAND2   gate15993  (.A(II26512), .B(II26528), .Z(II26536) ) ;
NAND2   gate15994  (.A(II26512), .B(II26536), .Z(II26537) ) ;
NAND2   gate15995  (.A(II26528), .B(II26536), .Z(II26538) ) ;
NAND2   gate15996  (.A(WX8760), .B(WX8437), .Z(II26545) ) ;
NAND2   gate15997  (.A(WX8760), .B(II26545), .Z(II26546) ) ;
NAND2   gate15998  (.A(WX8437), .B(II26545), .Z(II26547) ) ;
NAND2   gate15999  (.A(II26546), .B(II26547), .Z(II26544) ) ;
NAND2   gate16000  (.A(WX8501), .B(II26544), .Z(II26552) ) ;
NAND2   gate16001  (.A(WX8501), .B(II26552), .Z(II26553) ) ;
NAND2   gate16002  (.A(II26544), .B(II26552), .Z(II26554) ) ;
NAND2   gate16003  (.A(II26553), .B(II26554), .Z(II26543) ) ;
NAND2   gate16004  (.A(WX8565), .B(WX8629), .Z(II26560) ) ;
NAND2   gate16005  (.A(WX8565), .B(II26560), .Z(II26561) ) ;
NAND2   gate16006  (.A(WX8629), .B(II26560), .Z(II26562) ) ;
NAND2   gate16007  (.A(II26561), .B(II26562), .Z(II26559) ) ;
NAND2   gate16008  (.A(II26543), .B(II26559), .Z(II26567) ) ;
NAND2   gate16009  (.A(II26543), .B(II26567), .Z(II26568) ) ;
NAND2   gate16010  (.A(II26559), .B(II26567), .Z(II26569) ) ;
NAND2   gate16011  (.A(WX8760), .B(WX8439), .Z(II26576) ) ;
NAND2   gate16012  (.A(WX8760), .B(II26576), .Z(II26577) ) ;
NAND2   gate16013  (.A(WX8439), .B(II26576), .Z(II26578) ) ;
NAND2   gate16014  (.A(II26577), .B(II26578), .Z(II26575) ) ;
NAND2   gate16015  (.A(WX8503), .B(II26575), .Z(II26583) ) ;
NAND2   gate16016  (.A(WX8503), .B(II26583), .Z(II26584) ) ;
NAND2   gate16017  (.A(II26575), .B(II26583), .Z(II26585) ) ;
NAND2   gate16018  (.A(II26584), .B(II26585), .Z(II26574) ) ;
NAND2   gate16019  (.A(WX8567), .B(WX8631), .Z(II26591) ) ;
NAND2   gate16020  (.A(WX8567), .B(II26591), .Z(II26592) ) ;
NAND2   gate16021  (.A(WX8631), .B(II26591), .Z(II26593) ) ;
NAND2   gate16022  (.A(II26592), .B(II26593), .Z(II26590) ) ;
NAND2   gate16023  (.A(II26574), .B(II26590), .Z(II26598) ) ;
NAND2   gate16024  (.A(II26574), .B(II26598), .Z(II26599) ) ;
NAND2   gate16025  (.A(II26590), .B(II26598), .Z(II26600) ) ;
NAND2   gate16026  (.A(WX8760), .B(WX8441), .Z(II26607) ) ;
NAND2   gate16027  (.A(WX8760), .B(II26607), .Z(II26608) ) ;
NAND2   gate16028  (.A(WX8441), .B(II26607), .Z(II26609) ) ;
NAND2   gate16029  (.A(II26608), .B(II26609), .Z(II26606) ) ;
NAND2   gate16030  (.A(WX8505), .B(II26606), .Z(II26614) ) ;
NAND2   gate16031  (.A(WX8505), .B(II26614), .Z(II26615) ) ;
NAND2   gate16032  (.A(II26606), .B(II26614), .Z(II26616) ) ;
NAND2   gate16033  (.A(II26615), .B(II26616), .Z(II26605) ) ;
NAND2   gate16034  (.A(WX8569), .B(WX8633), .Z(II26622) ) ;
NAND2   gate16035  (.A(WX8569), .B(II26622), .Z(II26623) ) ;
NAND2   gate16036  (.A(WX8633), .B(II26622), .Z(II26624) ) ;
NAND2   gate16037  (.A(II26623), .B(II26624), .Z(II26621) ) ;
NAND2   gate16038  (.A(II26605), .B(II26621), .Z(II26629) ) ;
NAND2   gate16039  (.A(II26605), .B(II26629), .Z(II26630) ) ;
NAND2   gate16040  (.A(II26621), .B(II26629), .Z(II26631) ) ;
NAND2   gate16041  (.A(WX8760), .B(WX8443), .Z(II26638) ) ;
NAND2   gate16042  (.A(WX8760), .B(II26638), .Z(II26639) ) ;
NAND2   gate16043  (.A(WX8443), .B(II26638), .Z(II26640) ) ;
NAND2   gate16044  (.A(II26639), .B(II26640), .Z(II26637) ) ;
NAND2   gate16045  (.A(WX8507), .B(II26637), .Z(II26645) ) ;
NAND2   gate16046  (.A(WX8507), .B(II26645), .Z(II26646) ) ;
NAND2   gate16047  (.A(II26637), .B(II26645), .Z(II26647) ) ;
NAND2   gate16048  (.A(II26646), .B(II26647), .Z(II26636) ) ;
NAND2   gate16049  (.A(WX8571), .B(WX8635), .Z(II26653) ) ;
NAND2   gate16050  (.A(WX8571), .B(II26653), .Z(II26654) ) ;
NAND2   gate16051  (.A(WX8635), .B(II26653), .Z(II26655) ) ;
NAND2   gate16052  (.A(II26654), .B(II26655), .Z(II26652) ) ;
NAND2   gate16053  (.A(II26636), .B(II26652), .Z(II26660) ) ;
NAND2   gate16054  (.A(II26636), .B(II26660), .Z(II26661) ) ;
NAND2   gate16055  (.A(II26652), .B(II26660), .Z(II26662) ) ;
NAND2   gate16056  (.A(WX8760), .B(WX8445), .Z(II26669) ) ;
NAND2   gate16057  (.A(WX8760), .B(II26669), .Z(II26670) ) ;
NAND2   gate16058  (.A(WX8445), .B(II26669), .Z(II26671) ) ;
NAND2   gate16059  (.A(II26670), .B(II26671), .Z(II26668) ) ;
NAND2   gate16060  (.A(WX8509), .B(II26668), .Z(II26676) ) ;
NAND2   gate16061  (.A(WX8509), .B(II26676), .Z(II26677) ) ;
NAND2   gate16062  (.A(II26668), .B(II26676), .Z(II26678) ) ;
NAND2   gate16063  (.A(II26677), .B(II26678), .Z(II26667) ) ;
NAND2   gate16064  (.A(WX8573), .B(WX8637), .Z(II26684) ) ;
NAND2   gate16065  (.A(WX8573), .B(II26684), .Z(II26685) ) ;
NAND2   gate16066  (.A(WX8637), .B(II26684), .Z(II26686) ) ;
NAND2   gate16067  (.A(II26685), .B(II26686), .Z(II26683) ) ;
NAND2   gate16068  (.A(II26667), .B(II26683), .Z(II26691) ) ;
NAND2   gate16069  (.A(II26667), .B(II26691), .Z(II26692) ) ;
NAND2   gate16070  (.A(II26683), .B(II26691), .Z(II26693) ) ;
NAND2   gate16071  (.A(WX8760), .B(WX8447), .Z(II26700) ) ;
NAND2   gate16072  (.A(WX8760), .B(II26700), .Z(II26701) ) ;
NAND2   gate16073  (.A(WX8447), .B(II26700), .Z(II26702) ) ;
NAND2   gate16074  (.A(II26701), .B(II26702), .Z(II26699) ) ;
NAND2   gate16075  (.A(WX8511), .B(II26699), .Z(II26707) ) ;
NAND2   gate16076  (.A(WX8511), .B(II26707), .Z(II26708) ) ;
NAND2   gate16077  (.A(II26699), .B(II26707), .Z(II26709) ) ;
NAND2   gate16078  (.A(II26708), .B(II26709), .Z(II26698) ) ;
NAND2   gate16079  (.A(WX8575), .B(WX8639), .Z(II26715) ) ;
NAND2   gate16080  (.A(WX8575), .B(II26715), .Z(II26716) ) ;
NAND2   gate16081  (.A(WX8639), .B(II26715), .Z(II26717) ) ;
NAND2   gate16082  (.A(II26716), .B(II26717), .Z(II26714) ) ;
NAND2   gate16083  (.A(II26698), .B(II26714), .Z(II26722) ) ;
NAND2   gate16084  (.A(II26698), .B(II26722), .Z(II26723) ) ;
NAND2   gate16085  (.A(II26714), .B(II26722), .Z(II26724) ) ;
NAND2   gate16086  (.A(WX8760), .B(WX8449), .Z(II26731) ) ;
NAND2   gate16087  (.A(WX8760), .B(II26731), .Z(II26732) ) ;
NAND2   gate16088  (.A(WX8449), .B(II26731), .Z(II26733) ) ;
NAND2   gate16089  (.A(II26732), .B(II26733), .Z(II26730) ) ;
NAND2   gate16090  (.A(WX8513), .B(II26730), .Z(II26738) ) ;
NAND2   gate16091  (.A(WX8513), .B(II26738), .Z(II26739) ) ;
NAND2   gate16092  (.A(II26730), .B(II26738), .Z(II26740) ) ;
NAND2   gate16093  (.A(II26739), .B(II26740), .Z(II26729) ) ;
NAND2   gate16094  (.A(WX8577), .B(WX8641), .Z(II26746) ) ;
NAND2   gate16095  (.A(WX8577), .B(II26746), .Z(II26747) ) ;
NAND2   gate16096  (.A(WX8641), .B(II26746), .Z(II26748) ) ;
NAND2   gate16097  (.A(II26747), .B(II26748), .Z(II26745) ) ;
NAND2   gate16098  (.A(II26729), .B(II26745), .Z(II26753) ) ;
NAND2   gate16099  (.A(II26729), .B(II26753), .Z(II26754) ) ;
NAND2   gate16100  (.A(II26745), .B(II26753), .Z(II26755) ) ;
NAND2   gate16101  (.A(WX8760), .B(WX8451), .Z(II26762) ) ;
NAND2   gate16102  (.A(WX8760), .B(II26762), .Z(II26763) ) ;
NAND2   gate16103  (.A(WX8451), .B(II26762), .Z(II26764) ) ;
NAND2   gate16104  (.A(II26763), .B(II26764), .Z(II26761) ) ;
NAND2   gate16105  (.A(WX8515), .B(II26761), .Z(II26769) ) ;
NAND2   gate16106  (.A(WX8515), .B(II26769), .Z(II26770) ) ;
NAND2   gate16107  (.A(II26761), .B(II26769), .Z(II26771) ) ;
NAND2   gate16108  (.A(II26770), .B(II26771), .Z(II26760) ) ;
NAND2   gate16109  (.A(WX8579), .B(WX8643), .Z(II26777) ) ;
NAND2   gate16110  (.A(WX8579), .B(II26777), .Z(II26778) ) ;
NAND2   gate16111  (.A(WX8643), .B(II26777), .Z(II26779) ) ;
NAND2   gate16112  (.A(II26778), .B(II26779), .Z(II26776) ) ;
NAND2   gate16113  (.A(II26760), .B(II26776), .Z(II26784) ) ;
NAND2   gate16114  (.A(II26760), .B(II26784), .Z(II26785) ) ;
NAND2   gate16115  (.A(II26776), .B(II26784), .Z(II26786) ) ;
NAND2   gate16116  (.A(WX8760), .B(WX8453), .Z(II26793) ) ;
NAND2   gate16117  (.A(WX8760), .B(II26793), .Z(II26794) ) ;
NAND2   gate16118  (.A(WX8453), .B(II26793), .Z(II26795) ) ;
NAND2   gate16119  (.A(II26794), .B(II26795), .Z(II26792) ) ;
NAND2   gate16120  (.A(WX8517), .B(II26792), .Z(II26800) ) ;
NAND2   gate16121  (.A(WX8517), .B(II26800), .Z(II26801) ) ;
NAND2   gate16122  (.A(II26792), .B(II26800), .Z(II26802) ) ;
NAND2   gate16123  (.A(II26801), .B(II26802), .Z(II26791) ) ;
NAND2   gate16124  (.A(WX8581), .B(WX8645), .Z(II26808) ) ;
NAND2   gate16125  (.A(WX8581), .B(II26808), .Z(II26809) ) ;
NAND2   gate16126  (.A(WX8645), .B(II26808), .Z(II26810) ) ;
NAND2   gate16127  (.A(II26809), .B(II26810), .Z(II26807) ) ;
NAND2   gate16128  (.A(II26791), .B(II26807), .Z(II26815) ) ;
NAND2   gate16129  (.A(II26791), .B(II26815), .Z(II26816) ) ;
NAND2   gate16130  (.A(II26807), .B(II26815), .Z(II26817) ) ;
NAND2   gate16131  (.A(WX8760), .B(WX8455), .Z(II26824) ) ;
NAND2   gate16132  (.A(WX8760), .B(II26824), .Z(II26825) ) ;
NAND2   gate16133  (.A(WX8455), .B(II26824), .Z(II26826) ) ;
NAND2   gate16134  (.A(II26825), .B(II26826), .Z(II26823) ) ;
NAND2   gate16135  (.A(WX8519), .B(II26823), .Z(II26831) ) ;
NAND2   gate16136  (.A(WX8519), .B(II26831), .Z(II26832) ) ;
NAND2   gate16137  (.A(II26823), .B(II26831), .Z(II26833) ) ;
NAND2   gate16138  (.A(II26832), .B(II26833), .Z(II26822) ) ;
NAND2   gate16139  (.A(WX8583), .B(WX8647), .Z(II26839) ) ;
NAND2   gate16140  (.A(WX8583), .B(II26839), .Z(II26840) ) ;
NAND2   gate16141  (.A(WX8647), .B(II26839), .Z(II26841) ) ;
NAND2   gate16142  (.A(II26840), .B(II26841), .Z(II26838) ) ;
NAND2   gate16143  (.A(II26822), .B(II26838), .Z(II26846) ) ;
NAND2   gate16144  (.A(II26822), .B(II26846), .Z(II26847) ) ;
NAND2   gate16145  (.A(II26838), .B(II26846), .Z(II26848) ) ;
NAND2   gate16146  (.A(WX8760), .B(WX8457), .Z(II26855) ) ;
NAND2   gate16147  (.A(WX8760), .B(II26855), .Z(II26856) ) ;
NAND2   gate16148  (.A(WX8457), .B(II26855), .Z(II26857) ) ;
NAND2   gate16149  (.A(II26856), .B(II26857), .Z(II26854) ) ;
NAND2   gate16150  (.A(WX8521), .B(II26854), .Z(II26862) ) ;
NAND2   gate16151  (.A(WX8521), .B(II26862), .Z(II26863) ) ;
NAND2   gate16152  (.A(II26854), .B(II26862), .Z(II26864) ) ;
NAND2   gate16153  (.A(II26863), .B(II26864), .Z(II26853) ) ;
NAND2   gate16154  (.A(WX8585), .B(WX8649), .Z(II26870) ) ;
NAND2   gate16155  (.A(WX8585), .B(II26870), .Z(II26871) ) ;
NAND2   gate16156  (.A(WX8649), .B(II26870), .Z(II26872) ) ;
NAND2   gate16157  (.A(II26871), .B(II26872), .Z(II26869) ) ;
NAND2   gate16158  (.A(II26853), .B(II26869), .Z(II26877) ) ;
NAND2   gate16159  (.A(II26853), .B(II26877), .Z(II26878) ) ;
NAND2   gate16160  (.A(II26869), .B(II26877), .Z(II26879) ) ;
NAND2   gate16161  (.A(WX8760), .B(WX8459), .Z(II26886) ) ;
NAND2   gate16162  (.A(WX8760), .B(II26886), .Z(II26887) ) ;
NAND2   gate16163  (.A(WX8459), .B(II26886), .Z(II26888) ) ;
NAND2   gate16164  (.A(II26887), .B(II26888), .Z(II26885) ) ;
NAND2   gate16165  (.A(WX8523), .B(II26885), .Z(II26893) ) ;
NAND2   gate16166  (.A(WX8523), .B(II26893), .Z(II26894) ) ;
NAND2   gate16167  (.A(II26885), .B(II26893), .Z(II26895) ) ;
NAND2   gate16168  (.A(II26894), .B(II26895), .Z(II26884) ) ;
NAND2   gate16169  (.A(WX8587), .B(WX8651), .Z(II26901) ) ;
NAND2   gate16170  (.A(WX8587), .B(II26901), .Z(II26902) ) ;
NAND2   gate16171  (.A(WX8651), .B(II26901), .Z(II26903) ) ;
NAND2   gate16172  (.A(II26902), .B(II26903), .Z(II26900) ) ;
NAND2   gate16173  (.A(II26884), .B(II26900), .Z(II26908) ) ;
NAND2   gate16174  (.A(II26884), .B(II26908), .Z(II26909) ) ;
NAND2   gate16175  (.A(II26900), .B(II26908), .Z(II26910) ) ;
NAND2   gate16176  (.A(WX8760), .B(WX8461), .Z(II26917) ) ;
NAND2   gate16177  (.A(WX8760), .B(II26917), .Z(II26918) ) ;
NAND2   gate16178  (.A(WX8461), .B(II26917), .Z(II26919) ) ;
NAND2   gate16179  (.A(II26918), .B(II26919), .Z(II26916) ) ;
NAND2   gate16180  (.A(WX8525), .B(II26916), .Z(II26924) ) ;
NAND2   gate16181  (.A(WX8525), .B(II26924), .Z(II26925) ) ;
NAND2   gate16182  (.A(II26916), .B(II26924), .Z(II26926) ) ;
NAND2   gate16183  (.A(II26925), .B(II26926), .Z(II26915) ) ;
NAND2   gate16184  (.A(WX8589), .B(WX8653), .Z(II26932) ) ;
NAND2   gate16185  (.A(WX8589), .B(II26932), .Z(II26933) ) ;
NAND2   gate16186  (.A(WX8653), .B(II26932), .Z(II26934) ) ;
NAND2   gate16187  (.A(II26933), .B(II26934), .Z(II26931) ) ;
NAND2   gate16188  (.A(II26915), .B(II26931), .Z(II26939) ) ;
NAND2   gate16189  (.A(II26915), .B(II26939), .Z(II26940) ) ;
NAND2   gate16190  (.A(II26931), .B(II26939), .Z(II26941) ) ;
NAND2   gate16191  (.A(WX8760), .B(WX8463), .Z(II26948) ) ;
NAND2   gate16192  (.A(WX8760), .B(II26948), .Z(II26949) ) ;
NAND2   gate16193  (.A(WX8463), .B(II26948), .Z(II26950) ) ;
NAND2   gate16194  (.A(II26949), .B(II26950), .Z(II26947) ) ;
NAND2   gate16195  (.A(WX8527), .B(II26947), .Z(II26955) ) ;
NAND2   gate16196  (.A(WX8527), .B(II26955), .Z(II26956) ) ;
NAND2   gate16197  (.A(II26947), .B(II26955), .Z(II26957) ) ;
NAND2   gate16198  (.A(II26956), .B(II26957), .Z(II26946) ) ;
NAND2   gate16199  (.A(WX8591), .B(WX8655), .Z(II26963) ) ;
NAND2   gate16200  (.A(WX8591), .B(II26963), .Z(II26964) ) ;
NAND2   gate16201  (.A(WX8655), .B(II26963), .Z(II26965) ) ;
NAND2   gate16202  (.A(II26964), .B(II26965), .Z(II26962) ) ;
NAND2   gate16203  (.A(II26946), .B(II26962), .Z(II26970) ) ;
NAND2   gate16204  (.A(II26946), .B(II26970), .Z(II26971) ) ;
NAND2   gate16205  (.A(II26962), .B(II26970), .Z(II26972) ) ;
NAND2   gate16206  (.A(WX8760), .B(WX8465), .Z(II26979) ) ;
NAND2   gate16207  (.A(WX8760), .B(II26979), .Z(II26980) ) ;
NAND2   gate16208  (.A(WX8465), .B(II26979), .Z(II26981) ) ;
NAND2   gate16209  (.A(II26980), .B(II26981), .Z(II26978) ) ;
NAND2   gate16210  (.A(WX8529), .B(II26978), .Z(II26986) ) ;
NAND2   gate16211  (.A(WX8529), .B(II26986), .Z(II26987) ) ;
NAND2   gate16212  (.A(II26978), .B(II26986), .Z(II26988) ) ;
NAND2   gate16213  (.A(II26987), .B(II26988), .Z(II26977) ) ;
NAND2   gate16214  (.A(WX8593), .B(WX8657), .Z(II26994) ) ;
NAND2   gate16215  (.A(WX8593), .B(II26994), .Z(II26995) ) ;
NAND2   gate16216  (.A(WX8657), .B(II26994), .Z(II26996) ) ;
NAND2   gate16217  (.A(II26995), .B(II26996), .Z(II26993) ) ;
NAND2   gate16218  (.A(II26977), .B(II26993), .Z(II27001) ) ;
NAND2   gate16219  (.A(II26977), .B(II27001), .Z(II27002) ) ;
NAND2   gate16220  (.A(II26993), .B(II27001), .Z(II27003) ) ;
NAND2   gate16221  (.A(WX8338), .B(WX8243), .Z(II27082) ) ;
NAND2   gate16222  (.A(WX8338), .B(II27082), .Z(II27083) ) ;
NAND2   gate16223  (.A(WX8243), .B(II27082), .Z(II27084) ) ;
NAND2   gate16224  (.A(WX8339), .B(WX8245), .Z(II27095) ) ;
NAND2   gate16225  (.A(WX8339), .B(II27095), .Z(II27096) ) ;
NAND2   gate16226  (.A(WX8245), .B(II27095), .Z(II27097) ) ;
NAND2   gate16227  (.A(WX8340), .B(WX8247), .Z(II27108) ) ;
NAND2   gate16228  (.A(WX8340), .B(II27108), .Z(II27109) ) ;
NAND2   gate16229  (.A(WX8247), .B(II27108), .Z(II27110) ) ;
NAND2   gate16230  (.A(WX8341), .B(WX8249), .Z(II27121) ) ;
NAND2   gate16231  (.A(WX8341), .B(II27121), .Z(II27122) ) ;
NAND2   gate16232  (.A(WX8249), .B(II27121), .Z(II27123) ) ;
NAND2   gate16233  (.A(WX8342), .B(WX8251), .Z(II27134) ) ;
NAND2   gate16234  (.A(WX8342), .B(II27134), .Z(II27135) ) ;
NAND2   gate16235  (.A(WX8251), .B(II27134), .Z(II27136) ) ;
NAND2   gate16236  (.A(WX8343), .B(WX8253), .Z(II27147) ) ;
NAND2   gate16237  (.A(WX8343), .B(II27147), .Z(II27148) ) ;
NAND2   gate16238  (.A(WX8253), .B(II27147), .Z(II27149) ) ;
NAND2   gate16239  (.A(WX8344), .B(WX8255), .Z(II27160) ) ;
NAND2   gate16240  (.A(WX8344), .B(II27160), .Z(II27161) ) ;
NAND2   gate16241  (.A(WX8255), .B(II27160), .Z(II27162) ) ;
NAND2   gate16242  (.A(WX8345), .B(WX8257), .Z(II27173) ) ;
NAND2   gate16243  (.A(WX8345), .B(II27173), .Z(II27174) ) ;
NAND2   gate16244  (.A(WX8257), .B(II27173), .Z(II27175) ) ;
NAND2   gate16245  (.A(WX8346), .B(WX8259), .Z(II27186) ) ;
NAND2   gate16246  (.A(WX8346), .B(II27186), .Z(II27187) ) ;
NAND2   gate16247  (.A(WX8259), .B(II27186), .Z(II27188) ) ;
NAND2   gate16248  (.A(WX8347), .B(WX8261), .Z(II27199) ) ;
NAND2   gate16249  (.A(WX8347), .B(II27199), .Z(II27200) ) ;
NAND2   gate16250  (.A(WX8261), .B(II27199), .Z(II27201) ) ;
NAND2   gate16251  (.A(WX8348), .B(WX8263), .Z(II27212) ) ;
NAND2   gate16252  (.A(WX8348), .B(II27212), .Z(II27213) ) ;
NAND2   gate16253  (.A(WX8263), .B(II27212), .Z(II27214) ) ;
NAND2   gate16254  (.A(WX8349), .B(WX8265), .Z(II27225) ) ;
NAND2   gate16255  (.A(WX8349), .B(II27225), .Z(II27226) ) ;
NAND2   gate16256  (.A(WX8265), .B(II27225), .Z(II27227) ) ;
NAND2   gate16257  (.A(WX8350), .B(WX8267), .Z(II27238) ) ;
NAND2   gate16258  (.A(WX8350), .B(II27238), .Z(II27239) ) ;
NAND2   gate16259  (.A(WX8267), .B(II27238), .Z(II27240) ) ;
NAND2   gate16260  (.A(WX8351), .B(WX8269), .Z(II27251) ) ;
NAND2   gate16261  (.A(WX8351), .B(II27251), .Z(II27252) ) ;
NAND2   gate16262  (.A(WX8269), .B(II27251), .Z(II27253) ) ;
NAND2   gate16263  (.A(WX8352), .B(WX8271), .Z(II27264) ) ;
NAND2   gate16264  (.A(WX8352), .B(II27264), .Z(II27265) ) ;
NAND2   gate16265  (.A(WX8271), .B(II27264), .Z(II27266) ) ;
NAND2   gate16266  (.A(WX8353), .B(WX8273), .Z(II27277) ) ;
NAND2   gate16267  (.A(WX8353), .B(II27277), .Z(II27278) ) ;
NAND2   gate16268  (.A(WX8273), .B(II27277), .Z(II27279) ) ;
NAND2   gate16269  (.A(WX8354), .B(WX8275), .Z(II27290) ) ;
NAND2   gate16270  (.A(WX8354), .B(II27290), .Z(II27291) ) ;
NAND2   gate16271  (.A(WX8275), .B(II27290), .Z(II27292) ) ;
NAND2   gate16272  (.A(WX8355), .B(WX8277), .Z(II27303) ) ;
NAND2   gate16273  (.A(WX8355), .B(II27303), .Z(II27304) ) ;
NAND2   gate16274  (.A(WX8277), .B(II27303), .Z(II27305) ) ;
NAND2   gate16275  (.A(WX8356), .B(WX8279), .Z(II27316) ) ;
NAND2   gate16276  (.A(WX8356), .B(II27316), .Z(II27317) ) ;
NAND2   gate16277  (.A(WX8279), .B(II27316), .Z(II27318) ) ;
NAND2   gate16278  (.A(WX8357), .B(WX8281), .Z(II27329) ) ;
NAND2   gate16279  (.A(WX8357), .B(II27329), .Z(II27330) ) ;
NAND2   gate16280  (.A(WX8281), .B(II27329), .Z(II27331) ) ;
NAND2   gate16281  (.A(WX8358), .B(WX8283), .Z(II27342) ) ;
NAND2   gate16282  (.A(WX8358), .B(II27342), .Z(II27343) ) ;
NAND2   gate16283  (.A(WX8283), .B(II27342), .Z(II27344) ) ;
NAND2   gate16284  (.A(WX8359), .B(WX8285), .Z(II27355) ) ;
NAND2   gate16285  (.A(WX8359), .B(II27355), .Z(II27356) ) ;
NAND2   gate16286  (.A(WX8285), .B(II27355), .Z(II27357) ) ;
NAND2   gate16287  (.A(WX8360), .B(WX8287), .Z(II27368) ) ;
NAND2   gate16288  (.A(WX8360), .B(II27368), .Z(II27369) ) ;
NAND2   gate16289  (.A(WX8287), .B(II27368), .Z(II27370) ) ;
NAND2   gate16290  (.A(WX8361), .B(WX8289), .Z(II27381) ) ;
NAND2   gate16291  (.A(WX8361), .B(II27381), .Z(II27382) ) ;
NAND2   gate16292  (.A(WX8289), .B(II27381), .Z(II27383) ) ;
NAND2   gate16293  (.A(WX8362), .B(WX8291), .Z(II27394) ) ;
NAND2   gate16294  (.A(WX8362), .B(II27394), .Z(II27395) ) ;
NAND2   gate16295  (.A(WX8291), .B(II27394), .Z(II27396) ) ;
NAND2   gate16296  (.A(WX8363), .B(WX8293), .Z(II27407) ) ;
NAND2   gate16297  (.A(WX8363), .B(II27407), .Z(II27408) ) ;
NAND2   gate16298  (.A(WX8293), .B(II27407), .Z(II27409) ) ;
NAND2   gate16299  (.A(WX8364), .B(WX8295), .Z(II27420) ) ;
NAND2   gate16300  (.A(WX8364), .B(II27420), .Z(II27421) ) ;
NAND2   gate16301  (.A(WX8295), .B(II27420), .Z(II27422) ) ;
NAND2   gate16302  (.A(WX8365), .B(WX8297), .Z(II27433) ) ;
NAND2   gate16303  (.A(WX8365), .B(II27433), .Z(II27434) ) ;
NAND2   gate16304  (.A(WX8297), .B(II27433), .Z(II27435) ) ;
NAND2   gate16305  (.A(WX8366), .B(WX8299), .Z(II27446) ) ;
NAND2   gate16306  (.A(WX8366), .B(II27446), .Z(II27447) ) ;
NAND2   gate16307  (.A(WX8299), .B(II27446), .Z(II27448) ) ;
NAND2   gate16308  (.A(WX8367), .B(WX8301), .Z(II27459) ) ;
NAND2   gate16309  (.A(WX8367), .B(II27459), .Z(II27460) ) ;
NAND2   gate16310  (.A(WX8301), .B(II27459), .Z(II27461) ) ;
NAND2   gate16311  (.A(WX8368), .B(WX8303), .Z(II27472) ) ;
NAND2   gate16312  (.A(WX8368), .B(II27472), .Z(II27473) ) ;
NAND2   gate16313  (.A(WX8303), .B(II27472), .Z(II27474) ) ;
NAND2   gate16314  (.A(WX8369), .B(WX8305), .Z(II27485) ) ;
NAND2   gate16315  (.A(WX8369), .B(II27485), .Z(II27486) ) ;
NAND2   gate16316  (.A(WX8305), .B(II27485), .Z(II27487) ) ;
NAND2   gate16317  (.A(WX8385), .B(CRC_OUT_3_31), .Z(II27500) ) ;
NAND2   gate16318  (.A(WX8385), .B(II27500), .Z(II27501) ) ;
NAND2   gate16319  (.A(CRC_OUT_3_31), .B(II27500), .Z(II27502) ) ;
NAND2   gate16320  (.A(II27501), .B(II27502), .Z(II27499) ) ;
NAND2   gate16321  (.A(CRC_OUT_3_15), .B(II27499), .Z(II27507) ) ;
NAND2   gate16322  (.A(CRC_OUT_3_15), .B(II27507), .Z(II27508) ) ;
NAND2   gate16323  (.A(II27499), .B(II27507), .Z(II27509) ) ;
NAND2   gate16324  (.A(WX8390), .B(CRC_OUT_3_31), .Z(II27515) ) ;
NAND2   gate16325  (.A(WX8390), .B(II27515), .Z(II27516) ) ;
NAND2   gate16326  (.A(CRC_OUT_3_31), .B(II27515), .Z(II27517) ) ;
NAND2   gate16327  (.A(II27516), .B(II27517), .Z(II27514) ) ;
NAND2   gate16328  (.A(CRC_OUT_3_10), .B(II27514), .Z(II27522) ) ;
NAND2   gate16329  (.A(CRC_OUT_3_10), .B(II27522), .Z(II27523) ) ;
NAND2   gate16330  (.A(II27514), .B(II27522), .Z(II27524) ) ;
NAND2   gate16331  (.A(WX8397), .B(CRC_OUT_3_31), .Z(II27530) ) ;
NAND2   gate16332  (.A(WX8397), .B(II27530), .Z(II27531) ) ;
NAND2   gate16333  (.A(CRC_OUT_3_31), .B(II27530), .Z(II27532) ) ;
NAND2   gate16334  (.A(II27531), .B(II27532), .Z(II27529) ) ;
NAND2   gate16335  (.A(CRC_OUT_3_3), .B(II27529), .Z(II27537) ) ;
NAND2   gate16336  (.A(CRC_OUT_3_3), .B(II27537), .Z(II27538) ) ;
NAND2   gate16337  (.A(II27529), .B(II27537), .Z(II27539) ) ;
NAND2   gate16338  (.A(WX8401), .B(CRC_OUT_3_31), .Z(II27544) ) ;
NAND2   gate16339  (.A(WX8401), .B(II27544), .Z(II27545) ) ;
NAND2   gate16340  (.A(CRC_OUT_3_31), .B(II27544), .Z(II27546) ) ;
NAND2   gate16341  (.A(WX8370), .B(CRC_OUT_3_30), .Z(II27551) ) ;
NAND2   gate16342  (.A(WX8370), .B(II27551), .Z(II27552) ) ;
NAND2   gate16343  (.A(CRC_OUT_3_30), .B(II27551), .Z(II27553) ) ;
NAND2   gate16344  (.A(WX8371), .B(CRC_OUT_3_29), .Z(II27558) ) ;
NAND2   gate16345  (.A(WX8371), .B(II27558), .Z(II27559) ) ;
NAND2   gate16346  (.A(CRC_OUT_3_29), .B(II27558), .Z(II27560) ) ;
NAND2   gate16347  (.A(WX8372), .B(CRC_OUT_3_28), .Z(II27565) ) ;
NAND2   gate16348  (.A(WX8372), .B(II27565), .Z(II27566) ) ;
NAND2   gate16349  (.A(CRC_OUT_3_28), .B(II27565), .Z(II27567) ) ;
NAND2   gate16350  (.A(WX8373), .B(CRC_OUT_3_27), .Z(II27572) ) ;
NAND2   gate16351  (.A(WX8373), .B(II27572), .Z(II27573) ) ;
NAND2   gate16352  (.A(CRC_OUT_3_27), .B(II27572), .Z(II27574) ) ;
NAND2   gate16353  (.A(WX8374), .B(CRC_OUT_3_26), .Z(II27579) ) ;
NAND2   gate16354  (.A(WX8374), .B(II27579), .Z(II27580) ) ;
NAND2   gate16355  (.A(CRC_OUT_3_26), .B(II27579), .Z(II27581) ) ;
NAND2   gate16356  (.A(WX8375), .B(CRC_OUT_3_25), .Z(II27586) ) ;
NAND2   gate16357  (.A(WX8375), .B(II27586), .Z(II27587) ) ;
NAND2   gate16358  (.A(CRC_OUT_3_25), .B(II27586), .Z(II27588) ) ;
NAND2   gate16359  (.A(WX8376), .B(CRC_OUT_3_24), .Z(II27593) ) ;
NAND2   gate16360  (.A(WX8376), .B(II27593), .Z(II27594) ) ;
NAND2   gate16361  (.A(CRC_OUT_3_24), .B(II27593), .Z(II27595) ) ;
NAND2   gate16362  (.A(WX8377), .B(CRC_OUT_3_23), .Z(II27600) ) ;
NAND2   gate16363  (.A(WX8377), .B(II27600), .Z(II27601) ) ;
NAND2   gate16364  (.A(CRC_OUT_3_23), .B(II27600), .Z(II27602) ) ;
NAND2   gate16365  (.A(WX8378), .B(CRC_OUT_3_22), .Z(II27607) ) ;
NAND2   gate16366  (.A(WX8378), .B(II27607), .Z(II27608) ) ;
NAND2   gate16367  (.A(CRC_OUT_3_22), .B(II27607), .Z(II27609) ) ;
NAND2   gate16368  (.A(WX8379), .B(CRC_OUT_3_21), .Z(II27614) ) ;
NAND2   gate16369  (.A(WX8379), .B(II27614), .Z(II27615) ) ;
NAND2   gate16370  (.A(CRC_OUT_3_21), .B(II27614), .Z(II27616) ) ;
NAND2   gate16371  (.A(WX8380), .B(CRC_OUT_3_20), .Z(II27621) ) ;
NAND2   gate16372  (.A(WX8380), .B(II27621), .Z(II27622) ) ;
NAND2   gate16373  (.A(CRC_OUT_3_20), .B(II27621), .Z(II27623) ) ;
NAND2   gate16374  (.A(WX8381), .B(CRC_OUT_3_19), .Z(II27628) ) ;
NAND2   gate16375  (.A(WX8381), .B(II27628), .Z(II27629) ) ;
NAND2   gate16376  (.A(CRC_OUT_3_19), .B(II27628), .Z(II27630) ) ;
NAND2   gate16377  (.A(WX8382), .B(CRC_OUT_3_18), .Z(II27635) ) ;
NAND2   gate16378  (.A(WX8382), .B(II27635), .Z(II27636) ) ;
NAND2   gate16379  (.A(CRC_OUT_3_18), .B(II27635), .Z(II27637) ) ;
NAND2   gate16380  (.A(WX8383), .B(CRC_OUT_3_17), .Z(II27642) ) ;
NAND2   gate16381  (.A(WX8383), .B(II27642), .Z(II27643) ) ;
NAND2   gate16382  (.A(CRC_OUT_3_17), .B(II27642), .Z(II27644) ) ;
NAND2   gate16383  (.A(WX8384), .B(CRC_OUT_3_16), .Z(II27649) ) ;
NAND2   gate16384  (.A(WX8384), .B(II27649), .Z(II27650) ) ;
NAND2   gate16385  (.A(CRC_OUT_3_16), .B(II27649), .Z(II27651) ) ;
NAND2   gate16386  (.A(WX8386), .B(CRC_OUT_3_14), .Z(II27656) ) ;
NAND2   gate16387  (.A(WX8386), .B(II27656), .Z(II27657) ) ;
NAND2   gate16388  (.A(CRC_OUT_3_14), .B(II27656), .Z(II27658) ) ;
NAND2   gate16389  (.A(WX8387), .B(CRC_OUT_3_13), .Z(II27663) ) ;
NAND2   gate16390  (.A(WX8387), .B(II27663), .Z(II27664) ) ;
NAND2   gate16391  (.A(CRC_OUT_3_13), .B(II27663), .Z(II27665) ) ;
NAND2   gate16392  (.A(WX8388), .B(CRC_OUT_3_12), .Z(II27670) ) ;
NAND2   gate16393  (.A(WX8388), .B(II27670), .Z(II27671) ) ;
NAND2   gate16394  (.A(CRC_OUT_3_12), .B(II27670), .Z(II27672) ) ;
NAND2   gate16395  (.A(WX8389), .B(CRC_OUT_3_11), .Z(II27677) ) ;
NAND2   gate16396  (.A(WX8389), .B(II27677), .Z(II27678) ) ;
NAND2   gate16397  (.A(CRC_OUT_3_11), .B(II27677), .Z(II27679) ) ;
NAND2   gate16398  (.A(WX8391), .B(CRC_OUT_3_9), .Z(II27684) ) ;
NAND2   gate16399  (.A(WX8391), .B(II27684), .Z(II27685) ) ;
NAND2   gate16400  (.A(CRC_OUT_3_9), .B(II27684), .Z(II27686) ) ;
NAND2   gate16401  (.A(WX8392), .B(CRC_OUT_3_8), .Z(II27691) ) ;
NAND2   gate16402  (.A(WX8392), .B(II27691), .Z(II27692) ) ;
NAND2   gate16403  (.A(CRC_OUT_3_8), .B(II27691), .Z(II27693) ) ;
NAND2   gate16404  (.A(WX8393), .B(CRC_OUT_3_7), .Z(II27698) ) ;
NAND2   gate16405  (.A(WX8393), .B(II27698), .Z(II27699) ) ;
NAND2   gate16406  (.A(CRC_OUT_3_7), .B(II27698), .Z(II27700) ) ;
NAND2   gate16407  (.A(WX8394), .B(CRC_OUT_3_6), .Z(II27705) ) ;
NAND2   gate16408  (.A(WX8394), .B(II27705), .Z(II27706) ) ;
NAND2   gate16409  (.A(CRC_OUT_3_6), .B(II27705), .Z(II27707) ) ;
NAND2   gate16410  (.A(WX8395), .B(CRC_OUT_3_5), .Z(II27712) ) ;
NAND2   gate16411  (.A(WX8395), .B(II27712), .Z(II27713) ) ;
NAND2   gate16412  (.A(CRC_OUT_3_5), .B(II27712), .Z(II27714) ) ;
NAND2   gate16413  (.A(WX8396), .B(CRC_OUT_3_4), .Z(II27719) ) ;
NAND2   gate16414  (.A(WX8396), .B(II27719), .Z(II27720) ) ;
NAND2   gate16415  (.A(CRC_OUT_3_4), .B(II27719), .Z(II27721) ) ;
NAND2   gate16416  (.A(WX8398), .B(CRC_OUT_3_2), .Z(II27726) ) ;
NAND2   gate16417  (.A(WX8398), .B(II27726), .Z(II27727) ) ;
NAND2   gate16418  (.A(CRC_OUT_3_2), .B(II27726), .Z(II27728) ) ;
NAND2   gate16419  (.A(WX8399), .B(CRC_OUT_3_1), .Z(II27733) ) ;
NAND2   gate16420  (.A(WX8399), .B(II27733), .Z(II27734) ) ;
NAND2   gate16421  (.A(CRC_OUT_3_1), .B(II27733), .Z(II27735) ) ;
NAND2   gate16422  (.A(WX8400), .B(CRC_OUT_3_0), .Z(II27740) ) ;
NAND2   gate16423  (.A(WX8400), .B(II27740), .Z(II27741) ) ;
NAND2   gate16424  (.A(CRC_OUT_3_0), .B(II27740), .Z(II27742) ) ;
NAND2   gate16425  (.A(WX10052), .B(WX9696), .Z(II30023) ) ;
NAND2   gate16426  (.A(WX10052), .B(II30023), .Z(II30024) ) ;
NAND2   gate16427  (.A(WX9696), .B(II30023), .Z(II30025) ) ;
NAND2   gate16428  (.A(II30024), .B(II30025), .Z(II30022) ) ;
NAND2   gate16429  (.A(WX9760), .B(II30022), .Z(II30030) ) ;
NAND2   gate16430  (.A(WX9760), .B(II30030), .Z(II30031) ) ;
NAND2   gate16431  (.A(II30022), .B(II30030), .Z(II30032) ) ;
NAND2   gate16432  (.A(II30031), .B(II30032), .Z(II30021) ) ;
NAND2   gate16433  (.A(WX9824), .B(WX9888), .Z(II30038) ) ;
NAND2   gate16434  (.A(WX9824), .B(II30038), .Z(II30039) ) ;
NAND2   gate16435  (.A(WX9888), .B(II30038), .Z(II30040) ) ;
NAND2   gate16436  (.A(II30039), .B(II30040), .Z(II30037) ) ;
NAND2   gate16437  (.A(II30021), .B(II30037), .Z(II30045) ) ;
NAND2   gate16438  (.A(II30021), .B(II30045), .Z(II30046) ) ;
NAND2   gate16439  (.A(II30037), .B(II30045), .Z(II30047) ) ;
NAND2   gate16440  (.A(WX10052), .B(WX9698), .Z(II30054) ) ;
NAND2   gate16441  (.A(WX10052), .B(II30054), .Z(II30055) ) ;
NAND2   gate16442  (.A(WX9698), .B(II30054), .Z(II30056) ) ;
NAND2   gate16443  (.A(II30055), .B(II30056), .Z(II30053) ) ;
NAND2   gate16444  (.A(WX9762), .B(II30053), .Z(II30061) ) ;
NAND2   gate16445  (.A(WX9762), .B(II30061), .Z(II30062) ) ;
NAND2   gate16446  (.A(II30053), .B(II30061), .Z(II30063) ) ;
NAND2   gate16447  (.A(II30062), .B(II30063), .Z(II30052) ) ;
NAND2   gate16448  (.A(WX9826), .B(WX9890), .Z(II30069) ) ;
NAND2   gate16449  (.A(WX9826), .B(II30069), .Z(II30070) ) ;
NAND2   gate16450  (.A(WX9890), .B(II30069), .Z(II30071) ) ;
NAND2   gate16451  (.A(II30070), .B(II30071), .Z(II30068) ) ;
NAND2   gate16452  (.A(II30052), .B(II30068), .Z(II30076) ) ;
NAND2   gate16453  (.A(II30052), .B(II30076), .Z(II30077) ) ;
NAND2   gate16454  (.A(II30068), .B(II30076), .Z(II30078) ) ;
NAND2   gate16455  (.A(WX10052), .B(WX9700), .Z(II30085) ) ;
NAND2   gate16456  (.A(WX10052), .B(II30085), .Z(II30086) ) ;
NAND2   gate16457  (.A(WX9700), .B(II30085), .Z(II30087) ) ;
NAND2   gate16458  (.A(II30086), .B(II30087), .Z(II30084) ) ;
NAND2   gate16459  (.A(WX9764), .B(II30084), .Z(II30092) ) ;
NAND2   gate16460  (.A(WX9764), .B(II30092), .Z(II30093) ) ;
NAND2   gate16461  (.A(II30084), .B(II30092), .Z(II30094) ) ;
NAND2   gate16462  (.A(II30093), .B(II30094), .Z(II30083) ) ;
NAND2   gate16463  (.A(WX9828), .B(WX9892), .Z(II30100) ) ;
NAND2   gate16464  (.A(WX9828), .B(II30100), .Z(II30101) ) ;
NAND2   gate16465  (.A(WX9892), .B(II30100), .Z(II30102) ) ;
NAND2   gate16466  (.A(II30101), .B(II30102), .Z(II30099) ) ;
NAND2   gate16467  (.A(II30083), .B(II30099), .Z(II30107) ) ;
NAND2   gate16468  (.A(II30083), .B(II30107), .Z(II30108) ) ;
NAND2   gate16469  (.A(II30099), .B(II30107), .Z(II30109) ) ;
NAND2   gate16470  (.A(WX10052), .B(WX9702), .Z(II30116) ) ;
NAND2   gate16471  (.A(WX10052), .B(II30116), .Z(II30117) ) ;
NAND2   gate16472  (.A(WX9702), .B(II30116), .Z(II30118) ) ;
NAND2   gate16473  (.A(II30117), .B(II30118), .Z(II30115) ) ;
NAND2   gate16474  (.A(WX9766), .B(II30115), .Z(II30123) ) ;
NAND2   gate16475  (.A(WX9766), .B(II30123), .Z(II30124) ) ;
NAND2   gate16476  (.A(II30115), .B(II30123), .Z(II30125) ) ;
NAND2   gate16477  (.A(II30124), .B(II30125), .Z(II30114) ) ;
NAND2   gate16478  (.A(WX9830), .B(WX9894), .Z(II30131) ) ;
NAND2   gate16479  (.A(WX9830), .B(II30131), .Z(II30132) ) ;
NAND2   gate16480  (.A(WX9894), .B(II30131), .Z(II30133) ) ;
NAND2   gate16481  (.A(II30132), .B(II30133), .Z(II30130) ) ;
NAND2   gate16482  (.A(II30114), .B(II30130), .Z(II30138) ) ;
NAND2   gate16483  (.A(II30114), .B(II30138), .Z(II30139) ) ;
NAND2   gate16484  (.A(II30130), .B(II30138), .Z(II30140) ) ;
NAND2   gate16485  (.A(WX10052), .B(WX9704), .Z(II30147) ) ;
NAND2   gate16486  (.A(WX10052), .B(II30147), .Z(II30148) ) ;
NAND2   gate16487  (.A(WX9704), .B(II30147), .Z(II30149) ) ;
NAND2   gate16488  (.A(II30148), .B(II30149), .Z(II30146) ) ;
NAND2   gate16489  (.A(WX9768), .B(II30146), .Z(II30154) ) ;
NAND2   gate16490  (.A(WX9768), .B(II30154), .Z(II30155) ) ;
NAND2   gate16491  (.A(II30146), .B(II30154), .Z(II30156) ) ;
NAND2   gate16492  (.A(II30155), .B(II30156), .Z(II30145) ) ;
NAND2   gate16493  (.A(WX9832), .B(WX9896), .Z(II30162) ) ;
NAND2   gate16494  (.A(WX9832), .B(II30162), .Z(II30163) ) ;
NAND2   gate16495  (.A(WX9896), .B(II30162), .Z(II30164) ) ;
NAND2   gate16496  (.A(II30163), .B(II30164), .Z(II30161) ) ;
NAND2   gate16497  (.A(II30145), .B(II30161), .Z(II30169) ) ;
NAND2   gate16498  (.A(II30145), .B(II30169), .Z(II30170) ) ;
NAND2   gate16499  (.A(II30161), .B(II30169), .Z(II30171) ) ;
NAND2   gate16500  (.A(WX10052), .B(WX9706), .Z(II30178) ) ;
NAND2   gate16501  (.A(WX10052), .B(II30178), .Z(II30179) ) ;
NAND2   gate16502  (.A(WX9706), .B(II30178), .Z(II30180) ) ;
NAND2   gate16503  (.A(II30179), .B(II30180), .Z(II30177) ) ;
NAND2   gate16504  (.A(WX9770), .B(II30177), .Z(II30185) ) ;
NAND2   gate16505  (.A(WX9770), .B(II30185), .Z(II30186) ) ;
NAND2   gate16506  (.A(II30177), .B(II30185), .Z(II30187) ) ;
NAND2   gate16507  (.A(II30186), .B(II30187), .Z(II30176) ) ;
NAND2   gate16508  (.A(WX9834), .B(WX9898), .Z(II30193) ) ;
NAND2   gate16509  (.A(WX9834), .B(II30193), .Z(II30194) ) ;
NAND2   gate16510  (.A(WX9898), .B(II30193), .Z(II30195) ) ;
NAND2   gate16511  (.A(II30194), .B(II30195), .Z(II30192) ) ;
NAND2   gate16512  (.A(II30176), .B(II30192), .Z(II30200) ) ;
NAND2   gate16513  (.A(II30176), .B(II30200), .Z(II30201) ) ;
NAND2   gate16514  (.A(II30192), .B(II30200), .Z(II30202) ) ;
NAND2   gate16515  (.A(WX10052), .B(WX9708), .Z(II30209) ) ;
NAND2   gate16516  (.A(WX10052), .B(II30209), .Z(II30210) ) ;
NAND2   gate16517  (.A(WX9708), .B(II30209), .Z(II30211) ) ;
NAND2   gate16518  (.A(II30210), .B(II30211), .Z(II30208) ) ;
NAND2   gate16519  (.A(WX9772), .B(II30208), .Z(II30216) ) ;
NAND2   gate16520  (.A(WX9772), .B(II30216), .Z(II30217) ) ;
NAND2   gate16521  (.A(II30208), .B(II30216), .Z(II30218) ) ;
NAND2   gate16522  (.A(II30217), .B(II30218), .Z(II30207) ) ;
NAND2   gate16523  (.A(WX9836), .B(WX9900), .Z(II30224) ) ;
NAND2   gate16524  (.A(WX9836), .B(II30224), .Z(II30225) ) ;
NAND2   gate16525  (.A(WX9900), .B(II30224), .Z(II30226) ) ;
NAND2   gate16526  (.A(II30225), .B(II30226), .Z(II30223) ) ;
NAND2   gate16527  (.A(II30207), .B(II30223), .Z(II30231) ) ;
NAND2   gate16528  (.A(II30207), .B(II30231), .Z(II30232) ) ;
NAND2   gate16529  (.A(II30223), .B(II30231), .Z(II30233) ) ;
NAND2   gate16530  (.A(WX10052), .B(WX9710), .Z(II30240) ) ;
NAND2   gate16531  (.A(WX10052), .B(II30240), .Z(II30241) ) ;
NAND2   gate16532  (.A(WX9710), .B(II30240), .Z(II30242) ) ;
NAND2   gate16533  (.A(II30241), .B(II30242), .Z(II30239) ) ;
NAND2   gate16534  (.A(WX9774), .B(II30239), .Z(II30247) ) ;
NAND2   gate16535  (.A(WX9774), .B(II30247), .Z(II30248) ) ;
NAND2   gate16536  (.A(II30239), .B(II30247), .Z(II30249) ) ;
NAND2   gate16537  (.A(II30248), .B(II30249), .Z(II30238) ) ;
NAND2   gate16538  (.A(WX9838), .B(WX9902), .Z(II30255) ) ;
NAND2   gate16539  (.A(WX9838), .B(II30255), .Z(II30256) ) ;
NAND2   gate16540  (.A(WX9902), .B(II30255), .Z(II30257) ) ;
NAND2   gate16541  (.A(II30256), .B(II30257), .Z(II30254) ) ;
NAND2   gate16542  (.A(II30238), .B(II30254), .Z(II30262) ) ;
NAND2   gate16543  (.A(II30238), .B(II30262), .Z(II30263) ) ;
NAND2   gate16544  (.A(II30254), .B(II30262), .Z(II30264) ) ;
NAND2   gate16545  (.A(WX10052), .B(WX9712), .Z(II30271) ) ;
NAND2   gate16546  (.A(WX10052), .B(II30271), .Z(II30272) ) ;
NAND2   gate16547  (.A(WX9712), .B(II30271), .Z(II30273) ) ;
NAND2   gate16548  (.A(II30272), .B(II30273), .Z(II30270) ) ;
NAND2   gate16549  (.A(WX9776), .B(II30270), .Z(II30278) ) ;
NAND2   gate16550  (.A(WX9776), .B(II30278), .Z(II30279) ) ;
NAND2   gate16551  (.A(II30270), .B(II30278), .Z(II30280) ) ;
NAND2   gate16552  (.A(II30279), .B(II30280), .Z(II30269) ) ;
NAND2   gate16553  (.A(WX9840), .B(WX9904), .Z(II30286) ) ;
NAND2   gate16554  (.A(WX9840), .B(II30286), .Z(II30287) ) ;
NAND2   gate16555  (.A(WX9904), .B(II30286), .Z(II30288) ) ;
NAND2   gate16556  (.A(II30287), .B(II30288), .Z(II30285) ) ;
NAND2   gate16557  (.A(II30269), .B(II30285), .Z(II30293) ) ;
NAND2   gate16558  (.A(II30269), .B(II30293), .Z(II30294) ) ;
NAND2   gate16559  (.A(II30285), .B(II30293), .Z(II30295) ) ;
NAND2   gate16560  (.A(WX10052), .B(WX9714), .Z(II30302) ) ;
NAND2   gate16561  (.A(WX10052), .B(II30302), .Z(II30303) ) ;
NAND2   gate16562  (.A(WX9714), .B(II30302), .Z(II30304) ) ;
NAND2   gate16563  (.A(II30303), .B(II30304), .Z(II30301) ) ;
NAND2   gate16564  (.A(WX9778), .B(II30301), .Z(II30309) ) ;
NAND2   gate16565  (.A(WX9778), .B(II30309), .Z(II30310) ) ;
NAND2   gate16566  (.A(II30301), .B(II30309), .Z(II30311) ) ;
NAND2   gate16567  (.A(II30310), .B(II30311), .Z(II30300) ) ;
NAND2   gate16568  (.A(WX9842), .B(WX9906), .Z(II30317) ) ;
NAND2   gate16569  (.A(WX9842), .B(II30317), .Z(II30318) ) ;
NAND2   gate16570  (.A(WX9906), .B(II30317), .Z(II30319) ) ;
NAND2   gate16571  (.A(II30318), .B(II30319), .Z(II30316) ) ;
NAND2   gate16572  (.A(II30300), .B(II30316), .Z(II30324) ) ;
NAND2   gate16573  (.A(II30300), .B(II30324), .Z(II30325) ) ;
NAND2   gate16574  (.A(II30316), .B(II30324), .Z(II30326) ) ;
NAND2   gate16575  (.A(WX10052), .B(WX9716), .Z(II30333) ) ;
NAND2   gate16576  (.A(WX10052), .B(II30333), .Z(II30334) ) ;
NAND2   gate16577  (.A(WX9716), .B(II30333), .Z(II30335) ) ;
NAND2   gate16578  (.A(II30334), .B(II30335), .Z(II30332) ) ;
NAND2   gate16579  (.A(WX9780), .B(II30332), .Z(II30340) ) ;
NAND2   gate16580  (.A(WX9780), .B(II30340), .Z(II30341) ) ;
NAND2   gate16581  (.A(II30332), .B(II30340), .Z(II30342) ) ;
NAND2   gate16582  (.A(II30341), .B(II30342), .Z(II30331) ) ;
NAND2   gate16583  (.A(WX9844), .B(WX9908), .Z(II30348) ) ;
NAND2   gate16584  (.A(WX9844), .B(II30348), .Z(II30349) ) ;
NAND2   gate16585  (.A(WX9908), .B(II30348), .Z(II30350) ) ;
NAND2   gate16586  (.A(II30349), .B(II30350), .Z(II30347) ) ;
NAND2   gate16587  (.A(II30331), .B(II30347), .Z(II30355) ) ;
NAND2   gate16588  (.A(II30331), .B(II30355), .Z(II30356) ) ;
NAND2   gate16589  (.A(II30347), .B(II30355), .Z(II30357) ) ;
NAND2   gate16590  (.A(WX10052), .B(WX9718), .Z(II30364) ) ;
NAND2   gate16591  (.A(WX10052), .B(II30364), .Z(II30365) ) ;
NAND2   gate16592  (.A(WX9718), .B(II30364), .Z(II30366) ) ;
NAND2   gate16593  (.A(II30365), .B(II30366), .Z(II30363) ) ;
NAND2   gate16594  (.A(WX9782), .B(II30363), .Z(II30371) ) ;
NAND2   gate16595  (.A(WX9782), .B(II30371), .Z(II30372) ) ;
NAND2   gate16596  (.A(II30363), .B(II30371), .Z(II30373) ) ;
NAND2   gate16597  (.A(II30372), .B(II30373), .Z(II30362) ) ;
NAND2   gate16598  (.A(WX9846), .B(WX9910), .Z(II30379) ) ;
NAND2   gate16599  (.A(WX9846), .B(II30379), .Z(II30380) ) ;
NAND2   gate16600  (.A(WX9910), .B(II30379), .Z(II30381) ) ;
NAND2   gate16601  (.A(II30380), .B(II30381), .Z(II30378) ) ;
NAND2   gate16602  (.A(II30362), .B(II30378), .Z(II30386) ) ;
NAND2   gate16603  (.A(II30362), .B(II30386), .Z(II30387) ) ;
NAND2   gate16604  (.A(II30378), .B(II30386), .Z(II30388) ) ;
NAND2   gate16605  (.A(WX10052), .B(WX9720), .Z(II30395) ) ;
NAND2   gate16606  (.A(WX10052), .B(II30395), .Z(II30396) ) ;
NAND2   gate16607  (.A(WX9720), .B(II30395), .Z(II30397) ) ;
NAND2   gate16608  (.A(II30396), .B(II30397), .Z(II30394) ) ;
NAND2   gate16609  (.A(WX9784), .B(II30394), .Z(II30402) ) ;
NAND2   gate16610  (.A(WX9784), .B(II30402), .Z(II30403) ) ;
NAND2   gate16611  (.A(II30394), .B(II30402), .Z(II30404) ) ;
NAND2   gate16612  (.A(II30403), .B(II30404), .Z(II30393) ) ;
NAND2   gate16613  (.A(WX9848), .B(WX9912), .Z(II30410) ) ;
NAND2   gate16614  (.A(WX9848), .B(II30410), .Z(II30411) ) ;
NAND2   gate16615  (.A(WX9912), .B(II30410), .Z(II30412) ) ;
NAND2   gate16616  (.A(II30411), .B(II30412), .Z(II30409) ) ;
NAND2   gate16617  (.A(II30393), .B(II30409), .Z(II30417) ) ;
NAND2   gate16618  (.A(II30393), .B(II30417), .Z(II30418) ) ;
NAND2   gate16619  (.A(II30409), .B(II30417), .Z(II30419) ) ;
NAND2   gate16620  (.A(WX10052), .B(WX9722), .Z(II30426) ) ;
NAND2   gate16621  (.A(WX10052), .B(II30426), .Z(II30427) ) ;
NAND2   gate16622  (.A(WX9722), .B(II30426), .Z(II30428) ) ;
NAND2   gate16623  (.A(II30427), .B(II30428), .Z(II30425) ) ;
NAND2   gate16624  (.A(WX9786), .B(II30425), .Z(II30433) ) ;
NAND2   gate16625  (.A(WX9786), .B(II30433), .Z(II30434) ) ;
NAND2   gate16626  (.A(II30425), .B(II30433), .Z(II30435) ) ;
NAND2   gate16627  (.A(II30434), .B(II30435), .Z(II30424) ) ;
NAND2   gate16628  (.A(WX9850), .B(WX9914), .Z(II30441) ) ;
NAND2   gate16629  (.A(WX9850), .B(II30441), .Z(II30442) ) ;
NAND2   gate16630  (.A(WX9914), .B(II30441), .Z(II30443) ) ;
NAND2   gate16631  (.A(II30442), .B(II30443), .Z(II30440) ) ;
NAND2   gate16632  (.A(II30424), .B(II30440), .Z(II30448) ) ;
NAND2   gate16633  (.A(II30424), .B(II30448), .Z(II30449) ) ;
NAND2   gate16634  (.A(II30440), .B(II30448), .Z(II30450) ) ;
NAND2   gate16635  (.A(WX10052), .B(WX9724), .Z(II30457) ) ;
NAND2   gate16636  (.A(WX10052), .B(II30457), .Z(II30458) ) ;
NAND2   gate16637  (.A(WX9724), .B(II30457), .Z(II30459) ) ;
NAND2   gate16638  (.A(II30458), .B(II30459), .Z(II30456) ) ;
NAND2   gate16639  (.A(WX9788), .B(II30456), .Z(II30464) ) ;
NAND2   gate16640  (.A(WX9788), .B(II30464), .Z(II30465) ) ;
NAND2   gate16641  (.A(II30456), .B(II30464), .Z(II30466) ) ;
NAND2   gate16642  (.A(II30465), .B(II30466), .Z(II30455) ) ;
NAND2   gate16643  (.A(WX9852), .B(WX9916), .Z(II30472) ) ;
NAND2   gate16644  (.A(WX9852), .B(II30472), .Z(II30473) ) ;
NAND2   gate16645  (.A(WX9916), .B(II30472), .Z(II30474) ) ;
NAND2   gate16646  (.A(II30473), .B(II30474), .Z(II30471) ) ;
NAND2   gate16647  (.A(II30455), .B(II30471), .Z(II30479) ) ;
NAND2   gate16648  (.A(II30455), .B(II30479), .Z(II30480) ) ;
NAND2   gate16649  (.A(II30471), .B(II30479), .Z(II30481) ) ;
NAND2   gate16650  (.A(WX10052), .B(WX9726), .Z(II30488) ) ;
NAND2   gate16651  (.A(WX10052), .B(II30488), .Z(II30489) ) ;
NAND2   gate16652  (.A(WX9726), .B(II30488), .Z(II30490) ) ;
NAND2   gate16653  (.A(II30489), .B(II30490), .Z(II30487) ) ;
NAND2   gate16654  (.A(WX9790), .B(II30487), .Z(II30495) ) ;
NAND2   gate16655  (.A(WX9790), .B(II30495), .Z(II30496) ) ;
NAND2   gate16656  (.A(II30487), .B(II30495), .Z(II30497) ) ;
NAND2   gate16657  (.A(II30496), .B(II30497), .Z(II30486) ) ;
NAND2   gate16658  (.A(WX9854), .B(WX9918), .Z(II30503) ) ;
NAND2   gate16659  (.A(WX9854), .B(II30503), .Z(II30504) ) ;
NAND2   gate16660  (.A(WX9918), .B(II30503), .Z(II30505) ) ;
NAND2   gate16661  (.A(II30504), .B(II30505), .Z(II30502) ) ;
NAND2   gate16662  (.A(II30486), .B(II30502), .Z(II30510) ) ;
NAND2   gate16663  (.A(II30486), .B(II30510), .Z(II30511) ) ;
NAND2   gate16664  (.A(II30502), .B(II30510), .Z(II30512) ) ;
NAND2   gate16665  (.A(WX10053), .B(WX9728), .Z(II30519) ) ;
NAND2   gate16666  (.A(WX10053), .B(II30519), .Z(II30520) ) ;
NAND2   gate16667  (.A(WX9728), .B(II30519), .Z(II30521) ) ;
NAND2   gate16668  (.A(II30520), .B(II30521), .Z(II30518) ) ;
NAND2   gate16669  (.A(WX9792), .B(II30518), .Z(II30526) ) ;
NAND2   gate16670  (.A(WX9792), .B(II30526), .Z(II30527) ) ;
NAND2   gate16671  (.A(II30518), .B(II30526), .Z(II30528) ) ;
NAND2   gate16672  (.A(II30527), .B(II30528), .Z(II30517) ) ;
NAND2   gate16673  (.A(WX9856), .B(WX9920), .Z(II30534) ) ;
NAND2   gate16674  (.A(WX9856), .B(II30534), .Z(II30535) ) ;
NAND2   gate16675  (.A(WX9920), .B(II30534), .Z(II30536) ) ;
NAND2   gate16676  (.A(II30535), .B(II30536), .Z(II30533) ) ;
NAND2   gate16677  (.A(II30517), .B(II30533), .Z(II30541) ) ;
NAND2   gate16678  (.A(II30517), .B(II30541), .Z(II30542) ) ;
NAND2   gate16679  (.A(II30533), .B(II30541), .Z(II30543) ) ;
NAND2   gate16680  (.A(WX10053), .B(WX9730), .Z(II30550) ) ;
NAND2   gate16681  (.A(WX10053), .B(II30550), .Z(II30551) ) ;
NAND2   gate16682  (.A(WX9730), .B(II30550), .Z(II30552) ) ;
NAND2   gate16683  (.A(II30551), .B(II30552), .Z(II30549) ) ;
NAND2   gate16684  (.A(WX9794), .B(II30549), .Z(II30557) ) ;
NAND2   gate16685  (.A(WX9794), .B(II30557), .Z(II30558) ) ;
NAND2   gate16686  (.A(II30549), .B(II30557), .Z(II30559) ) ;
NAND2   gate16687  (.A(II30558), .B(II30559), .Z(II30548) ) ;
NAND2   gate16688  (.A(WX9858), .B(WX9922), .Z(II30565) ) ;
NAND2   gate16689  (.A(WX9858), .B(II30565), .Z(II30566) ) ;
NAND2   gate16690  (.A(WX9922), .B(II30565), .Z(II30567) ) ;
NAND2   gate16691  (.A(II30566), .B(II30567), .Z(II30564) ) ;
NAND2   gate16692  (.A(II30548), .B(II30564), .Z(II30572) ) ;
NAND2   gate16693  (.A(II30548), .B(II30572), .Z(II30573) ) ;
NAND2   gate16694  (.A(II30564), .B(II30572), .Z(II30574) ) ;
NAND2   gate16695  (.A(WX10053), .B(WX9732), .Z(II30581) ) ;
NAND2   gate16696  (.A(WX10053), .B(II30581), .Z(II30582) ) ;
NAND2   gate16697  (.A(WX9732), .B(II30581), .Z(II30583) ) ;
NAND2   gate16698  (.A(II30582), .B(II30583), .Z(II30580) ) ;
NAND2   gate16699  (.A(WX9796), .B(II30580), .Z(II30588) ) ;
NAND2   gate16700  (.A(WX9796), .B(II30588), .Z(II30589) ) ;
NAND2   gate16701  (.A(II30580), .B(II30588), .Z(II30590) ) ;
NAND2   gate16702  (.A(II30589), .B(II30590), .Z(II30579) ) ;
NAND2   gate16703  (.A(WX9860), .B(WX9924), .Z(II30596) ) ;
NAND2   gate16704  (.A(WX9860), .B(II30596), .Z(II30597) ) ;
NAND2   gate16705  (.A(WX9924), .B(II30596), .Z(II30598) ) ;
NAND2   gate16706  (.A(II30597), .B(II30598), .Z(II30595) ) ;
NAND2   gate16707  (.A(II30579), .B(II30595), .Z(II30603) ) ;
NAND2   gate16708  (.A(II30579), .B(II30603), .Z(II30604) ) ;
NAND2   gate16709  (.A(II30595), .B(II30603), .Z(II30605) ) ;
NAND2   gate16710  (.A(WX10053), .B(WX9734), .Z(II30612) ) ;
NAND2   gate16711  (.A(WX10053), .B(II30612), .Z(II30613) ) ;
NAND2   gate16712  (.A(WX9734), .B(II30612), .Z(II30614) ) ;
NAND2   gate16713  (.A(II30613), .B(II30614), .Z(II30611) ) ;
NAND2   gate16714  (.A(WX9798), .B(II30611), .Z(II30619) ) ;
NAND2   gate16715  (.A(WX9798), .B(II30619), .Z(II30620) ) ;
NAND2   gate16716  (.A(II30611), .B(II30619), .Z(II30621) ) ;
NAND2   gate16717  (.A(II30620), .B(II30621), .Z(II30610) ) ;
NAND2   gate16718  (.A(WX9862), .B(WX9926), .Z(II30627) ) ;
NAND2   gate16719  (.A(WX9862), .B(II30627), .Z(II30628) ) ;
NAND2   gate16720  (.A(WX9926), .B(II30627), .Z(II30629) ) ;
NAND2   gate16721  (.A(II30628), .B(II30629), .Z(II30626) ) ;
NAND2   gate16722  (.A(II30610), .B(II30626), .Z(II30634) ) ;
NAND2   gate16723  (.A(II30610), .B(II30634), .Z(II30635) ) ;
NAND2   gate16724  (.A(II30626), .B(II30634), .Z(II30636) ) ;
NAND2   gate16725  (.A(WX10053), .B(WX9736), .Z(II30643) ) ;
NAND2   gate16726  (.A(WX10053), .B(II30643), .Z(II30644) ) ;
NAND2   gate16727  (.A(WX9736), .B(II30643), .Z(II30645) ) ;
NAND2   gate16728  (.A(II30644), .B(II30645), .Z(II30642) ) ;
NAND2   gate16729  (.A(WX9800), .B(II30642), .Z(II30650) ) ;
NAND2   gate16730  (.A(WX9800), .B(II30650), .Z(II30651) ) ;
NAND2   gate16731  (.A(II30642), .B(II30650), .Z(II30652) ) ;
NAND2   gate16732  (.A(II30651), .B(II30652), .Z(II30641) ) ;
NAND2   gate16733  (.A(WX9864), .B(WX9928), .Z(II30658) ) ;
NAND2   gate16734  (.A(WX9864), .B(II30658), .Z(II30659) ) ;
NAND2   gate16735  (.A(WX9928), .B(II30658), .Z(II30660) ) ;
NAND2   gate16736  (.A(II30659), .B(II30660), .Z(II30657) ) ;
NAND2   gate16737  (.A(II30641), .B(II30657), .Z(II30665) ) ;
NAND2   gate16738  (.A(II30641), .B(II30665), .Z(II30666) ) ;
NAND2   gate16739  (.A(II30657), .B(II30665), .Z(II30667) ) ;
NAND2   gate16740  (.A(WX10053), .B(WX9738), .Z(II30674) ) ;
NAND2   gate16741  (.A(WX10053), .B(II30674), .Z(II30675) ) ;
NAND2   gate16742  (.A(WX9738), .B(II30674), .Z(II30676) ) ;
NAND2   gate16743  (.A(II30675), .B(II30676), .Z(II30673) ) ;
NAND2   gate16744  (.A(WX9802), .B(II30673), .Z(II30681) ) ;
NAND2   gate16745  (.A(WX9802), .B(II30681), .Z(II30682) ) ;
NAND2   gate16746  (.A(II30673), .B(II30681), .Z(II30683) ) ;
NAND2   gate16747  (.A(II30682), .B(II30683), .Z(II30672) ) ;
NAND2   gate16748  (.A(WX9866), .B(WX9930), .Z(II30689) ) ;
NAND2   gate16749  (.A(WX9866), .B(II30689), .Z(II30690) ) ;
NAND2   gate16750  (.A(WX9930), .B(II30689), .Z(II30691) ) ;
NAND2   gate16751  (.A(II30690), .B(II30691), .Z(II30688) ) ;
NAND2   gate16752  (.A(II30672), .B(II30688), .Z(II30696) ) ;
NAND2   gate16753  (.A(II30672), .B(II30696), .Z(II30697) ) ;
NAND2   gate16754  (.A(II30688), .B(II30696), .Z(II30698) ) ;
NAND2   gate16755  (.A(WX10053), .B(WX9740), .Z(II30705) ) ;
NAND2   gate16756  (.A(WX10053), .B(II30705), .Z(II30706) ) ;
NAND2   gate16757  (.A(WX9740), .B(II30705), .Z(II30707) ) ;
NAND2   gate16758  (.A(II30706), .B(II30707), .Z(II30704) ) ;
NAND2   gate16759  (.A(WX9804), .B(II30704), .Z(II30712) ) ;
NAND2   gate16760  (.A(WX9804), .B(II30712), .Z(II30713) ) ;
NAND2   gate16761  (.A(II30704), .B(II30712), .Z(II30714) ) ;
NAND2   gate16762  (.A(II30713), .B(II30714), .Z(II30703) ) ;
NAND2   gate16763  (.A(WX9868), .B(WX9932), .Z(II30720) ) ;
NAND2   gate16764  (.A(WX9868), .B(II30720), .Z(II30721) ) ;
NAND2   gate16765  (.A(WX9932), .B(II30720), .Z(II30722) ) ;
NAND2   gate16766  (.A(II30721), .B(II30722), .Z(II30719) ) ;
NAND2   gate16767  (.A(II30703), .B(II30719), .Z(II30727) ) ;
NAND2   gate16768  (.A(II30703), .B(II30727), .Z(II30728) ) ;
NAND2   gate16769  (.A(II30719), .B(II30727), .Z(II30729) ) ;
NAND2   gate16770  (.A(WX10053), .B(WX9742), .Z(II30736) ) ;
NAND2   gate16771  (.A(WX10053), .B(II30736), .Z(II30737) ) ;
NAND2   gate16772  (.A(WX9742), .B(II30736), .Z(II30738) ) ;
NAND2   gate16773  (.A(II30737), .B(II30738), .Z(II30735) ) ;
NAND2   gate16774  (.A(WX9806), .B(II30735), .Z(II30743) ) ;
NAND2   gate16775  (.A(WX9806), .B(II30743), .Z(II30744) ) ;
NAND2   gate16776  (.A(II30735), .B(II30743), .Z(II30745) ) ;
NAND2   gate16777  (.A(II30744), .B(II30745), .Z(II30734) ) ;
NAND2   gate16778  (.A(WX9870), .B(WX9934), .Z(II30751) ) ;
NAND2   gate16779  (.A(WX9870), .B(II30751), .Z(II30752) ) ;
NAND2   gate16780  (.A(WX9934), .B(II30751), .Z(II30753) ) ;
NAND2   gate16781  (.A(II30752), .B(II30753), .Z(II30750) ) ;
NAND2   gate16782  (.A(II30734), .B(II30750), .Z(II30758) ) ;
NAND2   gate16783  (.A(II30734), .B(II30758), .Z(II30759) ) ;
NAND2   gate16784  (.A(II30750), .B(II30758), .Z(II30760) ) ;
NAND2   gate16785  (.A(WX10053), .B(WX9744), .Z(II30767) ) ;
NAND2   gate16786  (.A(WX10053), .B(II30767), .Z(II30768) ) ;
NAND2   gate16787  (.A(WX9744), .B(II30767), .Z(II30769) ) ;
NAND2   gate16788  (.A(II30768), .B(II30769), .Z(II30766) ) ;
NAND2   gate16789  (.A(WX9808), .B(II30766), .Z(II30774) ) ;
NAND2   gate16790  (.A(WX9808), .B(II30774), .Z(II30775) ) ;
NAND2   gate16791  (.A(II30766), .B(II30774), .Z(II30776) ) ;
NAND2   gate16792  (.A(II30775), .B(II30776), .Z(II30765) ) ;
NAND2   gate16793  (.A(WX9872), .B(WX9936), .Z(II30782) ) ;
NAND2   gate16794  (.A(WX9872), .B(II30782), .Z(II30783) ) ;
NAND2   gate16795  (.A(WX9936), .B(II30782), .Z(II30784) ) ;
NAND2   gate16796  (.A(II30783), .B(II30784), .Z(II30781) ) ;
NAND2   gate16797  (.A(II30765), .B(II30781), .Z(II30789) ) ;
NAND2   gate16798  (.A(II30765), .B(II30789), .Z(II30790) ) ;
NAND2   gate16799  (.A(II30781), .B(II30789), .Z(II30791) ) ;
NAND2   gate16800  (.A(WX10053), .B(WX9746), .Z(II30798) ) ;
NAND2   gate16801  (.A(WX10053), .B(II30798), .Z(II30799) ) ;
NAND2   gate16802  (.A(WX9746), .B(II30798), .Z(II30800) ) ;
NAND2   gate16803  (.A(II30799), .B(II30800), .Z(II30797) ) ;
NAND2   gate16804  (.A(WX9810), .B(II30797), .Z(II30805) ) ;
NAND2   gate16805  (.A(WX9810), .B(II30805), .Z(II30806) ) ;
NAND2   gate16806  (.A(II30797), .B(II30805), .Z(II30807) ) ;
NAND2   gate16807  (.A(II30806), .B(II30807), .Z(II30796) ) ;
NAND2   gate16808  (.A(WX9874), .B(WX9938), .Z(II30813) ) ;
NAND2   gate16809  (.A(WX9874), .B(II30813), .Z(II30814) ) ;
NAND2   gate16810  (.A(WX9938), .B(II30813), .Z(II30815) ) ;
NAND2   gate16811  (.A(II30814), .B(II30815), .Z(II30812) ) ;
NAND2   gate16812  (.A(II30796), .B(II30812), .Z(II30820) ) ;
NAND2   gate16813  (.A(II30796), .B(II30820), .Z(II30821) ) ;
NAND2   gate16814  (.A(II30812), .B(II30820), .Z(II30822) ) ;
NAND2   gate16815  (.A(WX10053), .B(WX9748), .Z(II30829) ) ;
NAND2   gate16816  (.A(WX10053), .B(II30829), .Z(II30830) ) ;
NAND2   gate16817  (.A(WX9748), .B(II30829), .Z(II30831) ) ;
NAND2   gate16818  (.A(II30830), .B(II30831), .Z(II30828) ) ;
NAND2   gate16819  (.A(WX9812), .B(II30828), .Z(II30836) ) ;
NAND2   gate16820  (.A(WX9812), .B(II30836), .Z(II30837) ) ;
NAND2   gate16821  (.A(II30828), .B(II30836), .Z(II30838) ) ;
NAND2   gate16822  (.A(II30837), .B(II30838), .Z(II30827) ) ;
NAND2   gate16823  (.A(WX9876), .B(WX9940), .Z(II30844) ) ;
NAND2   gate16824  (.A(WX9876), .B(II30844), .Z(II30845) ) ;
NAND2   gate16825  (.A(WX9940), .B(II30844), .Z(II30846) ) ;
NAND2   gate16826  (.A(II30845), .B(II30846), .Z(II30843) ) ;
NAND2   gate16827  (.A(II30827), .B(II30843), .Z(II30851) ) ;
NAND2   gate16828  (.A(II30827), .B(II30851), .Z(II30852) ) ;
NAND2   gate16829  (.A(II30843), .B(II30851), .Z(II30853) ) ;
NAND2   gate16830  (.A(WX10053), .B(WX9750), .Z(II30860) ) ;
NAND2   gate16831  (.A(WX10053), .B(II30860), .Z(II30861) ) ;
NAND2   gate16832  (.A(WX9750), .B(II30860), .Z(II30862) ) ;
NAND2   gate16833  (.A(II30861), .B(II30862), .Z(II30859) ) ;
NAND2   gate16834  (.A(WX9814), .B(II30859), .Z(II30867) ) ;
NAND2   gate16835  (.A(WX9814), .B(II30867), .Z(II30868) ) ;
NAND2   gate16836  (.A(II30859), .B(II30867), .Z(II30869) ) ;
NAND2   gate16837  (.A(II30868), .B(II30869), .Z(II30858) ) ;
NAND2   gate16838  (.A(WX9878), .B(WX9942), .Z(II30875) ) ;
NAND2   gate16839  (.A(WX9878), .B(II30875), .Z(II30876) ) ;
NAND2   gate16840  (.A(WX9942), .B(II30875), .Z(II30877) ) ;
NAND2   gate16841  (.A(II30876), .B(II30877), .Z(II30874) ) ;
NAND2   gate16842  (.A(II30858), .B(II30874), .Z(II30882) ) ;
NAND2   gate16843  (.A(II30858), .B(II30882), .Z(II30883) ) ;
NAND2   gate16844  (.A(II30874), .B(II30882), .Z(II30884) ) ;
NAND2   gate16845  (.A(WX10053), .B(WX9752), .Z(II30891) ) ;
NAND2   gate16846  (.A(WX10053), .B(II30891), .Z(II30892) ) ;
NAND2   gate16847  (.A(WX9752), .B(II30891), .Z(II30893) ) ;
NAND2   gate16848  (.A(II30892), .B(II30893), .Z(II30890) ) ;
NAND2   gate16849  (.A(WX9816), .B(II30890), .Z(II30898) ) ;
NAND2   gate16850  (.A(WX9816), .B(II30898), .Z(II30899) ) ;
NAND2   gate16851  (.A(II30890), .B(II30898), .Z(II30900) ) ;
NAND2   gate16852  (.A(II30899), .B(II30900), .Z(II30889) ) ;
NAND2   gate16853  (.A(WX9880), .B(WX9944), .Z(II30906) ) ;
NAND2   gate16854  (.A(WX9880), .B(II30906), .Z(II30907) ) ;
NAND2   gate16855  (.A(WX9944), .B(II30906), .Z(II30908) ) ;
NAND2   gate16856  (.A(II30907), .B(II30908), .Z(II30905) ) ;
NAND2   gate16857  (.A(II30889), .B(II30905), .Z(II30913) ) ;
NAND2   gate16858  (.A(II30889), .B(II30913), .Z(II30914) ) ;
NAND2   gate16859  (.A(II30905), .B(II30913), .Z(II30915) ) ;
NAND2   gate16860  (.A(WX10053), .B(WX9754), .Z(II30922) ) ;
NAND2   gate16861  (.A(WX10053), .B(II30922), .Z(II30923) ) ;
NAND2   gate16862  (.A(WX9754), .B(II30922), .Z(II30924) ) ;
NAND2   gate16863  (.A(II30923), .B(II30924), .Z(II30921) ) ;
NAND2   gate16864  (.A(WX9818), .B(II30921), .Z(II30929) ) ;
NAND2   gate16865  (.A(WX9818), .B(II30929), .Z(II30930) ) ;
NAND2   gate16866  (.A(II30921), .B(II30929), .Z(II30931) ) ;
NAND2   gate16867  (.A(II30930), .B(II30931), .Z(II30920) ) ;
NAND2   gate16868  (.A(WX9882), .B(WX9946), .Z(II30937) ) ;
NAND2   gate16869  (.A(WX9882), .B(II30937), .Z(II30938) ) ;
NAND2   gate16870  (.A(WX9946), .B(II30937), .Z(II30939) ) ;
NAND2   gate16871  (.A(II30938), .B(II30939), .Z(II30936) ) ;
NAND2   gate16872  (.A(II30920), .B(II30936), .Z(II30944) ) ;
NAND2   gate16873  (.A(II30920), .B(II30944), .Z(II30945) ) ;
NAND2   gate16874  (.A(II30936), .B(II30944), .Z(II30946) ) ;
NAND2   gate16875  (.A(WX10053), .B(WX9756), .Z(II30953) ) ;
NAND2   gate16876  (.A(WX10053), .B(II30953), .Z(II30954) ) ;
NAND2   gate16877  (.A(WX9756), .B(II30953), .Z(II30955) ) ;
NAND2   gate16878  (.A(II30954), .B(II30955), .Z(II30952) ) ;
NAND2   gate16879  (.A(WX9820), .B(II30952), .Z(II30960) ) ;
NAND2   gate16880  (.A(WX9820), .B(II30960), .Z(II30961) ) ;
NAND2   gate16881  (.A(II30952), .B(II30960), .Z(II30962) ) ;
NAND2   gate16882  (.A(II30961), .B(II30962), .Z(II30951) ) ;
NAND2   gate16883  (.A(WX9884), .B(WX9948), .Z(II30968) ) ;
NAND2   gate16884  (.A(WX9884), .B(II30968), .Z(II30969) ) ;
NAND2   gate16885  (.A(WX9948), .B(II30968), .Z(II30970) ) ;
NAND2   gate16886  (.A(II30969), .B(II30970), .Z(II30967) ) ;
NAND2   gate16887  (.A(II30951), .B(II30967), .Z(II30975) ) ;
NAND2   gate16888  (.A(II30951), .B(II30975), .Z(II30976) ) ;
NAND2   gate16889  (.A(II30967), .B(II30975), .Z(II30977) ) ;
NAND2   gate16890  (.A(WX10053), .B(WX9758), .Z(II30984) ) ;
NAND2   gate16891  (.A(WX10053), .B(II30984), .Z(II30985) ) ;
NAND2   gate16892  (.A(WX9758), .B(II30984), .Z(II30986) ) ;
NAND2   gate16893  (.A(II30985), .B(II30986), .Z(II30983) ) ;
NAND2   gate16894  (.A(WX9822), .B(II30983), .Z(II30991) ) ;
NAND2   gate16895  (.A(WX9822), .B(II30991), .Z(II30992) ) ;
NAND2   gate16896  (.A(II30983), .B(II30991), .Z(II30993) ) ;
NAND2   gate16897  (.A(II30992), .B(II30993), .Z(II30982) ) ;
NAND2   gate16898  (.A(WX9886), .B(WX9950), .Z(II30999) ) ;
NAND2   gate16899  (.A(WX9886), .B(II30999), .Z(II31000) ) ;
NAND2   gate16900  (.A(WX9950), .B(II30999), .Z(II31001) ) ;
NAND2   gate16901  (.A(II31000), .B(II31001), .Z(II30998) ) ;
NAND2   gate16902  (.A(II30982), .B(II30998), .Z(II31006) ) ;
NAND2   gate16903  (.A(II30982), .B(II31006), .Z(II31007) ) ;
NAND2   gate16904  (.A(II30998), .B(II31006), .Z(II31008) ) ;
NAND2   gate16905  (.A(WX9631), .B(WX9536), .Z(II31087) ) ;
NAND2   gate16906  (.A(WX9631), .B(II31087), .Z(II31088) ) ;
NAND2   gate16907  (.A(WX9536), .B(II31087), .Z(II31089) ) ;
NAND2   gate16908  (.A(WX9632), .B(WX9538), .Z(II31100) ) ;
NAND2   gate16909  (.A(WX9632), .B(II31100), .Z(II31101) ) ;
NAND2   gate16910  (.A(WX9538), .B(II31100), .Z(II31102) ) ;
NAND2   gate16911  (.A(WX9633), .B(WX9540), .Z(II31113) ) ;
NAND2   gate16912  (.A(WX9633), .B(II31113), .Z(II31114) ) ;
NAND2   gate16913  (.A(WX9540), .B(II31113), .Z(II31115) ) ;
NAND2   gate16914  (.A(WX9634), .B(WX9542), .Z(II31126) ) ;
NAND2   gate16915  (.A(WX9634), .B(II31126), .Z(II31127) ) ;
NAND2   gate16916  (.A(WX9542), .B(II31126), .Z(II31128) ) ;
NAND2   gate16917  (.A(WX9635), .B(WX9544), .Z(II31139) ) ;
NAND2   gate16918  (.A(WX9635), .B(II31139), .Z(II31140) ) ;
NAND2   gate16919  (.A(WX9544), .B(II31139), .Z(II31141) ) ;
NAND2   gate16920  (.A(WX9636), .B(WX9546), .Z(II31152) ) ;
NAND2   gate16921  (.A(WX9636), .B(II31152), .Z(II31153) ) ;
NAND2   gate16922  (.A(WX9546), .B(II31152), .Z(II31154) ) ;
NAND2   gate16923  (.A(WX9637), .B(WX9548), .Z(II31165) ) ;
NAND2   gate16924  (.A(WX9637), .B(II31165), .Z(II31166) ) ;
NAND2   gate16925  (.A(WX9548), .B(II31165), .Z(II31167) ) ;
NAND2   gate16926  (.A(WX9638), .B(WX9550), .Z(II31178) ) ;
NAND2   gate16927  (.A(WX9638), .B(II31178), .Z(II31179) ) ;
NAND2   gate16928  (.A(WX9550), .B(II31178), .Z(II31180) ) ;
NAND2   gate16929  (.A(WX9639), .B(WX9552), .Z(II31191) ) ;
NAND2   gate16930  (.A(WX9639), .B(II31191), .Z(II31192) ) ;
NAND2   gate16931  (.A(WX9552), .B(II31191), .Z(II31193) ) ;
NAND2   gate16932  (.A(WX9640), .B(WX9554), .Z(II31204) ) ;
NAND2   gate16933  (.A(WX9640), .B(II31204), .Z(II31205) ) ;
NAND2   gate16934  (.A(WX9554), .B(II31204), .Z(II31206) ) ;
NAND2   gate16935  (.A(WX9641), .B(WX9556), .Z(II31217) ) ;
NAND2   gate16936  (.A(WX9641), .B(II31217), .Z(II31218) ) ;
NAND2   gate16937  (.A(WX9556), .B(II31217), .Z(II31219) ) ;
NAND2   gate16938  (.A(WX9642), .B(WX9558), .Z(II31230) ) ;
NAND2   gate16939  (.A(WX9642), .B(II31230), .Z(II31231) ) ;
NAND2   gate16940  (.A(WX9558), .B(II31230), .Z(II31232) ) ;
NAND2   gate16941  (.A(WX9643), .B(WX9560), .Z(II31243) ) ;
NAND2   gate16942  (.A(WX9643), .B(II31243), .Z(II31244) ) ;
NAND2   gate16943  (.A(WX9560), .B(II31243), .Z(II31245) ) ;
NAND2   gate16944  (.A(WX9644), .B(WX9562), .Z(II31256) ) ;
NAND2   gate16945  (.A(WX9644), .B(II31256), .Z(II31257) ) ;
NAND2   gate16946  (.A(WX9562), .B(II31256), .Z(II31258) ) ;
NAND2   gate16947  (.A(WX9645), .B(WX9564), .Z(II31269) ) ;
NAND2   gate16948  (.A(WX9645), .B(II31269), .Z(II31270) ) ;
NAND2   gate16949  (.A(WX9564), .B(II31269), .Z(II31271) ) ;
NAND2   gate16950  (.A(WX9646), .B(WX9566), .Z(II31282) ) ;
NAND2   gate16951  (.A(WX9646), .B(II31282), .Z(II31283) ) ;
NAND2   gate16952  (.A(WX9566), .B(II31282), .Z(II31284) ) ;
NAND2   gate16953  (.A(WX9647), .B(WX9568), .Z(II31295) ) ;
NAND2   gate16954  (.A(WX9647), .B(II31295), .Z(II31296) ) ;
NAND2   gate16955  (.A(WX9568), .B(II31295), .Z(II31297) ) ;
NAND2   gate16956  (.A(WX9648), .B(WX9570), .Z(II31308) ) ;
NAND2   gate16957  (.A(WX9648), .B(II31308), .Z(II31309) ) ;
NAND2   gate16958  (.A(WX9570), .B(II31308), .Z(II31310) ) ;
NAND2   gate16959  (.A(WX9649), .B(WX9572), .Z(II31321) ) ;
NAND2   gate16960  (.A(WX9649), .B(II31321), .Z(II31322) ) ;
NAND2   gate16961  (.A(WX9572), .B(II31321), .Z(II31323) ) ;
NAND2   gate16962  (.A(WX9650), .B(WX9574), .Z(II31334) ) ;
NAND2   gate16963  (.A(WX9650), .B(II31334), .Z(II31335) ) ;
NAND2   gate16964  (.A(WX9574), .B(II31334), .Z(II31336) ) ;
NAND2   gate16965  (.A(WX9651), .B(WX9576), .Z(II31347) ) ;
NAND2   gate16966  (.A(WX9651), .B(II31347), .Z(II31348) ) ;
NAND2   gate16967  (.A(WX9576), .B(II31347), .Z(II31349) ) ;
NAND2   gate16968  (.A(WX9652), .B(WX9578), .Z(II31360) ) ;
NAND2   gate16969  (.A(WX9652), .B(II31360), .Z(II31361) ) ;
NAND2   gate16970  (.A(WX9578), .B(II31360), .Z(II31362) ) ;
NAND2   gate16971  (.A(WX9653), .B(WX9580), .Z(II31373) ) ;
NAND2   gate16972  (.A(WX9653), .B(II31373), .Z(II31374) ) ;
NAND2   gate16973  (.A(WX9580), .B(II31373), .Z(II31375) ) ;
NAND2   gate16974  (.A(WX9654), .B(WX9582), .Z(II31386) ) ;
NAND2   gate16975  (.A(WX9654), .B(II31386), .Z(II31387) ) ;
NAND2   gate16976  (.A(WX9582), .B(II31386), .Z(II31388) ) ;
NAND2   gate16977  (.A(WX9655), .B(WX9584), .Z(II31399) ) ;
NAND2   gate16978  (.A(WX9655), .B(II31399), .Z(II31400) ) ;
NAND2   gate16979  (.A(WX9584), .B(II31399), .Z(II31401) ) ;
NAND2   gate16980  (.A(WX9656), .B(WX9586), .Z(II31412) ) ;
NAND2   gate16981  (.A(WX9656), .B(II31412), .Z(II31413) ) ;
NAND2   gate16982  (.A(WX9586), .B(II31412), .Z(II31414) ) ;
NAND2   gate16983  (.A(WX9657), .B(WX9588), .Z(II31425) ) ;
NAND2   gate16984  (.A(WX9657), .B(II31425), .Z(II31426) ) ;
NAND2   gate16985  (.A(WX9588), .B(II31425), .Z(II31427) ) ;
NAND2   gate16986  (.A(WX9658), .B(WX9590), .Z(II31438) ) ;
NAND2   gate16987  (.A(WX9658), .B(II31438), .Z(II31439) ) ;
NAND2   gate16988  (.A(WX9590), .B(II31438), .Z(II31440) ) ;
NAND2   gate16989  (.A(WX9659), .B(WX9592), .Z(II31451) ) ;
NAND2   gate16990  (.A(WX9659), .B(II31451), .Z(II31452) ) ;
NAND2   gate16991  (.A(WX9592), .B(II31451), .Z(II31453) ) ;
NAND2   gate16992  (.A(WX9660), .B(WX9594), .Z(II31464) ) ;
NAND2   gate16993  (.A(WX9660), .B(II31464), .Z(II31465) ) ;
NAND2   gate16994  (.A(WX9594), .B(II31464), .Z(II31466) ) ;
NAND2   gate16995  (.A(WX9661), .B(WX9596), .Z(II31477) ) ;
NAND2   gate16996  (.A(WX9661), .B(II31477), .Z(II31478) ) ;
NAND2   gate16997  (.A(WX9596), .B(II31477), .Z(II31479) ) ;
NAND2   gate16998  (.A(WX9662), .B(WX9598), .Z(II31490) ) ;
NAND2   gate16999  (.A(WX9662), .B(II31490), .Z(II31491) ) ;
NAND2   gate17000  (.A(WX9598), .B(II31490), .Z(II31492) ) ;
NAND2   gate17001  (.A(WX9678), .B(CRC_OUT_2_31), .Z(II31505) ) ;
NAND2   gate17002  (.A(WX9678), .B(II31505), .Z(II31506) ) ;
NAND2   gate17003  (.A(CRC_OUT_2_31), .B(II31505), .Z(II31507) ) ;
NAND2   gate17004  (.A(II31506), .B(II31507), .Z(II31504) ) ;
NAND2   gate17005  (.A(CRC_OUT_2_15), .B(II31504), .Z(II31512) ) ;
NAND2   gate17006  (.A(CRC_OUT_2_15), .B(II31512), .Z(II31513) ) ;
NAND2   gate17007  (.A(II31504), .B(II31512), .Z(II31514) ) ;
NAND2   gate17008  (.A(WX9683), .B(CRC_OUT_2_31), .Z(II31520) ) ;
NAND2   gate17009  (.A(WX9683), .B(II31520), .Z(II31521) ) ;
NAND2   gate17010  (.A(CRC_OUT_2_31), .B(II31520), .Z(II31522) ) ;
NAND2   gate17011  (.A(II31521), .B(II31522), .Z(II31519) ) ;
NAND2   gate17012  (.A(CRC_OUT_2_10), .B(II31519), .Z(II31527) ) ;
NAND2   gate17013  (.A(CRC_OUT_2_10), .B(II31527), .Z(II31528) ) ;
NAND2   gate17014  (.A(II31519), .B(II31527), .Z(II31529) ) ;
NAND2   gate17015  (.A(WX9690), .B(CRC_OUT_2_31), .Z(II31535) ) ;
NAND2   gate17016  (.A(WX9690), .B(II31535), .Z(II31536) ) ;
NAND2   gate17017  (.A(CRC_OUT_2_31), .B(II31535), .Z(II31537) ) ;
NAND2   gate17018  (.A(II31536), .B(II31537), .Z(II31534) ) ;
NAND2   gate17019  (.A(CRC_OUT_2_3), .B(II31534), .Z(II31542) ) ;
NAND2   gate17020  (.A(CRC_OUT_2_3), .B(II31542), .Z(II31543) ) ;
NAND2   gate17021  (.A(II31534), .B(II31542), .Z(II31544) ) ;
NAND2   gate17022  (.A(WX9694), .B(CRC_OUT_2_31), .Z(II31549) ) ;
NAND2   gate17023  (.A(WX9694), .B(II31549), .Z(II31550) ) ;
NAND2   gate17024  (.A(CRC_OUT_2_31), .B(II31549), .Z(II31551) ) ;
NAND2   gate17025  (.A(WX9663), .B(CRC_OUT_2_30), .Z(II31556) ) ;
NAND2   gate17026  (.A(WX9663), .B(II31556), .Z(II31557) ) ;
NAND2   gate17027  (.A(CRC_OUT_2_30), .B(II31556), .Z(II31558) ) ;
NAND2   gate17028  (.A(WX9664), .B(CRC_OUT_2_29), .Z(II31563) ) ;
NAND2   gate17029  (.A(WX9664), .B(II31563), .Z(II31564) ) ;
NAND2   gate17030  (.A(CRC_OUT_2_29), .B(II31563), .Z(II31565) ) ;
NAND2   gate17031  (.A(WX9665), .B(CRC_OUT_2_28), .Z(II31570) ) ;
NAND2   gate17032  (.A(WX9665), .B(II31570), .Z(II31571) ) ;
NAND2   gate17033  (.A(CRC_OUT_2_28), .B(II31570), .Z(II31572) ) ;
NAND2   gate17034  (.A(WX9666), .B(CRC_OUT_2_27), .Z(II31577) ) ;
NAND2   gate17035  (.A(WX9666), .B(II31577), .Z(II31578) ) ;
NAND2   gate17036  (.A(CRC_OUT_2_27), .B(II31577), .Z(II31579) ) ;
NAND2   gate17037  (.A(WX9667), .B(CRC_OUT_2_26), .Z(II31584) ) ;
NAND2   gate17038  (.A(WX9667), .B(II31584), .Z(II31585) ) ;
NAND2   gate17039  (.A(CRC_OUT_2_26), .B(II31584), .Z(II31586) ) ;
NAND2   gate17040  (.A(WX9668), .B(CRC_OUT_2_25), .Z(II31591) ) ;
NAND2   gate17041  (.A(WX9668), .B(II31591), .Z(II31592) ) ;
NAND2   gate17042  (.A(CRC_OUT_2_25), .B(II31591), .Z(II31593) ) ;
NAND2   gate17043  (.A(WX9669), .B(CRC_OUT_2_24), .Z(II31598) ) ;
NAND2   gate17044  (.A(WX9669), .B(II31598), .Z(II31599) ) ;
NAND2   gate17045  (.A(CRC_OUT_2_24), .B(II31598), .Z(II31600) ) ;
NAND2   gate17046  (.A(WX9670), .B(CRC_OUT_2_23), .Z(II31605) ) ;
NAND2   gate17047  (.A(WX9670), .B(II31605), .Z(II31606) ) ;
NAND2   gate17048  (.A(CRC_OUT_2_23), .B(II31605), .Z(II31607) ) ;
NAND2   gate17049  (.A(WX9671), .B(CRC_OUT_2_22), .Z(II31612) ) ;
NAND2   gate17050  (.A(WX9671), .B(II31612), .Z(II31613) ) ;
NAND2   gate17051  (.A(CRC_OUT_2_22), .B(II31612), .Z(II31614) ) ;
NAND2   gate17052  (.A(WX9672), .B(CRC_OUT_2_21), .Z(II31619) ) ;
NAND2   gate17053  (.A(WX9672), .B(II31619), .Z(II31620) ) ;
NAND2   gate17054  (.A(CRC_OUT_2_21), .B(II31619), .Z(II31621) ) ;
NAND2   gate17055  (.A(WX9673), .B(CRC_OUT_2_20), .Z(II31626) ) ;
NAND2   gate17056  (.A(WX9673), .B(II31626), .Z(II31627) ) ;
NAND2   gate17057  (.A(CRC_OUT_2_20), .B(II31626), .Z(II31628) ) ;
NAND2   gate17058  (.A(WX9674), .B(CRC_OUT_2_19), .Z(II31633) ) ;
NAND2   gate17059  (.A(WX9674), .B(II31633), .Z(II31634) ) ;
NAND2   gate17060  (.A(CRC_OUT_2_19), .B(II31633), .Z(II31635) ) ;
NAND2   gate17061  (.A(WX9675), .B(CRC_OUT_2_18), .Z(II31640) ) ;
NAND2   gate17062  (.A(WX9675), .B(II31640), .Z(II31641) ) ;
NAND2   gate17063  (.A(CRC_OUT_2_18), .B(II31640), .Z(II31642) ) ;
NAND2   gate17064  (.A(WX9676), .B(CRC_OUT_2_17), .Z(II31647) ) ;
NAND2   gate17065  (.A(WX9676), .B(II31647), .Z(II31648) ) ;
NAND2   gate17066  (.A(CRC_OUT_2_17), .B(II31647), .Z(II31649) ) ;
NAND2   gate17067  (.A(WX9677), .B(CRC_OUT_2_16), .Z(II31654) ) ;
NAND2   gate17068  (.A(WX9677), .B(II31654), .Z(II31655) ) ;
NAND2   gate17069  (.A(CRC_OUT_2_16), .B(II31654), .Z(II31656) ) ;
NAND2   gate17070  (.A(WX9679), .B(CRC_OUT_2_14), .Z(II31661) ) ;
NAND2   gate17071  (.A(WX9679), .B(II31661), .Z(II31662) ) ;
NAND2   gate17072  (.A(CRC_OUT_2_14), .B(II31661), .Z(II31663) ) ;
NAND2   gate17073  (.A(WX9680), .B(CRC_OUT_2_13), .Z(II31668) ) ;
NAND2   gate17074  (.A(WX9680), .B(II31668), .Z(II31669) ) ;
NAND2   gate17075  (.A(CRC_OUT_2_13), .B(II31668), .Z(II31670) ) ;
NAND2   gate17076  (.A(WX9681), .B(CRC_OUT_2_12), .Z(II31675) ) ;
NAND2   gate17077  (.A(WX9681), .B(II31675), .Z(II31676) ) ;
NAND2   gate17078  (.A(CRC_OUT_2_12), .B(II31675), .Z(II31677) ) ;
NAND2   gate17079  (.A(WX9682), .B(CRC_OUT_2_11), .Z(II31682) ) ;
NAND2   gate17080  (.A(WX9682), .B(II31682), .Z(II31683) ) ;
NAND2   gate17081  (.A(CRC_OUT_2_11), .B(II31682), .Z(II31684) ) ;
NAND2   gate17082  (.A(WX9684), .B(CRC_OUT_2_9), .Z(II31689) ) ;
NAND2   gate17083  (.A(WX9684), .B(II31689), .Z(II31690) ) ;
NAND2   gate17084  (.A(CRC_OUT_2_9), .B(II31689), .Z(II31691) ) ;
NAND2   gate17085  (.A(WX9685), .B(CRC_OUT_2_8), .Z(II31696) ) ;
NAND2   gate17086  (.A(WX9685), .B(II31696), .Z(II31697) ) ;
NAND2   gate17087  (.A(CRC_OUT_2_8), .B(II31696), .Z(II31698) ) ;
NAND2   gate17088  (.A(WX9686), .B(CRC_OUT_2_7), .Z(II31703) ) ;
NAND2   gate17089  (.A(WX9686), .B(II31703), .Z(II31704) ) ;
NAND2   gate17090  (.A(CRC_OUT_2_7), .B(II31703), .Z(II31705) ) ;
NAND2   gate17091  (.A(WX9687), .B(CRC_OUT_2_6), .Z(II31710) ) ;
NAND2   gate17092  (.A(WX9687), .B(II31710), .Z(II31711) ) ;
NAND2   gate17093  (.A(CRC_OUT_2_6), .B(II31710), .Z(II31712) ) ;
NAND2   gate17094  (.A(WX9688), .B(CRC_OUT_2_5), .Z(II31717) ) ;
NAND2   gate17095  (.A(WX9688), .B(II31717), .Z(II31718) ) ;
NAND2   gate17096  (.A(CRC_OUT_2_5), .B(II31717), .Z(II31719) ) ;
NAND2   gate17097  (.A(WX9689), .B(CRC_OUT_2_4), .Z(II31724) ) ;
NAND2   gate17098  (.A(WX9689), .B(II31724), .Z(II31725) ) ;
NAND2   gate17099  (.A(CRC_OUT_2_4), .B(II31724), .Z(II31726) ) ;
NAND2   gate17100  (.A(WX9691), .B(CRC_OUT_2_2), .Z(II31731) ) ;
NAND2   gate17101  (.A(WX9691), .B(II31731), .Z(II31732) ) ;
NAND2   gate17102  (.A(CRC_OUT_2_2), .B(II31731), .Z(II31733) ) ;
NAND2   gate17103  (.A(WX9692), .B(CRC_OUT_2_1), .Z(II31738) ) ;
NAND2   gate17104  (.A(WX9692), .B(II31738), .Z(II31739) ) ;
NAND2   gate17105  (.A(CRC_OUT_2_1), .B(II31738), .Z(II31740) ) ;
NAND2   gate17106  (.A(WX9693), .B(CRC_OUT_2_0), .Z(II31745) ) ;
NAND2   gate17107  (.A(WX9693), .B(II31745), .Z(II31746) ) ;
NAND2   gate17108  (.A(CRC_OUT_2_0), .B(II31745), .Z(II31747) ) ;
NAND2   gate17109  (.A(WX11345), .B(WX10989), .Z(II34028) ) ;
NAND2   gate17110  (.A(WX11345), .B(II34028), .Z(II34029) ) ;
NAND2   gate17111  (.A(WX10989), .B(II34028), .Z(II34030) ) ;
NAND2   gate17112  (.A(II34029), .B(II34030), .Z(II34027) ) ;
NAND2   gate17113  (.A(WX11053), .B(II34027), .Z(II34035) ) ;
NAND2   gate17114  (.A(WX11053), .B(II34035), .Z(II34036) ) ;
NAND2   gate17115  (.A(II34027), .B(II34035), .Z(II34037) ) ;
NAND2   gate17116  (.A(II34036), .B(II34037), .Z(II34026) ) ;
NAND2   gate17117  (.A(WX11117), .B(WX11181), .Z(II34043) ) ;
NAND2   gate17118  (.A(WX11117), .B(II34043), .Z(II34044) ) ;
NAND2   gate17119  (.A(WX11181), .B(II34043), .Z(II34045) ) ;
NAND2   gate17120  (.A(II34044), .B(II34045), .Z(II34042) ) ;
NAND2   gate17121  (.A(II34026), .B(II34042), .Z(II34050) ) ;
NAND2   gate17122  (.A(II34026), .B(II34050), .Z(II34051) ) ;
NAND2   gate17123  (.A(II34042), .B(II34050), .Z(II34052) ) ;
NAND2   gate17124  (.A(WX11345), .B(WX10991), .Z(II34059) ) ;
NAND2   gate17125  (.A(WX11345), .B(II34059), .Z(II34060) ) ;
NAND2   gate17126  (.A(WX10991), .B(II34059), .Z(II34061) ) ;
NAND2   gate17127  (.A(II34060), .B(II34061), .Z(II34058) ) ;
NAND2   gate17128  (.A(WX11055), .B(II34058), .Z(II34066) ) ;
NAND2   gate17129  (.A(WX11055), .B(II34066), .Z(II34067) ) ;
NAND2   gate17130  (.A(II34058), .B(II34066), .Z(II34068) ) ;
NAND2   gate17131  (.A(II34067), .B(II34068), .Z(II34057) ) ;
NAND2   gate17132  (.A(WX11119), .B(WX11183), .Z(II34074) ) ;
NAND2   gate17133  (.A(WX11119), .B(II34074), .Z(II34075) ) ;
NAND2   gate17134  (.A(WX11183), .B(II34074), .Z(II34076) ) ;
NAND2   gate17135  (.A(II34075), .B(II34076), .Z(II34073) ) ;
NAND2   gate17136  (.A(II34057), .B(II34073), .Z(II34081) ) ;
NAND2   gate17137  (.A(II34057), .B(II34081), .Z(II34082) ) ;
NAND2   gate17138  (.A(II34073), .B(II34081), .Z(II34083) ) ;
NAND2   gate17139  (.A(WX11345), .B(WX10993), .Z(II34090) ) ;
NAND2   gate17140  (.A(WX11345), .B(II34090), .Z(II34091) ) ;
NAND2   gate17141  (.A(WX10993), .B(II34090), .Z(II34092) ) ;
NAND2   gate17142  (.A(II34091), .B(II34092), .Z(II34089) ) ;
NAND2   gate17143  (.A(WX11057), .B(II34089), .Z(II34097) ) ;
NAND2   gate17144  (.A(WX11057), .B(II34097), .Z(II34098) ) ;
NAND2   gate17145  (.A(II34089), .B(II34097), .Z(II34099) ) ;
NAND2   gate17146  (.A(II34098), .B(II34099), .Z(II34088) ) ;
NAND2   gate17147  (.A(WX11121), .B(WX11185), .Z(II34105) ) ;
NAND2   gate17148  (.A(WX11121), .B(II34105), .Z(II34106) ) ;
NAND2   gate17149  (.A(WX11185), .B(II34105), .Z(II34107) ) ;
NAND2   gate17150  (.A(II34106), .B(II34107), .Z(II34104) ) ;
NAND2   gate17151  (.A(II34088), .B(II34104), .Z(II34112) ) ;
NAND2   gate17152  (.A(II34088), .B(II34112), .Z(II34113) ) ;
NAND2   gate17153  (.A(II34104), .B(II34112), .Z(II34114) ) ;
NAND2   gate17154  (.A(WX11345), .B(WX10995), .Z(II34121) ) ;
NAND2   gate17155  (.A(WX11345), .B(II34121), .Z(II34122) ) ;
NAND2   gate17156  (.A(WX10995), .B(II34121), .Z(II34123) ) ;
NAND2   gate17157  (.A(II34122), .B(II34123), .Z(II34120) ) ;
NAND2   gate17158  (.A(WX11059), .B(II34120), .Z(II34128) ) ;
NAND2   gate17159  (.A(WX11059), .B(II34128), .Z(II34129) ) ;
NAND2   gate17160  (.A(II34120), .B(II34128), .Z(II34130) ) ;
NAND2   gate17161  (.A(II34129), .B(II34130), .Z(II34119) ) ;
NAND2   gate17162  (.A(WX11123), .B(WX11187), .Z(II34136) ) ;
NAND2   gate17163  (.A(WX11123), .B(II34136), .Z(II34137) ) ;
NAND2   gate17164  (.A(WX11187), .B(II34136), .Z(II34138) ) ;
NAND2   gate17165  (.A(II34137), .B(II34138), .Z(II34135) ) ;
NAND2   gate17166  (.A(II34119), .B(II34135), .Z(II34143) ) ;
NAND2   gate17167  (.A(II34119), .B(II34143), .Z(II34144) ) ;
NAND2   gate17168  (.A(II34135), .B(II34143), .Z(II34145) ) ;
NAND2   gate17169  (.A(WX11345), .B(WX10997), .Z(II34152) ) ;
NAND2   gate17170  (.A(WX11345), .B(II34152), .Z(II34153) ) ;
NAND2   gate17171  (.A(WX10997), .B(II34152), .Z(II34154) ) ;
NAND2   gate17172  (.A(II34153), .B(II34154), .Z(II34151) ) ;
NAND2   gate17173  (.A(WX11061), .B(II34151), .Z(II34159) ) ;
NAND2   gate17174  (.A(WX11061), .B(II34159), .Z(II34160) ) ;
NAND2   gate17175  (.A(II34151), .B(II34159), .Z(II34161) ) ;
NAND2   gate17176  (.A(II34160), .B(II34161), .Z(II34150) ) ;
NAND2   gate17177  (.A(WX11125), .B(WX11189), .Z(II34167) ) ;
NAND2   gate17178  (.A(WX11125), .B(II34167), .Z(II34168) ) ;
NAND2   gate17179  (.A(WX11189), .B(II34167), .Z(II34169) ) ;
NAND2   gate17180  (.A(II34168), .B(II34169), .Z(II34166) ) ;
NAND2   gate17181  (.A(II34150), .B(II34166), .Z(II34174) ) ;
NAND2   gate17182  (.A(II34150), .B(II34174), .Z(II34175) ) ;
NAND2   gate17183  (.A(II34166), .B(II34174), .Z(II34176) ) ;
NAND2   gate17184  (.A(WX11345), .B(WX10999), .Z(II34183) ) ;
NAND2   gate17185  (.A(WX11345), .B(II34183), .Z(II34184) ) ;
NAND2   gate17186  (.A(WX10999), .B(II34183), .Z(II34185) ) ;
NAND2   gate17187  (.A(II34184), .B(II34185), .Z(II34182) ) ;
NAND2   gate17188  (.A(WX11063), .B(II34182), .Z(II34190) ) ;
NAND2   gate17189  (.A(WX11063), .B(II34190), .Z(II34191) ) ;
NAND2   gate17190  (.A(II34182), .B(II34190), .Z(II34192) ) ;
NAND2   gate17191  (.A(II34191), .B(II34192), .Z(II34181) ) ;
NAND2   gate17192  (.A(WX11127), .B(WX11191), .Z(II34198) ) ;
NAND2   gate17193  (.A(WX11127), .B(II34198), .Z(II34199) ) ;
NAND2   gate17194  (.A(WX11191), .B(II34198), .Z(II34200) ) ;
NAND2   gate17195  (.A(II34199), .B(II34200), .Z(II34197) ) ;
NAND2   gate17196  (.A(II34181), .B(II34197), .Z(II34205) ) ;
NAND2   gate17197  (.A(II34181), .B(II34205), .Z(II34206) ) ;
NAND2   gate17198  (.A(II34197), .B(II34205), .Z(II34207) ) ;
NAND2   gate17199  (.A(WX11345), .B(WX11001), .Z(II34214) ) ;
NAND2   gate17200  (.A(WX11345), .B(II34214), .Z(II34215) ) ;
NAND2   gate17201  (.A(WX11001), .B(II34214), .Z(II34216) ) ;
NAND2   gate17202  (.A(II34215), .B(II34216), .Z(II34213) ) ;
NAND2   gate17203  (.A(WX11065), .B(II34213), .Z(II34221) ) ;
NAND2   gate17204  (.A(WX11065), .B(II34221), .Z(II34222) ) ;
NAND2   gate17205  (.A(II34213), .B(II34221), .Z(II34223) ) ;
NAND2   gate17206  (.A(II34222), .B(II34223), .Z(II34212) ) ;
NAND2   gate17207  (.A(WX11129), .B(WX11193), .Z(II34229) ) ;
NAND2   gate17208  (.A(WX11129), .B(II34229), .Z(II34230) ) ;
NAND2   gate17209  (.A(WX11193), .B(II34229), .Z(II34231) ) ;
NAND2   gate17210  (.A(II34230), .B(II34231), .Z(II34228) ) ;
NAND2   gate17211  (.A(II34212), .B(II34228), .Z(II34236) ) ;
NAND2   gate17212  (.A(II34212), .B(II34236), .Z(II34237) ) ;
NAND2   gate17213  (.A(II34228), .B(II34236), .Z(II34238) ) ;
NAND2   gate17214  (.A(WX11345), .B(WX11003), .Z(II34245) ) ;
NAND2   gate17215  (.A(WX11345), .B(II34245), .Z(II34246) ) ;
NAND2   gate17216  (.A(WX11003), .B(II34245), .Z(II34247) ) ;
NAND2   gate17217  (.A(II34246), .B(II34247), .Z(II34244) ) ;
NAND2   gate17218  (.A(WX11067), .B(II34244), .Z(II34252) ) ;
NAND2   gate17219  (.A(WX11067), .B(II34252), .Z(II34253) ) ;
NAND2   gate17220  (.A(II34244), .B(II34252), .Z(II34254) ) ;
NAND2   gate17221  (.A(II34253), .B(II34254), .Z(II34243) ) ;
NAND2   gate17222  (.A(WX11131), .B(WX11195), .Z(II34260) ) ;
NAND2   gate17223  (.A(WX11131), .B(II34260), .Z(II34261) ) ;
NAND2   gate17224  (.A(WX11195), .B(II34260), .Z(II34262) ) ;
NAND2   gate17225  (.A(II34261), .B(II34262), .Z(II34259) ) ;
NAND2   gate17226  (.A(II34243), .B(II34259), .Z(II34267) ) ;
NAND2   gate17227  (.A(II34243), .B(II34267), .Z(II34268) ) ;
NAND2   gate17228  (.A(II34259), .B(II34267), .Z(II34269) ) ;
NAND2   gate17229  (.A(WX11345), .B(WX11005), .Z(II34276) ) ;
NAND2   gate17230  (.A(WX11345), .B(II34276), .Z(II34277) ) ;
NAND2   gate17231  (.A(WX11005), .B(II34276), .Z(II34278) ) ;
NAND2   gate17232  (.A(II34277), .B(II34278), .Z(II34275) ) ;
NAND2   gate17233  (.A(WX11069), .B(II34275), .Z(II34283) ) ;
NAND2   gate17234  (.A(WX11069), .B(II34283), .Z(II34284) ) ;
NAND2   gate17235  (.A(II34275), .B(II34283), .Z(II34285) ) ;
NAND2   gate17236  (.A(II34284), .B(II34285), .Z(II34274) ) ;
NAND2   gate17237  (.A(WX11133), .B(WX11197), .Z(II34291) ) ;
NAND2   gate17238  (.A(WX11133), .B(II34291), .Z(II34292) ) ;
NAND2   gate17239  (.A(WX11197), .B(II34291), .Z(II34293) ) ;
NAND2   gate17240  (.A(II34292), .B(II34293), .Z(II34290) ) ;
NAND2   gate17241  (.A(II34274), .B(II34290), .Z(II34298) ) ;
NAND2   gate17242  (.A(II34274), .B(II34298), .Z(II34299) ) ;
NAND2   gate17243  (.A(II34290), .B(II34298), .Z(II34300) ) ;
NAND2   gate17244  (.A(WX11345), .B(WX11007), .Z(II34307) ) ;
NAND2   gate17245  (.A(WX11345), .B(II34307), .Z(II34308) ) ;
NAND2   gate17246  (.A(WX11007), .B(II34307), .Z(II34309) ) ;
NAND2   gate17247  (.A(II34308), .B(II34309), .Z(II34306) ) ;
NAND2   gate17248  (.A(WX11071), .B(II34306), .Z(II34314) ) ;
NAND2   gate17249  (.A(WX11071), .B(II34314), .Z(II34315) ) ;
NAND2   gate17250  (.A(II34306), .B(II34314), .Z(II34316) ) ;
NAND2   gate17251  (.A(II34315), .B(II34316), .Z(II34305) ) ;
NAND2   gate17252  (.A(WX11135), .B(WX11199), .Z(II34322) ) ;
NAND2   gate17253  (.A(WX11135), .B(II34322), .Z(II34323) ) ;
NAND2   gate17254  (.A(WX11199), .B(II34322), .Z(II34324) ) ;
NAND2   gate17255  (.A(II34323), .B(II34324), .Z(II34321) ) ;
NAND2   gate17256  (.A(II34305), .B(II34321), .Z(II34329) ) ;
NAND2   gate17257  (.A(II34305), .B(II34329), .Z(II34330) ) ;
NAND2   gate17258  (.A(II34321), .B(II34329), .Z(II34331) ) ;
NAND2   gate17259  (.A(WX11345), .B(WX11009), .Z(II34338) ) ;
NAND2   gate17260  (.A(WX11345), .B(II34338), .Z(II34339) ) ;
NAND2   gate17261  (.A(WX11009), .B(II34338), .Z(II34340) ) ;
NAND2   gate17262  (.A(II34339), .B(II34340), .Z(II34337) ) ;
NAND2   gate17263  (.A(WX11073), .B(II34337), .Z(II34345) ) ;
NAND2   gate17264  (.A(WX11073), .B(II34345), .Z(II34346) ) ;
NAND2   gate17265  (.A(II34337), .B(II34345), .Z(II34347) ) ;
NAND2   gate17266  (.A(II34346), .B(II34347), .Z(II34336) ) ;
NAND2   gate17267  (.A(WX11137), .B(WX11201), .Z(II34353) ) ;
NAND2   gate17268  (.A(WX11137), .B(II34353), .Z(II34354) ) ;
NAND2   gate17269  (.A(WX11201), .B(II34353), .Z(II34355) ) ;
NAND2   gate17270  (.A(II34354), .B(II34355), .Z(II34352) ) ;
NAND2   gate17271  (.A(II34336), .B(II34352), .Z(II34360) ) ;
NAND2   gate17272  (.A(II34336), .B(II34360), .Z(II34361) ) ;
NAND2   gate17273  (.A(II34352), .B(II34360), .Z(II34362) ) ;
NAND2   gate17274  (.A(WX11345), .B(WX11011), .Z(II34369) ) ;
NAND2   gate17275  (.A(WX11345), .B(II34369), .Z(II34370) ) ;
NAND2   gate17276  (.A(WX11011), .B(II34369), .Z(II34371) ) ;
NAND2   gate17277  (.A(II34370), .B(II34371), .Z(II34368) ) ;
NAND2   gate17278  (.A(WX11075), .B(II34368), .Z(II34376) ) ;
NAND2   gate17279  (.A(WX11075), .B(II34376), .Z(II34377) ) ;
NAND2   gate17280  (.A(II34368), .B(II34376), .Z(II34378) ) ;
NAND2   gate17281  (.A(II34377), .B(II34378), .Z(II34367) ) ;
NAND2   gate17282  (.A(WX11139), .B(WX11203), .Z(II34384) ) ;
NAND2   gate17283  (.A(WX11139), .B(II34384), .Z(II34385) ) ;
NAND2   gate17284  (.A(WX11203), .B(II34384), .Z(II34386) ) ;
NAND2   gate17285  (.A(II34385), .B(II34386), .Z(II34383) ) ;
NAND2   gate17286  (.A(II34367), .B(II34383), .Z(II34391) ) ;
NAND2   gate17287  (.A(II34367), .B(II34391), .Z(II34392) ) ;
NAND2   gate17288  (.A(II34383), .B(II34391), .Z(II34393) ) ;
NAND2   gate17289  (.A(WX11345), .B(WX11013), .Z(II34400) ) ;
NAND2   gate17290  (.A(WX11345), .B(II34400), .Z(II34401) ) ;
NAND2   gate17291  (.A(WX11013), .B(II34400), .Z(II34402) ) ;
NAND2   gate17292  (.A(II34401), .B(II34402), .Z(II34399) ) ;
NAND2   gate17293  (.A(WX11077), .B(II34399), .Z(II34407) ) ;
NAND2   gate17294  (.A(WX11077), .B(II34407), .Z(II34408) ) ;
NAND2   gate17295  (.A(II34399), .B(II34407), .Z(II34409) ) ;
NAND2   gate17296  (.A(II34408), .B(II34409), .Z(II34398) ) ;
NAND2   gate17297  (.A(WX11141), .B(WX11205), .Z(II34415) ) ;
NAND2   gate17298  (.A(WX11141), .B(II34415), .Z(II34416) ) ;
NAND2   gate17299  (.A(WX11205), .B(II34415), .Z(II34417) ) ;
NAND2   gate17300  (.A(II34416), .B(II34417), .Z(II34414) ) ;
NAND2   gate17301  (.A(II34398), .B(II34414), .Z(II34422) ) ;
NAND2   gate17302  (.A(II34398), .B(II34422), .Z(II34423) ) ;
NAND2   gate17303  (.A(II34414), .B(II34422), .Z(II34424) ) ;
NAND2   gate17304  (.A(WX11345), .B(WX11015), .Z(II34431) ) ;
NAND2   gate17305  (.A(WX11345), .B(II34431), .Z(II34432) ) ;
NAND2   gate17306  (.A(WX11015), .B(II34431), .Z(II34433) ) ;
NAND2   gate17307  (.A(II34432), .B(II34433), .Z(II34430) ) ;
NAND2   gate17308  (.A(WX11079), .B(II34430), .Z(II34438) ) ;
NAND2   gate17309  (.A(WX11079), .B(II34438), .Z(II34439) ) ;
NAND2   gate17310  (.A(II34430), .B(II34438), .Z(II34440) ) ;
NAND2   gate17311  (.A(II34439), .B(II34440), .Z(II34429) ) ;
NAND2   gate17312  (.A(WX11143), .B(WX11207), .Z(II34446) ) ;
NAND2   gate17313  (.A(WX11143), .B(II34446), .Z(II34447) ) ;
NAND2   gate17314  (.A(WX11207), .B(II34446), .Z(II34448) ) ;
NAND2   gate17315  (.A(II34447), .B(II34448), .Z(II34445) ) ;
NAND2   gate17316  (.A(II34429), .B(II34445), .Z(II34453) ) ;
NAND2   gate17317  (.A(II34429), .B(II34453), .Z(II34454) ) ;
NAND2   gate17318  (.A(II34445), .B(II34453), .Z(II34455) ) ;
NAND2   gate17319  (.A(WX11345), .B(WX11017), .Z(II34462) ) ;
NAND2   gate17320  (.A(WX11345), .B(II34462), .Z(II34463) ) ;
NAND2   gate17321  (.A(WX11017), .B(II34462), .Z(II34464) ) ;
NAND2   gate17322  (.A(II34463), .B(II34464), .Z(II34461) ) ;
NAND2   gate17323  (.A(WX11081), .B(II34461), .Z(II34469) ) ;
NAND2   gate17324  (.A(WX11081), .B(II34469), .Z(II34470) ) ;
NAND2   gate17325  (.A(II34461), .B(II34469), .Z(II34471) ) ;
NAND2   gate17326  (.A(II34470), .B(II34471), .Z(II34460) ) ;
NAND2   gate17327  (.A(WX11145), .B(WX11209), .Z(II34477) ) ;
NAND2   gate17328  (.A(WX11145), .B(II34477), .Z(II34478) ) ;
NAND2   gate17329  (.A(WX11209), .B(II34477), .Z(II34479) ) ;
NAND2   gate17330  (.A(II34478), .B(II34479), .Z(II34476) ) ;
NAND2   gate17331  (.A(II34460), .B(II34476), .Z(II34484) ) ;
NAND2   gate17332  (.A(II34460), .B(II34484), .Z(II34485) ) ;
NAND2   gate17333  (.A(II34476), .B(II34484), .Z(II34486) ) ;
NAND2   gate17334  (.A(WX11345), .B(WX11019), .Z(II34493) ) ;
NAND2   gate17335  (.A(WX11345), .B(II34493), .Z(II34494) ) ;
NAND2   gate17336  (.A(WX11019), .B(II34493), .Z(II34495) ) ;
NAND2   gate17337  (.A(II34494), .B(II34495), .Z(II34492) ) ;
NAND2   gate17338  (.A(WX11083), .B(II34492), .Z(II34500) ) ;
NAND2   gate17339  (.A(WX11083), .B(II34500), .Z(II34501) ) ;
NAND2   gate17340  (.A(II34492), .B(II34500), .Z(II34502) ) ;
NAND2   gate17341  (.A(II34501), .B(II34502), .Z(II34491) ) ;
NAND2   gate17342  (.A(WX11147), .B(WX11211), .Z(II34508) ) ;
NAND2   gate17343  (.A(WX11147), .B(II34508), .Z(II34509) ) ;
NAND2   gate17344  (.A(WX11211), .B(II34508), .Z(II34510) ) ;
NAND2   gate17345  (.A(II34509), .B(II34510), .Z(II34507) ) ;
NAND2   gate17346  (.A(II34491), .B(II34507), .Z(II34515) ) ;
NAND2   gate17347  (.A(II34491), .B(II34515), .Z(II34516) ) ;
NAND2   gate17348  (.A(II34507), .B(II34515), .Z(II34517) ) ;
NAND2   gate17349  (.A(WX11346), .B(WX11021), .Z(II34524) ) ;
NAND2   gate17350  (.A(WX11346), .B(II34524), .Z(II34525) ) ;
NAND2   gate17351  (.A(WX11021), .B(II34524), .Z(II34526) ) ;
NAND2   gate17352  (.A(II34525), .B(II34526), .Z(II34523) ) ;
NAND2   gate17353  (.A(WX11085), .B(II34523), .Z(II34531) ) ;
NAND2   gate17354  (.A(WX11085), .B(II34531), .Z(II34532) ) ;
NAND2   gate17355  (.A(II34523), .B(II34531), .Z(II34533) ) ;
NAND2   gate17356  (.A(II34532), .B(II34533), .Z(II34522) ) ;
NAND2   gate17357  (.A(WX11149), .B(WX11213), .Z(II34539) ) ;
NAND2   gate17358  (.A(WX11149), .B(II34539), .Z(II34540) ) ;
NAND2   gate17359  (.A(WX11213), .B(II34539), .Z(II34541) ) ;
NAND2   gate17360  (.A(II34540), .B(II34541), .Z(II34538) ) ;
NAND2   gate17361  (.A(II34522), .B(II34538), .Z(II34546) ) ;
NAND2   gate17362  (.A(II34522), .B(II34546), .Z(II34547) ) ;
NAND2   gate17363  (.A(II34538), .B(II34546), .Z(II34548) ) ;
NAND2   gate17364  (.A(WX11346), .B(WX11023), .Z(II34555) ) ;
NAND2   gate17365  (.A(WX11346), .B(II34555), .Z(II34556) ) ;
NAND2   gate17366  (.A(WX11023), .B(II34555), .Z(II34557) ) ;
NAND2   gate17367  (.A(II34556), .B(II34557), .Z(II34554) ) ;
NAND2   gate17368  (.A(WX11087), .B(II34554), .Z(II34562) ) ;
NAND2   gate17369  (.A(WX11087), .B(II34562), .Z(II34563) ) ;
NAND2   gate17370  (.A(II34554), .B(II34562), .Z(II34564) ) ;
NAND2   gate17371  (.A(II34563), .B(II34564), .Z(II34553) ) ;
NAND2   gate17372  (.A(WX11151), .B(WX11215), .Z(II34570) ) ;
NAND2   gate17373  (.A(WX11151), .B(II34570), .Z(II34571) ) ;
NAND2   gate17374  (.A(WX11215), .B(II34570), .Z(II34572) ) ;
NAND2   gate17375  (.A(II34571), .B(II34572), .Z(II34569) ) ;
NAND2   gate17376  (.A(II34553), .B(II34569), .Z(II34577) ) ;
NAND2   gate17377  (.A(II34553), .B(II34577), .Z(II34578) ) ;
NAND2   gate17378  (.A(II34569), .B(II34577), .Z(II34579) ) ;
NAND2   gate17379  (.A(WX11346), .B(WX11025), .Z(II34586) ) ;
NAND2   gate17380  (.A(WX11346), .B(II34586), .Z(II34587) ) ;
NAND2   gate17381  (.A(WX11025), .B(II34586), .Z(II34588) ) ;
NAND2   gate17382  (.A(II34587), .B(II34588), .Z(II34585) ) ;
NAND2   gate17383  (.A(WX11089), .B(II34585), .Z(II34593) ) ;
NAND2   gate17384  (.A(WX11089), .B(II34593), .Z(II34594) ) ;
NAND2   gate17385  (.A(II34585), .B(II34593), .Z(II34595) ) ;
NAND2   gate17386  (.A(II34594), .B(II34595), .Z(II34584) ) ;
NAND2   gate17387  (.A(WX11153), .B(WX11217), .Z(II34601) ) ;
NAND2   gate17388  (.A(WX11153), .B(II34601), .Z(II34602) ) ;
NAND2   gate17389  (.A(WX11217), .B(II34601), .Z(II34603) ) ;
NAND2   gate17390  (.A(II34602), .B(II34603), .Z(II34600) ) ;
NAND2   gate17391  (.A(II34584), .B(II34600), .Z(II34608) ) ;
NAND2   gate17392  (.A(II34584), .B(II34608), .Z(II34609) ) ;
NAND2   gate17393  (.A(II34600), .B(II34608), .Z(II34610) ) ;
NAND2   gate17394  (.A(WX11346), .B(WX11027), .Z(II34617) ) ;
NAND2   gate17395  (.A(WX11346), .B(II34617), .Z(II34618) ) ;
NAND2   gate17396  (.A(WX11027), .B(II34617), .Z(II34619) ) ;
NAND2   gate17397  (.A(II34618), .B(II34619), .Z(II34616) ) ;
NAND2   gate17398  (.A(WX11091), .B(II34616), .Z(II34624) ) ;
NAND2   gate17399  (.A(WX11091), .B(II34624), .Z(II34625) ) ;
NAND2   gate17400  (.A(II34616), .B(II34624), .Z(II34626) ) ;
NAND2   gate17401  (.A(II34625), .B(II34626), .Z(II34615) ) ;
NAND2   gate17402  (.A(WX11155), .B(WX11219), .Z(II34632) ) ;
NAND2   gate17403  (.A(WX11155), .B(II34632), .Z(II34633) ) ;
NAND2   gate17404  (.A(WX11219), .B(II34632), .Z(II34634) ) ;
NAND2   gate17405  (.A(II34633), .B(II34634), .Z(II34631) ) ;
NAND2   gate17406  (.A(II34615), .B(II34631), .Z(II34639) ) ;
NAND2   gate17407  (.A(II34615), .B(II34639), .Z(II34640) ) ;
NAND2   gate17408  (.A(II34631), .B(II34639), .Z(II34641) ) ;
NAND2   gate17409  (.A(WX11346), .B(WX11029), .Z(II34648) ) ;
NAND2   gate17410  (.A(WX11346), .B(II34648), .Z(II34649) ) ;
NAND2   gate17411  (.A(WX11029), .B(II34648), .Z(II34650) ) ;
NAND2   gate17412  (.A(II34649), .B(II34650), .Z(II34647) ) ;
NAND2   gate17413  (.A(WX11093), .B(II34647), .Z(II34655) ) ;
NAND2   gate17414  (.A(WX11093), .B(II34655), .Z(II34656) ) ;
NAND2   gate17415  (.A(II34647), .B(II34655), .Z(II34657) ) ;
NAND2   gate17416  (.A(II34656), .B(II34657), .Z(II34646) ) ;
NAND2   gate17417  (.A(WX11157), .B(WX11221), .Z(II34663) ) ;
NAND2   gate17418  (.A(WX11157), .B(II34663), .Z(II34664) ) ;
NAND2   gate17419  (.A(WX11221), .B(II34663), .Z(II34665) ) ;
NAND2   gate17420  (.A(II34664), .B(II34665), .Z(II34662) ) ;
NAND2   gate17421  (.A(II34646), .B(II34662), .Z(II34670) ) ;
NAND2   gate17422  (.A(II34646), .B(II34670), .Z(II34671) ) ;
NAND2   gate17423  (.A(II34662), .B(II34670), .Z(II34672) ) ;
NAND2   gate17424  (.A(WX11346), .B(WX11031), .Z(II34679) ) ;
NAND2   gate17425  (.A(WX11346), .B(II34679), .Z(II34680) ) ;
NAND2   gate17426  (.A(WX11031), .B(II34679), .Z(II34681) ) ;
NAND2   gate17427  (.A(II34680), .B(II34681), .Z(II34678) ) ;
NAND2   gate17428  (.A(WX11095), .B(II34678), .Z(II34686) ) ;
NAND2   gate17429  (.A(WX11095), .B(II34686), .Z(II34687) ) ;
NAND2   gate17430  (.A(II34678), .B(II34686), .Z(II34688) ) ;
NAND2   gate17431  (.A(II34687), .B(II34688), .Z(II34677) ) ;
NAND2   gate17432  (.A(WX11159), .B(WX11223), .Z(II34694) ) ;
NAND2   gate17433  (.A(WX11159), .B(II34694), .Z(II34695) ) ;
NAND2   gate17434  (.A(WX11223), .B(II34694), .Z(II34696) ) ;
NAND2   gate17435  (.A(II34695), .B(II34696), .Z(II34693) ) ;
NAND2   gate17436  (.A(II34677), .B(II34693), .Z(II34701) ) ;
NAND2   gate17437  (.A(II34677), .B(II34701), .Z(II34702) ) ;
NAND2   gate17438  (.A(II34693), .B(II34701), .Z(II34703) ) ;
NAND2   gate17439  (.A(WX11346), .B(WX11033), .Z(II34710) ) ;
NAND2   gate17440  (.A(WX11346), .B(II34710), .Z(II34711) ) ;
NAND2   gate17441  (.A(WX11033), .B(II34710), .Z(II34712) ) ;
NAND2   gate17442  (.A(II34711), .B(II34712), .Z(II34709) ) ;
NAND2   gate17443  (.A(WX11097), .B(II34709), .Z(II34717) ) ;
NAND2   gate17444  (.A(WX11097), .B(II34717), .Z(II34718) ) ;
NAND2   gate17445  (.A(II34709), .B(II34717), .Z(II34719) ) ;
NAND2   gate17446  (.A(II34718), .B(II34719), .Z(II34708) ) ;
NAND2   gate17447  (.A(WX11161), .B(WX11225), .Z(II34725) ) ;
NAND2   gate17448  (.A(WX11161), .B(II34725), .Z(II34726) ) ;
NAND2   gate17449  (.A(WX11225), .B(II34725), .Z(II34727) ) ;
NAND2   gate17450  (.A(II34726), .B(II34727), .Z(II34724) ) ;
NAND2   gate17451  (.A(II34708), .B(II34724), .Z(II34732) ) ;
NAND2   gate17452  (.A(II34708), .B(II34732), .Z(II34733) ) ;
NAND2   gate17453  (.A(II34724), .B(II34732), .Z(II34734) ) ;
NAND2   gate17454  (.A(WX11346), .B(WX11035), .Z(II34741) ) ;
NAND2   gate17455  (.A(WX11346), .B(II34741), .Z(II34742) ) ;
NAND2   gate17456  (.A(WX11035), .B(II34741), .Z(II34743) ) ;
NAND2   gate17457  (.A(II34742), .B(II34743), .Z(II34740) ) ;
NAND2   gate17458  (.A(WX11099), .B(II34740), .Z(II34748) ) ;
NAND2   gate17459  (.A(WX11099), .B(II34748), .Z(II34749) ) ;
NAND2   gate17460  (.A(II34740), .B(II34748), .Z(II34750) ) ;
NAND2   gate17461  (.A(II34749), .B(II34750), .Z(II34739) ) ;
NAND2   gate17462  (.A(WX11163), .B(WX11227), .Z(II34756) ) ;
NAND2   gate17463  (.A(WX11163), .B(II34756), .Z(II34757) ) ;
NAND2   gate17464  (.A(WX11227), .B(II34756), .Z(II34758) ) ;
NAND2   gate17465  (.A(II34757), .B(II34758), .Z(II34755) ) ;
NAND2   gate17466  (.A(II34739), .B(II34755), .Z(II34763) ) ;
NAND2   gate17467  (.A(II34739), .B(II34763), .Z(II34764) ) ;
NAND2   gate17468  (.A(II34755), .B(II34763), .Z(II34765) ) ;
NAND2   gate17469  (.A(WX11346), .B(WX11037), .Z(II34772) ) ;
NAND2   gate17470  (.A(WX11346), .B(II34772), .Z(II34773) ) ;
NAND2   gate17471  (.A(WX11037), .B(II34772), .Z(II34774) ) ;
NAND2   gate17472  (.A(II34773), .B(II34774), .Z(II34771) ) ;
NAND2   gate17473  (.A(WX11101), .B(II34771), .Z(II34779) ) ;
NAND2   gate17474  (.A(WX11101), .B(II34779), .Z(II34780) ) ;
NAND2   gate17475  (.A(II34771), .B(II34779), .Z(II34781) ) ;
NAND2   gate17476  (.A(II34780), .B(II34781), .Z(II34770) ) ;
NAND2   gate17477  (.A(WX11165), .B(WX11229), .Z(II34787) ) ;
NAND2   gate17478  (.A(WX11165), .B(II34787), .Z(II34788) ) ;
NAND2   gate17479  (.A(WX11229), .B(II34787), .Z(II34789) ) ;
NAND2   gate17480  (.A(II34788), .B(II34789), .Z(II34786) ) ;
NAND2   gate17481  (.A(II34770), .B(II34786), .Z(II34794) ) ;
NAND2   gate17482  (.A(II34770), .B(II34794), .Z(II34795) ) ;
NAND2   gate17483  (.A(II34786), .B(II34794), .Z(II34796) ) ;
NAND2   gate17484  (.A(WX11346), .B(WX11039), .Z(II34803) ) ;
NAND2   gate17485  (.A(WX11346), .B(II34803), .Z(II34804) ) ;
NAND2   gate17486  (.A(WX11039), .B(II34803), .Z(II34805) ) ;
NAND2   gate17487  (.A(II34804), .B(II34805), .Z(II34802) ) ;
NAND2   gate17488  (.A(WX11103), .B(II34802), .Z(II34810) ) ;
NAND2   gate17489  (.A(WX11103), .B(II34810), .Z(II34811) ) ;
NAND2   gate17490  (.A(II34802), .B(II34810), .Z(II34812) ) ;
NAND2   gate17491  (.A(II34811), .B(II34812), .Z(II34801) ) ;
NAND2   gate17492  (.A(WX11167), .B(WX11231), .Z(II34818) ) ;
NAND2   gate17493  (.A(WX11167), .B(II34818), .Z(II34819) ) ;
NAND2   gate17494  (.A(WX11231), .B(II34818), .Z(II34820) ) ;
NAND2   gate17495  (.A(II34819), .B(II34820), .Z(II34817) ) ;
NAND2   gate17496  (.A(II34801), .B(II34817), .Z(II34825) ) ;
NAND2   gate17497  (.A(II34801), .B(II34825), .Z(II34826) ) ;
NAND2   gate17498  (.A(II34817), .B(II34825), .Z(II34827) ) ;
NAND2   gate17499  (.A(WX11346), .B(WX11041), .Z(II34834) ) ;
NAND2   gate17500  (.A(WX11346), .B(II34834), .Z(II34835) ) ;
NAND2   gate17501  (.A(WX11041), .B(II34834), .Z(II34836) ) ;
NAND2   gate17502  (.A(II34835), .B(II34836), .Z(II34833) ) ;
NAND2   gate17503  (.A(WX11105), .B(II34833), .Z(II34841) ) ;
NAND2   gate17504  (.A(WX11105), .B(II34841), .Z(II34842) ) ;
NAND2   gate17505  (.A(II34833), .B(II34841), .Z(II34843) ) ;
NAND2   gate17506  (.A(II34842), .B(II34843), .Z(II34832) ) ;
NAND2   gate17507  (.A(WX11169), .B(WX11233), .Z(II34849) ) ;
NAND2   gate17508  (.A(WX11169), .B(II34849), .Z(II34850) ) ;
NAND2   gate17509  (.A(WX11233), .B(II34849), .Z(II34851) ) ;
NAND2   gate17510  (.A(II34850), .B(II34851), .Z(II34848) ) ;
NAND2   gate17511  (.A(II34832), .B(II34848), .Z(II34856) ) ;
NAND2   gate17512  (.A(II34832), .B(II34856), .Z(II34857) ) ;
NAND2   gate17513  (.A(II34848), .B(II34856), .Z(II34858) ) ;
NAND2   gate17514  (.A(WX11346), .B(WX11043), .Z(II34865) ) ;
NAND2   gate17515  (.A(WX11346), .B(II34865), .Z(II34866) ) ;
NAND2   gate17516  (.A(WX11043), .B(II34865), .Z(II34867) ) ;
NAND2   gate17517  (.A(II34866), .B(II34867), .Z(II34864) ) ;
NAND2   gate17518  (.A(WX11107), .B(II34864), .Z(II34872) ) ;
NAND2   gate17519  (.A(WX11107), .B(II34872), .Z(II34873) ) ;
NAND2   gate17520  (.A(II34864), .B(II34872), .Z(II34874) ) ;
NAND2   gate17521  (.A(II34873), .B(II34874), .Z(II34863) ) ;
NAND2   gate17522  (.A(WX11171), .B(WX11235), .Z(II34880) ) ;
NAND2   gate17523  (.A(WX11171), .B(II34880), .Z(II34881) ) ;
NAND2   gate17524  (.A(WX11235), .B(II34880), .Z(II34882) ) ;
NAND2   gate17525  (.A(II34881), .B(II34882), .Z(II34879) ) ;
NAND2   gate17526  (.A(II34863), .B(II34879), .Z(II34887) ) ;
NAND2   gate17527  (.A(II34863), .B(II34887), .Z(II34888) ) ;
NAND2   gate17528  (.A(II34879), .B(II34887), .Z(II34889) ) ;
NAND2   gate17529  (.A(WX11346), .B(WX11045), .Z(II34896) ) ;
NAND2   gate17530  (.A(WX11346), .B(II34896), .Z(II34897) ) ;
NAND2   gate17531  (.A(WX11045), .B(II34896), .Z(II34898) ) ;
NAND2   gate17532  (.A(II34897), .B(II34898), .Z(II34895) ) ;
NAND2   gate17533  (.A(WX11109), .B(II34895), .Z(II34903) ) ;
NAND2   gate17534  (.A(WX11109), .B(II34903), .Z(II34904) ) ;
NAND2   gate17535  (.A(II34895), .B(II34903), .Z(II34905) ) ;
NAND2   gate17536  (.A(II34904), .B(II34905), .Z(II34894) ) ;
NAND2   gate17537  (.A(WX11173), .B(WX11237), .Z(II34911) ) ;
NAND2   gate17538  (.A(WX11173), .B(II34911), .Z(II34912) ) ;
NAND2   gate17539  (.A(WX11237), .B(II34911), .Z(II34913) ) ;
NAND2   gate17540  (.A(II34912), .B(II34913), .Z(II34910) ) ;
NAND2   gate17541  (.A(II34894), .B(II34910), .Z(II34918) ) ;
NAND2   gate17542  (.A(II34894), .B(II34918), .Z(II34919) ) ;
NAND2   gate17543  (.A(II34910), .B(II34918), .Z(II34920) ) ;
NAND2   gate17544  (.A(WX11346), .B(WX11047), .Z(II34927) ) ;
NAND2   gate17545  (.A(WX11346), .B(II34927), .Z(II34928) ) ;
NAND2   gate17546  (.A(WX11047), .B(II34927), .Z(II34929) ) ;
NAND2   gate17547  (.A(II34928), .B(II34929), .Z(II34926) ) ;
NAND2   gate17548  (.A(WX11111), .B(II34926), .Z(II34934) ) ;
NAND2   gate17549  (.A(WX11111), .B(II34934), .Z(II34935) ) ;
NAND2   gate17550  (.A(II34926), .B(II34934), .Z(II34936) ) ;
NAND2   gate17551  (.A(II34935), .B(II34936), .Z(II34925) ) ;
NAND2   gate17552  (.A(WX11175), .B(WX11239), .Z(II34942) ) ;
NAND2   gate17553  (.A(WX11175), .B(II34942), .Z(II34943) ) ;
NAND2   gate17554  (.A(WX11239), .B(II34942), .Z(II34944) ) ;
NAND2   gate17555  (.A(II34943), .B(II34944), .Z(II34941) ) ;
NAND2   gate17556  (.A(II34925), .B(II34941), .Z(II34949) ) ;
NAND2   gate17557  (.A(II34925), .B(II34949), .Z(II34950) ) ;
NAND2   gate17558  (.A(II34941), .B(II34949), .Z(II34951) ) ;
NAND2   gate17559  (.A(WX11346), .B(WX11049), .Z(II34958) ) ;
NAND2   gate17560  (.A(WX11346), .B(II34958), .Z(II34959) ) ;
NAND2   gate17561  (.A(WX11049), .B(II34958), .Z(II34960) ) ;
NAND2   gate17562  (.A(II34959), .B(II34960), .Z(II34957) ) ;
NAND2   gate17563  (.A(WX11113), .B(II34957), .Z(II34965) ) ;
NAND2   gate17564  (.A(WX11113), .B(II34965), .Z(II34966) ) ;
NAND2   gate17565  (.A(II34957), .B(II34965), .Z(II34967) ) ;
NAND2   gate17566  (.A(II34966), .B(II34967), .Z(II34956) ) ;
NAND2   gate17567  (.A(WX11177), .B(WX11241), .Z(II34973) ) ;
NAND2   gate17568  (.A(WX11177), .B(II34973), .Z(II34974) ) ;
NAND2   gate17569  (.A(WX11241), .B(II34973), .Z(II34975) ) ;
NAND2   gate17570  (.A(II34974), .B(II34975), .Z(II34972) ) ;
NAND2   gate17571  (.A(II34956), .B(II34972), .Z(II34980) ) ;
NAND2   gate17572  (.A(II34956), .B(II34980), .Z(II34981) ) ;
NAND2   gate17573  (.A(II34972), .B(II34980), .Z(II34982) ) ;
NAND2   gate17574  (.A(WX11346), .B(WX11051), .Z(II34989) ) ;
NAND2   gate17575  (.A(WX11346), .B(II34989), .Z(II34990) ) ;
NAND2   gate17576  (.A(WX11051), .B(II34989), .Z(II34991) ) ;
NAND2   gate17577  (.A(II34990), .B(II34991), .Z(II34988) ) ;
NAND2   gate17578  (.A(WX11115), .B(II34988), .Z(II34996) ) ;
NAND2   gate17579  (.A(WX11115), .B(II34996), .Z(II34997) ) ;
NAND2   gate17580  (.A(II34988), .B(II34996), .Z(II34998) ) ;
NAND2   gate17581  (.A(II34997), .B(II34998), .Z(II34987) ) ;
NAND2   gate17582  (.A(WX11179), .B(WX11243), .Z(II35004) ) ;
NAND2   gate17583  (.A(WX11179), .B(II35004), .Z(II35005) ) ;
NAND2   gate17584  (.A(WX11243), .B(II35004), .Z(II35006) ) ;
NAND2   gate17585  (.A(II35005), .B(II35006), .Z(II35003) ) ;
NAND2   gate17586  (.A(II34987), .B(II35003), .Z(II35011) ) ;
NAND2   gate17587  (.A(II34987), .B(II35011), .Z(II35012) ) ;
NAND2   gate17588  (.A(II35003), .B(II35011), .Z(II35013) ) ;
NAND2   gate17589  (.A(WX10924), .B(WX10829), .Z(II35092) ) ;
NAND2   gate17590  (.A(WX10924), .B(II35092), .Z(II35093) ) ;
NAND2   gate17591  (.A(WX10829), .B(II35092), .Z(II35094) ) ;
NAND2   gate17592  (.A(WX10925), .B(WX10831), .Z(II35105) ) ;
NAND2   gate17593  (.A(WX10925), .B(II35105), .Z(II35106) ) ;
NAND2   gate17594  (.A(WX10831), .B(II35105), .Z(II35107) ) ;
NAND2   gate17595  (.A(WX10926), .B(WX10833), .Z(II35118) ) ;
NAND2   gate17596  (.A(WX10926), .B(II35118), .Z(II35119) ) ;
NAND2   gate17597  (.A(WX10833), .B(II35118), .Z(II35120) ) ;
NAND2   gate17598  (.A(WX10927), .B(WX10835), .Z(II35131) ) ;
NAND2   gate17599  (.A(WX10927), .B(II35131), .Z(II35132) ) ;
NAND2   gate17600  (.A(WX10835), .B(II35131), .Z(II35133) ) ;
NAND2   gate17601  (.A(WX10928), .B(WX10837), .Z(II35144) ) ;
NAND2   gate17602  (.A(WX10928), .B(II35144), .Z(II35145) ) ;
NAND2   gate17603  (.A(WX10837), .B(II35144), .Z(II35146) ) ;
NAND2   gate17604  (.A(WX10929), .B(WX10839), .Z(II35157) ) ;
NAND2   gate17605  (.A(WX10929), .B(II35157), .Z(II35158) ) ;
NAND2   gate17606  (.A(WX10839), .B(II35157), .Z(II35159) ) ;
NAND2   gate17607  (.A(WX10930), .B(WX10841), .Z(II35170) ) ;
NAND2   gate17608  (.A(WX10930), .B(II35170), .Z(II35171) ) ;
NAND2   gate17609  (.A(WX10841), .B(II35170), .Z(II35172) ) ;
NAND2   gate17610  (.A(WX10931), .B(WX10843), .Z(II35183) ) ;
NAND2   gate17611  (.A(WX10931), .B(II35183), .Z(II35184) ) ;
NAND2   gate17612  (.A(WX10843), .B(II35183), .Z(II35185) ) ;
NAND2   gate17613  (.A(WX10932), .B(WX10845), .Z(II35196) ) ;
NAND2   gate17614  (.A(WX10932), .B(II35196), .Z(II35197) ) ;
NAND2   gate17615  (.A(WX10845), .B(II35196), .Z(II35198) ) ;
NAND2   gate17616  (.A(WX10933), .B(WX10847), .Z(II35209) ) ;
NAND2   gate17617  (.A(WX10933), .B(II35209), .Z(II35210) ) ;
NAND2   gate17618  (.A(WX10847), .B(II35209), .Z(II35211) ) ;
NAND2   gate17619  (.A(WX10934), .B(WX10849), .Z(II35222) ) ;
NAND2   gate17620  (.A(WX10934), .B(II35222), .Z(II35223) ) ;
NAND2   gate17621  (.A(WX10849), .B(II35222), .Z(II35224) ) ;
NAND2   gate17622  (.A(WX10935), .B(WX10851), .Z(II35235) ) ;
NAND2   gate17623  (.A(WX10935), .B(II35235), .Z(II35236) ) ;
NAND2   gate17624  (.A(WX10851), .B(II35235), .Z(II35237) ) ;
NAND2   gate17625  (.A(WX10936), .B(WX10853), .Z(II35248) ) ;
NAND2   gate17626  (.A(WX10936), .B(II35248), .Z(II35249) ) ;
NAND2   gate17627  (.A(WX10853), .B(II35248), .Z(II35250) ) ;
NAND2   gate17628  (.A(WX10937), .B(WX10855), .Z(II35261) ) ;
NAND2   gate17629  (.A(WX10937), .B(II35261), .Z(II35262) ) ;
NAND2   gate17630  (.A(WX10855), .B(II35261), .Z(II35263) ) ;
NAND2   gate17631  (.A(WX10938), .B(WX10857), .Z(II35274) ) ;
NAND2   gate17632  (.A(WX10938), .B(II35274), .Z(II35275) ) ;
NAND2   gate17633  (.A(WX10857), .B(II35274), .Z(II35276) ) ;
NAND2   gate17634  (.A(WX10939), .B(WX10859), .Z(II35287) ) ;
NAND2   gate17635  (.A(WX10939), .B(II35287), .Z(II35288) ) ;
NAND2   gate17636  (.A(WX10859), .B(II35287), .Z(II35289) ) ;
NAND2   gate17637  (.A(WX10940), .B(WX10861), .Z(II35300) ) ;
NAND2   gate17638  (.A(WX10940), .B(II35300), .Z(II35301) ) ;
NAND2   gate17639  (.A(WX10861), .B(II35300), .Z(II35302) ) ;
NAND2   gate17640  (.A(WX10941), .B(WX10863), .Z(II35313) ) ;
NAND2   gate17641  (.A(WX10941), .B(II35313), .Z(II35314) ) ;
NAND2   gate17642  (.A(WX10863), .B(II35313), .Z(II35315) ) ;
NAND2   gate17643  (.A(WX10942), .B(WX10865), .Z(II35326) ) ;
NAND2   gate17644  (.A(WX10942), .B(II35326), .Z(II35327) ) ;
NAND2   gate17645  (.A(WX10865), .B(II35326), .Z(II35328) ) ;
NAND2   gate17646  (.A(WX10943), .B(WX10867), .Z(II35339) ) ;
NAND2   gate17647  (.A(WX10943), .B(II35339), .Z(II35340) ) ;
NAND2   gate17648  (.A(WX10867), .B(II35339), .Z(II35341) ) ;
NAND2   gate17649  (.A(WX10944), .B(WX10869), .Z(II35352) ) ;
NAND2   gate17650  (.A(WX10944), .B(II35352), .Z(II35353) ) ;
NAND2   gate17651  (.A(WX10869), .B(II35352), .Z(II35354) ) ;
NAND2   gate17652  (.A(WX10945), .B(WX10871), .Z(II35365) ) ;
NAND2   gate17653  (.A(WX10945), .B(II35365), .Z(II35366) ) ;
NAND2   gate17654  (.A(WX10871), .B(II35365), .Z(II35367) ) ;
NAND2   gate17655  (.A(WX10946), .B(WX10873), .Z(II35378) ) ;
NAND2   gate17656  (.A(WX10946), .B(II35378), .Z(II35379) ) ;
NAND2   gate17657  (.A(WX10873), .B(II35378), .Z(II35380) ) ;
NAND2   gate17658  (.A(WX10947), .B(WX10875), .Z(II35391) ) ;
NAND2   gate17659  (.A(WX10947), .B(II35391), .Z(II35392) ) ;
NAND2   gate17660  (.A(WX10875), .B(II35391), .Z(II35393) ) ;
NAND2   gate17661  (.A(WX10948), .B(WX10877), .Z(II35404) ) ;
NAND2   gate17662  (.A(WX10948), .B(II35404), .Z(II35405) ) ;
NAND2   gate17663  (.A(WX10877), .B(II35404), .Z(II35406) ) ;
NAND2   gate17664  (.A(WX10949), .B(WX10879), .Z(II35417) ) ;
NAND2   gate17665  (.A(WX10949), .B(II35417), .Z(II35418) ) ;
NAND2   gate17666  (.A(WX10879), .B(II35417), .Z(II35419) ) ;
NAND2   gate17667  (.A(WX10950), .B(WX10881), .Z(II35430) ) ;
NAND2   gate17668  (.A(WX10950), .B(II35430), .Z(II35431) ) ;
NAND2   gate17669  (.A(WX10881), .B(II35430), .Z(II35432) ) ;
NAND2   gate17670  (.A(WX10951), .B(WX10883), .Z(II35443) ) ;
NAND2   gate17671  (.A(WX10951), .B(II35443), .Z(II35444) ) ;
NAND2   gate17672  (.A(WX10883), .B(II35443), .Z(II35445) ) ;
NAND2   gate17673  (.A(WX10952), .B(WX10885), .Z(II35456) ) ;
NAND2   gate17674  (.A(WX10952), .B(II35456), .Z(II35457) ) ;
NAND2   gate17675  (.A(WX10885), .B(II35456), .Z(II35458) ) ;
NAND2   gate17676  (.A(WX10953), .B(WX10887), .Z(II35469) ) ;
NAND2   gate17677  (.A(WX10953), .B(II35469), .Z(II35470) ) ;
NAND2   gate17678  (.A(WX10887), .B(II35469), .Z(II35471) ) ;
NAND2   gate17679  (.A(WX10954), .B(WX10889), .Z(II35482) ) ;
NAND2   gate17680  (.A(WX10954), .B(II35482), .Z(II35483) ) ;
NAND2   gate17681  (.A(WX10889), .B(II35482), .Z(II35484) ) ;
NAND2   gate17682  (.A(WX10955), .B(WX10891), .Z(II35495) ) ;
NAND2   gate17683  (.A(WX10955), .B(II35495), .Z(II35496) ) ;
NAND2   gate17684  (.A(WX10891), .B(II35495), .Z(II35497) ) ;
NAND2   gate17685  (.A(WX10971), .B(CRC_OUT_1_31), .Z(II35510) ) ;
NAND2   gate17686  (.A(WX10971), .B(II35510), .Z(II35511) ) ;
NAND2   gate17687  (.A(CRC_OUT_1_31), .B(II35510), .Z(II35512) ) ;
NAND2   gate17688  (.A(II35511), .B(II35512), .Z(II35509) ) ;
NAND2   gate17689  (.A(CRC_OUT_1_15), .B(II35509), .Z(II35517) ) ;
NAND2   gate17690  (.A(CRC_OUT_1_15), .B(II35517), .Z(II35518) ) ;
NAND2   gate17691  (.A(II35509), .B(II35517), .Z(II35519) ) ;
NAND2   gate17692  (.A(WX10976), .B(CRC_OUT_1_31), .Z(II35525) ) ;
NAND2   gate17693  (.A(WX10976), .B(II35525), .Z(II35526) ) ;
NAND2   gate17694  (.A(CRC_OUT_1_31), .B(II35525), .Z(II35527) ) ;
NAND2   gate17695  (.A(II35526), .B(II35527), .Z(II35524) ) ;
NAND2   gate17696  (.A(CRC_OUT_1_10), .B(II35524), .Z(II35532) ) ;
NAND2   gate17697  (.A(CRC_OUT_1_10), .B(II35532), .Z(II35533) ) ;
NAND2   gate17698  (.A(II35524), .B(II35532), .Z(II35534) ) ;
NAND2   gate17699  (.A(WX10983), .B(CRC_OUT_1_31), .Z(II35540) ) ;
NAND2   gate17700  (.A(WX10983), .B(II35540), .Z(II35541) ) ;
NAND2   gate17701  (.A(CRC_OUT_1_31), .B(II35540), .Z(II35542) ) ;
NAND2   gate17702  (.A(II35541), .B(II35542), .Z(II35539) ) ;
NAND2   gate17703  (.A(CRC_OUT_1_3), .B(II35539), .Z(II35547) ) ;
NAND2   gate17704  (.A(CRC_OUT_1_3), .B(II35547), .Z(II35548) ) ;
NAND2   gate17705  (.A(II35539), .B(II35547), .Z(II35549) ) ;
NAND2   gate17706  (.A(WX10987), .B(CRC_OUT_1_31), .Z(II35554) ) ;
NAND2   gate17707  (.A(WX10987), .B(II35554), .Z(II35555) ) ;
NAND2   gate17708  (.A(CRC_OUT_1_31), .B(II35554), .Z(II35556) ) ;
NAND2   gate17709  (.A(WX10956), .B(CRC_OUT_1_30), .Z(II35561) ) ;
NAND2   gate17710  (.A(WX10956), .B(II35561), .Z(II35562) ) ;
NAND2   gate17711  (.A(CRC_OUT_1_30), .B(II35561), .Z(II35563) ) ;
NAND2   gate17712  (.A(WX10957), .B(CRC_OUT_1_29), .Z(II35568) ) ;
NAND2   gate17713  (.A(WX10957), .B(II35568), .Z(II35569) ) ;
NAND2   gate17714  (.A(CRC_OUT_1_29), .B(II35568), .Z(II35570) ) ;
NAND2   gate17715  (.A(WX10958), .B(CRC_OUT_1_28), .Z(II35575) ) ;
NAND2   gate17716  (.A(WX10958), .B(II35575), .Z(II35576) ) ;
NAND2   gate17717  (.A(CRC_OUT_1_28), .B(II35575), .Z(II35577) ) ;
NAND2   gate17718  (.A(WX10959), .B(CRC_OUT_1_27), .Z(II35582) ) ;
NAND2   gate17719  (.A(WX10959), .B(II35582), .Z(II35583) ) ;
NAND2   gate17720  (.A(CRC_OUT_1_27), .B(II35582), .Z(II35584) ) ;
NAND2   gate17721  (.A(WX10960), .B(CRC_OUT_1_26), .Z(II35589) ) ;
NAND2   gate17722  (.A(WX10960), .B(II35589), .Z(II35590) ) ;
NAND2   gate17723  (.A(CRC_OUT_1_26), .B(II35589), .Z(II35591) ) ;
NAND2   gate17724  (.A(WX10961), .B(CRC_OUT_1_25), .Z(II35596) ) ;
NAND2   gate17725  (.A(WX10961), .B(II35596), .Z(II35597) ) ;
NAND2   gate17726  (.A(CRC_OUT_1_25), .B(II35596), .Z(II35598) ) ;
NAND2   gate17727  (.A(WX10962), .B(CRC_OUT_1_24), .Z(II35603) ) ;
NAND2   gate17728  (.A(WX10962), .B(II35603), .Z(II35604) ) ;
NAND2   gate17729  (.A(CRC_OUT_1_24), .B(II35603), .Z(II35605) ) ;
NAND2   gate17730  (.A(WX10963), .B(CRC_OUT_1_23), .Z(II35610) ) ;
NAND2   gate17731  (.A(WX10963), .B(II35610), .Z(II35611) ) ;
NAND2   gate17732  (.A(CRC_OUT_1_23), .B(II35610), .Z(II35612) ) ;
NAND2   gate17733  (.A(WX10964), .B(CRC_OUT_1_22), .Z(II35617) ) ;
NAND2   gate17734  (.A(WX10964), .B(II35617), .Z(II35618) ) ;
NAND2   gate17735  (.A(CRC_OUT_1_22), .B(II35617), .Z(II35619) ) ;
NAND2   gate17736  (.A(WX10965), .B(CRC_OUT_1_21), .Z(II35624) ) ;
NAND2   gate17737  (.A(WX10965), .B(II35624), .Z(II35625) ) ;
NAND2   gate17738  (.A(CRC_OUT_1_21), .B(II35624), .Z(II35626) ) ;
NAND2   gate17739  (.A(WX10966), .B(CRC_OUT_1_20), .Z(II35631) ) ;
NAND2   gate17740  (.A(WX10966), .B(II35631), .Z(II35632) ) ;
NAND2   gate17741  (.A(CRC_OUT_1_20), .B(II35631), .Z(II35633) ) ;
NAND2   gate17742  (.A(WX10967), .B(CRC_OUT_1_19), .Z(II35638) ) ;
NAND2   gate17743  (.A(WX10967), .B(II35638), .Z(II35639) ) ;
NAND2   gate17744  (.A(CRC_OUT_1_19), .B(II35638), .Z(II35640) ) ;
NAND2   gate17745  (.A(WX10968), .B(CRC_OUT_1_18), .Z(II35645) ) ;
NAND2   gate17746  (.A(WX10968), .B(II35645), .Z(II35646) ) ;
NAND2   gate17747  (.A(CRC_OUT_1_18), .B(II35645), .Z(II35647) ) ;
NAND2   gate17748  (.A(WX10969), .B(CRC_OUT_1_17), .Z(II35652) ) ;
NAND2   gate17749  (.A(WX10969), .B(II35652), .Z(II35653) ) ;
NAND2   gate17750  (.A(CRC_OUT_1_17), .B(II35652), .Z(II35654) ) ;
NAND2   gate17751  (.A(WX10970), .B(CRC_OUT_1_16), .Z(II35659) ) ;
NAND2   gate17752  (.A(WX10970), .B(II35659), .Z(II35660) ) ;
NAND2   gate17753  (.A(CRC_OUT_1_16), .B(II35659), .Z(II35661) ) ;
NAND2   gate17754  (.A(WX10972), .B(CRC_OUT_1_14), .Z(II35666) ) ;
NAND2   gate17755  (.A(WX10972), .B(II35666), .Z(II35667) ) ;
NAND2   gate17756  (.A(CRC_OUT_1_14), .B(II35666), .Z(II35668) ) ;
NAND2   gate17757  (.A(WX10973), .B(CRC_OUT_1_13), .Z(II35673) ) ;
NAND2   gate17758  (.A(WX10973), .B(II35673), .Z(II35674) ) ;
NAND2   gate17759  (.A(CRC_OUT_1_13), .B(II35673), .Z(II35675) ) ;
NAND2   gate17760  (.A(WX10974), .B(CRC_OUT_1_12), .Z(II35680) ) ;
NAND2   gate17761  (.A(WX10974), .B(II35680), .Z(II35681) ) ;
NAND2   gate17762  (.A(CRC_OUT_1_12), .B(II35680), .Z(II35682) ) ;
NAND2   gate17763  (.A(WX10975), .B(CRC_OUT_1_11), .Z(II35687) ) ;
NAND2   gate17764  (.A(WX10975), .B(II35687), .Z(II35688) ) ;
NAND2   gate17765  (.A(CRC_OUT_1_11), .B(II35687), .Z(II35689) ) ;
NAND2   gate17766  (.A(WX10977), .B(CRC_OUT_1_9), .Z(II35694) ) ;
NAND2   gate17767  (.A(WX10977), .B(II35694), .Z(II35695) ) ;
NAND2   gate17768  (.A(CRC_OUT_1_9), .B(II35694), .Z(II35696) ) ;
NAND2   gate17769  (.A(WX10978), .B(CRC_OUT_1_8), .Z(II35701) ) ;
NAND2   gate17770  (.A(WX10978), .B(II35701), .Z(II35702) ) ;
NAND2   gate17771  (.A(CRC_OUT_1_8), .B(II35701), .Z(II35703) ) ;
NAND2   gate17772  (.A(WX10979), .B(CRC_OUT_1_7), .Z(II35708) ) ;
NAND2   gate17773  (.A(WX10979), .B(II35708), .Z(II35709) ) ;
NAND2   gate17774  (.A(CRC_OUT_1_7), .B(II35708), .Z(II35710) ) ;
NAND2   gate17775  (.A(WX10980), .B(CRC_OUT_1_6), .Z(II35715) ) ;
NAND2   gate17776  (.A(WX10980), .B(II35715), .Z(II35716) ) ;
NAND2   gate17777  (.A(CRC_OUT_1_6), .B(II35715), .Z(II35717) ) ;
NAND2   gate17778  (.A(WX10981), .B(CRC_OUT_1_5), .Z(II35722) ) ;
NAND2   gate17779  (.A(WX10981), .B(II35722), .Z(II35723) ) ;
NAND2   gate17780  (.A(CRC_OUT_1_5), .B(II35722), .Z(II35724) ) ;
NAND2   gate17781  (.A(WX10982), .B(CRC_OUT_1_4), .Z(II35729) ) ;
NAND2   gate17782  (.A(WX10982), .B(II35729), .Z(II35730) ) ;
NAND2   gate17783  (.A(CRC_OUT_1_4), .B(II35729), .Z(II35731) ) ;
NAND2   gate17784  (.A(WX10984), .B(CRC_OUT_1_2), .Z(II35736) ) ;
NAND2   gate17785  (.A(WX10984), .B(II35736), .Z(II35737) ) ;
NAND2   gate17786  (.A(CRC_OUT_1_2), .B(II35736), .Z(II35738) ) ;
NAND2   gate17787  (.A(WX10985), .B(CRC_OUT_1_1), .Z(II35743) ) ;
NAND2   gate17788  (.A(WX10985), .B(II35743), .Z(II35744) ) ;
NAND2   gate17789  (.A(CRC_OUT_1_1), .B(II35743), .Z(II35745) ) ;
NAND2   gate17790  (.A(WX10986), .B(CRC_OUT_1_0), .Z(II35750) ) ;
NAND2   gate17791  (.A(WX10986), .B(II35750), .Z(II35751) ) ;
NAND2   gate17792  (.A(CRC_OUT_1_0), .B(II35750), .Z(II35752) ) ;

endmodule
