module s9234 (g89, g94, g98, g102, g107
    , g301, g306, g310, g314, g319
    , g557, g558, g559, g560, g561
    , g562, g563, g564, g705, CLK
    , g2584, g3222, g3600, g4307, g4321
    , g4422, g4809, g5137, g5468, g5469
    , g5692, g6282, g6284, g6360, g6362
    , g6364, g6366, g6368, g6370, g6372
    , g6374, g6728) ;

input   g89, g94, g98, g102, g107
    , g301, g306, g310, g314, g319
    , g557, g558, g559, g560, g561
    , g562, g563, g564, g705, CLK ;

output  g2584, g3222, g3600, g4307, g4321
    , g4422, g4809, g5137, g5468, g5469
    , g5692, g6282, g6284, g6360, g6362
    , g6364, g6366, g6368, g6370, g6372
    , g6374, g6728 ;

INV     gate0  (.A(II3705), .Z(g2584) ) ;
INV     gate1  (.A(II4465), .Z(g3222) ) ;
INV     gate2  (.A(II4791), .Z(g3600) ) ;
INV     gate3  (.A(II5774), .Z(g4307) ) ;
INV     gate4  (.A(II5790), .Z(g4321) ) ;
INV     gate5  (.A(g4111), .Z(g4422) ) ;
INV     gate6  (.A(II6485), .Z(g4809) ) ;
INV     gate7  (.A(II6789), .Z(g5137) ) ;
INV     gate8  (.A(II7150), .Z(g5468) ) ;
INV     gate9  (.A(II7153), .Z(g5469) ) ;
INV     gate10  (.A(II7451), .Z(g5692) ) ;
INV     gate11  (.A(II7996), .Z(g6282) ) ;
INV     gate12  (.A(II8002), .Z(g6284) ) ;
INV     gate13  (.A(II8144), .Z(g6360) ) ;
INV     gate14  (.A(II8150), .Z(g6362) ) ;
INV     gate15  (.A(II8156), .Z(g6364) ) ;
INV     gate16  (.A(II8162), .Z(g6366) ) ;
INV     gate17  (.A(II8168), .Z(g6368) ) ;
INV     gate18  (.A(II8174), .Z(g6370) ) ;
INV     gate19  (.A(II8180), .Z(g6372) ) ;
INV     gate20  (.A(II8186), .Z(g6374) ) ;
INV     gate21  (.A(II8878), .Z(g6728) ) ;
INV     gate22  (.A(II5409), .Z(g4109) ) ;
DFF     gate23  (.D(g4109), .CP(CLK), .Q(g46) ) ;
INV     gate24  (.A(II5406), .Z(g4108) ) ;
DFF     gate25  (.D(g4108), .CP(CLK), .Q(g45) ) ;
INV     gate26  (.A(II5403), .Z(g4107) ) ;
DFF     gate27  (.D(g4107), .CP(CLK), .Q(g44) ) ;
INV     gate28  (.A(II5400), .Z(g4106) ) ;
DFF     gate29  (.D(g4106), .CP(CLK), .Q(g42) ) ;
INV     gate30  (.A(II5397), .Z(g4105) ) ;
DFF     gate31  (.D(g4105), .CP(CLK), .Q(g40) ) ;
INV     gate32  (.A(II5391), .Z(g4103) ) ;
DFF     gate33  (.D(g4103), .CP(CLK), .Q(g39) ) ;
INV     gate34  (.A(II5388), .Z(g4102) ) ;
DFF     gate35  (.D(g4102), .CP(CLK), .Q(g38) ) ;
INV     gate36  (.A(II5385), .Z(g4101) ) ;
DFF     gate37  (.D(g4101), .CP(CLK), .Q(g37) ) ;
INV     gate38  (.A(II5382), .Z(g4100) ) ;
DFF     gate39  (.D(g4100), .CP(CLK), .Q(g36) ) ;
INV     gate40  (.A(II5379), .Z(g4099) ) ;
DFF     gate41  (.D(g4099), .CP(CLK), .Q(g32) ) ;
INV     gate42  (.A(II8875), .Z(g6727) ) ;
DFF     gate43  (.D(g6727), .CP(CLK), .Q(g28) ) ;
INV     gate44  (.A(II8872), .Z(g6726) ) ;
DFF     gate45  (.D(g6726), .CP(CLK), .Q(g24) ) ;
INV     gate46  (.A(II8869), .Z(g6725) ) ;
DFF     gate47  (.D(g6725), .CP(CLK), .Q(g18) ) ;
INV     gate48  (.A(II8866), .Z(g6724) ) ;
DFF     gate49  (.D(g6724), .CP(CLK), .Q(g14) ) ;
INV     gate50  (.A(II8863), .Z(g6723) ) ;
DFF     gate51  (.D(g6723), .CP(CLK), .Q(g10) ) ;
INV     gate52  (.A(II8860), .Z(g6722) ) ;
DFF     gate53  (.D(g6722), .CP(CLK), .Q(g6) ) ;
INV     gate54  (.A(II8857), .Z(g6721) ) ;
DFF     gate55  (.D(g6721), .CP(CLK), .Q(g2) ) ;
INV     gate56  (.A(II8854), .Z(g6720) ) ;
DFF     gate57  (.D(g6720), .CP(CLK), .Q(g1) ) ;
INV     gate58  (.A(II8881), .Z(g6729) ) ;
DFF     gate59  (.D(g6729), .CP(CLK), .Q(g48) ) ;
INV     gate60  (.A(II5418), .Z(g4112) ) ;
DFF     gate61  (.D(g4112), .CP(CLK), .Q(g47) ) ;
INV     gate62  (.A(II5412), .Z(g4110) ) ;
DFF     gate63  (.D(g4110), .CP(CLK), .Q(g41) ) ;
INV     gate64  (.A(II5394), .Z(g4104) ) ;
DFF     gate65  (.D(g4104), .CP(CLK), .Q(g22) ) ;
INV     gate66  (.A(II5376), .Z(g4098) ) ;
DFF     gate67  (.D(g4098), .CP(CLK), .Q(g23) ) ;
INV     gate68  (.A(II4471), .Z(g3224) ) ;
DFF     gate69  (.D(g3224), .CP(CLK), .Q(g284) ) ;
INV     gate70  (.A(II4474), .Z(g3225) ) ;
DFF     gate71  (.D(g3225), .CP(CLK), .Q(g285) ) ;
INV     gate72  (.A(II4477), .Z(g3226) ) ;
DFF     gate73  (.D(g3226), .CP(CLK), .Q(g286) ) ;
INV     gate74  (.A(II4480), .Z(g3227) ) ;
DFF     gate75  (.D(g3227), .CP(CLK), .Q(g287) ) ;
INV     gate76  (.A(II4483), .Z(g3228) ) ;
DFF     gate77  (.D(g3228), .CP(CLK), .Q(g288) ) ;
INV     gate78  (.A(II4486), .Z(g3229) ) ;
DFF     gate79  (.D(g3229), .CP(CLK), .Q(g289) ) ;
INV     gate80  (.A(II4489), .Z(g3230) ) ;
DFF     gate81  (.D(g3230), .CP(CLK), .Q(g290) ) ;
INV     gate82  (.A(II4492), .Z(g3231) ) ;
DFF     gate83  (.D(g3231), .CP(CLK), .Q(g291) ) ;
INV     gate84  (.A(II4495), .Z(g3232) ) ;
DFF     gate85  (.D(g3232), .CP(CLK), .Q(g292) ) ;
INV     gate86  (.A(II7161), .Z(g5475) ) ;
DFF     gate87  (.D(g5475), .CP(CLK), .Q(g338) ) ;
INV     gate88  (.A(II7164), .Z(g5476) ) ;
DFF     gate89  (.D(g5476), .CP(CLK), .Q(g341) ) ;
INV     gate90  (.A(II7167), .Z(g5477) ) ;
DFF     gate91  (.D(g5477), .CP(CLK), .Q(g345) ) ;
INV     gate92  (.A(II7170), .Z(g5478) ) ;
DFF     gate93  (.D(g5478), .CP(CLK), .Q(g349) ) ;
INV     gate94  (.A(II7173), .Z(g5479) ) ;
DFF     gate95  (.D(g5479), .CP(CLK), .Q(g353) ) ;
INV     gate96  (.A(II7176), .Z(g5480) ) ;
DFF     gate97  (.D(g5480), .CP(CLK), .Q(g357) ) ;
INV     gate98  (.A(II8614), .Z(g6582) ) ;
DFF     gate99  (.D(g6582), .CP(CLK), .Q(g361) ) ;
INV     gate100  (.A(II8617), .Z(g6583) ) ;
DFF     gate101  (.D(g6583), .CP(CLK), .Q(g49) ) ;
INV     gate102  (.A(II8620), .Z(g6584) ) ;
DFF     gate103  (.D(g6584), .CP(CLK), .Q(g54) ) ;
INV     gate104  (.A(II8623), .Z(g6585) ) ;
DFF     gate105  (.D(g6585), .CP(CLK), .Q(g59) ) ;
INV     gate106  (.A(II8626), .Z(g6586) ) ;
DFF     gate107  (.D(g6586), .CP(CLK), .Q(g64) ) ;
INV     gate108  (.A(II8629), .Z(g6587) ) ;
DFF     gate109  (.D(g6587), .CP(CLK), .Q(g69) ) ;
INV     gate110  (.A(II8632), .Z(g6588) ) ;
DFF     gate111  (.D(g6588), .CP(CLK), .Q(g74) ) ;
INV     gate112  (.A(II8635), .Z(g6589) ) ;
DFF     gate113  (.D(g6589), .CP(CLK), .Q(g79) ) ;
INV     gate114  (.A(II8638), .Z(g6590) ) ;
DFF     gate115  (.D(g6590), .CP(CLK), .Q(g84) ) ;
INV     gate116  (.A(II7966), .Z(g6278) ) ;
DFF     gate117  (.D(g6278), .CP(CLK), .Q(g366) ) ;
OR2     gate118  (.A(g5632), .B(g5481), .Z(g5693) ) ;
DFF     gate119  (.D(g5693), .CP(CLK), .Q(g370) ) ;
OR2     gate120  (.A(g5633), .B(g5482), .Z(g5694) ) ;
DFF     gate121  (.D(g5694), .CP(CLK), .Q(g374) ) ;
OR2     gate122  (.A(g5635), .B(g5483), .Z(g5695) ) ;
DFF     gate123  (.D(g5695), .CP(CLK), .Q(g378) ) ;
OR2     gate124  (.A(g5637), .B(g5484), .Z(g5696) ) ;
DFF     gate125  (.D(g5696), .CP(CLK), .Q(g382) ) ;
OR2     gate126  (.A(g5646), .B(g5485), .Z(g5697) ) ;
DFF     gate127  (.D(g5697), .CP(CLK), .Q(g386) ) ;
OR2     gate128  (.A(g5648), .B(g5486), .Z(g5698) ) ;
DFF     gate129  (.D(g5698), .CP(CLK), .Q(g390) ) ;
OR2     gate130  (.A(g5660), .B(g5487), .Z(g5699) ) ;
DFF     gate131  (.D(g5699), .CP(CLK), .Q(g394) ) ;
OR2     gate132  (.A(g5663), .B(g5488), .Z(g5700) ) ;
DFF     gate133  (.D(g5700), .CP(CLK), .Q(g398) ) ;
INV     gate134  (.A(II6528), .Z(g4840) ) ;
DFF     gate135  (.D(g4840), .CP(CLK), .Q(g326) ) ;
INV     gate136  (.A(II5433), .Z(g4117) ) ;
DFF     gate137  (.D(g4117), .CP(CLK), .Q(g327) ) ;
INV     gate138  (.A(II5436), .Z(g4118) ) ;
DFF     gate139  (.D(g4118), .CP(CLK), .Q(g328) ) ;
INV     gate140  (.A(II5439), .Z(g4119) ) ;
DFF     gate141  (.D(g4119), .CP(CLK), .Q(g331) ) ;
INV     gate142  (.A(II5442), .Z(g4120) ) ;
DFF     gate143  (.D(g4120), .CP(CLK), .Q(g323) ) ;
INV     gate144  (.A(II9002), .Z(g6823) ) ;
DFF     gate145  (.D(g6823), .CP(CLK), .Q(g332) ) ;
INV     gate146  (.A(II9208), .Z(g6925) ) ;
DFF     gate147  (.D(g6925), .CP(CLK), .Q(g336) ) ;
INV     gate148  (.A(II3708), .Z(g2585) ) ;
DFF     gate149  (.D(g2585), .CP(CLK), .Q(g337) ) ;
INV     gate150  (.A(II6792), .Z(g5138) ) ;
DFF     gate151  (.D(g5138), .CP(CLK), .Q(g128) ) ;
INV     gate152  (.A(II6795), .Z(g5139) ) ;
DFF     gate153  (.D(g5139), .CP(CLK), .Q(g131) ) ;
INV     gate154  (.A(II6798), .Z(g5140) ) ;
DFF     gate155  (.D(g5140), .CP(CLK), .Q(g135) ) ;
INV     gate156  (.A(II6801), .Z(g5141) ) ;
DFF     gate157  (.D(g5141), .CP(CLK), .Q(g139) ) ;
INV     gate158  (.A(II8217), .Z(g6401) ) ;
DFF     gate159  (.D(g6401), .CP(CLK), .Q(g143) ) ;
INV     gate160  (.A(II8220), .Z(g6402) ) ;
DFF     gate161  (.D(g6402), .CP(CLK), .Q(g152) ) ;
INV     gate162  (.A(II8223), .Z(g6403) ) ;
DFF     gate163  (.D(g6403), .CP(CLK), .Q(g161) ) ;
INV     gate164  (.A(II8226), .Z(g6404) ) ;
DFF     gate165  (.D(g6404), .CP(CLK), .Q(g170) ) ;
INV     gate166  (.A(II8229), .Z(g6405) ) ;
DFF     gate167  (.D(g6405), .CP(CLK), .Q(g179) ) ;
INV     gate168  (.A(II8232), .Z(g6406) ) ;
DFF     gate169  (.D(g6406), .CP(CLK), .Q(g188) ) ;
INV     gate170  (.A(II7634), .Z(g5874) ) ;
DFF     gate171  (.D(g5874), .CP(CLK), .Q(g148) ) ;
OR2     gate172  (.A(g5359), .B(g5142), .Z(g5470) ) ;
DFF     gate173  (.D(g5470), .CP(CLK), .Q(g157) ) ;
OR2     gate174  (.A(g5360), .B(g5143), .Z(g5471) ) ;
DFF     gate175  (.D(g5471), .CP(CLK), .Q(g166) ) ;
OR2     gate176  (.A(g5361), .B(g5144), .Z(g5472) ) ;
DFF     gate177  (.D(g5472), .CP(CLK), .Q(g175) ) ;
OR2     gate178  (.A(g5362), .B(g5145), .Z(g5473) ) ;
DFF     gate179  (.D(g5473), .CP(CLK), .Q(g184) ) ;
OR2     gate180  (.A(g5363), .B(g5146), .Z(g5474) ) ;
DFF     gate181  (.D(g5474), .CP(CLK), .Q(g193) ) ;
INV     gate182  (.A(II6525), .Z(g4839) ) ;
DFF     gate183  (.D(g4839), .CP(CLK), .Q(g117) ) ;
INV     gate184  (.A(II5421), .Z(g4113) ) ;
DFF     gate185  (.D(g4113), .CP(CLK), .Q(g118) ) ;
INV     gate186  (.A(II5424), .Z(g4114) ) ;
DFF     gate187  (.D(g4114), .CP(CLK), .Q(g119) ) ;
INV     gate188  (.A(II5427), .Z(g4115) ) ;
DFF     gate189  (.D(g4115), .CP(CLK), .Q(g122) ) ;
INV     gate190  (.A(II5430), .Z(g4116) ) ;
DFF     gate191  (.D(g4116), .CP(CLK), .Q(g114) ) ;
INV     gate192  (.A(II9233), .Z(g6940) ) ;
DFF     gate193  (.D(g6940), .CP(CLK), .Q(g123) ) ;
INV     gate194  (.A(II7963), .Z(g6277) ) ;
DFF     gate195  (.D(g6277), .CP(CLK), .Q(g111) ) ;
INV     gate196  (.A(II9236), .Z(g6941) ) ;
DFF     gate197  (.D(g6941), .CP(CLK), .Q(g127) ) ;
INV     gate198  (.A(II7643), .Z(g5877) ) ;
DFF     gate199  (.D(g5877), .CP(CLK), .Q(g276) ) ;
INV     gate200  (.A(II7808), .Z(g6104) ) ;
DFF     gate201  (.D(g6104), .CP(CLK), .Q(g277) ) ;
INV     gate202  (.A(II7811), .Z(g6105) ) ;
DFF     gate203  (.D(g6105), .CP(CLK), .Q(g278) ) ;
INV     gate204  (.A(II7814), .Z(g6106) ) ;
DFF     gate205  (.D(g6106), .CP(CLK), .Q(g279) ) ;
INV     gate206  (.A(II7646), .Z(g5878) ) ;
DFF     gate207  (.D(g5878), .CP(CLK), .Q(g280) ) ;
INV     gate208  (.A(II7817), .Z(g6107) ) ;
DFF     gate209  (.D(g6107), .CP(CLK), .Q(g281) ) ;
INV     gate210  (.A(II9044), .Z(g6841) ) ;
DFF     gate211  (.D(g6841), .CP(CLK), .Q(g282) ) ;
INV     gate212  (.A(II9047), .Z(g6842) ) ;
DFF     gate213  (.D(g6842), .CP(CLK), .Q(g283) ) ;
INV     gate214  (.A(II7637), .Z(g5875) ) ;
DFF     gate215  (.D(g5875), .CP(CLK), .Q(g204) ) ;
INV     gate216  (.A(II7796), .Z(g6100) ) ;
DFF     gate217  (.D(g6100), .CP(CLK), .Q(g205) ) ;
INV     gate218  (.A(II7799), .Z(g6101) ) ;
DFF     gate219  (.D(g6101), .CP(CLK), .Q(g206) ) ;
INV     gate220  (.A(II7802), .Z(g6102) ) ;
DFF     gate221  (.D(g6102), .CP(CLK), .Q(g207) ) ;
INV     gate222  (.A(II7640), .Z(g5876) ) ;
DFF     gate223  (.D(g5876), .CP(CLK), .Q(g208) ) ;
INV     gate224  (.A(II7805), .Z(g6103) ) ;
DFF     gate225  (.D(g6103), .CP(CLK), .Q(g209) ) ;
INV     gate226  (.A(II9038), .Z(g6839) ) ;
DFF     gate227  (.D(g6839), .CP(CLK), .Q(g210) ) ;
INV     gate228  (.A(II9041), .Z(g6840) ) ;
DFF     gate229  (.D(g6840), .CP(CLK), .Q(g211) ) ;
INV     gate230  (.A(II4498), .Z(g3233) ) ;
DFF     gate231  (.D(g3233), .CP(CLK), .Q(g212) ) ;
INV     gate232  (.A(II4501), .Z(g3234) ) ;
DFF     gate233  (.D(g3234), .CP(CLK), .Q(g218) ) ;
INV     gate234  (.A(II4504), .Z(g3235) ) ;
DFF     gate235  (.D(g3235), .CP(CLK), .Q(g224) ) ;
INV     gate236  (.A(II4507), .Z(g3236) ) ;
DFF     gate237  (.D(g3236), .CP(CLK), .Q(g230) ) ;
INV     gate238  (.A(II4510), .Z(g3237) ) ;
DFF     gate239  (.D(g3237), .CP(CLK), .Q(g236) ) ;
INV     gate240  (.A(II4513), .Z(g3238) ) ;
DFF     gate241  (.D(g3238), .CP(CLK), .Q(g242) ) ;
INV     gate242  (.A(II4516), .Z(g3239) ) ;
DFF     gate243  (.D(g3239), .CP(CLK), .Q(g248) ) ;
INV     gate244  (.A(II4519), .Z(g3240) ) ;
DFF     gate245  (.D(g3240), .CP(CLK), .Q(g254) ) ;
INV     gate246  (.A(II4522), .Z(g3241) ) ;
DFF     gate247  (.D(g3241), .CP(CLK), .Q(g260) ) ;
INV     gate248  (.A(II5445), .Z(g4121) ) ;
DFF     gate249  (.D(g4121), .CP(CLK), .Q(g567) ) ;
INV     gate250  (.A(II5448), .Z(g4122) ) ;
DFF     gate251  (.D(g4122), .CP(CLK), .Q(g598) ) ;
INV     gate252  (.A(II5923), .Z(g4424) ) ;
DFF     gate253  (.D(g4424), .CP(CLK), .Q(g634) ) ;
INV     gate254  (.A(II6247), .Z(g4658) ) ;
DFF     gate255  (.D(g4658), .CP(CLK), .Q(g642) ) ;
INV     gate256  (.A(II6579), .Z(g4857) ) ;
DFF     gate257  (.D(g4857), .CP(CLK), .Q(g606) ) ;
INV     gate258  (.A(II6812), .Z(g5148) ) ;
DFF     gate259  (.D(g5148), .CP(CLK), .Q(g646) ) ;
INV     gate260  (.A(II6989), .Z(g5329) ) ;
DFF     gate261  (.D(g5329), .CP(CLK), .Q(g650) ) ;
INV     gate262  (.A(II7190), .Z(g5490) ) ;
DFF     gate263  (.D(g5490), .CP(CLK), .Q(g654) ) ;
INV     gate264  (.A(II7336), .Z(g5580) ) ;
DFF     gate265  (.D(g5580), .CP(CLK), .Q(g571) ) ;
INV     gate266  (.A(II8644), .Z(g6592) ) ;
DFF     gate267  (.D(g6592), .CP(CLK), .Q(g578) ) ;
INV     gate268  (.A(II8647), .Z(g6593) ) ;
DFF     gate269  (.D(g6593), .CP(CLK), .Q(g582) ) ;
INV     gate270  (.A(II8650), .Z(g6594) ) ;
DFF     gate271  (.D(g6594), .CP(CLK), .Q(g586) ) ;
INV     gate272  (.A(II8641), .Z(g6591) ) ;
DFF     gate273  (.D(g6591), .CP(CLK), .Q(g574) ) ;
INV     gate274  (.A(II8653), .Z(g6595) ) ;
DFF     gate275  (.D(g6595), .CP(CLK), .Q(g590) ) ;
INV     gate276  (.A(II8656), .Z(g6596) ) ;
DFF     gate277  (.D(g6596), .CP(CLK), .Q(g594) ) ;
INV     gate278  (.A(II5451), .Z(g4123) ) ;
DFF     gate279  (.D(g4123), .CP(CLK), .Q(g602) ) ;
INV     gate280  (.A(II5454), .Z(g4124) ) ;
DFF     gate281  (.D(g4124), .CP(CLK), .Q(g610) ) ;
INV     gate282  (.A(II5920), .Z(g4423) ) ;
DFF     gate283  (.D(g4423), .CP(CLK), .Q(g613) ) ;
INV     gate284  (.A(II6244), .Z(g4657) ) ;
DFF     gate285  (.D(g4657), .CP(CLK), .Q(g616) ) ;
INV     gate286  (.A(II6582), .Z(g4858) ) ;
DFF     gate287  (.D(g4858), .CP(CLK), .Q(g619) ) ;
INV     gate288  (.A(II6809), .Z(g5147) ) ;
DFF     gate289  (.D(g5147), .CP(CLK), .Q(g622) ) ;
INV     gate290  (.A(II6986), .Z(g5328) ) ;
DFF     gate291  (.D(g5328), .CP(CLK), .Q(g625) ) ;
INV     gate292  (.A(II7187), .Z(g5489) ) ;
DFF     gate293  (.D(g5489), .CP(CLK), .Q(g628) ) ;
INV     gate294  (.A(II7339), .Z(g5581) ) ;
DFF     gate295  (.D(g5581), .CP(CLK), .Q(g631) ) ;
INV     gate296  (.A(II8235), .Z(g6407) ) ;
DFF     gate297  (.D(g6407), .CP(CLK), .Q(g43) ) ;
INV     gate298  (.A(II6250), .Z(g4659) ) ;
DFF     gate299  (.D(g4659), .CP(CLK), .Q(g266) ) ;
INV     gate300  (.A(II5926), .Z(g4425) ) ;
DFF     gate301  (.D(g4425), .CP(CLK), .Q(g658) ) ;
INV     gate302  (.A(II5463), .Z(g4127) ) ;
DFF     gate303  (.D(g4127), .CP(CLK), .Q(g667) ) ;
INV     gate304  (.A(II5466), .Z(g4128) ) ;
DFF     gate305  (.D(g4128), .CP(CLK), .Q(g666) ) ;
INV     gate306  (.A(II2907), .Z(g1831) ) ;
DFF     gate307  (.D(g1831), .CP(CLK), .Q(g662) ) ;
INV     gate308  (.A(II5457), .Z(g4125) ) ;
DFF     gate309  (.D(g4125), .CP(CLK), .Q(g663) ) ;
INV     gate310  (.A(II2269), .Z(g1288) ) ;
DFF     gate311  (.D(g1288), .CP(CLK), .Q(g664) ) ;
INV     gate312  (.A(II2278), .Z(g1291) ) ;
DFF     gate313  (.D(g1291), .CP(CLK), .Q(g471) ) ;
INV     gate314  (.A(II5460), .Z(g4126) ) ;
DFF     gate315  (.D(g4126), .CP(CLK), .Q(g665) ) ;
INV     gate316  (.A(II2281), .Z(g1292) ) ;
DFF     gate317  (.D(g1292), .CP(CLK), .Q(g478) ) ;
INV     gate318  (.A(II2272), .Z(g1289) ) ;
DFF     gate319  (.D(g1289), .CP(CLK), .Q(g638) ) ;
INV     gate320  (.A(II2275), .Z(g1290) ) ;
DFF     gate321  (.D(g1290), .CP(CLK), .Q(g639) ) ;
INV     gate322  (.A(II5929), .Z(g4426) ) ;
DFF     gate323  (.D(g4426), .CP(CLK), .Q(g699) ) ;
INV     gate324  (.A(II2284), .Z(g1293) ) ;
DFF     gate325  (.D(g1293), .CP(CLK), .Q(g702) ) ;
INV     gate326  (.A(II2287), .Z(g1294) ) ;
DFF     gate327  (.D(g1294), .CP(CLK), .Q(g675) ) ;
INV     gate328  (.A(II7342), .Z(g5582) ) ;
DFF     gate329  (.D(g5582), .CP(CLK), .Q(g669) ) ;
INV     gate330  (.A(II6992), .Z(g5330) ) ;
DFF     gate331  (.D(g5330), .CP(CLK), .Q(g676) ) ;
INV     gate332  (.A(II7193), .Z(g5491) ) ;
DFF     gate333  (.D(g5491), .CP(CLK), .Q(g672) ) ;
INV     gate334  (.A(II8659), .Z(g6597) ) ;
DFF     gate335  (.D(g6597), .CP(CLK), .Q(g3) ) ;
INV     gate336  (.A(II8662), .Z(g6598) ) ;
DFF     gate337  (.D(g6598), .CP(CLK), .Q(g7) ) ;
INV     gate338  (.A(II8665), .Z(g6599) ) ;
DFF     gate339  (.D(g6599), .CP(CLK), .Q(g11) ) ;
INV     gate340  (.A(II8674), .Z(g6602) ) ;
DFF     gate341  (.D(g6602), .CP(CLK), .Q(g15) ) ;
INV     gate342  (.A(II8668), .Z(g6600) ) ;
DFF     gate343  (.D(g6600), .CP(CLK), .Q(g19) ) ;
INV     gate344  (.A(II8671), .Z(g6601) ) ;
DFF     gate345  (.D(g6601), .CP(CLK), .Q(g25) ) ;
INV     gate346  (.A(II9082), .Z(g6853) ) ;
DFF     gate347  (.D(g6853), .CP(CLK), .Q(g29) ) ;
INV     gate348  (.A(II9085), .Z(g6854) ) ;
DFF     gate349  (.D(g6854), .CP(CLK), .Q(g33) ) ;
INV     gate350  (.A(II5508), .Z(g4142) ) ;
DFF     gate351  (.D(g4142), .CP(CLK), .Q(g690) ) ;
INV     gate352  (.A(II5511), .Z(g4143) ) ;
DFF     gate353  (.D(g4143), .CP(CLK), .Q(g691) ) ;
INV     gate354  (.A(II5514), .Z(g4144) ) ;
DFF     gate355  (.D(g4144), .CP(CLK), .Q(g692) ) ;
INV     gate356  (.A(II5517), .Z(g4145) ) ;
DFF     gate357  (.D(g4145), .CP(CLK), .Q(g693) ) ;
INV     gate358  (.A(II5520), .Z(g4146) ) ;
DFF     gate359  (.D(g4146), .CP(CLK), .Q(g694) ) ;
INV     gate360  (.A(II5523), .Z(g4147) ) ;
DFF     gate361  (.D(g4147), .CP(CLK), .Q(g695) ) ;
INV     gate362  (.A(II5526), .Z(g4148) ) ;
DFF     gate363  (.D(g4148), .CP(CLK), .Q(g696) ) ;
INV     gate364  (.A(II5529), .Z(g4149) ) ;
DFF     gate365  (.D(g4149), .CP(CLK), .Q(g697) ) ;
INV     gate366  (.A(II5469), .Z(g4129) ) ;
DFF     gate367  (.D(g4129), .CP(CLK), .Q(g677) ) ;
INV     gate368  (.A(II5472), .Z(g4130) ) ;
DFF     gate369  (.D(g4130), .CP(CLK), .Q(g678) ) ;
INV     gate370  (.A(II5475), .Z(g4131) ) ;
DFF     gate371  (.D(g4131), .CP(CLK), .Q(g679) ) ;
INV     gate372  (.A(II5478), .Z(g4132) ) ;
DFF     gate373  (.D(g4132), .CP(CLK), .Q(g680) ) ;
INV     gate374  (.A(II5481), .Z(g4133) ) ;
DFF     gate375  (.D(g4133), .CP(CLK), .Q(g681) ) ;
INV     gate376  (.A(II5484), .Z(g4134) ) ;
DFF     gate377  (.D(g4134), .CP(CLK), .Q(g682) ) ;
INV     gate378  (.A(II5487), .Z(g4135) ) ;
DFF     gate379  (.D(g4135), .CP(CLK), .Q(g683) ) ;
INV     gate380  (.A(II5490), .Z(g4136) ) ;
DFF     gate381  (.D(g4136), .CP(CLK), .Q(g684) ) ;
INV     gate382  (.A(II5493), .Z(g4137) ) ;
DFF     gate383  (.D(g4137), .CP(CLK), .Q(g685) ) ;
INV     gate384  (.A(II5496), .Z(g4138) ) ;
DFF     gate385  (.D(g4138), .CP(CLK), .Q(g686) ) ;
INV     gate386  (.A(II5499), .Z(g4139) ) ;
DFF     gate387  (.D(g4139), .CP(CLK), .Q(g687) ) ;
INV     gate388  (.A(II5502), .Z(g4140) ) ;
DFF     gate389  (.D(g4140), .CP(CLK), .Q(g688) ) ;
INV     gate390  (.A(II5505), .Z(g4141) ) ;
DFF     gate391  (.D(g4141), .CP(CLK), .Q(g689) ) ;
INV     gate392  (.A(II5532), .Z(g4150) ) ;
DFF     gate393  (.D(g4150), .CP(CLK), .Q(g698) ) ;
INV     gate394  (.A(II8966), .Z(g6800) ) ;
DFF     gate395  (.D(g6800), .CP(CLK), .Q(g668) ) ;
INV     gate396  (.A(II8969), .Z(g6801) ) ;
DFF     gate397  (.D(g6801), .CP(CLK), .Q(g485) ) ;
INV     gate398  (.A(II6555), .Z(g4849) ) ;
DFF     gate399  (.D(g4849), .CP(CLK), .Q(g402) ) ;
INV     gate400  (.A(II6558), .Z(g4850) ) ;
DFF     gate401  (.D(g4850), .CP(CLK), .Q(g406) ) ;
INV     gate402  (.A(II6561), .Z(g4851) ) ;
DFF     gate403  (.D(g4851), .CP(CLK), .Q(g410) ) ;
INV     gate404  (.A(II6564), .Z(g4852) ) ;
DFF     gate405  (.D(g4852), .CP(CLK), .Q(g414) ) ;
INV     gate406  (.A(II6567), .Z(g4853) ) ;
DFF     gate407  (.D(g4853), .CP(CLK), .Q(g418) ) ;
INV     gate408  (.A(II6570), .Z(g4854) ) ;
DFF     gate409  (.D(g4854), .CP(CLK), .Q(g422) ) ;
INV     gate410  (.A(II6573), .Z(g4855) ) ;
DFF     gate411  (.D(g4855), .CP(CLK), .Q(g426) ) ;
INV     gate412  (.A(II6576), .Z(g4856) ) ;
DFF     gate413  (.D(g4856), .CP(CLK), .Q(g430) ) ;
INV     gate414  (.A(II6531), .Z(g4841) ) ;
DFF     gate415  (.D(g4841), .CP(CLK), .Q(g461) ) ;
INV     gate416  (.A(II6534), .Z(g4842) ) ;
DFF     gate417  (.D(g4842), .CP(CLK), .Q(g457) ) ;
INV     gate418  (.A(II6537), .Z(g4843) ) ;
DFF     gate419  (.D(g4843), .CP(CLK), .Q(g453) ) ;
INV     gate420  (.A(II6540), .Z(g4844) ) ;
DFF     gate421  (.D(g4844), .CP(CLK), .Q(g449) ) ;
INV     gate422  (.A(II6543), .Z(g4845) ) ;
DFF     gate423  (.D(g4845), .CP(CLK), .Q(g445) ) ;
INV     gate424  (.A(II6546), .Z(g4846) ) ;
DFF     gate425  (.D(g4846), .CP(CLK), .Q(g441) ) ;
INV     gate426  (.A(II6549), .Z(g4847) ) ;
DFF     gate427  (.D(g4847), .CP(CLK), .Q(g437) ) ;
INV     gate428  (.A(II6552), .Z(g4848) ) ;
DFF     gate429  (.D(g4848), .CP(CLK), .Q(g434) ) ;
INV     gate430  (.A(II9005), .Z(g6824) ) ;
DFF     gate431  (.D(g6824), .CP(CLK), .Q(g545) ) ;
INV     gate432  (.A(II9008), .Z(g6825) ) ;
DFF     gate433  (.D(g6825), .CP(CLK), .Q(g548) ) ;
INV     gate434  (.A(II9011), .Z(g6826) ) ;
DFF     gate435  (.D(g6826), .CP(CLK), .Q(g551) ) ;
INV     gate436  (.A(II9014), .Z(g6827) ) ;
DFF     gate437  (.D(g6827), .CP(CLK), .Q(g554) ) ;
INV     gate438  (.A(II8447), .Z(g6509) ) ;
DFF     gate439  (.D(g6509), .CP(CLK), .Q(g197) ) ;
INV     gate440  (.A(II8450), .Z(g6510) ) ;
DFF     gate441  (.D(g6510), .CP(CLK), .Q(g269) ) ;
INV     gate442  (.A(II8453), .Z(g6511) ) ;
DFF     gate443  (.D(g6511), .CP(CLK), .Q(g293) ) ;
INV     gate444  (.A(II8456), .Z(g6512) ) ;
DFF     gate445  (.D(g6512), .CP(CLK), .Q(g297) ) ;
INV     gate446  (.A(II8411), .Z(g6497) ) ;
DFF     gate447  (.D(g6497), .CP(CLK), .Q(g500) ) ;
INV     gate448  (.A(II8414), .Z(g6498) ) ;
DFF     gate449  (.D(g6498), .CP(CLK), .Q(g504) ) ;
INV     gate450  (.A(II8417), .Z(g6499) ) ;
DFF     gate451  (.D(g6499), .CP(CLK), .Q(g508) ) ;
INV     gate452  (.A(II8420), .Z(g6500) ) ;
DFF     gate453  (.D(g6500), .CP(CLK), .Q(g512) ) ;
INV     gate454  (.A(II8423), .Z(g6501) ) ;
DFF     gate455  (.D(g6501), .CP(CLK), .Q(g516) ) ;
INV     gate456  (.A(II8426), .Z(g6502) ) ;
DFF     gate457  (.D(g6502), .CP(CLK), .Q(g520) ) ;
INV     gate458  (.A(II8429), .Z(g6503) ) ;
DFF     gate459  (.D(g6503), .CP(CLK), .Q(g524) ) ;
INV     gate460  (.A(II8432), .Z(g6504) ) ;
DFF     gate461  (.D(g6504), .CP(CLK), .Q(g528) ) ;
INV     gate462  (.A(II8444), .Z(g6508) ) ;
DFF     gate463  (.D(g6508), .CP(CLK), .Q(g532) ) ;
INV     gate464  (.A(II8441), .Z(g6507) ) ;
DFF     gate465  (.D(g6507), .CP(CLK), .Q(g465) ) ;
INV     gate466  (.A(II8438), .Z(g6506) ) ;
DFF     gate467  (.D(g6506), .CP(CLK), .Q(g536) ) ;
INV     gate468  (.A(II8435), .Z(g6505) ) ;
DFF     gate469  (.D(g6505), .CP(CLK), .Q(g541) ) ;
INV     gate470  (.A(II3711), .Z(g2586) ) ;
DFF     gate471  (.D(g2586), .CP(CLK), .Q(g486) ) ;
INV     gate472  (.A(II3714), .Z(g2587) ) ;
DFF     gate473  (.D(g2587), .CP(CLK), .Q(g489) ) ;
INV     gate474  (.A(II8913), .Z(g6745) ) ;
DFF     gate475  (.D(g6745), .CP(CLK), .Q(g496) ) ;
INV     gate476  (.A(II8910), .Z(g6744) ) ;
DFF     gate477  (.D(g6744), .CP(CLK), .Q(g492) ) ;
INV     gate478  (.A(g361), .Z(II1825) ) ;
INV     gate479  (.A(II1825), .Z(g706) ) ;
INV     gate480  (.A(g114), .Z(g709) ) ;
INV     gate481  (.A(g128), .Z(g710) ) ;
INV     gate482  (.A(g131), .Z(g714) ) ;
INV     gate483  (.A(g135), .Z(g715) ) ;
INV     gate484  (.A(g143), .Z(II1832) ) ;
INV     gate485  (.A(II1832), .Z(g716) ) ;
INV     gate486  (.A(g205), .Z(II1835) ) ;
INV     gate487  (.A(II1835), .Z(g719) ) ;
INV     gate488  (.A(g206), .Z(II1838) ) ;
INV     gate489  (.A(II1838), .Z(g729) ) ;
INV     gate490  (.A(g207), .Z(II1841) ) ;
INV     gate491  (.A(II1841), .Z(g736) ) ;
INV     gate492  (.A(g208), .Z(II1844) ) ;
INV     gate493  (.A(II1844), .Z(g743) ) ;
INV     gate494  (.A(g209), .Z(II1847) ) ;
INV     gate495  (.A(II1847), .Z(g749) ) ;
INV     gate496  (.A(g210), .Z(II1850) ) ;
INV     gate497  (.A(II1850), .Z(g754) ) ;
INV     gate498  (.A(g211), .Z(II1853) ) ;
INV     gate499  (.A(II1853), .Z(g760) ) ;
INV     gate500  (.A(g204), .Z(II1856) ) ;
INV     gate501  (.A(II1856), .Z(g766) ) ;
INV     gate502  (.A(g277), .Z(II1859) ) ;
INV     gate503  (.A(II1859), .Z(g774) ) ;
INV     gate504  (.A(g278), .Z(II1862) ) ;
INV     gate505  (.A(II1862), .Z(g784) ) ;
INV     gate506  (.A(g279), .Z(II1865) ) ;
INV     gate507  (.A(II1865), .Z(g791) ) ;
INV     gate508  (.A(g280), .Z(II1868) ) ;
INV     gate509  (.A(II1868), .Z(g798) ) ;
INV     gate510  (.A(g281), .Z(II1871) ) ;
INV     gate511  (.A(II1871), .Z(g804) ) ;
INV     gate512  (.A(g282), .Z(II1874) ) ;
INV     gate513  (.A(II1874), .Z(g809) ) ;
INV     gate514  (.A(g283), .Z(II1877) ) ;
INV     gate515  (.A(II1877), .Z(g815) ) ;
INV     gate516  (.A(g276), .Z(II1880) ) ;
INV     gate517  (.A(II1880), .Z(g821) ) ;
INV     gate518  (.A(g323), .Z(g829) ) ;
INV     gate519  (.A(g338), .Z(g830) ) ;
INV     gate520  (.A(g341), .Z(g834) ) ;
INV     gate521  (.A(g345), .Z(g835) ) ;
INV     gate522  (.A(g349), .Z(g836) ) ;
INV     gate523  (.A(g353), .Z(g837) ) ;
INV     gate524  (.A(g564), .Z(g838) ) ;
INV     gate525  (.A(g567), .Z(g839) ) ;
INV     gate526  (.A(g571), .Z(g842) ) ;
INV     gate527  (.A(g574), .Z(g843) ) ;
INV     gate528  (.A(g578), .Z(g844) ) ;
INV     gate529  (.A(g582), .Z(g845) ) ;
INV     gate530  (.A(g586), .Z(g846) ) ;
INV     gate531  (.A(g590), .Z(g847) ) ;
INV     gate532  (.A(g594), .Z(g848) ) ;
INV     gate533  (.A(g598), .Z(g849) ) ;
INV     gate534  (.A(g602), .Z(g850) ) ;
INV     gate535  (.A(g606), .Z(g851) ) ;
INV     gate536  (.A(g634), .Z(g852) ) ;
INV     gate537  (.A(g642), .Z(g853) ) ;
INV     gate538  (.A(g646), .Z(g854) ) ;
INV     gate539  (.A(g650), .Z(g855) ) ;
INV     gate540  (.A(g654), .Z(g856) ) ;
INV     gate541  (.A(g170), .Z(g857) ) ;
INV     gate542  (.A(g301), .Z(g858) ) ;
INV     gate543  (.A(g179), .Z(g861) ) ;
INV     gate544  (.A(g319), .Z(g862) ) ;
INV     gate545  (.A(g188), .Z(g865) ) ;
INV     gate546  (.A(g314), .Z(g866) ) ;
INV     gate547  (.A(g143), .Z(g872) ) ;
INV     gate548  (.A(g306), .Z(g873) ) ;
INV     gate549  (.A(g639), .Z(g878) ) ;
INV     gate550  (.A(g310), .Z(g889) ) ;
INV     gate551  (.A(g23), .Z(g893) ) ;
INV     gate552  (.A(g48), .Z(II1917) ) ;
INV     gate553  (.A(II1917), .Z(g894) ) ;
INV     gate554  (.A(g139), .Z(g895) ) ;
INV     gate555  (.A(g22), .Z(g896) ) ;
INV     gate556  (.A(g41), .Z(g897) ) ;
INV     gate557  (.A(g47), .Z(g898) ) ;
INV     gate558  (.A(g663), .Z(II1924) ) ;
INV     gate559  (.A(II1924), .Z(g899) ) ;
INV     gate560  (.A(g665), .Z(II1927) ) ;
INV     gate561  (.A(II1927), .Z(g900) ) ;
INV     gate562  (.A(g667), .Z(II1932) ) ;
INV     gate563  (.A(II1932), .Z(g908) ) ;
INV     gate564  (.A(g666), .Z(II1935) ) ;
INV     gate565  (.A(II1935), .Z(g909) ) ;
INV     gate566  (.A(g332), .Z(II1938) ) ;
INV     gate567  (.A(II1938), .Z(g910) ) ;
INV     gate568  (.A(g658), .Z(g913) ) ;
INV     gate569  (.A(g664), .Z(II1942) ) ;
INV     gate570  (.A(II1942), .Z(g917) ) ;
INV     gate571  (.A(g111), .Z(g921) ) ;
INV     gate572  (.A(g699), .Z(II1947) ) ;
INV     gate573  (.A(II1947), .Z(g922) ) ;
INV     gate574  (.A(g332), .Z(g923) ) ;
INV     gate575  (.A(g702), .Z(II1958) ) ;
INV     gate576  (.A(II1958), .Z(g927) ) ;
INV     gate577  (.A(g49), .Z(g929) ) ;
INV     gate578  (.A(g54), .Z(g931) ) ;
INV     gate579  (.A(g337), .Z(g932) ) ;
INV     gate580  (.A(g59), .Z(g938) ) ;
INV     gate581  (.A(g64), .Z(g940) ) ;
INV     gate582  (.A(g69), .Z(g942) ) ;
INV     gate583  (.A(g496), .Z(g943) ) ;
INV     gate584  (.A(g536), .Z(g945) ) ;
INV     gate585  (.A(g361), .Z(g946) ) ;
INV     gate586  (.A(g74), .Z(g947) ) ;
INV     gate587  (.A(g79), .Z(g949) ) ;
INV     gate588  (.A(g84), .Z(g951) ) ;
INV     gate589  (.A(g677), .Z(II2029) ) ;
INV     gate590  (.A(II2029), .Z(g952) ) ;
INV     gate591  (.A(g357), .Z(g964) ) ;
INV     gate592  (.A(g678), .Z(II2033) ) ;
INV     gate593  (.A(II2033), .Z(g965) ) ;
INV     gate594  (.A(g658), .Z(g971) ) ;
INV     gate595  (.A(g679), .Z(II2037) ) ;
INV     gate596  (.A(II2037), .Z(g980) ) ;
INV     gate597  (.A(g638), .Z(g985) ) ;
INV     gate598  (.A(g680), .Z(II2041) ) ;
INV     gate599  (.A(II2041), .Z(g996) ) ;
INV     gate600  (.A(g681), .Z(II2044) ) ;
INV     gate601  (.A(II2044), .Z(g1001) ) ;
INV     gate602  (.A(g682), .Z(II2047) ) ;
INV     gate603  (.A(II2047), .Z(g1006) ) ;
INV     gate604  (.A(g683), .Z(II2050) ) ;
INV     gate605  (.A(II2050), .Z(g1011) ) ;
INV     gate606  (.A(g684), .Z(II2053) ) ;
INV     gate607  (.A(II2053), .Z(g1017) ) ;
INV     gate608  (.A(g685), .Z(II2057) ) ;
INV     gate609  (.A(II2057), .Z(g1030) ) ;
INV     gate610  (.A(g686), .Z(II2067) ) ;
INV     gate611  (.A(II2067), .Z(g1037) ) ;
INV     gate612  (.A(g127), .Z(g1038) ) ;
INV     gate613  (.A(g662), .Z(g1039) ) ;
INV     gate614  (.A(g486), .Z(g1043) ) ;
INV     gate615  (.A(g699), .Z(g1045) ) ;
INV     gate616  (.A(g489), .Z(g1046) ) ;
INV     gate617  (.A(g492), .Z(g1048) ) ;
INV     gate618  (.A(g266), .Z(g1049) ) ;
INV     gate619  (.A(g668), .Z(g1052) ) ;
INV     gate620  (.A(g197), .Z(g1053) ) ;
INV     gate621  (.A(g485), .Z(g1054) ) ;
INV     gate622  (.A(g269), .Z(g1055) ) ;
INV     gate623  (.A(g89), .Z(g1056) ) ;
INV     gate624  (.A(g702), .Z(g1059) ) ;
INV     gate625  (.A(g107), .Z(g1060) ) ;
INV     gate626  (.A(g675), .Z(g1063) ) ;
INV     gate627  (.A(g102), .Z(g1064) ) ;
INV     gate628  (.A(g94), .Z(g1070) ) ;
INV     gate629  (.A(g687), .Z(II2115) ) ;
INV     gate630  (.A(II2115), .Z(g1076) ) ;
INV     gate631  (.A(g98), .Z(g1084) ) ;
INV     gate632  (.A(g688), .Z(II2119) ) ;
INV     gate633  (.A(II2119), .Z(g1088) ) ;
INV     gate634  (.A(g689), .Z(II2122) ) ;
INV     gate635  (.A(II2122), .Z(g1094) ) ;
INV     gate636  (.A(g698), .Z(II2125) ) ;
INV     gate637  (.A(II2125), .Z(g1101) ) ;
INV     gate638  (.A(g18), .Z(II2128) ) ;
INV     gate639  (.A(II2128), .Z(g1106) ) ;
INV     gate640  (.A(g24), .Z(II2131) ) ;
INV     gate641  (.A(II2131), .Z(g1107) ) ;
INV     gate642  (.A(g705), .Z(II2134) ) ;
INV     gate643  (.A(II2134), .Z(g1108) ) ;
INV     gate644  (.A(g1), .Z(II2137) ) ;
INV     gate645  (.A(II2137), .Z(g1109) ) ;
INV     gate646  (.A(g28), .Z(II2140) ) ;
INV     gate647  (.A(II2140), .Z(g1110) ) ;
INV     gate648  (.A(g2), .Z(II2143) ) ;
INV     gate649  (.A(II2143), .Z(g1111) ) ;
INV     gate650  (.A(g336), .Z(g1112) ) ;
INV     gate651  (.A(g6), .Z(II2147) ) ;
INV     gate652  (.A(II2147), .Z(g1113) ) ;
INV     gate653  (.A(g10), .Z(II2150) ) ;
INV     gate654  (.A(II2150), .Z(g1114) ) ;
INV     gate655  (.A(g40), .Z(g1115) ) ;
INV     gate656  (.A(g14), .Z(II2154) ) ;
INV     gate657  (.A(II2154), .Z(g1116) ) ;
INV     gate658  (.A(g32), .Z(g1117) ) ;
INV     gate659  (.A(g36), .Z(g1118) ) ;
INV     gate660  (.A(g465), .Z(II2159) ) ;
INV     gate661  (.A(II2159), .Z(g1119) ) ;
INV     gate662  (.A(g197), .Z(II2162) ) ;
INV     gate663  (.A(II2162), .Z(g1122) ) ;
INV     gate664  (.A(g690), .Z(II2165) ) ;
INV     gate665  (.A(II2165), .Z(g1123) ) ;
INV     gate666  (.A(g269), .Z(II2169) ) ;
INV     gate667  (.A(II2169), .Z(g1142) ) ;
INV     gate668  (.A(g691), .Z(II2172) ) ;
INV     gate669  (.A(II2172), .Z(g1143) ) ;
INV     gate670  (.A(g25), .Z(II2175) ) ;
INV     gate671  (.A(II2175), .Z(g1156) ) ;
INV     gate672  (.A(g293), .Z(II2179) ) ;
INV     gate673  (.A(II2179), .Z(g1160) ) ;
INV     gate674  (.A(g692), .Z(II2182) ) ;
INV     gate675  (.A(II2182), .Z(g1161) ) ;
INV     gate676  (.A(g29), .Z(II2185) ) ;
INV     gate677  (.A(II2185), .Z(g1173) ) ;
INV     gate678  (.A(g37), .Z(g1174) ) ;
INV     gate679  (.A(g42), .Z(g1175) ) ;
INV     gate680  (.A(g297), .Z(II2190) ) ;
INV     gate681  (.A(II2190), .Z(g1176) ) ;
INV     gate682  (.A(g693), .Z(II2193) ) ;
INV     gate683  (.A(II2193), .Z(g1177) ) ;
INV     gate684  (.A(g3), .Z(II2196) ) ;
INV     gate685  (.A(II2196), .Z(g1189) ) ;
INV     gate686  (.A(g33), .Z(II2199) ) ;
INV     gate687  (.A(II2199), .Z(g1190) ) ;
INV     gate688  (.A(g38), .Z(g1191) ) ;
INV     gate689  (.A(g44), .Z(g1192) ) ;
INV     gate690  (.A(g694), .Z(II2204) ) ;
INV     gate691  (.A(II2204), .Z(g1193) ) ;
INV     gate692  (.A(g7), .Z(II2207) ) ;
INV     gate693  (.A(II2207), .Z(g1203) ) ;
INV     gate694  (.A(g39), .Z(g1204) ) ;
INV     gate695  (.A(g45), .Z(g1205) ) ;
INV     gate696  (.A(g123), .Z(II2212) ) ;
INV     gate697  (.A(II2212), .Z(g1206) ) ;
INV     gate698  (.A(g695), .Z(II2215) ) ;
INV     gate699  (.A(II2215), .Z(g1209) ) ;
INV     gate700  (.A(g11), .Z(II2218) ) ;
INV     gate701  (.A(II2218), .Z(g1219) ) ;
INV     gate702  (.A(g43), .Z(II2221) ) ;
INV     gate703  (.A(II2221), .Z(g1220) ) ;
INV     gate704  (.A(g46), .Z(g1221) ) ;
INV     gate705  (.A(g696), .Z(II2225) ) ;
INV     gate706  (.A(II2225), .Z(g1222) ) ;
INV     gate707  (.A(g15), .Z(II2228) ) ;
INV     gate708  (.A(II2228), .Z(g1232) ) ;
INV     gate709  (.A(g465), .Z(II2231) ) ;
INV     gate710  (.A(II2231), .Z(g1233) ) ;
INV     gate711  (.A(g697), .Z(II2234) ) ;
INV     gate712  (.A(II2234), .Z(g1236) ) ;
INV     gate713  (.A(g465), .Z(II2237) ) ;
INV     gate714  (.A(II2237), .Z(g1246) ) ;
INV     gate715  (.A(g19), .Z(II2240) ) ;
INV     gate716  (.A(II2240), .Z(g1249) ) ;
INV     gate717  (.A(g123), .Z(g1250) ) ;
INV     gate718  (.A(g152), .Z(g1254) ) ;
INV     gate719  (.A(g161), .Z(g1255) ) ;
INV     gate720  (.A(g838), .Z(g1256) ) ;
INV     gate721  (.A(g845), .Z(g1257) ) ;
INV     gate722  (.A(g846), .Z(g1263) ) ;
INV     gate723  (.A(g843), .Z(g1267) ) ;
INV     gate724  (.A(g844), .Z(g1270) ) ;
INV     gate725  (.A(g839), .Z(g1273) ) ;
INV     gate726  (.A(g856), .Z(g1274) ) ;
INV     gate727  (.A(g842), .Z(g1275) ) ;
INV     gate728  (.A(g847), .Z(g1276) ) ;
INV     gate729  (.A(g848), .Z(g1279) ) ;
INV     gate730  (.A(g849), .Z(g1282) ) ;
INV     gate731  (.A(g853), .Z(g1283) ) ;
INV     gate732  (.A(g851), .Z(g1284) ) ;
INV     gate733  (.A(g852), .Z(g1285) ) ;
INV     gate734  (.A(g854), .Z(g1286) ) ;
INV     gate735  (.A(g855), .Z(g1287) ) ;
INV     gate736  (.A(g899), .Z(II2269) ) ;
INV     gate737  (.A(g908), .Z(II2272) ) ;
INV     gate738  (.A(g909), .Z(II2275) ) ;
INV     gate739  (.A(g917), .Z(II2278) ) ;
INV     gate740  (.A(g900), .Z(II2281) ) ;
INV     gate741  (.A(g922), .Z(II2284) ) ;
INV     gate742  (.A(g927), .Z(II2287) ) ;
INV     gate743  (.A(g971), .Z(II2290) ) ;
INV     gate744  (.A(II2290), .Z(g1295) ) ;
INV     gate745  (.A(g971), .Z(II2293) ) ;
INV     gate746  (.A(II2293), .Z(g1305) ) ;
INV     gate747  (.A(g893), .Z(II2296) ) ;
INV     gate748  (.A(II2296), .Z(g1315) ) ;
INV     gate749  (.A(g896), .Z(II2306) ) ;
INV     gate750  (.A(II2306), .Z(g1317) ) ;
INV     gate751  (.A(g1236), .Z(II2309) ) ;
INV     gate752  (.A(II2309), .Z(g1318) ) ;
INV     gate753  (.A(g897), .Z(II2312) ) ;
INV     gate754  (.A(II2312), .Z(g1319) ) ;
INV     gate755  (.A(g1222), .Z(II2315) ) ;
INV     gate756  (.A(II2315), .Z(g1320) ) ;
INV     gate757  (.A(g1236), .Z(II2318) ) ;
INV     gate758  (.A(II2318), .Z(g1321) ) ;
INV     gate759  (.A(g898), .Z(II2321) ) ;
INV     gate760  (.A(II2321), .Z(g1322) ) ;
INV     gate761  (.A(g1209), .Z(II2324) ) ;
INV     gate762  (.A(II2324), .Z(g1323) ) ;
INV     gate763  (.A(g1222), .Z(II2327) ) ;
INV     gate764  (.A(II2327), .Z(g1324) ) ;
INV     gate765  (.A(g1122), .Z(II2330) ) ;
INV     gate766  (.A(II2330), .Z(g1325) ) ;
INV     gate767  (.A(g894), .Z(g1326) ) ;
INV     gate768  (.A(g1193), .Z(II2334) ) ;
INV     gate769  (.A(II2334), .Z(g1327) ) ;
INV     gate770  (.A(g1209), .Z(II2337) ) ;
INV     gate771  (.A(II2337), .Z(g1328) ) ;
INV     gate772  (.A(g1142), .Z(II2340) ) ;
INV     gate773  (.A(II2340), .Z(g1329) ) ;
INV     gate774  (.A(g1177), .Z(II2343) ) ;
INV     gate775  (.A(II2343), .Z(g1330) ) ;
INV     gate776  (.A(g1193), .Z(II2346) ) ;
INV     gate777  (.A(II2346), .Z(g1331) ) ;
INV     gate778  (.A(g1160), .Z(II2349) ) ;
INV     gate779  (.A(II2349), .Z(g1332) ) ;
INV     gate780  (.A(g1161), .Z(II2352) ) ;
INV     gate781  (.A(II2352), .Z(g1333) ) ;
INV     gate782  (.A(g1177), .Z(II2355) ) ;
INV     gate783  (.A(II2355), .Z(g1334) ) ;
INV     gate784  (.A(g1176), .Z(II2358) ) ;
INV     gate785  (.A(II2358), .Z(g1335) ) ;
NAND2   gate786  (.A(II2109), .B(II2110), .Z(g1075) ) ;
INV     gate787  (.A(g1075), .Z(II2361) ) ;
INV     gate788  (.A(II2361), .Z(g1336) ) ;
INV     gate789  (.A(g1143), .Z(II2364) ) ;
INV     gate790  (.A(II2364), .Z(g1337) ) ;
INV     gate791  (.A(g1161), .Z(II2367) ) ;
INV     gate792  (.A(II2367), .Z(g1338) ) ;
INV     gate793  (.A(g1123), .Z(II2370) ) ;
INV     gate794  (.A(II2370), .Z(g1339) ) ;
INV     gate795  (.A(g1143), .Z(II2373) ) ;
INV     gate796  (.A(II2373), .Z(g1340) ) ;
INV     gate797  (.A(g729), .Z(II2376) ) ;
INV     gate798  (.A(II2376), .Z(g1341) ) ;
INV     gate799  (.A(g1123), .Z(II2379) ) ;
INV     gate800  (.A(II2379), .Z(g1344) ) ;
INV     gate801  (.A(g719), .Z(II2382) ) ;
INV     gate802  (.A(II2382), .Z(g1345) ) ;
INV     gate803  (.A(g784), .Z(II2385) ) ;
INV     gate804  (.A(II2385), .Z(g1348) ) ;
INV     gate805  (.A(g878), .Z(II2388) ) ;
INV     gate806  (.A(II2388), .Z(g1351) ) ;
INV     gate807  (.A(g774), .Z(II2391) ) ;
INV     gate808  (.A(II2391), .Z(g1352) ) ;
INV     gate809  (.A(g719), .Z(II2394) ) ;
INV     gate810  (.A(II2394), .Z(g1355) ) ;
INV     gate811  (.A(g1119), .Z(g1358) ) ;
INV     gate812  (.A(g729), .Z(II2399) ) ;
INV     gate813  (.A(II2399), .Z(g1363) ) ;
INV     gate814  (.A(g774), .Z(II2402) ) ;
INV     gate815  (.A(II2402), .Z(g1366) ) ;
INV     gate816  (.A(g1112), .Z(II2405) ) ;
INV     gate817  (.A(II2405), .Z(g1369) ) ;
INV     gate818  (.A(g719), .Z(II2408) ) ;
INV     gate819  (.A(II2408), .Z(g1372) ) ;
INV     gate820  (.A(g736), .Z(II2411) ) ;
INV     gate821  (.A(II2411), .Z(g1375) ) ;
INV     gate822  (.A(g784), .Z(II2414) ) ;
INV     gate823  (.A(II2414), .Z(g1378) ) ;
INV     gate824  (.A(g774), .Z(II2417) ) ;
INV     gate825  (.A(II2417), .Z(g1381) ) ;
INV     gate826  (.A(g791), .Z(II2420) ) ;
INV     gate827  (.A(II2420), .Z(g1384) ) ;
INV     gate828  (.A(g719), .Z(II2424) ) ;
INV     gate829  (.A(II2424), .Z(g1391) ) ;
INV     gate830  (.A(g1206), .Z(g1394) ) ;
INV     gate831  (.A(g774), .Z(II2428) ) ;
INV     gate832  (.A(II2428), .Z(g1395) ) ;
INV     gate833  (.A(g1233), .Z(g1410) ) ;
INV     gate834  (.A(g1246), .Z(g1415) ) ;
INV     gate835  (.A(g872), .Z(II2442) ) ;
INV     gate836  (.A(II2442), .Z(g1423) ) ;
INV     gate837  (.A(g971), .Z(II2445) ) ;
INV     gate838  (.A(II2445), .Z(g1426) ) ;
INV     gate839  (.A(g971), .Z(II2449) ) ;
INV     gate840  (.A(II2449), .Z(g1439) ) ;
INV     gate841  (.A(g952), .Z(II2453) ) ;
INV     gate842  (.A(II2453), .Z(g1450) ) ;
NAND2   gate843  (.A(II2245), .B(II2246), .Z(g1253) ) ;
INV     gate844  (.A(g1253), .Z(II2457) ) ;
INV     gate845  (.A(II2457), .Z(g1460) ) ;
INV     gate846  (.A(g952), .Z(II2460) ) ;
INV     gate847  (.A(II2460), .Z(g1461) ) ;
INV     gate848  (.A(g850), .Z(II2464) ) ;
INV     gate849  (.A(II2464), .Z(g1471) ) ;
INV     gate850  (.A(g952), .Z(g1472) ) ;
INV     gate851  (.A(g952), .Z(g1477) ) ;
INV     gate852  (.A(g985), .Z(g1480) ) ;
INV     gate853  (.A(g971), .Z(II2473) ) ;
INV     gate854  (.A(II2473), .Z(g1484) ) ;
INV     gate855  (.A(g971), .Z(II2476) ) ;
INV     gate856  (.A(II2476), .Z(g1491) ) ;
INV     gate857  (.A(g1049), .Z(II2479) ) ;
INV     gate858  (.A(II2479), .Z(g1498) ) ;
INV     gate859  (.A(g709), .Z(g1502) ) ;
INV     gate860  (.A(g878), .Z(g1503) ) ;
INV     gate861  (.A(g766), .Z(II2485) ) ;
INV     gate862  (.A(II2485), .Z(g1504) ) ;
INV     gate863  (.A(g878), .Z(g1513) ) ;
INV     gate864  (.A(g821), .Z(II2491) ) ;
INV     gate865  (.A(II2491), .Z(g1519) ) ;
INV     gate866  (.A(g878), .Z(g1528) ) ;
INV     gate867  (.A(g1076), .Z(g1529) ) ;
INV     gate868  (.A(g878), .Z(g1533) ) ;
INV     gate869  (.A(g1088), .Z(g1535) ) ;
INV     gate870  (.A(g878), .Z(g1539) ) ;
INV     gate871  (.A(g1094), .Z(g1541) ) ;
INV     gate872  (.A(g878), .Z(g1542) ) ;
INV     gate873  (.A(g1006), .Z(g1543) ) ;
INV     gate874  (.A(g1101), .Z(g1546) ) ;
INV     gate875  (.A(g878), .Z(g1549) ) ;
INV     gate876  (.A(g996), .Z(g1550) ) ;
INV     gate877  (.A(g1011), .Z(g1551) ) ;
INV     gate878  (.A(g1030), .Z(g1552) ) ;
INV     gate879  (.A(g1063), .Z(II2521) ) ;
INV     gate880  (.A(II2521), .Z(g1555) ) ;
INV     gate881  (.A(g878), .Z(g1556) ) ;
INV     gate882  (.A(g1017), .Z(g1557) ) ;
INV     gate883  (.A(g965), .Z(g1559) ) ;
INV     gate884  (.A(g1006), .Z(g1563) ) ;
INV     gate885  (.A(g1030), .Z(g1564) ) ;
INV     gate886  (.A(g971), .Z(II2537) ) ;
INV     gate887  (.A(II2537), .Z(g1567) ) ;
INV     gate888  (.A(g1001), .Z(g1577) ) ;
INV     gate889  (.A(g971), .Z(II2552) ) ;
INV     gate890  (.A(II2552), .Z(g1578) ) ;
INV     gate891  (.A(g910), .Z(g1581) ) ;
INV     gate892  (.A(g1001), .Z(g1583) ) ;
INV     gate893  (.A(g743), .Z(g1584) ) ;
INV     gate894  (.A(g1052), .Z(g1586) ) ;
INV     gate895  (.A(g1123), .Z(g1587) ) ;
INV     gate896  (.A(g798), .Z(g1588) ) ;
INV     gate897  (.A(g1054), .Z(g1593) ) ;
INV     gate898  (.A(g1143), .Z(g1594) ) ;
INV     gate899  (.A(g1222), .Z(II2570) ) ;
INV     gate900  (.A(II2570), .Z(g1608) ) ;
INV     gate901  (.A(g1209), .Z(II2578) ) ;
INV     gate902  (.A(II2578), .Z(g1623) ) ;
INV     gate903  (.A(g946), .Z(II2581) ) ;
INV     gate904  (.A(II2581), .Z(g1624) ) ;
INV     gate905  (.A(g839), .Z(II2584) ) ;
INV     gate906  (.A(II2584), .Z(g1627) ) ;
INV     gate907  (.A(g1193), .Z(II2588) ) ;
INV     gate908  (.A(II2588), .Z(g1631) ) ;
INV     gate909  (.A(g760), .Z(g1632) ) ;
INV     gate910  (.A(g1177), .Z(II2593) ) ;
INV     gate911  (.A(II2593), .Z(g1636) ) ;
INV     gate912  (.A(g985), .Z(II2596) ) ;
INV     gate913  (.A(II2596), .Z(g1637) ) ;
INV     gate914  (.A(g754), .Z(g1638) ) ;
INV     gate915  (.A(g815), .Z(g1639) ) ;
INV     gate916  (.A(g1161), .Z(II2601) ) ;
INV     gate917  (.A(II2601), .Z(g1640) ) ;
INV     gate918  (.A(g1222), .Z(II2604) ) ;
INV     gate919  (.A(II2604), .Z(g1641) ) ;
INV     gate920  (.A(g809), .Z(g1642) ) ;
INV     gate921  (.A(g1143), .Z(II2608) ) ;
INV     gate922  (.A(II2608), .Z(g1643) ) ;
INV     gate923  (.A(g1209), .Z(II2611) ) ;
INV     gate924  (.A(II2611), .Z(g1644) ) ;
INV     gate925  (.A(g1123), .Z(II2614) ) ;
INV     gate926  (.A(II2614), .Z(g1645) ) ;
INV     gate927  (.A(g1193), .Z(II2617) ) ;
INV     gate928  (.A(II2617), .Z(g1646) ) ;
INV     gate929  (.A(g1177), .Z(II2620) ) ;
INV     gate930  (.A(II2620), .Z(g1647) ) ;
INV     gate931  (.A(g1161), .Z(II2623) ) ;
INV     gate932  (.A(II2623), .Z(g1648) ) ;
INV     gate933  (.A(g985), .Z(g1649) ) ;
INV     gate934  (.A(g1053), .Z(II2627) ) ;
INV     gate935  (.A(II2627), .Z(g1650) ) ;
INV     gate936  (.A(g1143), .Z(II2630) ) ;
INV     gate937  (.A(II2630), .Z(g1653) ) ;
INV     gate938  (.A(g878), .Z(g1654) ) ;
INV     gate939  (.A(g985), .Z(g1655) ) ;
INV     gate940  (.A(g1055), .Z(II2635) ) ;
INV     gate941  (.A(II2635), .Z(g1656) ) ;
INV     gate942  (.A(g1123), .Z(II2638) ) ;
INV     gate943  (.A(II2638), .Z(g1659) ) ;
INV     gate944  (.A(g985), .Z(g1660) ) ;
INV     gate945  (.A(g1076), .Z(g1661) ) ;
INV     gate946  (.A(g965), .Z(II2643) ) ;
INV     gate947  (.A(II2643), .Z(g1664) ) ;
INV     gate948  (.A(g985), .Z(g1665) ) ;
INV     gate949  (.A(g1088), .Z(g1666) ) ;
INV     gate950  (.A(g980), .Z(II2648) ) ;
INV     gate951  (.A(II2648), .Z(g1670) ) ;
INV     gate952  (.A(g985), .Z(g1671) ) ;
INV     gate953  (.A(g1094), .Z(g1672) ) ;
INV     gate954  (.A(g996), .Z(II2653) ) ;
INV     gate955  (.A(II2653), .Z(g1673) ) ;
INV     gate956  (.A(g985), .Z(g1674) ) ;
INV     gate957  (.A(g1101), .Z(g1675) ) ;
INV     gate958  (.A(g1001), .Z(II2658) ) ;
INV     gate959  (.A(II2658), .Z(g1678) ) ;
INV     gate960  (.A(g985), .Z(g1679) ) ;
INV     gate961  (.A(g1011), .Z(g1680) ) ;
INV     gate962  (.A(g1006), .Z(II2663) ) ;
INV     gate963  (.A(II2663), .Z(g1681) ) ;
INV     gate964  (.A(g829), .Z(g1682) ) ;
INV     gate965  (.A(g1017), .Z(g1683) ) ;
INV     gate966  (.A(g1011), .Z(II2668) ) ;
INV     gate967  (.A(II2668), .Z(g1684) ) ;
INV     gate968  (.A(g1017), .Z(II2671) ) ;
INV     gate969  (.A(II2671), .Z(g1685) ) ;
INV     gate970  (.A(g1030), .Z(II2688) ) ;
INV     gate971  (.A(II2688), .Z(g1688) ) ;
INV     gate972  (.A(g1037), .Z(II2692) ) ;
INV     gate973  (.A(II2692), .Z(g1690) ) ;
INV     gate974  (.A(g1156), .Z(II2696) ) ;
INV     gate975  (.A(II2696), .Z(g1692) ) ;
INV     gate976  (.A(g1106), .Z(g1695) ) ;
INV     gate977  (.A(g1173), .Z(II2700) ) ;
INV     gate978  (.A(II2700), .Z(g1696) ) ;
INV     gate979  (.A(g1189), .Z(II2703) ) ;
INV     gate980  (.A(II2703), .Z(g1699) ) ;
INV     gate981  (.A(g1107), .Z(g1702) ) ;
INV     gate982  (.A(g1190), .Z(II2707) ) ;
INV     gate983  (.A(II2707), .Z(g1703) ) ;
INV     gate984  (.A(g1109), .Z(g1710) ) ;
INV     gate985  (.A(g1203), .Z(II2712) ) ;
INV     gate986  (.A(II2712), .Z(g1711) ) ;
INV     gate987  (.A(g1110), .Z(g1714) ) ;
INV     gate988  (.A(g1115), .Z(II2716) ) ;
INV     gate989  (.A(II2716), .Z(g1715) ) ;
INV     gate990  (.A(g1111), .Z(g1720) ) ;
INV     gate991  (.A(g1219), .Z(II2721) ) ;
INV     gate992  (.A(II2721), .Z(g1721) ) ;
INV     gate993  (.A(g1220), .Z(II2724) ) ;
INV     gate994  (.A(II2724), .Z(g1724) ) ;
INV     gate995  (.A(g1113), .Z(g1725) ) ;
INV     gate996  (.A(g1232), .Z(II2728) ) ;
INV     gate997  (.A(II2728), .Z(g1726) ) ;
INV     gate998  (.A(g1117), .Z(II2731) ) ;
INV     gate999  (.A(II2731), .Z(g1729) ) ;
INV     gate1000  (.A(g1114), .Z(g1730) ) ;
INV     gate1001  (.A(g1118), .Z(II2735) ) ;
INV     gate1002  (.A(II2735), .Z(g1731) ) ;
INV     gate1003  (.A(g1236), .Z(II2738) ) ;
INV     gate1004  (.A(II2738), .Z(g1732) ) ;
INV     gate1005  (.A(g1222), .Z(II2741) ) ;
INV     gate1006  (.A(II2741), .Z(g1733) ) ;
INV     gate1007  (.A(g952), .Z(g1734) ) ;
INV     gate1008  (.A(g1249), .Z(II2745) ) ;
INV     gate1009  (.A(II2745), .Z(g1735) ) ;
INV     gate1010  (.A(g1108), .Z(g1738) ) ;
INV     gate1011  (.A(g1209), .Z(II2749) ) ;
INV     gate1012  (.A(II2749), .Z(g1739) ) ;
INV     gate1013  (.A(g1116), .Z(g1740) ) ;
INV     gate1014  (.A(g1174), .Z(II2753) ) ;
INV     gate1015  (.A(II2753), .Z(g1741) ) ;
INV     gate1016  (.A(g1175), .Z(II2756) ) ;
INV     gate1017  (.A(II2756), .Z(g1742) ) ;
INV     gate1018  (.A(g1193), .Z(II2760) ) ;
INV     gate1019  (.A(II2760), .Z(g1747) ) ;
INV     gate1020  (.A(g1236), .Z(II2763) ) ;
INV     gate1021  (.A(II2763), .Z(g1748) ) ;
INV     gate1022  (.A(g1191), .Z(II2773) ) ;
INV     gate1023  (.A(II2773), .Z(g1754) ) ;
INV     gate1024  (.A(g1192), .Z(II2776) ) ;
INV     gate1025  (.A(II2776), .Z(g1755) ) ;
INV     gate1026  (.A(g1038), .Z(II2779) ) ;
INV     gate1027  (.A(II2779), .Z(g1756) ) ;
INV     gate1028  (.A(g1177), .Z(II2782) ) ;
INV     gate1029  (.A(II2782), .Z(g1759) ) ;
INV     gate1030  (.A(g1222), .Z(II2785) ) ;
INV     gate1031  (.A(II2785), .Z(g1760) ) ;
INV     gate1032  (.A(g1236), .Z(II2788) ) ;
INV     gate1033  (.A(II2788), .Z(g1761) ) ;
INV     gate1034  (.A(g1236), .Z(II2791) ) ;
INV     gate1035  (.A(II2791), .Z(g1762) ) ;
INV     gate1036  (.A(g1204), .Z(II2802) ) ;
INV     gate1037  (.A(II2802), .Z(g1769) ) ;
INV     gate1038  (.A(g1205), .Z(II2805) ) ;
INV     gate1039  (.A(II2805), .Z(g1770) ) ;
INV     gate1040  (.A(g1161), .Z(II2808) ) ;
INV     gate1041  (.A(II2808), .Z(g1771) ) ;
INV     gate1042  (.A(g1209), .Z(II2811) ) ;
INV     gate1043  (.A(II2811), .Z(g1772) ) ;
INV     gate1044  (.A(g1222), .Z(II2814) ) ;
INV     gate1045  (.A(II2814), .Z(g1773) ) ;
INV     gate1046  (.A(g1222), .Z(II2817) ) ;
INV     gate1047  (.A(II2817), .Z(g1774) ) ;
INV     gate1048  (.A(g952), .Z(g1775) ) ;
INV     gate1049  (.A(g1221), .Z(II2821) ) ;
INV     gate1050  (.A(II2821), .Z(g1776) ) ;
INV     gate1051  (.A(g1143), .Z(II2825) ) ;
INV     gate1052  (.A(II2825), .Z(g1781) ) ;
INV     gate1053  (.A(g1193), .Z(II2828) ) ;
INV     gate1054  (.A(II2828), .Z(g1782) ) ;
INV     gate1055  (.A(g1209), .Z(II2831) ) ;
INV     gate1056  (.A(II2831), .Z(g1783) ) ;
INV     gate1057  (.A(g1209), .Z(II2835) ) ;
INV     gate1058  (.A(II2835), .Z(g1787) ) ;
INV     gate1059  (.A(g985), .Z(g1788) ) ;
INV     gate1060  (.A(g1123), .Z(II2839) ) ;
INV     gate1061  (.A(II2839), .Z(g1789) ) ;
INV     gate1062  (.A(g1177), .Z(II2842) ) ;
INV     gate1063  (.A(II2842), .Z(g1790) ) ;
INV     gate1064  (.A(g1193), .Z(II2845) ) ;
INV     gate1065  (.A(II2845), .Z(g1791) ) ;
INV     gate1066  (.A(g1193), .Z(II2848) ) ;
INV     gate1067  (.A(II2848), .Z(g1792) ) ;
INV     gate1068  (.A(g1236), .Z(II2854) ) ;
INV     gate1069  (.A(II2854), .Z(g1805) ) ;
INV     gate1070  (.A(g1161), .Z(II2857) ) ;
INV     gate1071  (.A(II2857), .Z(g1806) ) ;
INV     gate1072  (.A(g1177), .Z(II2860) ) ;
INV     gate1073  (.A(II2860), .Z(g1807) ) ;
INV     gate1074  (.A(g1177), .Z(II2864) ) ;
INV     gate1075  (.A(II2864), .Z(g1811) ) ;
INV     gate1076  (.A(g1143), .Z(II2867) ) ;
INV     gate1077  (.A(II2867), .Z(g1812) ) ;
INV     gate1078  (.A(g1161), .Z(II2870) ) ;
INV     gate1079  (.A(II2870), .Z(g1813) ) ;
INV     gate1080  (.A(g1161), .Z(II2873) ) ;
INV     gate1081  (.A(II2873), .Z(g1814) ) ;
INV     gate1082  (.A(g1123), .Z(II2877) ) ;
INV     gate1083  (.A(II2877), .Z(g1819) ) ;
INV     gate1084  (.A(g1143), .Z(II2880) ) ;
INV     gate1085  (.A(II2880), .Z(g1820) ) ;
INV     gate1086  (.A(g1143), .Z(II2883) ) ;
INV     gate1087  (.A(II2883), .Z(g1821) ) ;
INV     gate1088  (.A(g1123), .Z(II2887) ) ;
INV     gate1089  (.A(II2887), .Z(g1823) ) ;
INV     gate1090  (.A(g1123), .Z(II2890) ) ;
INV     gate1091  (.A(II2890), .Z(g1824) ) ;
INV     gate1092  (.A(g1236), .Z(II2893) ) ;
INV     gate1093  (.A(II2893), .Z(g1825) ) ;
INV     gate1094  (.A(g1256), .Z(II2904) ) ;
INV     gate1095  (.A(II2904), .Z(g1830) ) ;
INV     gate1096  (.A(g1498), .Z(II2907) ) ;
INV     gate1097  (.A(g1645), .Z(II2910) ) ;
INV     gate1098  (.A(II2910), .Z(g1832) ) ;
INV     gate1099  (.A(g1792), .Z(II2913) ) ;
INV     gate1100  (.A(II2913), .Z(g1833) ) ;
INV     gate1101  (.A(g1643), .Z(II2916) ) ;
INV     gate1102  (.A(II2916), .Z(g1834) ) ;
INV     gate1103  (.A(g1787), .Z(II2919) ) ;
INV     gate1104  (.A(II2919), .Z(g1835) ) ;
INV     gate1105  (.A(g1774), .Z(II2922) ) ;
INV     gate1106  (.A(II2922), .Z(g1836) ) ;
INV     gate1107  (.A(g1762), .Z(II2925) ) ;
INV     gate1108  (.A(II2925), .Z(g1837) ) ;
AND4    gate1109  (.A(g729), .B(g719), .C(g766), .D(II2566), .Z(g1595) ) ;
INV     gate1110  (.A(g1595), .Z(g1838) ) ;
INV     gate1111  (.A(g1659), .Z(II2929) ) ;
INV     gate1112  (.A(II2929), .Z(g1841) ) ;
AND4    gate1113  (.A(g784), .B(g774), .C(g821), .D(II2574), .Z(g1612) ) ;
INV     gate1114  (.A(g1612), .Z(g1842) ) ;
INV     gate1115  (.A(g1653), .Z(II2940) ) ;
INV     gate1116  (.A(II2940), .Z(g1846) ) ;
INV     gate1117  (.A(g1715), .Z(II2943) ) ;
INV     gate1118  (.A(II2943), .Z(g1847) ) ;
INV     gate1119  (.A(g1587), .Z(II2946) ) ;
INV     gate1120  (.A(II2946), .Z(g1848) ) ;
INV     gate1121  (.A(g1263), .Z(II2949) ) ;
INV     gate1122  (.A(II2949), .Z(g1849) ) ;
INV     gate1123  (.A(g1594), .Z(II2952) ) ;
INV     gate1124  (.A(II2952), .Z(g1852) ) ;
INV     gate1125  (.A(g1729), .Z(II2955) ) ;
INV     gate1126  (.A(II2955), .Z(g1853) ) ;
INV     gate1127  (.A(g1257), .Z(II2958) ) ;
INV     gate1128  (.A(II2958), .Z(g1854) ) ;
INV     gate1129  (.A(g1731), .Z(II2961) ) ;
INV     gate1130  (.A(II2961), .Z(g1857) ) ;
INV     gate1131  (.A(g1257), .Z(II2964) ) ;
INV     gate1132  (.A(II2964), .Z(g1858) ) ;
INV     gate1133  (.A(g1682), .Z(II2967) ) ;
INV     gate1134  (.A(II2967), .Z(g1861) ) ;
INV     gate1135  (.A(g1504), .Z(II2970) ) ;
INV     gate1136  (.A(II2970), .Z(g1875) ) ;
NAND2   gate1137  (.A(II2682), .B(II2683), .Z(g1687) ) ;
INV     gate1138  (.A(g1687), .Z(II2973) ) ;
INV     gate1139  (.A(II2973), .Z(g1878) ) ;
NOR2    gate1140  (.A(g1039), .B(g658), .Z(g1603) ) ;
INV     gate1141  (.A(g1603), .Z(g1880) ) ;
NAND3   gate1142  (.A(g98), .B(g1064), .C(g1070), .Z(g1797) ) ;
INV     gate1143  (.A(g1797), .Z(g1883) ) ;
INV     gate1144  (.A(g1263), .Z(II2979) ) ;
INV     gate1145  (.A(II2979), .Z(g1884) ) ;
INV     gate1146  (.A(g1426), .Z(II2982) ) ;
INV     gate1147  (.A(II2982), .Z(g1887) ) ;
NAND2   gate1148  (.A(g866), .B(g306), .Z(g1359) ) ;
INV     gate1149  (.A(g1359), .Z(g1890) ) ;
INV     gate1150  (.A(g1504), .Z(II2986) ) ;
INV     gate1151  (.A(II2986), .Z(g1891) ) ;
INV     gate1152  (.A(g1519), .Z(II2989) ) ;
INV     gate1153  (.A(II2989), .Z(g1894) ) ;
INV     gate1154  (.A(g1741), .Z(II2992) ) ;
INV     gate1155  (.A(II2992), .Z(g1897) ) ;
INV     gate1156  (.A(g1742), .Z(II2995) ) ;
INV     gate1157  (.A(II2995), .Z(g1898) ) ;
INV     gate1158  (.A(g1257), .Z(II2998) ) ;
INV     gate1159  (.A(II2998), .Z(g1899) ) ;
INV     gate1160  (.A(g1267), .Z(II3001) ) ;
INV     gate1161  (.A(II3001), .Z(g1902) ) ;
INV     gate1162  (.A(g1426), .Z(II3004) ) ;
INV     gate1163  (.A(II3004), .Z(g1905) ) ;
INV     gate1164  (.A(g1439), .Z(II3007) ) ;
INV     gate1165  (.A(II3007), .Z(g1908) ) ;
INV     gate1166  (.A(g1504), .Z(II3010) ) ;
INV     gate1167  (.A(II3010), .Z(g1911) ) ;
INV     gate1168  (.A(g1519), .Z(II3013) ) ;
INV     gate1169  (.A(II3013), .Z(g1914) ) ;
INV     gate1170  (.A(g1754), .Z(II3016) ) ;
INV     gate1171  (.A(II3016), .Z(g1917) ) ;
INV     gate1172  (.A(g1755), .Z(II3019) ) ;
INV     gate1173  (.A(II3019), .Z(g1918) ) ;
INV     gate1174  (.A(g1426), .Z(II3022) ) ;
INV     gate1175  (.A(II3022), .Z(g1919) ) ;
INV     gate1176  (.A(g1439), .Z(II3025) ) ;
INV     gate1177  (.A(II3025), .Z(g1922) ) ;
INV     gate1178  (.A(g1504), .Z(II3028) ) ;
INV     gate1179  (.A(II3028), .Z(g1925) ) ;
INV     gate1180  (.A(g1504), .Z(II3031) ) ;
INV     gate1181  (.A(II3031), .Z(g1928) ) ;
INV     gate1182  (.A(g1519), .Z(II3034) ) ;
INV     gate1183  (.A(II3034), .Z(g1931) ) ;
INV     gate1184  (.A(g1769), .Z(II3037) ) ;
INV     gate1185  (.A(II3037), .Z(g1934) ) ;
INV     gate1186  (.A(g1770), .Z(II3040) ) ;
INV     gate1187  (.A(II3040), .Z(g1935) ) ;
INV     gate1188  (.A(g1756), .Z(g1936) ) ;
INV     gate1189  (.A(g1257), .Z(II3044) ) ;
INV     gate1190  (.A(II3044), .Z(g1937) ) ;
INV     gate1191  (.A(g1426), .Z(II3047) ) ;
INV     gate1192  (.A(II3047), .Z(g1940) ) ;
INV     gate1193  (.A(g1439), .Z(II3050) ) ;
INV     gate1194  (.A(II3050), .Z(g1943) ) ;
AND2    gate1195  (.A(g301), .B(g866), .Z(g1407) ) ;
INV     gate1196  (.A(g1407), .Z(II3053) ) ;
INV     gate1197  (.A(II3053), .Z(g1946) ) ;
INV     gate1198  (.A(g1519), .Z(II3056) ) ;
INV     gate1199  (.A(II3056), .Z(g1947) ) ;
INV     gate1200  (.A(g1519), .Z(II3059) ) ;
INV     gate1201  (.A(II3059), .Z(g1950) ) ;
INV     gate1202  (.A(g1776), .Z(II3062) ) ;
INV     gate1203  (.A(II3062), .Z(g1953) ) ;
INV     gate1204  (.A(g1426), .Z(II3065) ) ;
INV     gate1205  (.A(II3065), .Z(g1954) ) ;
INV     gate1206  (.A(g1439), .Z(II3068) ) ;
INV     gate1207  (.A(II3068), .Z(g1957) ) ;
INV     gate1208  (.A(g1504), .Z(II3071) ) ;
INV     gate1209  (.A(II3071), .Z(g1960) ) ;
INV     gate1210  (.A(g1426), .Z(II3074) ) ;
INV     gate1211  (.A(II3074), .Z(g1963) ) ;
INV     gate1212  (.A(g1439), .Z(II3077) ) ;
INV     gate1213  (.A(II3077), .Z(g1966) ) ;
INV     gate1214  (.A(g1519), .Z(II3080) ) ;
INV     gate1215  (.A(II3080), .Z(g1969) ) ;
INV     gate1216  (.A(g1426), .Z(II3083) ) ;
INV     gate1217  (.A(II3083), .Z(g1972) ) ;
INV     gate1218  (.A(g1439), .Z(II3086) ) ;
INV     gate1219  (.A(II3086), .Z(g1975) ) ;
NAND3   gate1220  (.A(g862), .B(g314), .C(g301), .Z(g1387) ) ;
INV     gate1221  (.A(g1387), .Z(g1978) ) ;
INV     gate1222  (.A(g1504), .Z(II3090) ) ;
INV     gate1223  (.A(II3090), .Z(g1979) ) ;
INV     gate1224  (.A(g1426), .Z(II3093) ) ;
INV     gate1225  (.A(II3093), .Z(g1982) ) ;
INV     gate1226  (.A(g1439), .Z(II3096) ) ;
INV     gate1227  (.A(II3096), .Z(g1985) ) ;
INV     gate1228  (.A(g1519), .Z(II3099) ) ;
INV     gate1229  (.A(II3099), .Z(g1988) ) ;
INV     gate1230  (.A(g1426), .Z(II3102) ) ;
INV     gate1231  (.A(II3102), .Z(g1991) ) ;
INV     gate1232  (.A(g1439), .Z(II3105) ) ;
INV     gate1233  (.A(II3105), .Z(g1994) ) ;
NAND2   gate1234  (.A(g306), .B(g889), .Z(g1398) ) ;
INV     gate1235  (.A(g1398), .Z(g1997) ) ;
INV     gate1236  (.A(g1504), .Z(II3109) ) ;
INV     gate1237  (.A(II3109), .Z(g1998) ) ;
INV     gate1238  (.A(g1439), .Z(II3112) ) ;
INV     gate1239  (.A(II3112), .Z(g2001) ) ;
INV     gate1240  (.A(g1519), .Z(II3115) ) ;
INV     gate1241  (.A(II3115), .Z(g2004) ) ;
NAND2   gate1242  (.A(g314), .B(g873), .Z(g1411) ) ;
INV     gate1243  (.A(g1411), .Z(g2007) ) ;
INV     gate1244  (.A(g1276), .Z(g2025) ) ;
INV     gate1245  (.A(g1336), .Z(II3134) ) ;
INV     gate1246  (.A(II3134), .Z(g2029) ) ;
INV     gate1247  (.A(g1315), .Z(II3137) ) ;
INV     gate1248  (.A(II3137), .Z(g2030) ) ;
INV     gate1249  (.A(g1317), .Z(II3140) ) ;
INV     gate1250  (.A(II3140), .Z(g2031) ) ;
NAND2   gate1251  (.A(II2767), .B(II2768), .Z(g1749) ) ;
INV     gate1252  (.A(g1749), .Z(g2032) ) ;
INV     gate1253  (.A(g1319), .Z(II3144) ) ;
INV     gate1254  (.A(II3144), .Z(g2035) ) ;
NAND2   gate1255  (.A(II2796), .B(II2797), .Z(g1764) ) ;
INV     gate1256  (.A(g1764), .Z(g2036) ) ;
INV     gate1257  (.A(g1595), .Z(II3148) ) ;
INV     gate1258  (.A(II3148), .Z(g2039) ) ;
INV     gate1259  (.A(g1738), .Z(g2040) ) ;
INV     gate1260  (.A(g1322), .Z(II3152) ) ;
INV     gate1261  (.A(II3152), .Z(g2041) ) ;
INV     gate1262  (.A(g1612), .Z(II3155) ) ;
INV     gate1263  (.A(II3155), .Z(g2042) ) ;
NAND2   gate1264  (.A(II2898), .B(II2899), .Z(g1829) ) ;
INV     gate1265  (.A(g1829), .Z(II3158) ) ;
INV     gate1266  (.A(II3158), .Z(g2043) ) ;
INV     gate1267  (.A(g1270), .Z(II3161) ) ;
INV     gate1268  (.A(II3161), .Z(g2044) ) ;
NAND3   gate1269  (.A(g310), .B(g866), .C(g873), .Z(g1402) ) ;
INV     gate1270  (.A(g1402), .Z(g2059) ) ;
INV     gate1271  (.A(g1369), .Z(g2060) ) ;
INV     gate1272  (.A(g1341), .Z(g2066) ) ;
INV     gate1273  (.A(g1345), .Z(g2078) ) ;
INV     gate1274  (.A(g1348), .Z(g2079) ) ;
INV     gate1275  (.A(g1819), .Z(II3198) ) ;
INV     gate1276  (.A(II3198), .Z(g2086) ) ;
INV     gate1277  (.A(g1352), .Z(g2087) ) ;
INV     gate1278  (.A(g1812), .Z(II3202) ) ;
INV     gate1279  (.A(II3202), .Z(g2088) ) ;
INV     gate1280  (.A(g1823), .Z(II3206) ) ;
INV     gate1281  (.A(II3206), .Z(g2090) ) ;
INV     gate1282  (.A(g1355), .Z(g2091) ) ;
INV     gate1283  (.A(g1806), .Z(II3212) ) ;
INV     gate1284  (.A(II3212), .Z(g2096) ) ;
INV     gate1285  (.A(g1820), .Z(II3215) ) ;
INV     gate1286  (.A(II3215), .Z(g2097) ) ;
INV     gate1287  (.A(g1363), .Z(g2098) ) ;
INV     gate1288  (.A(g1366), .Z(g2099) ) ;
INV     gate1289  (.A(g1790), .Z(II3222) ) ;
INV     gate1290  (.A(II3222), .Z(g2102) ) ;
INV     gate1291  (.A(g1813), .Z(II3225) ) ;
INV     gate1292  (.A(II3225), .Z(g2103) ) ;
INV     gate1293  (.A(g1372), .Z(g2104) ) ;
INV     gate1294  (.A(g1375), .Z(g2105) ) ;
INV     gate1295  (.A(g1378), .Z(g2106) ) ;
INV     gate1296  (.A(g1782), .Z(II3232) ) ;
INV     gate1297  (.A(II3232), .Z(g2108) ) ;
INV     gate1298  (.A(g1807), .Z(II3235) ) ;
INV     gate1299  (.A(II3235), .Z(g2109) ) ;
INV     gate1300  (.A(g1381), .Z(g2110) ) ;
INV     gate1301  (.A(g1384), .Z(g2111) ) ;
INV     gate1302  (.A(g1460), .Z(II3240) ) ;
INV     gate1303  (.A(II3240), .Z(g2112) ) ;
INV     gate1304  (.A(g1772), .Z(II3244) ) ;
INV     gate1305  (.A(II3244), .Z(g2117) ) ;
INV     gate1306  (.A(g1791), .Z(II3247) ) ;
INV     gate1307  (.A(II3247), .Z(g2118) ) ;
INV     gate1308  (.A(g1391), .Z(g2119) ) ;
INV     gate1309  (.A(g1471), .Z(II3251) ) ;
INV     gate1310  (.A(II3251), .Z(g2120) ) ;
INV     gate1311  (.A(g1650), .Z(II3255) ) ;
INV     gate1312  (.A(II3255), .Z(g2125) ) ;
INV     gate1313  (.A(g1760), .Z(II3258) ) ;
INV     gate1314  (.A(II3258), .Z(g2134) ) ;
INV     gate1315  (.A(g1783), .Z(II3261) ) ;
INV     gate1316  (.A(II3261), .Z(g2135) ) ;
INV     gate1317  (.A(g1395), .Z(g2136) ) ;
INV     gate1318  (.A(g1656), .Z(II3268) ) ;
INV     gate1319  (.A(II3268), .Z(g2145) ) ;
INV     gate1320  (.A(g1748), .Z(II3271) ) ;
INV     gate1321  (.A(II3271), .Z(g2154) ) ;
INV     gate1322  (.A(g1773), .Z(II3274) ) ;
INV     gate1323  (.A(II3274), .Z(g2155) ) ;
INV     gate1324  (.A(g1695), .Z(II3278) ) ;
INV     gate1325  (.A(II3278), .Z(g2157) ) ;
INV     gate1326  (.A(g1761), .Z(II3281) ) ;
INV     gate1327  (.A(II3281), .Z(g2158) ) ;
INV     gate1328  (.A(g1702), .Z(II3284) ) ;
INV     gate1329  (.A(II3284), .Z(g2159) ) ;
INV     gate1330  (.A(g1710), .Z(II3288) ) ;
INV     gate1331  (.A(II3288), .Z(g2163) ) ;
INV     gate1332  (.A(g1714), .Z(II3291) ) ;
INV     gate1333  (.A(II3291), .Z(g2164) ) ;
INV     gate1334  (.A(g1720), .Z(II3294) ) ;
INV     gate1335  (.A(II3294), .Z(g2165) ) ;
INV     gate1336  (.A(g1725), .Z(II3298) ) ;
INV     gate1337  (.A(II3298), .Z(g2169) ) ;
INV     gate1338  (.A(g1730), .Z(II3301) ) ;
INV     gate1339  (.A(II3301), .Z(g2170) ) ;
INV     gate1340  (.A(g1740), .Z(II3304) ) ;
INV     gate1341  (.A(II3304), .Z(g2171) ) ;
INV     gate1342  (.A(g1339), .Z(II3307) ) ;
INV     gate1343  (.A(II3307), .Z(g2172) ) ;
INV     gate1344  (.A(g1640), .Z(II3310) ) ;
INV     gate1345  (.A(II3310), .Z(g2173) ) ;
INV     gate1346  (.A(g1337), .Z(II3313) ) ;
INV     gate1347  (.A(II3313), .Z(g2174) ) ;
INV     gate1348  (.A(g1344), .Z(II3316) ) ;
INV     gate1349  (.A(II3316), .Z(g2175) ) ;
INV     gate1350  (.A(g1636), .Z(II3319) ) ;
INV     gate1351  (.A(II3319), .Z(g2176) ) ;
INV     gate1352  (.A(g1333), .Z(II3322) ) ;
INV     gate1353  (.A(II3322), .Z(g2177) ) ;
INV     gate1354  (.A(g1340), .Z(II3325) ) ;
INV     gate1355  (.A(II3325), .Z(g2178) ) ;
INV     gate1356  (.A(g1273), .Z(II3328) ) ;
INV     gate1357  (.A(II3328), .Z(g2179) ) ;
INV     gate1358  (.A(g1631), .Z(II3331) ) ;
INV     gate1359  (.A(II3331), .Z(g2194) ) ;
INV     gate1360  (.A(g1330), .Z(II3334) ) ;
INV     gate1361  (.A(II3334), .Z(g2195) ) ;
INV     gate1362  (.A(g1338), .Z(II3337) ) ;
INV     gate1363  (.A(II3337), .Z(g2196) ) ;
INV     gate1364  (.A(g1282), .Z(II3340) ) ;
INV     gate1365  (.A(II3340), .Z(g2197) ) ;
INV     gate1366  (.A(g1623), .Z(II3343) ) ;
INV     gate1367  (.A(II3343), .Z(g2212) ) ;
INV     gate1368  (.A(g1327), .Z(II3346) ) ;
INV     gate1369  (.A(II3346), .Z(g2213) ) ;
INV     gate1370  (.A(g1334), .Z(II3349) ) ;
INV     gate1371  (.A(II3349), .Z(g2214) ) ;
INV     gate1372  (.A(g1285), .Z(II3352) ) ;
INV     gate1373  (.A(II3352), .Z(g2215) ) ;
INV     gate1374  (.A(g1608), .Z(II3355) ) ;
INV     gate1375  (.A(II3355), .Z(g2230) ) ;
INV     gate1376  (.A(g1323), .Z(II3358) ) ;
INV     gate1377  (.A(II3358), .Z(g2231) ) ;
INV     gate1378  (.A(g1331), .Z(II3361) ) ;
INV     gate1379  (.A(II3361), .Z(g2232) ) ;
INV     gate1380  (.A(g1648), .Z(II3364) ) ;
INV     gate1381  (.A(II3364), .Z(g2233) ) ;
INV     gate1382  (.A(g1283), .Z(II3367) ) ;
INV     gate1383  (.A(II3367), .Z(g2234) ) ;
INV     gate1384  (.A(g1805), .Z(II3370) ) ;
INV     gate1385  (.A(II3370), .Z(g2241) ) ;
INV     gate1386  (.A(g1320), .Z(II3373) ) ;
INV     gate1387  (.A(II3373), .Z(g2242) ) ;
INV     gate1388  (.A(g1328), .Z(II3376) ) ;
INV     gate1389  (.A(II3376), .Z(g2243) ) ;
INV     gate1390  (.A(g1647), .Z(II3379) ) ;
INV     gate1391  (.A(II3379), .Z(g2244) ) ;
INV     gate1392  (.A(g1284), .Z(II3382) ) ;
INV     gate1393  (.A(II3382), .Z(g2245) ) ;
INV     gate1394  (.A(g1318), .Z(II3385) ) ;
INV     gate1395  (.A(II3385), .Z(g2252) ) ;
INV     gate1396  (.A(g1324), .Z(II3388) ) ;
INV     gate1397  (.A(II3388), .Z(g2253) ) ;
INV     gate1398  (.A(g1646), .Z(II3391) ) ;
INV     gate1399  (.A(II3391), .Z(g2254) ) ;
INV     gate1400  (.A(g1286), .Z(II3395) ) ;
INV     gate1401  (.A(II3395), .Z(g2256) ) ;
INV     gate1402  (.A(g1321), .Z(II3405) ) ;
INV     gate1403  (.A(II3405), .Z(g2264) ) ;
INV     gate1404  (.A(g1644), .Z(II3408) ) ;
INV     gate1405  (.A(II3408), .Z(g2265) ) ;
INV     gate1406  (.A(g1287), .Z(II3419) ) ;
INV     gate1407  (.A(II3419), .Z(g2268) ) ;
INV     gate1408  (.A(g1641), .Z(II3422) ) ;
INV     gate1409  (.A(II3422), .Z(g2275) ) ;
INV     gate1410  (.A(g1274), .Z(II3425) ) ;
INV     gate1411  (.A(II3425), .Z(g2276) ) ;
INV     gate1412  (.A(g1825), .Z(II3428) ) ;
INV     gate1413  (.A(II3428), .Z(g2283) ) ;
INV     gate1414  (.A(g1275), .Z(II3431) ) ;
INV     gate1415  (.A(II3431), .Z(g2284) ) ;
INV     gate1416  (.A(g1627), .Z(II3434) ) ;
INV     gate1417  (.A(II3434), .Z(g2291) ) ;
INV     gate1418  (.A(g1567), .Z(g2293) ) ;
INV     gate1419  (.A(g1578), .Z(g2295) ) ;
INV     gate1420  (.A(g1502), .Z(II3441) ) ;
INV     gate1421  (.A(II3441), .Z(g2296) ) ;
NAND2   gate1422  (.A(g1064), .B(g94), .Z(g1743) ) ;
INV     gate1423  (.A(g1743), .Z(g2306) ) ;
INV     gate1424  (.A(g1450), .Z(II3452) ) ;
INV     gate1425  (.A(II3452), .Z(g2308) ) ;
INV     gate1426  (.A(g1450), .Z(II3462) ) ;
INV     gate1427  (.A(II3462), .Z(g2312) ) ;
INV     gate1428  (.A(g1724), .Z(II3465) ) ;
INV     gate1429  (.A(II3465), .Z(g2315) ) ;
AND2    gate1430  (.A(g89), .B(g1064), .Z(g1802) ) ;
INV     gate1431  (.A(g1802), .Z(II3468) ) ;
INV     gate1432  (.A(II3468), .Z(g2316) ) ;
INV     gate1433  (.A(g1450), .Z(II3471) ) ;
INV     gate1434  (.A(II3471), .Z(g2317) ) ;
INV     gate1435  (.A(g1450), .Z(II3474) ) ;
INV     gate1436  (.A(II3474), .Z(g2320) ) ;
INV     gate1437  (.A(g1450), .Z(II3478) ) ;
INV     gate1438  (.A(II3478), .Z(g2324) ) ;
INV     gate1439  (.A(g1461), .Z(II3481) ) ;
INV     gate1440  (.A(II3481), .Z(g2327) ) ;
NAND3   gate1441  (.A(g1060), .B(g102), .C(g89), .Z(g1777) ) ;
INV     gate1442  (.A(g1777), .Z(g2330) ) ;
INV     gate1443  (.A(g1450), .Z(II3485) ) ;
INV     gate1444  (.A(II3485), .Z(g2333) ) ;
INV     gate1445  (.A(g1295), .Z(II3488) ) ;
INV     gate1446  (.A(II3488), .Z(g2336) ) ;
INV     gate1447  (.A(g1461), .Z(II3493) ) ;
INV     gate1448  (.A(II3493), .Z(g2343) ) ;
INV     gate1449  (.A(g1326), .Z(II3496) ) ;
INV     gate1450  (.A(II3496), .Z(g2346) ) ;
INV     gate1451  (.A(g1450), .Z(II3499) ) ;
INV     gate1452  (.A(II3499), .Z(g2347) ) ;
INV     gate1453  (.A(g1295), .Z(II3502) ) ;
INV     gate1454  (.A(II3502), .Z(g2350) ) ;
INV     gate1455  (.A(g1305), .Z(II3505) ) ;
INV     gate1456  (.A(II3505), .Z(g2353) ) ;
INV     gate1457  (.A(g1461), .Z(II3509) ) ;
INV     gate1458  (.A(II3509), .Z(g2357) ) ;
NAND2   gate1459  (.A(g94), .B(g1084), .Z(g1793) ) ;
INV     gate1460  (.A(g1793), .Z(g2360) ) ;
INV     gate1461  (.A(g1450), .Z(II3513) ) ;
INV     gate1462  (.A(II3513), .Z(g2361) ) ;
INV     gate1463  (.A(g1295), .Z(II3516) ) ;
INV     gate1464  (.A(II3516), .Z(g2364) ) ;
INV     gate1465  (.A(g1305), .Z(II3519) ) ;
INV     gate1466  (.A(II3519), .Z(g2367) ) ;
INV     gate1467  (.A(g1664), .Z(II3522) ) ;
INV     gate1468  (.A(II3522), .Z(g2370) ) ;
INV     gate1469  (.A(g1461), .Z(II3525) ) ;
INV     gate1470  (.A(II3525), .Z(g2378) ) ;
NOR2    gate1471  (.A(g1039), .B(g913), .Z(g1422) ) ;
INV     gate1472  (.A(g1422), .Z(II3528) ) ;
INV     gate1473  (.A(II3528), .Z(g2381) ) ;
INV     gate1474  (.A(g1593), .Z(II3531) ) ;
INV     gate1475  (.A(II3531), .Z(g2390) ) ;
INV     gate1476  (.A(g1295), .Z(II3534) ) ;
INV     gate1477  (.A(II3534), .Z(g2391) ) ;
INV     gate1478  (.A(g1305), .Z(II3537) ) ;
INV     gate1479  (.A(II3537), .Z(g2394) ) ;
INV     gate1480  (.A(g1670), .Z(II3540) ) ;
INV     gate1481  (.A(II3540), .Z(g2397) ) ;
INV     gate1482  (.A(g1461), .Z(II3543) ) ;
INV     gate1483  (.A(II3543), .Z(g2405) ) ;
INV     gate1484  (.A(g1586), .Z(II3546) ) ;
INV     gate1485  (.A(II3546), .Z(g2408) ) ;
NAND2   gate1486  (.A(g102), .B(g1070), .Z(g1815) ) ;
INV     gate1487  (.A(g1815), .Z(g2409) ) ;
INV     gate1488  (.A(g1295), .Z(II3550) ) ;
INV     gate1489  (.A(II3550), .Z(g2410) ) ;
INV     gate1490  (.A(g1305), .Z(II3553) ) ;
INV     gate1491  (.A(II3553), .Z(g2413) ) ;
INV     gate1492  (.A(g1484), .Z(II3556) ) ;
INV     gate1493  (.A(II3556), .Z(g2416) ) ;
INV     gate1494  (.A(g1673), .Z(II3560) ) ;
INV     gate1495  (.A(II3560), .Z(g2422) ) ;
INV     gate1496  (.A(g1461), .Z(II3563) ) ;
INV     gate1497  (.A(II3563), .Z(g2430) ) ;
INV     gate1498  (.A(g1789), .Z(II3569) ) ;
INV     gate1499  (.A(II3569), .Z(g2436) ) ;
INV     gate1500  (.A(g1295), .Z(II3572) ) ;
INV     gate1501  (.A(II3572), .Z(g2437) ) ;
INV     gate1502  (.A(g1305), .Z(II3575) ) ;
INV     gate1503  (.A(II3575), .Z(g2440) ) ;
INV     gate1504  (.A(g1484), .Z(II3578) ) ;
INV     gate1505  (.A(II3578), .Z(g2443) ) ;
INV     gate1506  (.A(g1491), .Z(II3581) ) ;
INV     gate1507  (.A(II3581), .Z(g2446) ) ;
INV     gate1508  (.A(g1678), .Z(II3584) ) ;
INV     gate1509  (.A(II3584), .Z(g2449) ) ;
INV     gate1510  (.A(g1461), .Z(II3587) ) ;
INV     gate1511  (.A(II3587), .Z(g2457) ) ;
INV     gate1512  (.A(g1781), .Z(II3590) ) ;
INV     gate1513  (.A(II3590), .Z(g2460) ) ;
INV     gate1514  (.A(g1295), .Z(II3593) ) ;
INV     gate1515  (.A(II3593), .Z(g2461) ) ;
INV     gate1516  (.A(g1305), .Z(II3596) ) ;
INV     gate1517  (.A(II3596), .Z(g2464) ) ;
INV     gate1518  (.A(g1484), .Z(II3599) ) ;
INV     gate1519  (.A(II3599), .Z(g2467) ) ;
INV     gate1520  (.A(g1491), .Z(II3602) ) ;
INV     gate1521  (.A(II3602), .Z(g2470) ) ;
INV     gate1522  (.A(g1681), .Z(II3605) ) ;
INV     gate1523  (.A(II3605), .Z(g2473) ) ;
INV     gate1524  (.A(g1461), .Z(II3608) ) ;
INV     gate1525  (.A(II3608), .Z(g2481) ) ;
INV     gate1526  (.A(g1771), .Z(II3611) ) ;
INV     gate1527  (.A(II3611), .Z(g2484) ) ;
INV     gate1528  (.A(g1295), .Z(II3614) ) ;
INV     gate1529  (.A(II3614), .Z(g2485) ) ;
INV     gate1530  (.A(g1305), .Z(II3617) ) ;
INV     gate1531  (.A(II3617), .Z(g2488) ) ;
INV     gate1532  (.A(g1484), .Z(II3620) ) ;
INV     gate1533  (.A(II3620), .Z(g2491) ) ;
INV     gate1534  (.A(g1491), .Z(II3623) ) ;
INV     gate1535  (.A(II3623), .Z(g2494) ) ;
INV     gate1536  (.A(g1684), .Z(II3626) ) ;
INV     gate1537  (.A(II3626), .Z(g2497) ) ;
INV     gate1538  (.A(g1759), .Z(II3629) ) ;
INV     gate1539  (.A(II3629), .Z(g2505) ) ;
INV     gate1540  (.A(g1295), .Z(II3632) ) ;
INV     gate1541  (.A(II3632), .Z(g2506) ) ;
INV     gate1542  (.A(g1305), .Z(II3635) ) ;
INV     gate1543  (.A(II3635), .Z(g2509) ) ;
INV     gate1544  (.A(g1484), .Z(II3638) ) ;
INV     gate1545  (.A(II3638), .Z(g2512) ) ;
INV     gate1546  (.A(g1491), .Z(II3641) ) ;
INV     gate1547  (.A(II3641), .Z(g2515) ) ;
INV     gate1548  (.A(g1685), .Z(II3644) ) ;
INV     gate1549  (.A(II3644), .Z(g2518) ) ;
INV     gate1550  (.A(g1747), .Z(II3647) ) ;
INV     gate1551  (.A(II3647), .Z(g2524) ) ;
INV     gate1552  (.A(g1650), .Z(II3650) ) ;
INV     gate1553  (.A(II3650), .Z(g2525) ) ;
INV     gate1554  (.A(g1305), .Z(II3653) ) ;
INV     gate1555  (.A(II3653), .Z(g2535) ) ;
INV     gate1556  (.A(g1484), .Z(II3656) ) ;
INV     gate1557  (.A(II3656), .Z(g2538) ) ;
INV     gate1558  (.A(g1491), .Z(II3659) ) ;
INV     gate1559  (.A(II3659), .Z(g2541) ) ;
INV     gate1560  (.A(g1688), .Z(II3662) ) ;
INV     gate1561  (.A(II3662), .Z(g2544) ) ;
INV     gate1562  (.A(g1824), .Z(II3665) ) ;
INV     gate1563  (.A(II3665), .Z(g2550) ) ;
INV     gate1564  (.A(g1739), .Z(II3669) ) ;
INV     gate1565  (.A(II3669), .Z(g2554) ) ;
INV     gate1566  (.A(g1656), .Z(II3672) ) ;
INV     gate1567  (.A(II3672), .Z(g2555) ) ;
INV     gate1568  (.A(g1491), .Z(II3675) ) ;
INV     gate1569  (.A(II3675), .Z(g2565) ) ;
INV     gate1570  (.A(g1690), .Z(II3678) ) ;
INV     gate1571  (.A(II3678), .Z(g2568) ) ;
INV     gate1572  (.A(g1821), .Z(II3681) ) ;
INV     gate1573  (.A(II3681), .Z(g2574) ) ;
INV     gate1574  (.A(g1733), .Z(II3684) ) ;
INV     gate1575  (.A(II3684), .Z(g2575) ) ;
INV     gate1576  (.A(g1814), .Z(II3687) ) ;
INV     gate1577  (.A(II3687), .Z(g2576) ) ;
INV     gate1578  (.A(g1732), .Z(II3691) ) ;
INV     gate1579  (.A(II3691), .Z(g2580) ) ;
INV     gate1580  (.A(g1811), .Z(II3694) ) ;
INV     gate1581  (.A(II3694), .Z(g2581) ) ;
INV     gate1582  (.A(g1830), .Z(g2583) ) ;
INV     gate1583  (.A(g2316), .Z(II3705) ) ;
INV     gate1584  (.A(g1946), .Z(II3708) ) ;
INV     gate1585  (.A(g1848), .Z(II3711) ) ;
INV     gate1586  (.A(g1852), .Z(II3714) ) ;
INV     gate1587  (.A(g2154), .Z(II3717) ) ;
INV     gate1588  (.A(II3717), .Z(g2588) ) ;
INV     gate1589  (.A(g2155), .Z(II3720) ) ;
INV     gate1590  (.A(II3720), .Z(g2591) ) ;
INV     gate1591  (.A(g2158), .Z(II3723) ) ;
INV     gate1592  (.A(II3723), .Z(g2594) ) ;
INV     gate1593  (.A(g2030), .Z(II3726) ) ;
INV     gate1594  (.A(II3726), .Z(g2598) ) ;
INV     gate1595  (.A(g2436), .Z(II3729) ) ;
INV     gate1596  (.A(II3729), .Z(g2599) ) ;
NAND2   gate1597  (.A(II3169), .B(II3170), .Z(g2061) ) ;
INV     gate1598  (.A(g2061), .Z(g2602) ) ;
INV     gate1599  (.A(g2031), .Z(II3733) ) ;
INV     gate1600  (.A(II3733), .Z(g2603) ) ;
INV     gate1601  (.A(g2460), .Z(II3736) ) ;
INV     gate1602  (.A(II3736), .Z(g2604) ) ;
INV     gate1603  (.A(g2035), .Z(II3746) ) ;
INV     gate1604  (.A(II3746), .Z(g2608) ) ;
INV     gate1605  (.A(g2484), .Z(II3749) ) ;
INV     gate1606  (.A(II3749), .Z(g2609) ) ;
INV     gate1607  (.A(g2044), .Z(II3752) ) ;
INV     gate1608  (.A(II3752), .Z(g2612) ) ;
INV     gate1609  (.A(g2125), .Z(II3755) ) ;
INV     gate1610  (.A(II3755), .Z(g2615) ) ;
INV     gate1611  (.A(g2041), .Z(II3758) ) ;
INV     gate1612  (.A(II3758), .Z(g2618) ) ;
INV     gate1613  (.A(g2505), .Z(II3761) ) ;
INV     gate1614  (.A(II3761), .Z(g2619) ) ;
INV     gate1615  (.A(g2044), .Z(II3764) ) ;
INV     gate1616  (.A(II3764), .Z(g2622) ) ;
INV     gate1617  (.A(g2125), .Z(II3767) ) ;
INV     gate1618  (.A(II3767), .Z(g2625) ) ;
INV     gate1619  (.A(g2145), .Z(II3770) ) ;
INV     gate1620  (.A(II3770), .Z(g2628) ) ;
INV     gate1621  (.A(g2524), .Z(II3773) ) ;
INV     gate1622  (.A(II3773), .Z(g2631) ) ;
INV     gate1623  (.A(g2044), .Z(II3776) ) ;
INV     gate1624  (.A(II3776), .Z(g2634) ) ;
INV     gate1625  (.A(g2125), .Z(II3779) ) ;
INV     gate1626  (.A(II3779), .Z(g2637) ) ;
INV     gate1627  (.A(g2145), .Z(II3782) ) ;
INV     gate1628  (.A(II3782), .Z(g2640) ) ;
INV     gate1629  (.A(g2346), .Z(II3785) ) ;
INV     gate1630  (.A(II3785), .Z(g2643) ) ;
INV     gate1631  (.A(g2554), .Z(II3788) ) ;
INV     gate1632  (.A(II3788), .Z(g2644) ) ;
INV     gate1633  (.A(g2044), .Z(II3791) ) ;
INV     gate1634  (.A(II3791), .Z(g2647) ) ;
INV     gate1635  (.A(g2044), .Z(II3794) ) ;
INV     gate1636  (.A(II3794), .Z(g2650) ) ;
INV     gate1637  (.A(g2125), .Z(II3797) ) ;
INV     gate1638  (.A(II3797), .Z(g2653) ) ;
INV     gate1639  (.A(g2145), .Z(II3800) ) ;
INV     gate1640  (.A(II3800), .Z(g2656) ) ;
INV     gate1641  (.A(g2575), .Z(II3804) ) ;
INV     gate1642  (.A(II3804), .Z(g2660) ) ;
INV     gate1643  (.A(g2308), .Z(g2663) ) ;
INV     gate1644  (.A(g2125), .Z(II3808) ) ;
INV     gate1645  (.A(II3808), .Z(g2664) ) ;
INV     gate1646  (.A(g2145), .Z(II3811) ) ;
INV     gate1647  (.A(II3811), .Z(g2667) ) ;
INV     gate1648  (.A(g2580), .Z(II3816) ) ;
INV     gate1649  (.A(II3816), .Z(g2672) ) ;
INV     gate1650  (.A(g2044), .Z(II3819) ) ;
INV     gate1651  (.A(II3819), .Z(g2675) ) ;
INV     gate1652  (.A(g2312), .Z(g2678) ) ;
INV     gate1653  (.A(g2125), .Z(II3823) ) ;
INV     gate1654  (.A(II3823), .Z(g2679) ) ;
INV     gate1655  (.A(g2145), .Z(II3826) ) ;
INV     gate1656  (.A(II3826), .Z(g2682) ) ;
INV     gate1657  (.A(g2179), .Z(II3830) ) ;
INV     gate1658  (.A(II3830), .Z(g2686) ) ;
NAND2   gate1659  (.A(II3412), .B(II3413), .Z(g2266) ) ;
INV     gate1660  (.A(g2266), .Z(II3833) ) ;
INV     gate1661  (.A(II3833), .Z(g2687) ) ;
INV     gate1662  (.A(g1832), .Z(II3836) ) ;
INV     gate1663  (.A(II3836), .Z(g2688) ) ;
INV     gate1664  (.A(g2317), .Z(g2691) ) ;
INV     gate1665  (.A(g2125), .Z(II3840) ) ;
INV     gate1666  (.A(II3840), .Z(g2692) ) ;
INV     gate1667  (.A(g2145), .Z(II3843) ) ;
INV     gate1668  (.A(II3843), .Z(g2695) ) ;
INV     gate1669  (.A(g2550), .Z(II3855) ) ;
INV     gate1670  (.A(II3855), .Z(g2701) ) ;
INV     gate1671  (.A(g2197), .Z(II3858) ) ;
INV     gate1672  (.A(II3858), .Z(g2705) ) ;
INV     gate1673  (.A(g1834), .Z(II3861) ) ;
INV     gate1674  (.A(II3861), .Z(g2706) ) ;
INV     gate1675  (.A(g2044), .Z(II3864) ) ;
INV     gate1676  (.A(II3864), .Z(g2709) ) ;
INV     gate1677  (.A(g2320), .Z(g2712) ) ;
INV     gate1678  (.A(g2125), .Z(II3868) ) ;
INV     gate1679  (.A(II3868), .Z(g2713) ) ;
INV     gate1680  (.A(g2145), .Z(II3871) ) ;
INV     gate1681  (.A(II3871), .Z(g2716) ) ;
INV     gate1682  (.A(g2574), .Z(II3883) ) ;
INV     gate1683  (.A(II3883), .Z(g2722) ) ;
INV     gate1684  (.A(g2215), .Z(II3886) ) ;
INV     gate1685  (.A(II3886), .Z(g2726) ) ;
INV     gate1686  (.A(g2324), .Z(g2727) ) ;
INV     gate1687  (.A(g2145), .Z(II3890) ) ;
INV     gate1688  (.A(II3890), .Z(g2728) ) ;
INV     gate1689  (.A(g2576), .Z(II3902) ) ;
INV     gate1690  (.A(II3902), .Z(g2734) ) ;
INV     gate1691  (.A(g2327), .Z(g2738) ) ;
INV     gate1692  (.A(g2234), .Z(II3906) ) ;
INV     gate1693  (.A(II3906), .Z(g2739) ) ;
INV     gate1694  (.A(g2044), .Z(II3909) ) ;
INV     gate1695  (.A(II3909), .Z(g2740) ) ;
INV     gate1696  (.A(g2333), .Z(g2743) ) ;
INV     gate1697  (.A(g2336), .Z(g2744) ) ;
INV     gate1698  (.A(g2581), .Z(II3923) ) ;
INV     gate1699  (.A(II3923), .Z(g2748) ) ;
INV     gate1700  (.A(g2343), .Z(g2752) ) ;
INV     gate1701  (.A(g2245), .Z(II3927) ) ;
INV     gate1702  (.A(II3927), .Z(g2753) ) ;
INV     gate1703  (.A(g2347), .Z(g2754) ) ;
INV     gate1704  (.A(g2350), .Z(g2755) ) ;
INV     gate1705  (.A(g2353), .Z(g2756) ) ;
INV     gate1706  (.A(g1833), .Z(II3942) ) ;
INV     gate1707  (.A(II3942), .Z(g2760) ) ;
INV     gate1708  (.A(g2357), .Z(g2764) ) ;
INV     gate1709  (.A(g2256), .Z(II3946) ) ;
INV     gate1710  (.A(II3946), .Z(g2765) ) ;
INV     gate1711  (.A(g2361), .Z(g2766) ) ;
INV     gate1712  (.A(g2364), .Z(g2767) ) ;
INV     gate1713  (.A(g2367), .Z(g2768) ) ;
INV     gate1714  (.A(g1835), .Z(II3961) ) ;
INV     gate1715  (.A(II3961), .Z(g2772) ) ;
INV     gate1716  (.A(g2378), .Z(g2776) ) ;
INV     gate1717  (.A(g2268), .Z(II3965) ) ;
INV     gate1718  (.A(II3965), .Z(g2777) ) ;
INV     gate1719  (.A(g2391), .Z(g2778) ) ;
INV     gate1720  (.A(g2394), .Z(g2779) ) ;
INV     gate1721  (.A(g1836), .Z(II3979) ) ;
INV     gate1722  (.A(II3979), .Z(g2783) ) ;
INV     gate1723  (.A(g2405), .Z(g2787) ) ;
INV     gate1724  (.A(g2276), .Z(II3983) ) ;
INV     gate1725  (.A(II3983), .Z(g2788) ) ;
INV     gate1726  (.A(g2410), .Z(g2789) ) ;
INV     gate1727  (.A(g2413), .Z(g2790) ) ;
INV     gate1728  (.A(g2416), .Z(g2792) ) ;
INV     gate1729  (.A(g1837), .Z(II3999) ) ;
INV     gate1730  (.A(II3999), .Z(g2796) ) ;
INV     gate1731  (.A(g2430), .Z(g2800) ) ;
INV     gate1732  (.A(g2284), .Z(II4003) ) ;
INV     gate1733  (.A(II4003), .Z(g2801) ) ;
INV     gate1734  (.A(g2437), .Z(g2802) ) ;
INV     gate1735  (.A(g2440), .Z(g2803) ) ;
INV     gate1736  (.A(g2443), .Z(g2805) ) ;
INV     gate1737  (.A(g2446), .Z(g2806) ) ;
INV     gate1738  (.A(g1841), .Z(II4019) ) ;
INV     gate1739  (.A(II4019), .Z(g2809) ) ;
INV     gate1740  (.A(g2457), .Z(g2813) ) ;
INV     gate1741  (.A(g2315), .Z(II4023) ) ;
INV     gate1742  (.A(II4023), .Z(g2814) ) ;
INV     gate1743  (.A(g2461), .Z(g2817) ) ;
INV     gate1744  (.A(g2464), .Z(g2818) ) ;
INV     gate1745  (.A(g2467), .Z(g2819) ) ;
INV     gate1746  (.A(g2470), .Z(g2820) ) ;
INV     gate1747  (.A(g1846), .Z(II4031) ) ;
INV     gate1748  (.A(II4031), .Z(g2822) ) ;
INV     gate1749  (.A(g2481), .Z(g2826) ) ;
INV     gate1750  (.A(g2485), .Z(g2827) ) ;
INV     gate1751  (.A(g2488), .Z(g2828) ) ;
INV     gate1752  (.A(g2491), .Z(g2829) ) ;
INV     gate1753  (.A(g2494), .Z(g2830) ) ;
INV     gate1754  (.A(g2506), .Z(g2835) ) ;
INV     gate1755  (.A(g2509), .Z(g2836) ) ;
INV     gate1756  (.A(g2512), .Z(g2837) ) ;
INV     gate1757  (.A(g2515), .Z(g2838) ) ;
INV     gate1758  (.A(g2535), .Z(g2839) ) ;
INV     gate1759  (.A(g2538), .Z(g2840) ) ;
INV     gate1760  (.A(g2541), .Z(g2841) ) ;
INV     gate1761  (.A(g2059), .Z(II4050) ) ;
INV     gate1762  (.A(II4050), .Z(g2842) ) ;
INV     gate1763  (.A(g2565), .Z(g2845) ) ;
AND4    gate1764  (.A(g1743), .B(g1797), .C(g1793), .D(g1138), .Z(g2577) ) ;
INV     gate1765  (.A(g2577), .Z(g2849) ) ;
NAND3   gate1766  (.A(g1473), .B(g1470), .C(g1459), .Z(g2010) ) ;
INV     gate1767  (.A(g2010), .Z(g2856) ) ;
INV     gate1768  (.A(g1878), .Z(II4059) ) ;
INV     gate1769  (.A(II4059), .Z(g2857) ) ;
NAND2   gate1770  (.A(II3698), .B(II3699), .Z(g2582) ) ;
INV     gate1771  (.A(g2582), .Z(II4066) ) ;
INV     gate1772  (.A(II4066), .Z(g2862) ) ;
INV     gate1773  (.A(g2296), .Z(g2863) ) ;
INV     gate1774  (.A(g1887), .Z(g2864) ) ;
INV     gate1775  (.A(g2296), .Z(g2865) ) ;
INV     gate1776  (.A(g1905), .Z(g2866) ) ;
INV     gate1777  (.A(g1908), .Z(g2867) ) ;
NOR2    gate1778  (.A(g1418), .B(g1449), .Z(g2433) ) ;
INV     gate1779  (.A(g2433), .Z(g2869) ) ;
INV     gate1780  (.A(g2296), .Z(g2870) ) ;
INV     gate1781  (.A(g1919), .Z(g2871) ) ;
INV     gate1782  (.A(g1922), .Z(g2872) ) ;
INV     gate1783  (.A(g1849), .Z(g2874) ) ;
INV     gate1784  (.A(g1940), .Z(g2875) ) ;
INV     gate1785  (.A(g1943), .Z(g2876) ) ;
NAND3   gate1786  (.A(g1064), .B(g1070), .C(g1620), .Z(g2434) ) ;
INV     gate1787  (.A(g2434), .Z(g2877) ) ;
INV     gate1788  (.A(g1854), .Z(g2882) ) ;
INV     gate1789  (.A(g1954), .Z(g2883) ) ;
INV     gate1790  (.A(g1957), .Z(g2884) ) ;
INV     gate1791  (.A(g1963), .Z(g2885) ) ;
INV     gate1792  (.A(g1966), .Z(g2886) ) ;
INV     gate1793  (.A(g1858), .Z(g2887) ) ;
INV     gate1794  (.A(g1972), .Z(g2888) ) ;
INV     gate1795  (.A(g1975), .Z(g2889) ) ;
INV     gate1796  (.A(g1875), .Z(g2890) ) ;
INV     gate1797  (.A(g1884), .Z(g2891) ) ;
INV     gate1798  (.A(g1982), .Z(g2892) ) ;
INV     gate1799  (.A(g1985), .Z(g2893) ) ;
INV     gate1800  (.A(g1891), .Z(g2894) ) ;
INV     gate1801  (.A(g1894), .Z(g2895) ) ;
INV     gate1802  (.A(g1899), .Z(g2902) ) ;
INV     gate1803  (.A(g1902), .Z(g2903) ) ;
INV     gate1804  (.A(g1991), .Z(g2904) ) ;
INV     gate1805  (.A(g1994), .Z(g2905) ) ;
INV     gate1806  (.A(g1911), .Z(g2906) ) ;
INV     gate1807  (.A(g1914), .Z(g2907) ) ;
INV     gate1808  (.A(g2001), .Z(g2912) ) ;
INV     gate1809  (.A(g1925), .Z(g2913) ) ;
INV     gate1810  (.A(g1928), .Z(g2914) ) ;
INV     gate1811  (.A(g1931), .Z(g2915) ) ;
INV     gate1812  (.A(g1937), .Z(g2919) ) ;
INV     gate1813  (.A(g1947), .Z(g2920) ) ;
INV     gate1814  (.A(g1950), .Z(g2921) ) ;
INV     gate1815  (.A(g1960), .Z(g2922) ) ;
INV     gate1816  (.A(g1969), .Z(g2923) ) ;
INV     gate1817  (.A(g1979), .Z(g2927) ) ;
INV     gate1818  (.A(g1988), .Z(g2931) ) ;
INV     gate1819  (.A(g1998), .Z(g2932) ) ;
INV     gate1820  (.A(g2043), .Z(II4123) ) ;
INV     gate1821  (.A(II4123), .Z(g2933) ) ;
INV     gate1822  (.A(g2004), .Z(g2934) ) ;
AND4    gate1823  (.A(g1359), .B(g1402), .C(g1398), .D(g901), .Z(g2026) ) ;
INV     gate1824  (.A(g2026), .Z(g2936) ) ;
INV     gate1825  (.A(g2040), .Z(II4133) ) ;
INV     gate1826  (.A(II4133), .Z(g2945) ) ;
INV     gate1827  (.A(g2296), .Z(g2946) ) ;
INV     gate1828  (.A(g2381), .Z(g2952) ) ;
INV     gate1829  (.A(g2381), .Z(g2954) ) ;
INV     gate1830  (.A(g1861), .Z(g2956) ) ;
INV     gate1831  (.A(g1861), .Z(g2957) ) ;
INV     gate1832  (.A(g1861), .Z(g2958) ) ;
INV     gate1833  (.A(g1861), .Z(g2959) ) ;
INV     gate1834  (.A(g1861), .Z(g2961) ) ;
NAND3   gate1835  (.A(g866), .B(g873), .C(g1784), .Z(g2008) ) ;
INV     gate1836  (.A(g2008), .Z(g2962) ) ;
INV     gate1837  (.A(g2390), .Z(II4166) ) ;
INV     gate1838  (.A(II4166), .Z(g2967) ) ;
INV     gate1839  (.A(g2179), .Z(g2968) ) ;
INV     gate1840  (.A(g2157), .Z(II4170) ) ;
INV     gate1841  (.A(II4170), .Z(g2973) ) ;
INV     gate1842  (.A(g2408), .Z(II4173) ) ;
INV     gate1843  (.A(II4173), .Z(g2974) ) ;
INV     gate1844  (.A(g2268), .Z(II4176) ) ;
INV     gate1845  (.A(II4176), .Z(g2975) ) ;
INV     gate1846  (.A(g2197), .Z(g2976) ) ;
INV     gate1847  (.A(g2179), .Z(g2981) ) ;
INV     gate1848  (.A(g2010), .Z(g2986) ) ;
INV     gate1849  (.A(g2159), .Z(II4189) ) ;
INV     gate1850  (.A(II4189), .Z(g2996) ) ;
INV     gate1851  (.A(g1847), .Z(II4192) ) ;
INV     gate1852  (.A(II4192), .Z(g2997) ) ;
INV     gate1853  (.A(g2173), .Z(II4195) ) ;
INV     gate1854  (.A(II4195), .Z(g2998) ) ;
INV     gate1855  (.A(g2276), .Z(II4198) ) ;
INV     gate1856  (.A(II4198), .Z(g3001) ) ;
INV     gate1857  (.A(g2215), .Z(g3002) ) ;
INV     gate1858  (.A(g2197), .Z(g3007) ) ;
INV     gate1859  (.A(g2163), .Z(II4217) ) ;
INV     gate1860  (.A(II4217), .Z(g3014) ) ;
INV     gate1861  (.A(g2164), .Z(II4220) ) ;
INV     gate1862  (.A(II4220), .Z(g3015) ) ;
INV     gate1863  (.A(g2176), .Z(II4223) ) ;
INV     gate1864  (.A(II4223), .Z(g3016) ) ;
INV     gate1865  (.A(g2525), .Z(II4226) ) ;
INV     gate1866  (.A(II4226), .Z(g3019) ) ;
INV     gate1867  (.A(g2284), .Z(II4229) ) ;
INV     gate1868  (.A(II4229), .Z(g3022) ) ;
INV     gate1869  (.A(g2215), .Z(g3023) ) ;
INV     gate1870  (.A(g2165), .Z(II4240) ) ;
INV     gate1871  (.A(II4240), .Z(g3029) ) ;
INV     gate1872  (.A(g1853), .Z(II4243) ) ;
INV     gate1873  (.A(II4243), .Z(g3030) ) ;
INV     gate1874  (.A(g2194), .Z(II4246) ) ;
INV     gate1875  (.A(II4246), .Z(g3031) ) ;
INV     gate1876  (.A(g2525), .Z(II4249) ) ;
INV     gate1877  (.A(II4249), .Z(g3034) ) ;
INV     gate1878  (.A(g2555), .Z(II4252) ) ;
INV     gate1879  (.A(II4252), .Z(g3037) ) ;
INV     gate1880  (.A(g2179), .Z(II4255) ) ;
INV     gate1881  (.A(II4255), .Z(g3040) ) ;
INV     gate1882  (.A(g2169), .Z(II4258) ) ;
INV     gate1883  (.A(II4258), .Z(g3041) ) ;
INV     gate1884  (.A(g1857), .Z(II4261) ) ;
INV     gate1885  (.A(II4261), .Z(g3042) ) ;
INV     gate1886  (.A(g2212), .Z(II4264) ) ;
INV     gate1887  (.A(II4264), .Z(g3043) ) ;
INV     gate1888  (.A(g2525), .Z(II4267) ) ;
INV     gate1889  (.A(II4267), .Z(g3046) ) ;
INV     gate1890  (.A(g2555), .Z(II4270) ) ;
INV     gate1891  (.A(II4270), .Z(g3049) ) ;
INV     gate1892  (.A(g2197), .Z(II4273) ) ;
INV     gate1893  (.A(II4273), .Z(g3052) ) ;
INV     gate1894  (.A(g2170), .Z(II4276) ) ;
INV     gate1895  (.A(II4276), .Z(g3053) ) ;
INV     gate1896  (.A(g2230), .Z(II4279) ) ;
INV     gate1897  (.A(II4279), .Z(g3054) ) ;
INV     gate1898  (.A(g2525), .Z(II4282) ) ;
INV     gate1899  (.A(II4282), .Z(g3057) ) ;
INV     gate1900  (.A(g2555), .Z(II4285) ) ;
INV     gate1901  (.A(II4285), .Z(g3060) ) ;
INV     gate1902  (.A(g2215), .Z(II4288) ) ;
INV     gate1903  (.A(II4288), .Z(g3063) ) ;
INV     gate1904  (.A(g2241), .Z(II4291) ) ;
INV     gate1905  (.A(II4291), .Z(g3064) ) ;
INV     gate1906  (.A(g2525), .Z(II4294) ) ;
INV     gate1907  (.A(II4294), .Z(g3067) ) ;
INV     gate1908  (.A(g2555), .Z(II4297) ) ;
INV     gate1909  (.A(II4297), .Z(g3070) ) ;
INV     gate1910  (.A(g2234), .Z(II4300) ) ;
INV     gate1911  (.A(II4300), .Z(g3073) ) ;
INV     gate1912  (.A(g1897), .Z(II4303) ) ;
INV     gate1913  (.A(II4303), .Z(g3074) ) ;
INV     gate1914  (.A(g1898), .Z(II4306) ) ;
INV     gate1915  (.A(II4306), .Z(g3075) ) ;
INV     gate1916  (.A(g2525), .Z(II4309) ) ;
INV     gate1917  (.A(II4309), .Z(g3076) ) ;
INV     gate1918  (.A(g2555), .Z(II4312) ) ;
INV     gate1919  (.A(II4312), .Z(g3079) ) ;
INV     gate1920  (.A(g2245), .Z(II4315) ) ;
INV     gate1921  (.A(II4315), .Z(g3082) ) ;
INV     gate1922  (.A(g2171), .Z(II4318) ) ;
INV     gate1923  (.A(II4318), .Z(g3083) ) ;
INV     gate1924  (.A(g1917), .Z(II4321) ) ;
INV     gate1925  (.A(II4321), .Z(g3084) ) ;
INV     gate1926  (.A(g1918), .Z(II4324) ) ;
INV     gate1927  (.A(II4324), .Z(g3085) ) ;
INV     gate1928  (.A(g2525), .Z(II4327) ) ;
INV     gate1929  (.A(II4327), .Z(g3086) ) ;
INV     gate1930  (.A(g2555), .Z(II4331) ) ;
INV     gate1931  (.A(II4331), .Z(g3090) ) ;
INV     gate1932  (.A(g2256), .Z(II4334) ) ;
INV     gate1933  (.A(II4334), .Z(g3093) ) ;
INV     gate1934  (.A(g1934), .Z(II4337) ) ;
INV     gate1935  (.A(II4337), .Z(g3094) ) ;
INV     gate1936  (.A(g1935), .Z(II4340) ) ;
INV     gate1937  (.A(II4340), .Z(g3095) ) ;
INV     gate1938  (.A(g2525), .Z(II4343) ) ;
INV     gate1939  (.A(II4343), .Z(g3096) ) ;
INV     gate1940  (.A(g2555), .Z(II4347) ) ;
INV     gate1941  (.A(II4347), .Z(g3100) ) ;
INV     gate1942  (.A(g2233), .Z(II4351) ) ;
INV     gate1943  (.A(II4351), .Z(g3104) ) ;
INV     gate1944  (.A(g1953), .Z(II4354) ) ;
INV     gate1945  (.A(II4354), .Z(g3108) ) ;
INV     gate1946  (.A(g2525), .Z(II4358) ) ;
INV     gate1947  (.A(II4358), .Z(g3110) ) ;
INV     gate1948  (.A(g2555), .Z(II4362) ) ;
INV     gate1949  (.A(II4362), .Z(g3114) ) ;
INV     gate1950  (.A(g2244), .Z(II4366) ) ;
INV     gate1951  (.A(II4366), .Z(g3118) ) ;
INV     gate1952  (.A(g2555), .Z(II4371) ) ;
INV     gate1953  (.A(II4371), .Z(g3124) ) ;
INV     gate1954  (.A(g2254), .Z(II4375) ) ;
INV     gate1955  (.A(II4375), .Z(g3128) ) ;
INV     gate1956  (.A(g2265), .Z(II4382) ) ;
INV     gate1957  (.A(II4382), .Z(g3136) ) ;
INV     gate1958  (.A(g2275), .Z(II4391) ) ;
INV     gate1959  (.A(II4391), .Z(g3150) ) ;
INV     gate1960  (.A(g2086), .Z(II4398) ) ;
INV     gate1961  (.A(II4398), .Z(g3158) ) ;
INV     gate1962  (.A(g2283), .Z(II4402) ) ;
INV     gate1963  (.A(II4402), .Z(g3162) ) ;
INV     gate1964  (.A(g2088), .Z(II4410) ) ;
INV     gate1965  (.A(II4410), .Z(g3173) ) ;
INV     gate1966  (.A(g2090), .Z(II4414) ) ;
INV     gate1967  (.A(II4414), .Z(g3177) ) ;
INV     gate1968  (.A(g2096), .Z(II4420) ) ;
INV     gate1969  (.A(II4420), .Z(g3183) ) ;
INV     gate1970  (.A(g2097), .Z(II4424) ) ;
INV     gate1971  (.A(II4424), .Z(g3187) ) ;
INV     gate1972  (.A(g2102), .Z(II4429) ) ;
INV     gate1973  (.A(II4429), .Z(g3192) ) ;
INV     gate1974  (.A(g2103), .Z(II4433) ) ;
INV     gate1975  (.A(II4433), .Z(g3196) ) ;
INV     gate1976  (.A(g1861), .Z(g3199) ) ;
INV     gate1977  (.A(g2108), .Z(II4437) ) ;
INV     gate1978  (.A(II4437), .Z(g3200) ) ;
INV     gate1979  (.A(g2109), .Z(II4441) ) ;
INV     gate1980  (.A(II4441), .Z(g3204) ) ;
INV     gate1981  (.A(g2117), .Z(II4452) ) ;
INV     gate1982  (.A(II4452), .Z(g3209) ) ;
INV     gate1983  (.A(g2118), .Z(II4455) ) ;
INV     gate1984  (.A(II4455), .Z(g3212) ) ;
INV     gate1985  (.A(g2134), .Z(II4459) ) ;
INV     gate1986  (.A(II4459), .Z(g3216) ) ;
INV     gate1987  (.A(g2135), .Z(II4462) ) ;
INV     gate1988  (.A(II4462), .Z(g3219) ) ;
INV     gate1989  (.A(g2945), .Z(II4465) ) ;
INV     gate1990  (.A(g2583), .Z(II4468) ) ;
INV     gate1991  (.A(II4468), .Z(g3223) ) ;
INV     gate1992  (.A(g3040), .Z(II4471) ) ;
INV     gate1993  (.A(g3052), .Z(II4474) ) ;
INV     gate1994  (.A(g3063), .Z(II4477) ) ;
INV     gate1995  (.A(g3073), .Z(II4480) ) ;
INV     gate1996  (.A(g3082), .Z(II4483) ) ;
INV     gate1997  (.A(g3093), .Z(II4486) ) ;
INV     gate1998  (.A(g2975), .Z(II4489) ) ;
INV     gate1999  (.A(g3001), .Z(II4492) ) ;
INV     gate2000  (.A(g3022), .Z(II4495) ) ;
INV     gate2001  (.A(g2686), .Z(II4498) ) ;
INV     gate2002  (.A(g2705), .Z(II4501) ) ;
INV     gate2003  (.A(g2726), .Z(II4504) ) ;
INV     gate2004  (.A(g2739), .Z(II4507) ) ;
INV     gate2005  (.A(g2753), .Z(II4510) ) ;
INV     gate2006  (.A(g2765), .Z(II4513) ) ;
INV     gate2007  (.A(g2777), .Z(II4516) ) ;
INV     gate2008  (.A(g2788), .Z(II4519) ) ;
INV     gate2009  (.A(g2801), .Z(II4522) ) ;
INV     gate2010  (.A(g3083), .Z(g3242) ) ;
INV     gate2011  (.A(g2973), .Z(g3247) ) ;
NAND2   gate2012  (.A(g1815), .B(g2577), .Z(g2858) ) ;
INV     gate2013  (.A(g2858), .Z(II4534) ) ;
INV     gate2014  (.A(II4534), .Z(g3251) ) ;
INV     gate2015  (.A(g2877), .Z(II4537) ) ;
INV     gate2016  (.A(II4537), .Z(g3258) ) ;
INV     gate2017  (.A(g2996), .Z(g3259) ) ;
INV     gate2018  (.A(g3015), .Z(g3263) ) ;
INV     gate2019  (.A(g3030), .Z(g3267) ) ;
INV     gate2020  (.A(g3042), .Z(g3271) ) ;
INV     gate2021  (.A(g3019), .Z(g3284) ) ;
INV     gate2022  (.A(g3034), .Z(g3289) ) ;
INV     gate2023  (.A(g3037), .Z(g3291) ) ;
INV     gate2024  (.A(g3046), .Z(g3297) ) ;
INV     gate2025  (.A(g3049), .Z(g3299) ) ;
INV     gate2026  (.A(g3057), .Z(g3306) ) ;
INV     gate2027  (.A(g3060), .Z(g3308) ) ;
INV     gate2028  (.A(g2962), .Z(II4587) ) ;
INV     gate2029  (.A(II4587), .Z(g3312) ) ;
NAND2   gate2030  (.A(II4160), .B(II4161), .Z(g2966) ) ;
INV     gate2031  (.A(g2966), .Z(II4593) ) ;
INV     gate2032  (.A(II4593), .Z(g3318) ) ;
INV     gate2033  (.A(g3067), .Z(g3320) ) ;
INV     gate2034  (.A(g3070), .Z(g3322) ) ;
INV     gate2035  (.A(g3076), .Z(g3331) ) ;
INV     gate2036  (.A(g3079), .Z(g3332) ) ;
INV     gate2037  (.A(g3086), .Z(g3342) ) ;
INV     gate2038  (.A(g3090), .Z(g3343) ) ;
INV     gate2039  (.A(g2962), .Z(II4623) ) ;
INV     gate2040  (.A(II4623), .Z(g3346) ) ;
INV     gate2041  (.A(g3096), .Z(g3354) ) ;
INV     gate2042  (.A(g3100), .Z(g3355) ) ;
INV     gate2043  (.A(g3110), .Z(g3363) ) ;
INV     gate2044  (.A(g3114), .Z(g3364) ) ;
INV     gate2045  (.A(g2602), .Z(II4646) ) ;
INV     gate2046  (.A(II4646), .Z(g3369) ) ;
INV     gate2047  (.A(g3124), .Z(g3370) ) ;
NAND3   gate2048  (.A(g2007), .B(g862), .C(g1784), .Z(g2831) ) ;
INV     gate2049  (.A(g2831), .Z(g3380) ) ;
AND4    gate2050  (.A(g1263), .B(g1257), .C(g1270), .D(II4040), .Z(g2834) ) ;
INV     gate2051  (.A(g2834), .Z(g3384) ) ;
OR2     gate2052  (.A(g2095), .B(g1573), .Z(g2924) ) ;
INV     gate2053  (.A(g2924), .Z(II4664) ) ;
INV     gate2054  (.A(II4664), .Z(g3387) ) ;
NOR3    gate2055  (.A(g536), .B(g2010), .C(g541), .Z(g2908) ) ;
INV     gate2056  (.A(g2908), .Z(II4667) ) ;
INV     gate2057  (.A(II4667), .Z(g3388) ) ;
OR2     gate2058  (.A(g2100), .B(g1582), .Z(g2928) ) ;
INV     gate2059  (.A(g2928), .Z(II4671) ) ;
INV     gate2060  (.A(II4671), .Z(g3424) ) ;
AND2    gate2061  (.A(g2029), .B(g1503), .Z(g2670) ) ;
INV     gate2062  (.A(g2670), .Z(II4678) ) ;
INV     gate2063  (.A(II4678), .Z(g3440) ) ;
NAND2   gate2064  (.A(g1411), .B(g2026), .Z(g2947) ) ;
INV     gate2065  (.A(g2947), .Z(II4681) ) ;
INV     gate2066  (.A(II4681), .Z(g3441) ) ;
INV     gate2067  (.A(g2687), .Z(II4684) ) ;
INV     gate2068  (.A(II4684), .Z(g3448) ) ;
NAND2   gate2069  (.A(II4445), .B(II4446), .Z(g3207) ) ;
INV     gate2070  (.A(g3207), .Z(II4688) ) ;
INV     gate2071  (.A(II4688), .Z(g3450) ) ;
INV     gate2072  (.A(g2615), .Z(g3451) ) ;
INV     gate2073  (.A(g2625), .Z(g3452) ) ;
INV     gate2074  (.A(g2628), .Z(g3453) ) ;
INV     gate2075  (.A(g2637), .Z(g3455) ) ;
INV     gate2076  (.A(g2640), .Z(g3456) ) ;
INV     gate2077  (.A(g2653), .Z(g3457) ) ;
INV     gate2078  (.A(g2656), .Z(g3458) ) ;
INV     gate2079  (.A(g2664), .Z(g3459) ) ;
INV     gate2080  (.A(g2667), .Z(g3460) ) ;
INV     gate2081  (.A(g2986), .Z(g3461) ) ;
INV     gate2082  (.A(g2679), .Z(g3462) ) ;
INV     gate2083  (.A(g2682), .Z(g3463) ) ;
INV     gate2084  (.A(g2986), .Z(g3465) ) ;
INV     gate2085  (.A(g2877), .Z(II4706) ) ;
INV     gate2086  (.A(II4706), .Z(g3466) ) ;
INV     gate2087  (.A(g2692), .Z(g3477) ) ;
INV     gate2088  (.A(g2695), .Z(g3478) ) ;
INV     gate2089  (.A(g2986), .Z(g3480) ) ;
INV     gate2090  (.A(g2612), .Z(g3481) ) ;
INV     gate2091  (.A(g2713), .Z(g3482) ) ;
INV     gate2092  (.A(g2716), .Z(g3483) ) ;
INV     gate2093  (.A(g2986), .Z(g3485) ) ;
INV     gate2094  (.A(g2869), .Z(g3486) ) ;
INV     gate2095  (.A(g2622), .Z(g3487) ) ;
INV     gate2096  (.A(g2728), .Z(g3488) ) ;
INV     gate2097  (.A(g2608), .Z(g3491) ) ;
INV     gate2098  (.A(g2634), .Z(g3498) ) ;
INV     gate2099  (.A(g2647), .Z(g3500) ) ;
INV     gate2100  (.A(g2650), .Z(g3501) ) ;
INV     gate2101  (.A(g2675), .Z(g3504) ) ;
INV     gate2102  (.A(g2709), .Z(g3510) ) ;
INV     gate2103  (.A(g2740), .Z(g3519) ) ;
INV     gate2104  (.A(g2594), .Z(II4743) ) ;
INV     gate2105  (.A(II4743), .Z(g3527) ) ;
AND2    gate2106  (.A(g2112), .B(g1649), .Z(g2859) ) ;
INV     gate2107  (.A(g2859), .Z(II4752) ) ;
INV     gate2108  (.A(II4752), .Z(g3534) ) ;
AND2    gate2109  (.A(g2120), .B(g1654), .Z(g2861) ) ;
INV     gate2110  (.A(g2861), .Z(II4757) ) ;
INV     gate2111  (.A(II4757), .Z(g3537) ) ;
INV     gate2112  (.A(g2862), .Z(II4762) ) ;
INV     gate2113  (.A(II4762), .Z(g3540) ) ;
INV     gate2114  (.A(g2643), .Z(g3541) ) ;
INV     gate2115  (.A(g3085), .Z(g3545) ) ;
INV     gate2116  (.A(g3095), .Z(g3546) ) ;
INV     gate2117  (.A(g2598), .Z(g3557) ) ;
INV     gate2118  (.A(g2603), .Z(g3559) ) ;
INV     gate2119  (.A(g2618), .Z(g3564) ) ;
INV     gate2120  (.A(g3074), .Z(g3567) ) ;
INV     gate2121  (.A(g3084), .Z(g3571) ) ;
INV     gate2122  (.A(g2962), .Z(II4777) ) ;
INV     gate2123  (.A(II4777), .Z(g3575) ) ;
INV     gate2124  (.A(g3094), .Z(g3589) ) ;
INV     gate2125  (.A(g2997), .Z(g3593) ) ;
INV     gate2126  (.A(g2814), .Z(II4791) ) ;
INV     gate2127  (.A(g2814), .Z(II4794) ) ;
INV     gate2128  (.A(II4794), .Z(g3601) ) ;
INV     gate2129  (.A(g2967), .Z(II4799) ) ;
INV     gate2130  (.A(II4799), .Z(g3604) ) ;
INV     gate2131  (.A(g2877), .Z(II4802) ) ;
INV     gate2132  (.A(II4802), .Z(g3605) ) ;
INV     gate2133  (.A(g2974), .Z(II4809) ) ;
INV     gate2134  (.A(II4809), .Z(g3612) ) ;
INV     gate2135  (.A(g2877), .Z(II4821) ) ;
INV     gate2136  (.A(II4821), .Z(g3622) ) ;
INV     gate2137  (.A(g3108), .Z(g3638) ) ;
INV     gate2138  (.A(g3075), .Z(g3673) ) ;
NAND3   gate2139  (.A(g2409), .B(g1060), .C(g1620), .Z(g3140) ) ;
INV     gate2140  (.A(g3140), .Z(g3677) ) ;
INV     gate2141  (.A(g3014), .Z(g3705) ) ;
INV     gate2142  (.A(g3029), .Z(g3710) ) ;
INV     gate2143  (.A(g3041), .Z(g3714) ) ;
INV     gate2144  (.A(g3053), .Z(g3719) ) ;
INV     gate2145  (.A(g3223), .Z(II4903) ) ;
INV     gate2146  (.A(II4903), .Z(g3723) ) ;
INV     gate2147  (.A(g3369), .Z(II4935) ) ;
INV     gate2148  (.A(II4935), .Z(g3752) ) ;
INV     gate2149  (.A(g3605), .Z(g3761) ) ;
INV     gate2150  (.A(g3673), .Z(II4955) ) ;
INV     gate2151  (.A(II4955), .Z(g3766) ) ;
INV     gate2152  (.A(g3622), .Z(g3769) ) ;
NAND2   gate2153  (.A(II4783), .B(II4784), .Z(g3597) ) ;
INV     gate2154  (.A(g3597), .Z(II4961) ) ;
INV     gate2155  (.A(II4961), .Z(g3770) ) ;
INV     gate2156  (.A(g3673), .Z(II4964) ) ;
INV     gate2157  (.A(II4964), .Z(g3771) ) ;
INV     gate2158  (.A(g3466), .Z(g3772) ) ;
INV     gate2159  (.A(g3466), .Z(g3773) ) ;
INV     gate2160  (.A(g3388), .Z(g3775) ) ;
INV     gate2161  (.A(g3466), .Z(g3776) ) ;
INV     gate2162  (.A(g3388), .Z(g3777) ) ;
INV     gate2163  (.A(g3388), .Z(g3778) ) ;
INV     gate2164  (.A(g3466), .Z(g3779) ) ;
INV     gate2165  (.A(g3575), .Z(II4976) ) ;
INV     gate2166  (.A(II4976), .Z(g3781) ) ;
INV     gate2167  (.A(g3388), .Z(g3782) ) ;
INV     gate2168  (.A(g3546), .Z(II4980) ) ;
INV     gate2169  (.A(II4980), .Z(g3783) ) ;
INV     gate2170  (.A(g3466), .Z(g3785) ) ;
INV     gate2171  (.A(g3388), .Z(g3786) ) ;
INV     gate2172  (.A(g3638), .Z(II4986) ) ;
INV     gate2173  (.A(II4986), .Z(g3787) ) ;
INV     gate2174  (.A(g3466), .Z(g3788) ) ;
INV     gate2175  (.A(g3388), .Z(g3789) ) ;
INV     gate2176  (.A(g3388), .Z(g3790) ) ;
INV     gate2177  (.A(g3388), .Z(g3791) ) ;
INV     gate2178  (.A(g3388), .Z(g3792) ) ;
INV     gate2179  (.A(g3491), .Z(g3793) ) ;
INV     gate2180  (.A(g3388), .Z(g3796) ) ;
INV     gate2181  (.A(g3388), .Z(g3797) ) ;
INV     gate2182  (.A(g3388), .Z(g3798) ) ;
INV     gate2183  (.A(g3388), .Z(g3799) ) ;
INV     gate2184  (.A(g3388), .Z(g3800) ) ;
INV     gate2185  (.A(g3388), .Z(g3801) ) ;
INV     gate2186  (.A(g3388), .Z(g3802) ) ;
INV     gate2187  (.A(g3612), .Z(II5002) ) ;
INV     gate2188  (.A(II5002), .Z(g3803) ) ;
INV     gate2189  (.A(g3604), .Z(II5006) ) ;
INV     gate2190  (.A(II5006), .Z(g3807) ) ;
INV     gate2191  (.A(g3258), .Z(g3813) ) ;
INV     gate2192  (.A(g3318), .Z(II5019) ) ;
INV     gate2193  (.A(II5019), .Z(g3830) ) ;
INV     gate2194  (.A(g3263), .Z(II5023) ) ;
INV     gate2195  (.A(II5023), .Z(g3832) ) ;
INV     gate2196  (.A(g3267), .Z(II5027) ) ;
INV     gate2197  (.A(II5027), .Z(g3834) ) ;
INV     gate2198  (.A(g3242), .Z(II5030) ) ;
INV     gate2199  (.A(II5030), .Z(g3835) ) ;
INV     gate2200  (.A(g3527), .Z(II5033) ) ;
INV     gate2201  (.A(II5033), .Z(g3836) ) ;
INV     gate2202  (.A(g3705), .Z(II5037) ) ;
INV     gate2203  (.A(II5037), .Z(g3838) ) ;
INV     gate2204  (.A(g3271), .Z(II5040) ) ;
INV     gate2205  (.A(II5040), .Z(g3839) ) ;
INV     gate2206  (.A(g3247), .Z(II5043) ) ;
INV     gate2207  (.A(II5043), .Z(g3840) ) ;
NAND2   gate2208  (.A(II4527), .B(II4528), .Z(g3246) ) ;
INV     gate2209  (.A(g3246), .Z(II5050) ) ;
INV     gate2210  (.A(II5050), .Z(g3845) ) ;
INV     gate2211  (.A(g3710), .Z(II5053) ) ;
INV     gate2212  (.A(II5053), .Z(g3846) ) ;
INV     gate2213  (.A(g3567), .Z(II5056) ) ;
INV     gate2214  (.A(II5056), .Z(g3847) ) ;
INV     gate2215  (.A(g3259), .Z(II5059) ) ;
INV     gate2216  (.A(II5059), .Z(g3848) ) ;
INV     gate2217  (.A(g3714), .Z(II5065) ) ;
INV     gate2218  (.A(II5065), .Z(g3852) ) ;
INV     gate2219  (.A(g3571), .Z(II5068) ) ;
INV     gate2220  (.A(II5068), .Z(g3853) ) ;
INV     gate2221  (.A(g3263), .Z(II5071) ) ;
INV     gate2222  (.A(II5071), .Z(g3854) ) ;
INV     gate2223  (.A(g3719), .Z(II5078) ) ;
INV     gate2224  (.A(II5078), .Z(g3859) ) ;
INV     gate2225  (.A(g3589), .Z(II5081) ) ;
INV     gate2226  (.A(II5081), .Z(g3860) ) ;
INV     gate2227  (.A(g3593), .Z(II5084) ) ;
INV     gate2228  (.A(II5084), .Z(g3861) ) ;
INV     gate2229  (.A(g3242), .Z(II5091) ) ;
INV     gate2230  (.A(II5091), .Z(g3866) ) ;
INV     gate2231  (.A(g3705), .Z(II5094) ) ;
INV     gate2232  (.A(II5094), .Z(g3867) ) ;
INV     gate2233  (.A(g3491), .Z(g3868) ) ;
INV     gate2234  (.A(g3312), .Z(g3872) ) ;
INV     gate2235  (.A(g3440), .Z(II5103) ) ;
INV     gate2236  (.A(II5103), .Z(g3874) ) ;
INV     gate2237  (.A(g3247), .Z(II5106) ) ;
INV     gate2238  (.A(II5106), .Z(g3875) ) ;
INV     gate2239  (.A(g3710), .Z(II5109) ) ;
INV     gate2240  (.A(II5109), .Z(g3876) ) ;
INV     gate2241  (.A(g3259), .Z(II5116) ) ;
INV     gate2242  (.A(II5116), .Z(g3881) ) ;
INV     gate2243  (.A(g3714), .Z(II5119) ) ;
INV     gate2244  (.A(II5119), .Z(g3882) ) ;
INV     gate2245  (.A(g3719), .Z(II5124) ) ;
INV     gate2246  (.A(II5124), .Z(g3885) ) ;
INV     gate2247  (.A(g3346), .Z(g3886) ) ;
INV     gate2248  (.A(g3575), .Z(g3889) ) ;
INV     gate2249  (.A(g3575), .Z(g3890) ) ;
INV     gate2250  (.A(g3575), .Z(g3892) ) ;
INV     gate2251  (.A(g3251), .Z(g3897) ) ;
INV     gate2252  (.A(g3575), .Z(g3898) ) ;
INV     gate2253  (.A(g3575), .Z(g3900) ) ;
INV     gate2254  (.A(g3575), .Z(g3901) ) ;
INV     gate2255  (.A(g3575), .Z(g3902) ) ;
INV     gate2256  (.A(g3575), .Z(g3904) ) ;
INV     gate2257  (.A(g3575), .Z(g3906) ) ;
INV     gate2258  (.A(g3450), .Z(II5148) ) ;
INV     gate2259  (.A(II5148), .Z(g3911) ) ;
AND2    gate2260  (.A(g2924), .B(g1749), .Z(g3505) ) ;
INV     gate2261  (.A(g3505), .Z(g3912) ) ;
NAND3   gate2262  (.A(g1815), .B(g1797), .C(g3109), .Z(g3330) ) ;
INV     gate2263  (.A(g3330), .Z(II5153) ) ;
INV     gate2264  (.A(II5153), .Z(g3914) ) ;
AND2    gate2265  (.A(g2928), .B(g1764), .Z(g3512) ) ;
INV     gate2266  (.A(g3512), .Z(g3921) ) ;
AND2    gate2267  (.A(g2933), .B(g1660), .Z(g3454) ) ;
INV     gate2268  (.A(g3454), .Z(II5157) ) ;
INV     gate2269  (.A(II5157), .Z(g3922) ) ;
INV     gate2270  (.A(g3593), .Z(II5169) ) ;
INV     gate2271  (.A(II5169), .Z(g3932) ) ;
INV     gate2272  (.A(g3267), .Z(II5177) ) ;
INV     gate2273  (.A(II5177), .Z(g3940) ) ;
INV     gate2274  (.A(g3271), .Z(II5182) ) ;
INV     gate2275  (.A(II5182), .Z(g3952) ) ;
INV     gate2276  (.A(g3534), .Z(II5204) ) ;
INV     gate2277  (.A(II5204), .Z(g3960) ) ;
INV     gate2278  (.A(g3567), .Z(II5214) ) ;
INV     gate2279  (.A(II5214), .Z(g3962) ) ;
INV     gate2280  (.A(g3673), .Z(II5217) ) ;
INV     gate2281  (.A(II5217), .Z(g3963) ) ;
INV     gate2282  (.A(g3537), .Z(II5223) ) ;
INV     gate2283  (.A(II5223), .Z(g3967) ) ;
INV     gate2284  (.A(g3571), .Z(II5233) ) ;
INV     gate2285  (.A(II5233), .Z(g3969) ) ;
INV     gate2286  (.A(g3545), .Z(II5236) ) ;
INV     gate2287  (.A(II5236), .Z(g3970) ) ;
INV     gate2288  (.A(g3589), .Z(II5249) ) ;
INV     gate2289  (.A(II5249), .Z(g3975) ) ;
INV     gate2290  (.A(g3546), .Z(II5252) ) ;
INV     gate2291  (.A(II5252), .Z(g3976) ) ;
INV     gate2292  (.A(g3638), .Z(II5264) ) ;
INV     gate2293  (.A(II5264), .Z(g3980) ) ;
INV     gate2294  (.A(g3564), .Z(g3984) ) ;
INV     gate2295  (.A(g3441), .Z(g4003) ) ;
INV     gate2296  (.A(g3601), .Z(g4010) ) ;
INV     gate2297  (.A(g3486), .Z(g4011) ) ;
INV     gate2298  (.A(g3557), .Z(II5316) ) ;
INV     gate2299  (.A(II5316), .Z(g4014) ) ;
INV     gate2300  (.A(g3559), .Z(II5320) ) ;
INV     gate2301  (.A(II5320), .Z(g4016) ) ;
INV     gate2302  (.A(g3466), .Z(II5324) ) ;
INV     gate2303  (.A(II5324), .Z(g4020) ) ;
NAND3   gate2304  (.A(g1411), .B(g1402), .C(g2795), .Z(g3502) ) ;
INV     gate2305  (.A(g3502), .Z(II5328) ) ;
INV     gate2306  (.A(II5328), .Z(g4022) ) ;
INV     gate2307  (.A(g3491), .Z(II5333) ) ;
INV     gate2308  (.A(II5333), .Z(g4034) ) ;
INV     gate2309  (.A(g3564), .Z(II5337) ) ;
INV     gate2310  (.A(II5337), .Z(g4036) ) ;
OR2     gate2311  (.A(g2935), .B(g1637), .Z(g3599) ) ;
INV     gate2312  (.A(g3599), .Z(II5343) ) ;
INV     gate2313  (.A(II5343), .Z(g4040) ) ;
INV     gate2314  (.A(g4014), .Z(II5376) ) ;
INV     gate2315  (.A(g3940), .Z(II5379) ) ;
INV     gate2316  (.A(g3952), .Z(II5382) ) ;
INV     gate2317  (.A(g3962), .Z(II5385) ) ;
INV     gate2318  (.A(g3969), .Z(II5388) ) ;
INV     gate2319  (.A(g3975), .Z(II5391) ) ;
INV     gate2320  (.A(g4016), .Z(II5394) ) ;
INV     gate2321  (.A(g3932), .Z(II5397) ) ;
INV     gate2322  (.A(g3963), .Z(II5400) ) ;
INV     gate2323  (.A(g3970), .Z(II5403) ) ;
INV     gate2324  (.A(g3976), .Z(II5406) ) ;
INV     gate2325  (.A(g3980), .Z(II5409) ) ;
INV     gate2326  (.A(g4034), .Z(II5412) ) ;
INV     gate2327  (.A(g3723), .Z(II5415) ) ;
INV     gate2328  (.A(II5415), .Z(g4111) ) ;
INV     gate2329  (.A(g4036), .Z(II5418) ) ;
AND2    gate2330  (.A(g117), .B(g3251), .Z(g3724) ) ;
INV     gate2331  (.A(g3724), .Z(II5421) ) ;
AND2    gate2332  (.A(g118), .B(g3251), .Z(g3725) ) ;
INV     gate2333  (.A(g3725), .Z(II5424) ) ;
AND2    gate2334  (.A(g119), .B(g3251), .Z(g3726) ) ;
INV     gate2335  (.A(g3726), .Z(II5427) ) ;
AND2    gate2336  (.A(g122), .B(g3251), .Z(g3727) ) ;
INV     gate2337  (.A(g3727), .Z(II5430) ) ;
AND2    gate2338  (.A(g326), .B(g3441), .Z(g3728) ) ;
INV     gate2339  (.A(g3728), .Z(II5433) ) ;
AND2    gate2340  (.A(g327), .B(g3441), .Z(g3729) ) ;
INV     gate2341  (.A(g3729), .Z(II5436) ) ;
AND2    gate2342  (.A(g328), .B(g3441), .Z(g3730) ) ;
INV     gate2343  (.A(g3730), .Z(II5439) ) ;
AND2    gate2344  (.A(g331), .B(g3441), .Z(g3731) ) ;
INV     gate2345  (.A(g3731), .Z(II5442) ) ;
INV     gate2346  (.A(g4040), .Z(II5445) ) ;
INV     gate2347  (.A(g3960), .Z(II5448) ) ;
INV     gate2348  (.A(g3967), .Z(II5451) ) ;
INV     gate2349  (.A(g3874), .Z(II5454) ) ;
INV     gate2350  (.A(g3766), .Z(II5457) ) ;
INV     gate2351  (.A(g3771), .Z(II5460) ) ;
INV     gate2352  (.A(g3783), .Z(II5463) ) ;
INV     gate2353  (.A(g3787), .Z(II5466) ) ;
INV     gate2354  (.A(g3838), .Z(II5469) ) ;
INV     gate2355  (.A(g3846), .Z(II5472) ) ;
INV     gate2356  (.A(g3852), .Z(II5475) ) ;
INV     gate2357  (.A(g3859), .Z(II5478) ) ;
INV     gate2358  (.A(g3866), .Z(II5481) ) ;
INV     gate2359  (.A(g3875), .Z(II5484) ) ;
INV     gate2360  (.A(g3881), .Z(II5487) ) ;
INV     gate2361  (.A(g3832), .Z(II5490) ) ;
INV     gate2362  (.A(g3834), .Z(II5493) ) ;
INV     gate2363  (.A(g3839), .Z(II5496) ) ;
INV     gate2364  (.A(g3847), .Z(II5499) ) ;
INV     gate2365  (.A(g3853), .Z(II5502) ) ;
INV     gate2366  (.A(g3860), .Z(II5505) ) ;
INV     gate2367  (.A(g3867), .Z(II5508) ) ;
INV     gate2368  (.A(g3876), .Z(II5511) ) ;
INV     gate2369  (.A(g3882), .Z(II5514) ) ;
INV     gate2370  (.A(g3885), .Z(II5517) ) ;
INV     gate2371  (.A(g3835), .Z(II5520) ) ;
INV     gate2372  (.A(g3840), .Z(II5523) ) ;
INV     gate2373  (.A(g3848), .Z(II5526) ) ;
INV     gate2374  (.A(g3854), .Z(II5529) ) ;
INV     gate2375  (.A(g3861), .Z(II5532) ) ;
INV     gate2376  (.A(g3984), .Z(II5542) ) ;
INV     gate2377  (.A(II5542), .Z(g4152) ) ;
AND2    gate2378  (.A(g913), .B(g3546), .Z(g3814) ) ;
INV     gate2379  (.A(g3814), .Z(II5545) ) ;
INV     gate2380  (.A(II5545), .Z(g4153) ) ;
OR2     gate2381  (.A(g3466), .B(g3425), .Z(g4059) ) ;
INV     gate2382  (.A(g4059), .Z(II5548) ) ;
INV     gate2383  (.A(II5548), .Z(g4154) ) ;
INV     gate2384  (.A(g4059), .Z(II5551) ) ;
INV     gate2385  (.A(II5551), .Z(g4155) ) ;
INV     gate2386  (.A(g4059), .Z(II5556) ) ;
INV     gate2387  (.A(II5556), .Z(g4158) ) ;
NAND2   gate2388  (.A(II5293), .B(II5294), .Z(g4002) ) ;
INV     gate2389  (.A(g4002), .Z(II5562) ) ;
INV     gate2390  (.A(II5562), .Z(g4162) ) ;
INV     gate2391  (.A(g3897), .Z(II5568) ) ;
INV     gate2392  (.A(II5568), .Z(g4166) ) ;
INV     gate2393  (.A(g4022), .Z(II5577) ) ;
INV     gate2394  (.A(II5577), .Z(g4173) ) ;
OR2     gate2395  (.A(g2951), .B(g3466), .Z(g3821) ) ;
INV     gate2396  (.A(g3821), .Z(II5591) ) ;
INV     gate2397  (.A(II5591), .Z(g4187) ) ;
INV     gate2398  (.A(g3821), .Z(II5594) ) ;
INV     gate2399  (.A(II5594), .Z(g4188) ) ;
INV     gate2400  (.A(g3821), .Z(II5597) ) ;
INV     gate2401  (.A(II5597), .Z(g4189) ) ;
INV     gate2402  (.A(g3821), .Z(II5600) ) ;
INV     gate2403  (.A(II5600), .Z(g4190) ) ;
NAND3   gate2404  (.A(g3664), .B(g3656), .C(g3647), .Z(g3893) ) ;
INV     gate2405  (.A(g3893), .Z(II5603) ) ;
INV     gate2406  (.A(II5603), .Z(g4191) ) ;
INV     gate2407  (.A(g3821), .Z(II5606) ) ;
INV     gate2408  (.A(II5606), .Z(g4192) ) ;
INV     gate2409  (.A(g3893), .Z(II5609) ) ;
INV     gate2410  (.A(II5609), .Z(g4193) ) ;
AND2    gate2411  (.A(g3546), .B(g1049), .Z(g3910) ) ;
INV     gate2412  (.A(g3910), .Z(II5612) ) ;
INV     gate2413  (.A(II5612), .Z(g4194) ) ;
INV     gate2414  (.A(g3914), .Z(II5615) ) ;
INV     gate2415  (.A(II5615), .Z(g4195) ) ;
INV     gate2416  (.A(g3821), .Z(II5618) ) ;
INV     gate2417  (.A(II5618), .Z(g4198) ) ;
INV     gate2418  (.A(g3914), .Z(II5622) ) ;
INV     gate2419  (.A(II5622), .Z(g4202) ) ;
INV     gate2420  (.A(g3914), .Z(II5626) ) ;
INV     gate2421  (.A(II5626), .Z(g4206) ) ;
INV     gate2422  (.A(g3914), .Z(II5630) ) ;
INV     gate2423  (.A(II5630), .Z(g4210) ) ;
AND2    gate2424  (.A(g3448), .B(g1528), .Z(g3768) ) ;
INV     gate2425  (.A(g3768), .Z(II5633) ) ;
INV     gate2426  (.A(II5633), .Z(g4213) ) ;
INV     gate2427  (.A(g3914), .Z(II5637) ) ;
INV     gate2428  (.A(II5637), .Z(g4215) ) ;
INV     gate2429  (.A(g3770), .Z(II5640) ) ;
INV     gate2430  (.A(II5640), .Z(g4218) ) ;
INV     gate2431  (.A(g4059), .Z(II5644) ) ;
INV     gate2432  (.A(II5644), .Z(g4220) ) ;
NAND2   gate2433  (.A(II4920), .B(II4921), .Z(g3742) ) ;
INV     gate2434  (.A(g3742), .Z(II5654) ) ;
INV     gate2435  (.A(II5654), .Z(g4222) ) ;
AND2    gate2436  (.A(II5351), .B(II5352), .Z(g4046) ) ;
INV     gate2437  (.A(g4046), .Z(g4224) ) ;
INV     gate2438  (.A(g4059), .Z(g4225) ) ;
AND2    gate2439  (.A(II5359), .B(II5360), .Z(g4050) ) ;
INV     gate2440  (.A(g4050), .Z(g4226) ) ;
INV     gate2441  (.A(g4059), .Z(g4227) ) ;
OR2     gate2442  (.A(g3304), .B(g1351), .Z(g3828) ) ;
INV     gate2443  (.A(g3828), .Z(II5668) ) ;
INV     gate2444  (.A(II5668), .Z(g4228) ) ;
INV     gate2445  (.A(g4059), .Z(g4229) ) ;
INV     gate2446  (.A(g4003), .Z(II5674) ) ;
INV     gate2447  (.A(II5674), .Z(g4232) ) ;
OR2     gate2448  (.A(g3215), .B(g3575), .Z(g3942) ) ;
INV     gate2449  (.A(g3942), .Z(II5686) ) ;
INV     gate2450  (.A(II5686), .Z(g4242) ) ;
INV     gate2451  (.A(g3942), .Z(II5692) ) ;
INV     gate2452  (.A(II5692), .Z(g4246) ) ;
INV     gate2453  (.A(g3942), .Z(II5696) ) ;
INV     gate2454  (.A(II5696), .Z(g4248) ) ;
AND2    gate2455  (.A(g3540), .B(g1665), .Z(g3844) ) ;
INV     gate2456  (.A(g3844), .Z(II5699) ) ;
INV     gate2457  (.A(II5699), .Z(g4249) ) ;
INV     gate2458  (.A(g3845), .Z(II5702) ) ;
INV     gate2459  (.A(II5702), .Z(g4250) ) ;
INV     gate2460  (.A(g3942), .Z(II5705) ) ;
INV     gate2461  (.A(II5705), .Z(g4251) ) ;
INV     gate2462  (.A(g3942), .Z(II5708) ) ;
INV     gate2463  (.A(II5708), .Z(g4252) ) ;
INV     gate2464  (.A(g4022), .Z(II5713) ) ;
INV     gate2465  (.A(II5713), .Z(g4262) ) ;
INV     gate2466  (.A(g3942), .Z(II5716) ) ;
INV     gate2467  (.A(II5716), .Z(g4265) ) ;
INV     gate2468  (.A(g4022), .Z(II5720) ) ;
INV     gate2469  (.A(II5720), .Z(g4267) ) ;
INV     gate2470  (.A(g3942), .Z(II5723) ) ;
INV     gate2471  (.A(II5723), .Z(g4270) ) ;
INV     gate2472  (.A(g4022), .Z(II5728) ) ;
INV     gate2473  (.A(II5728), .Z(g4273) ) ;
INV     gate2474  (.A(g3942), .Z(II5731) ) ;
INV     gate2475  (.A(II5731), .Z(g4276) ) ;
INV     gate2476  (.A(g4022), .Z(II5736) ) ;
INV     gate2477  (.A(II5736), .Z(g4281) ) ;
INV     gate2478  (.A(g3942), .Z(II5739) ) ;
INV     gate2479  (.A(II5739), .Z(g4284) ) ;
INV     gate2480  (.A(g4022), .Z(II5743) ) ;
INV     gate2481  (.A(II5743), .Z(g4286) ) ;
INV     gate2482  (.A(g4022), .Z(II5746) ) ;
INV     gate2483  (.A(II5746), .Z(g4289) ) ;
INV     gate2484  (.A(g4059), .Z(g4292) ) ;
INV     gate2485  (.A(g4022), .Z(II5750) ) ;
INV     gate2486  (.A(II5750), .Z(g4293) ) ;
INV     gate2487  (.A(g4022), .Z(II5753) ) ;
INV     gate2488  (.A(II5753), .Z(g4296) ) ;
INV     gate2489  (.A(g3922), .Z(II5756) ) ;
INV     gate2490  (.A(II5756), .Z(g4299) ) ;
OR2     gate2491  (.A(g3293), .B(g2685), .Z(g4068) ) ;
INV     gate2492  (.A(g4068), .Z(g4302) ) ;
INV     gate2493  (.A(g3807), .Z(II5774) ) ;
INV     gate2494  (.A(g3807), .Z(II5777) ) ;
INV     gate2495  (.A(II5777), .Z(g4308) ) ;
OR2     gate2496  (.A(g3301), .B(g2699), .Z(g4074) ) ;
INV     gate2497  (.A(g4074), .Z(g4309) ) ;
OR2     gate2498  (.A(g3302), .B(g2700), .Z(g4080) ) ;
INV     gate2499  (.A(g4080), .Z(g4314) ) ;
INV     gate2500  (.A(g4011), .Z(g4320) ) ;
INV     gate2501  (.A(g3803), .Z(II5790) ) ;
INV     gate2502  (.A(g3803), .Z(II5793) ) ;
INV     gate2503  (.A(II5793), .Z(g4322) ) ;
OR2     gate2504  (.A(g3310), .B(g2720), .Z(g4086) ) ;
INV     gate2505  (.A(g4086), .Z(g4323) ) ;
OR2     gate2506  (.A(g3311), .B(g2721), .Z(g4092) ) ;
INV     gate2507  (.A(g4092), .Z(g4328) ) ;
OR2     gate2508  (.A(g3325), .B(g2733), .Z(g3733) ) ;
INV     gate2509  (.A(g3733), .Z(g4334) ) ;
INV     gate2510  (.A(g4011), .Z(g4343) ) ;
INV     gate2511  (.A(g4010), .Z(g4350) ) ;
INV     gate2512  (.A(g3914), .Z(II5825) ) ;
INV     gate2513  (.A(II5825), .Z(g4364) ) ;
OR2     gate2514  (.A(g3670), .B(g3135), .Z(g3842) ) ;
INV     gate2515  (.A(g3842), .Z(II5831) ) ;
INV     gate2516  (.A(II5831), .Z(g4370) ) ;
OR2     gate2517  (.A(g3680), .B(g3145), .Z(g3850) ) ;
INV     gate2518  (.A(g3850), .Z(II5837) ) ;
INV     gate2519  (.A(II5837), .Z(g4374) ) ;
OR2     gate2520  (.A(g3324), .B(g2732), .Z(g3732) ) ;
INV     gate2521  (.A(g3732), .Z(II5840) ) ;
INV     gate2522  (.A(II5840), .Z(g4375) ) ;
OR2     gate2523  (.A(g3681), .B(g3146), .Z(g3851) ) ;
INV     gate2524  (.A(g3851), .Z(II5843) ) ;
INV     gate2525  (.A(II5843), .Z(g4376) ) ;
OR2     gate2526  (.A(g3686), .B(g3157), .Z(g3856) ) ;
INV     gate2527  (.A(g3856), .Z(II5848) ) ;
INV     gate2528  (.A(II5848), .Z(g4379) ) ;
OR2     gate2529  (.A(g3334), .B(g2746), .Z(g3739) ) ;
INV     gate2530  (.A(g3739), .Z(II5851) ) ;
INV     gate2531  (.A(II5851), .Z(g4380) ) ;
OR2     gate2532  (.A(g3687), .B(g3161), .Z(g3857) ) ;
INV     gate2533  (.A(g3857), .Z(II5854) ) ;
INV     gate2534  (.A(II5854), .Z(g4381) ) ;
OR2     gate2535  (.A(g3335), .B(g2747), .Z(g3740) ) ;
INV     gate2536  (.A(g3740), .Z(II5857) ) ;
INV     gate2537  (.A(II5857), .Z(g4382) ) ;
OR2     gate2538  (.A(g3692), .B(g3172), .Z(g3863) ) ;
INV     gate2539  (.A(g3863), .Z(II5862) ) ;
INV     gate2540  (.A(II5862), .Z(g4385) ) ;
OR2     gate2541  (.A(g3344), .B(g2758), .Z(g3743) ) ;
INV     gate2542  (.A(g3743), .Z(II5865) ) ;
INV     gate2543  (.A(II5865), .Z(g4386) ) ;
OR2     gate2544  (.A(g3693), .B(g3176), .Z(g3864) ) ;
INV     gate2545  (.A(g3864), .Z(II5868) ) ;
INV     gate2546  (.A(II5868), .Z(g4387) ) ;
OR2     gate2547  (.A(g3345), .B(g2759), .Z(g3744) ) ;
INV     gate2548  (.A(g3744), .Z(II5871) ) ;
INV     gate2549  (.A(II5871), .Z(g4388) ) ;
OR2     gate2550  (.A(g3700), .B(g3182), .Z(g3870) ) ;
INV     gate2551  (.A(g3870), .Z(II5876) ) ;
INV     gate2552  (.A(II5876), .Z(g4391) ) ;
OR2     gate2553  (.A(g3356), .B(g2770), .Z(g3745) ) ;
INV     gate2554  (.A(g3745), .Z(II5879) ) ;
INV     gate2555  (.A(II5879), .Z(g4392) ) ;
OR2     gate2556  (.A(g3701), .B(g3186), .Z(g3871) ) ;
INV     gate2557  (.A(g3871), .Z(II5882) ) ;
INV     gate2558  (.A(II5882), .Z(g4393) ) ;
OR2     gate2559  (.A(g3357), .B(g2771), .Z(g3746) ) ;
INV     gate2560  (.A(g3746), .Z(II5885) ) ;
INV     gate2561  (.A(II5885), .Z(g4394) ) ;
OR2     gate2562  (.A(g3703), .B(g3191), .Z(g3878) ) ;
INV     gate2563  (.A(g3878), .Z(II5890) ) ;
INV     gate2564  (.A(II5890), .Z(g4397) ) ;
OR2     gate2565  (.A(g3365), .B(g2781), .Z(g3747) ) ;
INV     gate2566  (.A(g3747), .Z(II5893) ) ;
INV     gate2567  (.A(II5893), .Z(g4398) ) ;
OR2     gate2568  (.A(g3704), .B(g3195), .Z(g3879) ) ;
INV     gate2569  (.A(g3879), .Z(II5896) ) ;
INV     gate2570  (.A(II5896), .Z(g4399) ) ;
OR2     gate2571  (.A(g3366), .B(g2782), .Z(g3748) ) ;
INV     gate2572  (.A(g3748), .Z(II5899) ) ;
INV     gate2573  (.A(II5899), .Z(g4400) ) ;
NAND2   gate2574  (.A(g107), .B(g3425), .Z(g4017) ) ;
INV     gate2575  (.A(g4017), .Z(g4402) ) ;
OR2     gate2576  (.A(g3371), .B(g2793), .Z(g3749) ) ;
INV     gate2577  (.A(g3749), .Z(II5904) ) ;
INV     gate2578  (.A(II5904), .Z(g4403) ) ;
OR2     gate2579  (.A(g3709), .B(g3203), .Z(g3883) ) ;
INV     gate2580  (.A(g3883), .Z(II5907) ) ;
INV     gate2581  (.A(II5907), .Z(g4404) ) ;
OR2     gate2582  (.A(g3372), .B(g2794), .Z(g3750) ) ;
INV     gate2583  (.A(g3750), .Z(II5910) ) ;
INV     gate2584  (.A(II5910), .Z(g4405) ) ;
OR2     gate2585  (.A(g3375), .B(g2807), .Z(g3751) ) ;
INV     gate2586  (.A(g3751), .Z(II5913) ) ;
INV     gate2587  (.A(II5913), .Z(g4406) ) ;
INV     gate2588  (.A(g4228), .Z(II5920) ) ;
INV     gate2589  (.A(g4299), .Z(II5923) ) ;
INV     gate2590  (.A(g4153), .Z(II5926) ) ;
INV     gate2591  (.A(g4152), .Z(II5929) ) ;
AND2    gate2592  (.A(g157), .B(g3773), .Z(g4346) ) ;
INV     gate2593  (.A(g4346), .Z(II5933) ) ;
INV     gate2594  (.A(II5933), .Z(g4428) ) ;
AND2    gate2595  (.A(g166), .B(g3776), .Z(g4351) ) ;
INV     gate2596  (.A(g4351), .Z(II5938) ) ;
INV     gate2597  (.A(II5938), .Z(g4431) ) ;
AND2    gate2598  (.A(g175), .B(g3779), .Z(g4356) ) ;
INV     gate2599  (.A(g4356), .Z(II5944) ) ;
INV     gate2600  (.A(II5944), .Z(g4435) ) ;
AND2    gate2601  (.A(g184), .B(g3785), .Z(g4360) ) ;
INV     gate2602  (.A(g4360), .Z(II5948) ) ;
INV     gate2603  (.A(II5948), .Z(g4437) ) ;
AND2    gate2604  (.A(g193), .B(g3788), .Z(g4367) ) ;
INV     gate2605  (.A(g4367), .Z(II5952) ) ;
INV     gate2606  (.A(II5952), .Z(g4439) ) ;
NAND2   gate2607  (.A(II5783), .B(II5784), .Z(g4319) ) ;
INV     gate2608  (.A(g4319), .Z(II5977) ) ;
INV     gate2609  (.A(II5977), .Z(g4462) ) ;
INV     gate2610  (.A(g4364), .Z(g4463) ) ;
INV     gate2611  (.A(g4224), .Z(II5987) ) ;
INV     gate2612  (.A(II5987), .Z(g4485) ) ;
INV     gate2613  (.A(g4226), .Z(II5991) ) ;
INV     gate2614  (.A(II5991), .Z(g4487) ) ;
AND2    gate2615  (.A(g3830), .B(g1533), .Z(g4157) ) ;
INV     gate2616  (.A(g4157), .Z(II5998) ) ;
INV     gate2617  (.A(II5998), .Z(g4492) ) ;
INV     gate2618  (.A(g4162), .Z(II6001) ) ;
INV     gate2619  (.A(II6001), .Z(g4493) ) ;
AND2    gate2620  (.A(g370), .B(g3890), .Z(g4159) ) ;
INV     gate2621  (.A(g4159), .Z(II6004) ) ;
INV     gate2622  (.A(II6004), .Z(g4494) ) ;
AND2    gate2623  (.A(g374), .B(g3892), .Z(g4163) ) ;
INV     gate2624  (.A(g4163), .Z(II6008) ) ;
INV     gate2625  (.A(II6008), .Z(g4496) ) ;
AND2    gate2626  (.A(g378), .B(g3898), .Z(g4167) ) ;
INV     gate2627  (.A(g4167), .Z(II6012) ) ;
INV     gate2628  (.A(II6012), .Z(g4498) ) ;
AND2    gate2629  (.A(g382), .B(g3900), .Z(g4170) ) ;
INV     gate2630  (.A(g4170), .Z(II6015) ) ;
INV     gate2631  (.A(II6015), .Z(g4499) ) ;
AND2    gate2632  (.A(g386), .B(g3901), .Z(g4176) ) ;
INV     gate2633  (.A(g4176), .Z(II6020) ) ;
INV     gate2634  (.A(II6020), .Z(g4502) ) ;
NAND2   gate2635  (.A(II5536), .B(II5537), .Z(g4151) ) ;
INV     gate2636  (.A(g4151), .Z(II6023) ) ;
INV     gate2637  (.A(II6023), .Z(g4503) ) ;
AND2    gate2638  (.A(g390), .B(g3902), .Z(g4179) ) ;
INV     gate2639  (.A(g4179), .Z(II6033) ) ;
INV     gate2640  (.A(II6033), .Z(g4507) ) ;
INV     gate2641  (.A(g4370), .Z(II6036) ) ;
INV     gate2642  (.A(II6036), .Z(g4508) ) ;
AND2    gate2643  (.A(g394), .B(g3904), .Z(g4182) ) ;
INV     gate2644  (.A(g4182), .Z(II6039) ) ;
INV     gate2645  (.A(II6039), .Z(g4509) ) ;
INV     gate2646  (.A(g4374), .Z(II6042) ) ;
INV     gate2647  (.A(II6042), .Z(g4510) ) ;
INV     gate2648  (.A(g4375), .Z(II6045) ) ;
INV     gate2649  (.A(II6045), .Z(g4511) ) ;
INV     gate2650  (.A(g4376), .Z(II6048) ) ;
INV     gate2651  (.A(II6048), .Z(g4512) ) ;
AND2    gate2652  (.A(g398), .B(g3906), .Z(g4185) ) ;
INV     gate2653  (.A(g4185), .Z(II6051) ) ;
INV     gate2654  (.A(II6051), .Z(g4513) ) ;
INV     gate2655  (.A(g4194), .Z(II6054) ) ;
INV     gate2656  (.A(II6054), .Z(g4514) ) ;
INV     gate2657  (.A(g4379), .Z(II6057) ) ;
INV     gate2658  (.A(II6057), .Z(g4515) ) ;
INV     gate2659  (.A(g4380), .Z(II6060) ) ;
INV     gate2660  (.A(II6060), .Z(g4516) ) ;
INV     gate2661  (.A(g4381), .Z(II6063) ) ;
INV     gate2662  (.A(II6063), .Z(g4517) ) ;
INV     gate2663  (.A(g4382), .Z(II6066) ) ;
INV     gate2664  (.A(II6066), .Z(g4518) ) ;
INV     gate2665  (.A(g4213), .Z(II6069) ) ;
INV     gate2666  (.A(II6069), .Z(g4519) ) ;
INV     gate2667  (.A(g4385), .Z(II6072) ) ;
INV     gate2668  (.A(II6072), .Z(g4520) ) ;
INV     gate2669  (.A(g4386), .Z(II6075) ) ;
INV     gate2670  (.A(II6075), .Z(g4521) ) ;
INV     gate2671  (.A(g4387), .Z(II6078) ) ;
INV     gate2672  (.A(II6078), .Z(g4522) ) ;
INV     gate2673  (.A(g4388), .Z(II6081) ) ;
INV     gate2674  (.A(II6081), .Z(g4523) ) ;
INV     gate2675  (.A(g4391), .Z(II6084) ) ;
INV     gate2676  (.A(II6084), .Z(g4524) ) ;
INV     gate2677  (.A(g4392), .Z(II6087) ) ;
INV     gate2678  (.A(II6087), .Z(g4525) ) ;
INV     gate2679  (.A(g4393), .Z(II6090) ) ;
INV     gate2680  (.A(II6090), .Z(g4526) ) ;
INV     gate2681  (.A(g4394), .Z(II6093) ) ;
INV     gate2682  (.A(II6093), .Z(g4527) ) ;
INV     gate2683  (.A(g4397), .Z(II6096) ) ;
INV     gate2684  (.A(II6096), .Z(g4528) ) ;
INV     gate2685  (.A(g4398), .Z(II6099) ) ;
INV     gate2686  (.A(II6099), .Z(g4529) ) ;
INV     gate2687  (.A(g4399), .Z(II6102) ) ;
INV     gate2688  (.A(II6102), .Z(g4530) ) ;
INV     gate2689  (.A(g4400), .Z(II6105) ) ;
INV     gate2690  (.A(II6105), .Z(g4531) ) ;
INV     gate2691  (.A(g4403), .Z(II6108) ) ;
INV     gate2692  (.A(II6108), .Z(g4532) ) ;
INV     gate2693  (.A(g4404), .Z(II6111) ) ;
INV     gate2694  (.A(II6111), .Z(g4533) ) ;
INV     gate2695  (.A(g4405), .Z(II6114) ) ;
INV     gate2696  (.A(II6114), .Z(g4534) ) ;
INV     gate2697  (.A(g4173), .Z(g4535) ) ;
INV     gate2698  (.A(g4406), .Z(II6118) ) ;
INV     gate2699  (.A(II6118), .Z(g4536) ) ;
AND2    gate2700  (.A(g3903), .B(g1474), .Z(g4410) ) ;
INV     gate2701  (.A(g4410), .Z(g4537) ) ;
AND2    gate2702  (.A(g3905), .B(g1481), .Z(g4416) ) ;
INV     gate2703  (.A(g4416), .Z(g4545) ) ;
NOR3    gate2704  (.A(g1589), .B(g1879), .C(g3793), .Z(g4240) ) ;
INV     gate2705  (.A(g4240), .Z(II6126) ) ;
INV     gate2706  (.A(II6126), .Z(g4550) ) ;
INV     gate2707  (.A(g4187), .Z(g4559) ) ;
INV     gate2708  (.A(g4188), .Z(g4560) ) ;
INV     gate2709  (.A(g4189), .Z(g4561) ) ;
AND2    gate2710  (.A(g3911), .B(g1655), .Z(g4219) ) ;
INV     gate2711  (.A(g4219), .Z(II6132) ) ;
INV     gate2712  (.A(II6132), .Z(g4562) ) ;
INV     gate2713  (.A(g4190), .Z(g4563) ) ;
INV     gate2714  (.A(g4192), .Z(g4564) ) ;
INV     gate2715  (.A(g4195), .Z(g4565) ) ;
INV     gate2716  (.A(g4198), .Z(g4566) ) ;
INV     gate2717  (.A(g4222), .Z(II6139) ) ;
INV     gate2718  (.A(II6139), .Z(g4567) ) ;
NAND2   gate2719  (.A(g4049), .B(g4017), .Z(g4237) ) ;
INV     gate2720  (.A(g4237), .Z(II6143) ) ;
INV     gate2721  (.A(II6143), .Z(g4569) ) ;
INV     gate2722  (.A(g4202), .Z(g4577) ) ;
INV     gate2723  (.A(g4206), .Z(g4579) ) ;
INV     gate2724  (.A(g4210), .Z(g4582) ) ;
INV     gate2725  (.A(g4215), .Z(g4587) ) ;
INV     gate2726  (.A(g4191), .Z(g4601) ) ;
INV     gate2727  (.A(g4343), .Z(II6170) ) ;
INV     gate2728  (.A(II6170), .Z(g4603) ) ;
INV     gate2729  (.A(g4193), .Z(g4606) ) ;
INV     gate2730  (.A(g4249), .Z(II6182) ) ;
INV     gate2731  (.A(II6182), .Z(g4609) ) ;
INV     gate2732  (.A(g4320), .Z(g4612) ) ;
INV     gate2733  (.A(g4308), .Z(g4614) ) ;
INV     gate2734  (.A(g4322), .Z(g4615) ) ;
INV     gate2735  (.A(g4242), .Z(g4617) ) ;
INV     gate2736  (.A(g4246), .Z(g4618) ) ;
INV     gate2737  (.A(g4248), .Z(g4619) ) ;
INV     gate2738  (.A(g4251), .Z(g4620) ) ;
INV     gate2739  (.A(g4252), .Z(g4622) ) ;
INV     gate2740  (.A(g4262), .Z(g4623) ) ;
INV     gate2741  (.A(g4265), .Z(g4624) ) ;
INV     gate2742  (.A(g4267), .Z(g4625) ) ;
INV     gate2743  (.A(g4270), .Z(g4626) ) ;
INV     gate2744  (.A(g4273), .Z(g4628) ) ;
INV     gate2745  (.A(g4276), .Z(g4629) ) ;
INV     gate2746  (.A(g4281), .Z(g4632) ) ;
INV     gate2747  (.A(g4284), .Z(g4633) ) ;
INV     gate2748  (.A(g4286), .Z(g4636) ) ;
INV     gate2749  (.A(g4289), .Z(g4639) ) ;
INV     gate2750  (.A(g4293), .Z(g4643) ) ;
INV     gate2751  (.A(g4350), .Z(II6231) ) ;
INV     gate2752  (.A(II6231), .Z(g4644) ) ;
INV     gate2753  (.A(g4296), .Z(g4647) ) ;
INV     gate2754  (.A(g4519), .Z(II6244) ) ;
INV     gate2755  (.A(g4609), .Z(II6247) ) ;
INV     gate2756  (.A(g4514), .Z(II6250) ) ;
NAND2   gate2757  (.A(II6176), .B(II6177), .Z(g4608) ) ;
INV     gate2758  (.A(g4608), .Z(II6253) ) ;
INV     gate2759  (.A(II6253), .Z(g4660) ) ;
NAND2   gate2760  (.A(g4402), .B(g1056), .Z(g4640) ) ;
INV     gate2761  (.A(g4640), .Z(g4662) ) ;
OR2     gate2762  (.A(g4368), .B(g3660), .Z(g4655) ) ;
INV     gate2763  (.A(g4655), .Z(II6269) ) ;
INV     gate2764  (.A(II6269), .Z(g4679) ) ;
OR2     gate2765  (.A(g4349), .B(g4015), .Z(g4430) ) ;
INV     gate2766  (.A(g4430), .Z(II6280) ) ;
INV     gate2767  (.A(II6280), .Z(g4692) ) ;
NAND2   gate2768  (.A(II6195), .B(II6196), .Z(g4613) ) ;
INV     gate2769  (.A(g4613), .Z(II6283) ) ;
INV     gate2770  (.A(II6283), .Z(g4693) ) ;
OR2     gate2771  (.A(g4354), .B(g4032), .Z(g4433) ) ;
INV     gate2772  (.A(g4433), .Z(II6289) ) ;
INV     gate2773  (.A(II6289), .Z(g4699) ) ;
OR2     gate2774  (.A(g4355), .B(g4033), .Z(g4434) ) ;
INV     gate2775  (.A(g4434), .Z(II6292) ) ;
INV     gate2776  (.A(II6292), .Z(g4700) ) ;
OR2     gate2777  (.A(g4359), .B(g4035), .Z(g4436) ) ;
INV     gate2778  (.A(g4436), .Z(II6296) ) ;
INV     gate2779  (.A(II6296), .Z(g4702) ) ;
OR2     gate2780  (.A(g4363), .B(g4037), .Z(g4438) ) ;
INV     gate2781  (.A(g4438), .Z(II6299) ) ;
INV     gate2782  (.A(II6299), .Z(g4703) ) ;
OR2     gate2783  (.A(g4371), .B(g4038), .Z(g4440) ) ;
INV     gate2784  (.A(g4440), .Z(II6302) ) ;
INV     gate2785  (.A(II6302), .Z(g4704) ) ;
OR2     gate2786  (.A(g4372), .B(g4039), .Z(g4441) ) ;
INV     gate2787  (.A(g4441), .Z(II6305) ) ;
INV     gate2788  (.A(II6305), .Z(g4705) ) ;
OR2     gate2789  (.A(g4377), .B(g4041), .Z(g4443) ) ;
INV     gate2790  (.A(g4443), .Z(II6308) ) ;
INV     gate2791  (.A(II6308), .Z(g4706) ) ;
OR2     gate2792  (.A(g4378), .B(g4042), .Z(g4444) ) ;
INV     gate2793  (.A(g4444), .Z(II6311) ) ;
INV     gate2794  (.A(II6311), .Z(g4707) ) ;
OR2     gate2795  (.A(g4383), .B(g4043), .Z(g4446) ) ;
INV     gate2796  (.A(g4446), .Z(II6315) ) ;
INV     gate2797  (.A(II6315), .Z(g4711) ) ;
OR2     gate2798  (.A(g4384), .B(g4044), .Z(g4447) ) ;
INV     gate2799  (.A(g4447), .Z(II6318) ) ;
INV     gate2800  (.A(II6318), .Z(g4712) ) ;
INV     gate2801  (.A(g4559), .Z(II6321) ) ;
INV     gate2802  (.A(II6321), .Z(g4713) ) ;
OR2     gate2803  (.A(g4389), .B(g4047), .Z(g4450) ) ;
INV     gate2804  (.A(g4450), .Z(II6324) ) ;
INV     gate2805  (.A(II6324), .Z(g4714) ) ;
OR2     gate2806  (.A(g4390), .B(g4048), .Z(g4451) ) ;
INV     gate2807  (.A(g4451), .Z(II6327) ) ;
INV     gate2808  (.A(II6327), .Z(g4715) ) ;
INV     gate2809  (.A(g4560), .Z(II6330) ) ;
INV     gate2810  (.A(II6330), .Z(g4716) ) ;
NAND2   gate2811  (.A(g319), .B(g4253), .Z(g4465) ) ;
INV     gate2812  (.A(g4465), .Z(g4717) ) ;
OR2     gate2813  (.A(g4395), .B(g4051), .Z(g4454) ) ;
INV     gate2814  (.A(g4454), .Z(II6334) ) ;
INV     gate2815  (.A(II6334), .Z(g4718) ) ;
OR2     gate2816  (.A(g4396), .B(g4052), .Z(g4455) ) ;
INV     gate2817  (.A(g4455), .Z(II6337) ) ;
INV     gate2818  (.A(II6337), .Z(g4719) ) ;
INV     gate2819  (.A(g4561), .Z(II6340) ) ;
INV     gate2820  (.A(II6340), .Z(g4720) ) ;
OR2     gate2821  (.A(g4401), .B(g4057), .Z(g4458) ) ;
INV     gate2822  (.A(g4458), .Z(II6343) ) ;
INV     gate2823  (.A(II6343), .Z(g4721) ) ;
INV     gate2824  (.A(g4563), .Z(II6346) ) ;
INV     gate2825  (.A(II6346), .Z(g4722) ) ;
INV     gate2826  (.A(g4569), .Z(II6349) ) ;
INV     gate2827  (.A(II6349), .Z(g4723) ) ;
INV     gate2828  (.A(g4564), .Z(II6352) ) ;
INV     gate2829  (.A(II6352), .Z(g4726) ) ;
INV     gate2830  (.A(g4569), .Z(II6355) ) ;
INV     gate2831  (.A(II6355), .Z(g4727) ) ;
INV     gate2832  (.A(g4566), .Z(II6359) ) ;
INV     gate2833  (.A(II6359), .Z(g4731) ) ;
INV     gate2834  (.A(g4569), .Z(II6362) ) ;
INV     gate2835  (.A(II6362), .Z(g4732) ) ;
INV     gate2836  (.A(g4569), .Z(II6366) ) ;
INV     gate2837  (.A(II6366), .Z(g4736) ) ;
INV     gate2838  (.A(g4569), .Z(II6371) ) ;
INV     gate2839  (.A(II6371), .Z(g4741) ) ;
INV     gate2840  (.A(g4569), .Z(II6377) ) ;
INV     gate2841  (.A(II6377), .Z(g4753) ) ;
AND2    gate2842  (.A(g4218), .B(g1539), .Z(g4460) ) ;
INV     gate2843  (.A(g4460), .Z(II6382) ) ;
INV     gate2844  (.A(II6382), .Z(g4758) ) ;
INV     gate2845  (.A(g4462), .Z(II6386) ) ;
INV     gate2846  (.A(II6386), .Z(g4760) ) ;
OR2     gate2847  (.A(g3575), .B(g4253), .Z(g4473) ) ;
INV     gate2848  (.A(g4473), .Z(II6397) ) ;
INV     gate2849  (.A(II6397), .Z(g4763) ) ;
INV     gate2850  (.A(g4473), .Z(II6400) ) ;
INV     gate2851  (.A(II6400), .Z(g4764) ) ;
INV     gate2852  (.A(g4492), .Z(II6403) ) ;
INV     gate2853  (.A(II6403), .Z(g4765) ) ;
INV     gate2854  (.A(g4473), .Z(II6406) ) ;
INV     gate2855  (.A(II6406), .Z(g4766) ) ;
INV     gate2856  (.A(g4601), .Z(g4767) ) ;
INV     gate2857  (.A(g4473), .Z(II6410) ) ;
INV     gate2858  (.A(II6410), .Z(g4768) ) ;
INV     gate2859  (.A(g4606), .Z(g4769) ) ;
OR2     gate2860  (.A(g4166), .B(g3784), .Z(g4497) ) ;
INV     gate2861  (.A(g4497), .Z(II6414) ) ;
INV     gate2862  (.A(II6414), .Z(g4770) ) ;
INV     gate2863  (.A(g4617), .Z(II6417) ) ;
INV     gate2864  (.A(II6417), .Z(g4771) ) ;
INV     gate2865  (.A(g4618), .Z(II6420) ) ;
INV     gate2866  (.A(II6420), .Z(g4772) ) ;
INV     gate2867  (.A(g4619), .Z(II6425) ) ;
INV     gate2868  (.A(II6425), .Z(g4775) ) ;
INV     gate2869  (.A(g4620), .Z(II6430) ) ;
INV     gate2870  (.A(II6430), .Z(g4778) ) ;
INV     gate2871  (.A(g4622), .Z(II6434) ) ;
INV     gate2872  (.A(II6434), .Z(g4780) ) ;
AND2    gate2873  (.A(g4250), .B(g1671), .Z(g4501) ) ;
INV     gate2874  (.A(g4501), .Z(II6437) ) ;
INV     gate2875  (.A(II6437), .Z(g4781) ) ;
INV     gate2876  (.A(g4624), .Z(II6441) ) ;
INV     gate2877  (.A(II6441), .Z(g4783) ) ;
INV     gate2878  (.A(g4503), .Z(II6444) ) ;
INV     gate2879  (.A(II6444), .Z(g4784) ) ;
INV     gate2880  (.A(g4626), .Z(II6448) ) ;
INV     gate2881  (.A(II6448), .Z(g4786) ) ;
INV     gate2882  (.A(g4629), .Z(II6452) ) ;
INV     gate2883  (.A(II6452), .Z(g4788) ) ;
INV     gate2884  (.A(g4633), .Z(II6456) ) ;
INV     gate2885  (.A(II6456), .Z(g4790) ) ;
INV     gate2886  (.A(g4562), .Z(II6464) ) ;
INV     gate2887  (.A(II6464), .Z(g4798) ) ;
INV     gate2888  (.A(g4485), .Z(g4799) ) ;
INV     gate2889  (.A(g4487), .Z(g4801) ) ;
INV     gate2890  (.A(g4473), .Z(II6470) ) ;
INV     gate2891  (.A(II6470), .Z(g4802) ) ;
INV     gate2892  (.A(g4473), .Z(g4804) ) ;
INV     gate2893  (.A(g4473), .Z(g4805) ) ;
INV     gate2894  (.A(g4473), .Z(g4806) ) ;
INV     gate2895  (.A(g4473), .Z(g4807) ) ;
INV     gate2896  (.A(g4473), .Z(g4808) ) ;
INV     gate2897  (.A(g4603), .Z(II6485) ) ;
INV     gate2898  (.A(g4603), .Z(II6488) ) ;
INV     gate2899  (.A(II6488), .Z(g4810) ) ;
OR2     gate2900  (.A(g4232), .B(g3899), .Z(g4607) ) ;
INV     gate2901  (.A(g4607), .Z(II6495) ) ;
INV     gate2902  (.A(II6495), .Z(g4815) ) ;
INV     gate2903  (.A(g4614), .Z(g4822) ) ;
INV     gate2904  (.A(g4644), .Z(II6507) ) ;
INV     gate2905  (.A(II6507), .Z(g4823) ) ;
INV     gate2906  (.A(g4615), .Z(g4824) ) ;
INV     gate2907  (.A(g4473), .Z(g4837) ) ;
INV     gate2908  (.A(g4770), .Z(II6525) ) ;
INV     gate2909  (.A(g4815), .Z(II6528) ) ;
INV     gate2910  (.A(g4704), .Z(II6531) ) ;
INV     gate2911  (.A(g4706), .Z(II6534) ) ;
INV     gate2912  (.A(g4711), .Z(II6537) ) ;
INV     gate2913  (.A(g4714), .Z(II6540) ) ;
INV     gate2914  (.A(g4718), .Z(II6543) ) ;
INV     gate2915  (.A(g4692), .Z(II6546) ) ;
INV     gate2916  (.A(g4699), .Z(II6549) ) ;
INV     gate2917  (.A(g4702), .Z(II6552) ) ;
INV     gate2918  (.A(g4703), .Z(II6555) ) ;
INV     gate2919  (.A(g4705), .Z(II6558) ) ;
INV     gate2920  (.A(g4707), .Z(II6561) ) ;
INV     gate2921  (.A(g4712), .Z(II6564) ) ;
INV     gate2922  (.A(g4715), .Z(II6567) ) ;
INV     gate2923  (.A(g4719), .Z(II6570) ) ;
INV     gate2924  (.A(g4721), .Z(II6573) ) ;
INV     gate2925  (.A(g4700), .Z(II6576) ) ;
INV     gate2926  (.A(g4798), .Z(II6579) ) ;
INV     gate2927  (.A(g4765), .Z(II6582) ) ;
NAND2   gate2928  (.A(II6474), .B(II6475), .Z(g4803) ) ;
INV     gate2929  (.A(g4803), .Z(II6587) ) ;
INV     gate2930  (.A(II6587), .Z(g4861) ) ;
INV     gate2931  (.A(g4662), .Z(g4869) ) ;
INV     gate2932  (.A(g4823), .Z(II6599) ) ;
INV     gate2933  (.A(II6599), .Z(g4871) ) ;
NAND4   gate2934  (.A(g4550), .B(g965), .C(g1560), .D(g2073), .Z(g4813) ) ;
INV     gate2935  (.A(g4813), .Z(g4894) ) ;
OR2     gate2936  (.A(g4468), .B(g4569), .Z(g4745) ) ;
INV     gate2937  (.A(g4745), .Z(II6607) ) ;
INV     gate2938  (.A(II6607), .Z(g4900) ) ;
NAND4   gate2939  (.A(g4550), .B(g1560), .C(g1559), .D(g2073), .Z(g4812) ) ;
INV     gate2940  (.A(g4812), .Z(g4904) ) ;
INV     gate2941  (.A(g4660), .Z(II6612) ) ;
INV     gate2942  (.A(II6612), .Z(g4910) ) ;
INV     gate2943  (.A(g4745), .Z(II6615) ) ;
INV     gate2944  (.A(II6615), .Z(g4911) ) ;
NAND4   gate2945  (.A(g996), .B(g4550), .C(g1518), .D(g2073), .Z(g4816) ) ;
INV     gate2946  (.A(g4816), .Z(g4914) ) ;
NAND4   gate2947  (.A(g4550), .B(g1017), .C(g1680), .D(g2897), .Z(g4669) ) ;
INV     gate2948  (.A(g4669), .Z(g4915) ) ;
INV     gate2949  (.A(g4745), .Z(II6621) ) ;
INV     gate2950  (.A(II6621), .Z(g4929) ) ;
INV     gate2951  (.A(g4745), .Z(II6625) ) ;
INV     gate2952  (.A(II6625), .Z(g4933) ) ;
INV     gate2953  (.A(g4745), .Z(II6630) ) ;
INV     gate2954  (.A(II6630), .Z(g4938) ) ;
INV     gate2955  (.A(g4745), .Z(II6635) ) ;
INV     gate2956  (.A(II6635), .Z(g4943) ) ;
NAND4   gate2957  (.A(g2897), .B(g2101), .C(g1514), .D(g4550), .Z(g4678) ) ;
INV     gate2958  (.A(g4678), .Z(g4980) ) ;
AND2    gate2959  (.A(g4493), .B(g1542), .Z(g4687) ) ;
INV     gate2960  (.A(g4687), .Z(II6646) ) ;
INV     gate2961  (.A(II6646), .Z(g5010) ) ;
INV     gate2962  (.A(g4693), .Z(II6649) ) ;
INV     gate2963  (.A(II6649), .Z(g5011) ) ;
OR2     gate2964  (.A(g4448), .B(g4154), .Z(g4740) ) ;
INV     gate2965  (.A(g4740), .Z(II6666) ) ;
INV     gate2966  (.A(II6666), .Z(g5022) ) ;
NAND4   gate2967  (.A(g4550), .B(g1575), .C(g1550), .D(g2073), .Z(g4814) ) ;
INV     gate2968  (.A(g4814), .Z(g5025) ) ;
OR2     gate2969  (.A(g4452), .B(g4155), .Z(g4752) ) ;
INV     gate2970  (.A(g4752), .Z(II6672) ) ;
INV     gate2971  (.A(II6672), .Z(g5042) ) ;
OR2     gate2972  (.A(g4456), .B(g4158), .Z(g4757) ) ;
INV     gate2973  (.A(g4757), .Z(II6677) ) ;
INV     gate2974  (.A(II6677), .Z(g5045) ) ;
INV     gate2975  (.A(g4713), .Z(II6680) ) ;
INV     gate2976  (.A(II6680), .Z(g5046) ) ;
INV     gate2977  (.A(g4716), .Z(II6685) ) ;
INV     gate2978  (.A(II6685), .Z(g5049) ) ;
INV     gate2979  (.A(g4758), .Z(II6689) ) ;
INV     gate2980  (.A(II6689), .Z(g5051) ) ;
INV     gate2981  (.A(g4720), .Z(II6692) ) ;
INV     gate2982  (.A(II6692), .Z(g5052) ) ;
INV     gate2983  (.A(g4816), .Z(g5054) ) ;
INV     gate2984  (.A(g4722), .Z(II6697) ) ;
INV     gate2985  (.A(II6697), .Z(g5059) ) ;
INV     gate2986  (.A(g4726), .Z(II6701) ) ;
INV     gate2987  (.A(II6701), .Z(g5061) ) ;
INV     gate2988  (.A(g4799), .Z(g5063) ) ;
INV     gate2989  (.A(g4731), .Z(II6706) ) ;
INV     gate2990  (.A(II6706), .Z(g5064) ) ;
INV     gate2991  (.A(g4801), .Z(g5067) ) ;
INV     gate2992  (.A(g4723), .Z(g5082) ) ;
INV     gate2993  (.A(g4727), .Z(g5084) ) ;
INV     gate2994  (.A(g4732), .Z(g5086) ) ;
INV     gate2995  (.A(g4736), .Z(g5087) ) ;
AND2    gate2996  (.A(g4567), .B(g1674), .Z(g4761) ) ;
INV     gate2997  (.A(g4761), .Z(II6723) ) ;
INV     gate2998  (.A(II6723), .Z(g5089) ) ;
INV     gate2999  (.A(g4741), .Z(g5090) ) ;
INV     gate3000  (.A(g4753), .Z(g5092) ) ;
OR2     gate3001  (.A(g4495), .B(g4220), .Z(g4773) ) ;
INV     gate3002  (.A(g4773), .Z(II6733) ) ;
INV     gate3003  (.A(II6733), .Z(g5097) ) ;
INV     gate3004  (.A(g4662), .Z(II6737) ) ;
INV     gate3005  (.A(II6737), .Z(g5099) ) ;
INV     gate3006  (.A(g4781), .Z(II6740) ) ;
INV     gate3007  (.A(II6740), .Z(g5110) ) ;
INV     gate3008  (.A(g4771), .Z(II6750) ) ;
INV     gate3009  (.A(II6750), .Z(g5112) ) ;
INV     gate3010  (.A(g4772), .Z(II6753) ) ;
INV     gate3011  (.A(II6753), .Z(g5113) ) ;
INV     gate3012  (.A(g4775), .Z(II6756) ) ;
INV     gate3013  (.A(II6756), .Z(g5114) ) ;
INV     gate3014  (.A(g4778), .Z(II6759) ) ;
INV     gate3015  (.A(II6759), .Z(g5115) ) ;
INV     gate3016  (.A(g4810), .Z(g5116) ) ;
INV     gate3017  (.A(g4780), .Z(II6763) ) ;
INV     gate3018  (.A(II6763), .Z(g5117) ) ;
INV     gate3019  (.A(g4783), .Z(II6766) ) ;
INV     gate3020  (.A(II6766), .Z(g5118) ) ;
INV     gate3021  (.A(g4786), .Z(II6769) ) ;
INV     gate3022  (.A(II6769), .Z(g5119) ) ;
INV     gate3023  (.A(g4788), .Z(II6772) ) ;
INV     gate3024  (.A(II6772), .Z(g5120) ) ;
INV     gate3025  (.A(g4790), .Z(II6775) ) ;
INV     gate3026  (.A(II6775), .Z(g5121) ) ;
NAND2   gate3027  (.A(g4472), .B(g4465), .Z(g4825) ) ;
INV     gate3028  (.A(g4825), .Z(II6780) ) ;
INV     gate3029  (.A(II6780), .Z(g5124) ) ;
INV     gate3030  (.A(g4822), .Z(II6783) ) ;
INV     gate3031  (.A(II6783), .Z(g5135) ) ;
INV     gate3032  (.A(g4824), .Z(II6786) ) ;
INV     gate3033  (.A(II6786), .Z(g5136) ) ;
INV     gate3034  (.A(g4871), .Z(II6789) ) ;
INV     gate3035  (.A(g5097), .Z(II6792) ) ;
INV     gate3036  (.A(g5022), .Z(II6795) ) ;
INV     gate3037  (.A(g5042), .Z(II6798) ) ;
INV     gate3038  (.A(g5045), .Z(II6801) ) ;
INV     gate3039  (.A(g5051), .Z(II6809) ) ;
INV     gate3040  (.A(g5110), .Z(II6812) ) ;
NAND2   gate3041  (.A(II6744), .B(II6745), .Z(g5111) ) ;
INV     gate3042  (.A(g5111), .Z(II6816) ) ;
INV     gate3043  (.A(II6816), .Z(g5150) ) ;
NAND2   gate3044  (.A(II6660), .B(II6661), .Z(g5019) ) ;
INV     gate3045  (.A(g5019), .Z(II6819) ) ;
INV     gate3046  (.A(II6819), .Z(g5151) ) ;
INV     gate3047  (.A(g5099), .Z(g5155) ) ;
INV     gate3048  (.A(g5099), .Z(g5160) ) ;
INV     gate3049  (.A(g5099), .Z(g5168) ) ;
INV     gate3050  (.A(g5099), .Z(g5174) ) ;
INV     gate3051  (.A(g5099), .Z(g5179) ) ;
INV     gate3052  (.A(g5082), .Z(II6867) ) ;
INV     gate3053  (.A(II6867), .Z(g5199) ) ;
INV     gate3054  (.A(g4861), .Z(II6874) ) ;
INV     gate3055  (.A(II6874), .Z(g5210) ) ;
AND2    gate3056  (.A(g4760), .B(g1549), .Z(g4872) ) ;
INV     gate3057  (.A(g4872), .Z(II6885) ) ;
INV     gate3058  (.A(II6885), .Z(g5219) ) ;
NAND2   gate3059  (.A(g4717), .B(g858), .Z(g4903) ) ;
INV     gate3060  (.A(g4903), .Z(g5220) ) ;
INV     gate3061  (.A(g5010), .Z(II6895) ) ;
INV     gate3062  (.A(II6895), .Z(g5230) ) ;
OR2     gate3063  (.A(g4688), .B(g4271), .Z(g5083) ) ;
INV     gate3064  (.A(g5083), .Z(g5237) ) ;
OR2     gate3065  (.A(g4694), .B(g4280), .Z(g5085) ) ;
INV     gate3066  (.A(g5085), .Z(g5242) ) ;
INV     gate3067  (.A(g4900), .Z(g5247) ) ;
INV     gate3068  (.A(g4911), .Z(g5248) ) ;
INV     gate3069  (.A(g4929), .Z(g5250) ) ;
OR2     gate3070  (.A(g1595), .B(g4688), .Z(g5069) ) ;
INV     gate3071  (.A(g5069), .Z(g5251) ) ;
INV     gate3072  (.A(g4933), .Z(g5255) ) ;
OR2     gate3073  (.A(g1612), .B(g4694), .Z(g5077) ) ;
INV     gate3074  (.A(g5077), .Z(g5256) ) ;
INV     gate3075  (.A(g4938), .Z(g5260) ) ;
INV     gate3076  (.A(g5124), .Z(II6918) ) ;
INV     gate3077  (.A(II6918), .Z(g5261) ) ;
INV     gate3078  (.A(g4943), .Z(g5264) ) ;
INV     gate3079  (.A(g5124), .Z(II6923) ) ;
INV     gate3080  (.A(II6923), .Z(g5266) ) ;
INV     gate3081  (.A(g5124), .Z(II6927) ) ;
INV     gate3082  (.A(II6927), .Z(g5270) ) ;
AND2    gate3083  (.A(g4784), .B(g1679), .Z(g5017) ) ;
INV     gate3084  (.A(g5017), .Z(II6930) ) ;
INV     gate3085  (.A(II6930), .Z(g5273) ) ;
INV     gate3086  (.A(g5124), .Z(II6933) ) ;
INV     gate3087  (.A(II6933), .Z(g5274) ) ;
INV     gate3088  (.A(g5124), .Z(II6937) ) ;
INV     gate3089  (.A(II6937), .Z(g5278) ) ;
INV     gate3090  (.A(g5124), .Z(II6942) ) ;
INV     gate3091  (.A(II6942), .Z(g5292) ) ;
INV     gate3092  (.A(g5124), .Z(II6946) ) ;
INV     gate3093  (.A(II6946), .Z(g5296) ) ;
AND2    gate3094  (.A(g4285), .B(g4807), .Z(g5050) ) ;
INV     gate3095  (.A(g5050), .Z(II6949) ) ;
INV     gate3096  (.A(II6949), .Z(g5299) ) ;
INV     gate3097  (.A(g5124), .Z(II6952) ) ;
INV     gate3098  (.A(II6952), .Z(g5300) ) ;
INV     gate3099  (.A(g5124), .Z(II6956) ) ;
INV     gate3100  (.A(II6956), .Z(g5304) ) ;
INV     gate3101  (.A(g5089), .Z(II6959) ) ;
INV     gate3102  (.A(II6959), .Z(g5307) ) ;
INV     gate3103  (.A(g5063), .Z(g5309) ) ;
INV     gate3104  (.A(g5067), .Z(g5310) ) ;
INV     gate3105  (.A(g5135), .Z(II6972) ) ;
INV     gate3106  (.A(II6972), .Z(g5314) ) ;
INV     gate3107  (.A(g5116), .Z(g5315) ) ;
INV     gate3108  (.A(g5136), .Z(II6976) ) ;
INV     gate3109  (.A(II6976), .Z(g5316) ) ;
INV     gate3110  (.A(g5230), .Z(II6986) ) ;
INV     gate3111  (.A(g5307), .Z(II6989) ) ;
INV     gate3112  (.A(g5151), .Z(II6992) ) ;
INV     gate3113  (.A(g5220), .Z(II6995) ) ;
INV     gate3114  (.A(II6995), .Z(g5331) ) ;
NAND2   gate3115  (.A(II6963), .B(II6964), .Z(g5308) ) ;
INV     gate3116  (.A(g5308), .Z(II7002) ) ;
INV     gate3117  (.A(II7002), .Z(g5352) ) ;
INV     gate3118  (.A(g5314), .Z(II7007) ) ;
INV     gate3119  (.A(II7007), .Z(g5355) ) ;
INV     gate3120  (.A(g5316), .Z(II7012) ) ;
INV     gate3121  (.A(II7012), .Z(g5358) ) ;
AND2    gate3122  (.A(g4910), .B(g1480), .Z(g5149) ) ;
INV     gate3123  (.A(g5149), .Z(II7029) ) ;
INV     gate3124  (.A(II7029), .Z(g5375) ) ;
INV     gate3125  (.A(g5150), .Z(II7035) ) ;
INV     gate3126  (.A(II7035), .Z(g5379) ) ;
INV     gate3127  (.A(g5309), .Z(II7039) ) ;
INV     gate3128  (.A(II7039), .Z(g5381) ) ;
INV     gate3129  (.A(g5310), .Z(II7042) ) ;
INV     gate3130  (.A(II7042), .Z(g5382) ) ;
AND2    gate3131  (.A(g5011), .B(g1556), .Z(g5167) ) ;
INV     gate3132  (.A(g5167), .Z(II7045) ) ;
INV     gate3133  (.A(II7045), .Z(g5383) ) ;
INV     gate3134  (.A(g5220), .Z(g5384) ) ;
INV     gate3135  (.A(g5219), .Z(II7051) ) ;
INV     gate3136  (.A(II7051), .Z(g5387) ) ;
NAND2   gate3137  (.A(g676), .B(g5060), .Z(g5318) ) ;
INV     gate3138  (.A(g5318), .Z(II7055) ) ;
INV     gate3139  (.A(II7055), .Z(g5391) ) ;
OR2     gate3140  (.A(g5074), .B(g5124), .Z(g5281) ) ;
INV     gate3141  (.A(g5281), .Z(II7058) ) ;
INV     gate3142  (.A(II7058), .Z(g5392) ) ;
INV     gate3143  (.A(g5281), .Z(II7061) ) ;
INV     gate3144  (.A(II7061), .Z(g5395) ) ;
INV     gate3145  (.A(g5281), .Z(II7065) ) ;
INV     gate3146  (.A(II7065), .Z(g5399) ) ;
INV     gate3147  (.A(g5281), .Z(II7069) ) ;
INV     gate3148  (.A(II7069), .Z(g5403) ) ;
INV     gate3149  (.A(g5281), .Z(II7073) ) ;
INV     gate3150  (.A(II7073), .Z(g5407) ) ;
INV     gate3151  (.A(g5281), .Z(II7077) ) ;
INV     gate3152  (.A(II7077), .Z(g5411) ) ;
INV     gate3153  (.A(g5281), .Z(II7081) ) ;
INV     gate3154  (.A(II7081), .Z(g5415) ) ;
INV     gate3155  (.A(g5281), .Z(II7086) ) ;
INV     gate3156  (.A(II7086), .Z(g5420) ) ;
INV     gate3157  (.A(g5281), .Z(II7091) ) ;
INV     gate3158  (.A(II7091), .Z(g5425) ) ;
INV     gate3159  (.A(g5273), .Z(II7104) ) ;
INV     gate3160  (.A(II7104), .Z(g5432) ) ;
OR2     gate3161  (.A(g5023), .B(g4763), .Z(g5277) ) ;
INV     gate3162  (.A(g5277), .Z(II7107) ) ;
INV     gate3163  (.A(II7107), .Z(g5433) ) ;
OR2     gate3164  (.A(g5043), .B(g4764), .Z(g5291) ) ;
INV     gate3165  (.A(g5291), .Z(II7110) ) ;
INV     gate3166  (.A(II7110), .Z(g5434) ) ;
OR2     gate3167  (.A(g5047), .B(g4766), .Z(g5295) ) ;
INV     gate3168  (.A(g5295), .Z(II7113) ) ;
INV     gate3169  (.A(II7113), .Z(g5435) ) ;
INV     gate3170  (.A(g5299), .Z(II7116) ) ;
INV     gate3171  (.A(II7116), .Z(g5436) ) ;
OR2     gate3172  (.A(g5053), .B(g4768), .Z(g5303) ) ;
INV     gate3173  (.A(g5303), .Z(II7119) ) ;
INV     gate3174  (.A(II7119), .Z(g5437) ) ;
INV     gate3175  (.A(g5261), .Z(g5439) ) ;
INV     gate3176  (.A(g5266), .Z(g5440) ) ;
INV     gate3177  (.A(g5270), .Z(g5442) ) ;
INV     gate3178  (.A(g5274), .Z(g5445) ) ;
INV     gate3179  (.A(g5278), .Z(g5448) ) ;
INV     gate3180  (.A(g5292), .Z(g5450) ) ;
INV     gate3181  (.A(g5296), .Z(g5453) ) ;
INV     gate3182  (.A(g5300), .Z(g5456) ) ;
INV     gate3183  (.A(g5304), .Z(g5457) ) ;
OR2     gate3184  (.A(g5098), .B(g4802), .Z(g5323) ) ;
INV     gate3185  (.A(g5323), .Z(II7143) ) ;
INV     gate3186  (.A(II7143), .Z(g5465) ) ;
OR2     gate3187  (.A(g5048), .B(g672), .Z(g5231) ) ;
INV     gate3188  (.A(g5231), .Z(II7146) ) ;
INV     gate3189  (.A(II7146), .Z(g5466) ) ;
INV     gate3190  (.A(g5355), .Z(II7150) ) ;
INV     gate3191  (.A(g5358), .Z(II7153) ) ;
INV     gate3192  (.A(g5465), .Z(II7161) ) ;
INV     gate3193  (.A(g5433), .Z(II7164) ) ;
INV     gate3194  (.A(g5434), .Z(II7167) ) ;
INV     gate3195  (.A(g5435), .Z(II7170) ) ;
INV     gate3196  (.A(g5436), .Z(II7173) ) ;
INV     gate3197  (.A(g5437), .Z(II7176) ) ;
INV     gate3198  (.A(g5387), .Z(II7187) ) ;
INV     gate3199  (.A(g5432), .Z(II7190) ) ;
INV     gate3200  (.A(g5466), .Z(II7193) ) ;
NAND2   gate3201  (.A(II7098), .B(II7099), .Z(g5431) ) ;
INV     gate3202  (.A(g5431), .Z(II7197) ) ;
INV     gate3203  (.A(II7197), .Z(g5493) ) ;
OR2     gate3204  (.A(g3466), .B(g5311), .Z(g5458) ) ;
INV     gate3205  (.A(g5458), .Z(II7251) ) ;
INV     gate3206  (.A(II7251), .Z(g5509) ) ;
INV     gate3207  (.A(g5458), .Z(II7254) ) ;
INV     gate3208  (.A(II7254), .Z(g5512) ) ;
INV     gate3209  (.A(g5458), .Z(II7258) ) ;
INV     gate3210  (.A(II7258), .Z(g5518) ) ;
INV     gate3211  (.A(g5458), .Z(II7261) ) ;
INV     gate3212  (.A(II7261), .Z(g5521) ) ;
INV     gate3213  (.A(g5458), .Z(II7264) ) ;
INV     gate3214  (.A(II7264), .Z(g5524) ) ;
INV     gate3215  (.A(g5458), .Z(II7267) ) ;
INV     gate3216  (.A(II7267), .Z(g5527) ) ;
INV     gate3217  (.A(g5352), .Z(II7270) ) ;
INV     gate3218  (.A(II7270), .Z(g5530) ) ;
INV     gate3219  (.A(g5375), .Z(II7276) ) ;
INV     gate3220  (.A(II7276), .Z(g5534) ) ;
OR3     gate3221  (.A(g3868), .B(g5318), .C(g3992), .Z(g5467) ) ;
INV     gate3222  (.A(g5467), .Z(g5536) ) ;
OR2     gate3223  (.A(g3992), .B(g5318), .Z(g5385) ) ;
INV     gate3224  (.A(g5385), .Z(g5537) ) ;
INV     gate3225  (.A(g5331), .Z(g5538) ) ;
INV     gate3226  (.A(g5331), .Z(g5539) ) ;
INV     gate3227  (.A(g5383), .Z(II7284) ) ;
INV     gate3228  (.A(II7284), .Z(g5540) ) ;
INV     gate3229  (.A(g5331), .Z(g5542) ) ;
INV     gate3230  (.A(g5331), .Z(g5543) ) ;
INV     gate3231  (.A(g5331), .Z(g5544) ) ;
INV     gate3232  (.A(g5331), .Z(g5545) ) ;
OR3     gate3233  (.A(g5318), .B(g1589), .C(g3491), .Z(g5388) ) ;
INV     gate3234  (.A(g5388), .Z(g5546) ) ;
INV     gate3235  (.A(g5331), .Z(g5549) ) ;
INV     gate3236  (.A(g5331), .Z(g5550) ) ;
INV     gate3237  (.A(g5439), .Z(II7295) ) ;
INV     gate3238  (.A(II7295), .Z(g5551) ) ;
NAND2   gate3239  (.A(g2330), .B(g5311), .Z(g5455) ) ;
INV     gate3240  (.A(g5455), .Z(g5554) ) ;
INV     gate3241  (.A(g5381), .Z(g5563) ) ;
INV     gate3242  (.A(g5382), .Z(g5564) ) ;
AND2    gate3243  (.A(g5315), .B(g4612), .Z(g5452) ) ;
INV     gate3244  (.A(g5452), .Z(II7318) ) ;
INV     gate3245  (.A(II7318), .Z(g5566) ) ;
NOR2    gate3246  (.A(g5162), .B(g5169), .Z(g5418) ) ;
INV     gate3247  (.A(g5418), .Z(g5567) ) ;
NOR2    gate3248  (.A(g5170), .B(g5175), .Z(g5423) ) ;
INV     gate3249  (.A(g5423), .Z(g5568) ) ;
INV     gate3250  (.A(g5392), .Z(g5570) ) ;
INV     gate3251  (.A(g5395), .Z(g5571) ) ;
INV     gate3252  (.A(g5399), .Z(g5572) ) ;
INV     gate3253  (.A(g5403), .Z(g5573) ) ;
INV     gate3254  (.A(g5407), .Z(g5574) ) ;
INV     gate3255  (.A(g5411), .Z(g5575) ) ;
INV     gate3256  (.A(g5415), .Z(g5576) ) ;
INV     gate3257  (.A(g5420), .Z(g5577) ) ;
INV     gate3258  (.A(g5425), .Z(g5578) ) ;
OR2     gate3259  (.A(g5227), .B(g669), .Z(g5386) ) ;
INV     gate3260  (.A(g5386), .Z(II7333) ) ;
INV     gate3261  (.A(II7333), .Z(g5579) ) ;
INV     gate3262  (.A(g5534), .Z(II7336) ) ;
INV     gate3263  (.A(g5540), .Z(II7339) ) ;
INV     gate3264  (.A(g5579), .Z(II7342) ) ;
OR2     gate3265  (.A(g5349), .B(g3275), .Z(g5531) ) ;
INV     gate3266  (.A(g5531), .Z(II7346) ) ;
INV     gate3267  (.A(II7346), .Z(g5584) ) ;
OR2     gate3268  (.A(g5350), .B(g3278), .Z(g5532) ) ;
INV     gate3269  (.A(g5532), .Z(II7349) ) ;
INV     gate3270  (.A(II7349), .Z(g5587) ) ;
OR2     gate3271  (.A(g5351), .B(g3290), .Z(g5533) ) ;
INV     gate3272  (.A(g5533), .Z(II7352) ) ;
INV     gate3273  (.A(II7352), .Z(g5590) ) ;
OR2     gate3274  (.A(g5353), .B(g3300), .Z(g5535) ) ;
INV     gate3275  (.A(g5535), .Z(II7355) ) ;
INV     gate3276  (.A(II7355), .Z(g5593) ) ;
NAND2   gate3277  (.A(II7312), .B(II7313), .Z(g5565) ) ;
INV     gate3278  (.A(g5565), .Z(II7358) ) ;
INV     gate3279  (.A(II7358), .Z(g5596) ) ;
INV     gate3280  (.A(g5566), .Z(II7361) ) ;
INV     gate3281  (.A(II7361), .Z(g5597) ) ;
INV     gate3282  (.A(g5493), .Z(II7372) ) ;
INV     gate3283  (.A(II7372), .Z(g5615) ) ;
INV     gate3284  (.A(g5536), .Z(g5631) ) ;
NOR4    gate3285  (.A(g5391), .B(g1589), .C(g3793), .D(g1880), .Z(g5561) ) ;
INV     gate3286  (.A(g5561), .Z(II7397) ) ;
INV     gate3287  (.A(II7397), .Z(g5638) ) ;
INV     gate3288  (.A(g5537), .Z(g5645) ) ;
INV     gate3289  (.A(g5509), .Z(g5647) ) ;
NOR2    gate3290  (.A(g5388), .B(g1880), .Z(g5541) ) ;
INV     gate3291  (.A(g5541), .Z(II7404) ) ;
INV     gate3292  (.A(II7404), .Z(g5649) ) ;
INV     gate3293  (.A(g5512), .Z(g5658) ) ;
INV     gate3294  (.A(g5518), .Z(g5661) ) ;
INV     gate3295  (.A(g5521), .Z(g5664) ) ;
INV     gate3296  (.A(g5524), .Z(g5667) ) ;
INV     gate3297  (.A(g5527), .Z(g5670) ) ;
NOR2    gate3298  (.A(g5354), .B(g5356), .Z(g5552) ) ;
INV     gate3299  (.A(g5552), .Z(g5685) ) ;
INV     gate3300  (.A(g5567), .Z(g5687) ) ;
INV     gate3301  (.A(g5568), .Z(g5691) ) ;
INV     gate3302  (.A(g5597), .Z(II7451) ) ;
OR2     gate3303  (.A(g5492), .B(g3277), .Z(g5622) ) ;
INV     gate3304  (.A(g5622), .Z(II7463) ) ;
INV     gate3305  (.A(II7463), .Z(g5702) ) ;
OR2     gate3306  (.A(g5494), .B(g3280), .Z(g5624) ) ;
INV     gate3307  (.A(g5624), .Z(II7466) ) ;
INV     gate3308  (.A(II7466), .Z(g5705) ) ;
OR2     gate3309  (.A(g5495), .B(g3281), .Z(g5625) ) ;
INV     gate3310  (.A(g5625), .Z(II7469) ) ;
INV     gate3311  (.A(II7469), .Z(g5708) ) ;
OR2     gate3312  (.A(g5496), .B(g3285), .Z(g5626) ) ;
INV     gate3313  (.A(g5626), .Z(II7472) ) ;
INV     gate3314  (.A(II7472), .Z(g5711) ) ;
OR2     gate3315  (.A(g5497), .B(g3286), .Z(g5627) ) ;
INV     gate3316  (.A(g5627), .Z(II7475) ) ;
INV     gate3317  (.A(II7475), .Z(g5714) ) ;
OR2     gate3318  (.A(g5498), .B(g3292), .Z(g5628) ) ;
INV     gate3319  (.A(g5628), .Z(II7478) ) ;
INV     gate3320  (.A(II7478), .Z(g5717) ) ;
OR2     gate3321  (.A(g5499), .B(g3298), .Z(g5629) ) ;
INV     gate3322  (.A(g5629), .Z(II7481) ) ;
INV     gate3323  (.A(II7481), .Z(g5720) ) ;
OR2     gate3324  (.A(g5501), .B(g3309), .Z(g5630) ) ;
INV     gate3325  (.A(g5630), .Z(II7484) ) ;
INV     gate3326  (.A(II7484), .Z(g5723) ) ;
NAND2   gate3327  (.A(II7440), .B(II7441), .Z(g5684) ) ;
INV     gate3328  (.A(g5684), .Z(II7487) ) ;
INV     gate3329  (.A(II7487), .Z(g5726) ) ;
OR2     gate3330  (.A(g5569), .B(g4020), .Z(g5583) ) ;
INV     gate3331  (.A(g5583), .Z(II7490) ) ;
INV     gate3332  (.A(II7490), .Z(g5727) ) ;
INV     gate3333  (.A(g5691), .Z(II7494) ) ;
INV     gate3334  (.A(II7494), .Z(g5729) ) ;
INV     gate3335  (.A(g5687), .Z(II7497) ) ;
INV     gate3336  (.A(II7497), .Z(g5730) ) ;
INV     gate3337  (.A(g5596), .Z(II7501) ) ;
INV     gate3338  (.A(II7501), .Z(g5740) ) ;
AND2    gate3339  (.A(g594), .B(g5515), .Z(g5602) ) ;
INV     gate3340  (.A(g5602), .Z(g5741) ) ;
NAND4   gate3341  (.A(g5546), .B(g1017), .C(g1551), .D(g2916), .Z(g5686) ) ;
INV     gate3342  (.A(g5686), .Z(g5742) ) ;
INV     gate3343  (.A(g5584), .Z(II7506) ) ;
INV     gate3344  (.A(II7506), .Z(g5751) ) ;
INV     gate3345  (.A(g5587), .Z(II7509) ) ;
INV     gate3346  (.A(II7509), .Z(g5752) ) ;
INV     gate3347  (.A(g5645), .Z(g5770) ) ;
INV     gate3348  (.A(g5590), .Z(II7514) ) ;
INV     gate3349  (.A(II7514), .Z(g5773) ) ;
INV     gate3350  (.A(g5593), .Z(II7517) ) ;
INV     gate3351  (.A(II7517), .Z(g5774) ) ;
OR2     gate3352  (.A(g3575), .B(g5500), .Z(g5605) ) ;
INV     gate3353  (.A(g5605), .Z(II7583) ) ;
INV     gate3354  (.A(II7583), .Z(g5784) ) ;
INV     gate3355  (.A(g5685), .Z(g5787) ) ;
INV     gate3356  (.A(g5605), .Z(II7587) ) ;
INV     gate3357  (.A(II7587), .Z(g5788) ) ;
INV     gate3358  (.A(g5605), .Z(II7590) ) ;
INV     gate3359  (.A(II7590), .Z(g5791) ) ;
INV     gate3360  (.A(g5605), .Z(II7593) ) ;
INV     gate3361  (.A(II7593), .Z(g5794) ) ;
INV     gate3362  (.A(g5605), .Z(II7596) ) ;
INV     gate3363  (.A(II7596), .Z(g5797) ) ;
INV     gate3364  (.A(g5605), .Z(II7600) ) ;
INV     gate3365  (.A(II7600), .Z(g5801) ) ;
INV     gate3366  (.A(g5605), .Z(II7604) ) ;
INV     gate3367  (.A(II7604), .Z(g5805) ) ;
INV     gate3368  (.A(g5605), .Z(II7608) ) ;
INV     gate3369  (.A(II7608), .Z(g5809) ) ;
INV     gate3370  (.A(g5605), .Z(II7612) ) ;
INV     gate3371  (.A(II7612), .Z(g5813) ) ;
INV     gate3372  (.A(g5631), .Z(g5824) ) ;
NAND2   gate3373  (.A(g5563), .B(g4767), .Z(g5634) ) ;
INV     gate3374  (.A(g5634), .Z(g5860) ) ;
NAND2   gate3375  (.A(g5564), .B(g4769), .Z(g5636) ) ;
INV     gate3376  (.A(g5636), .Z(g5861) ) ;
INV     gate3377  (.A(g5727), .Z(II7634) ) ;
INV     gate3378  (.A(g5751), .Z(II7637) ) ;
INV     gate3379  (.A(g5773), .Z(II7640) ) ;
INV     gate3380  (.A(g5752), .Z(II7643) ) ;
INV     gate3381  (.A(g5774), .Z(II7646) ) ;
INV     gate3382  (.A(g5770), .Z(g5879) ) ;
INV     gate3383  (.A(g5824), .Z(g5880) ) ;
NAND4   gate3384  (.A(g5649), .B(g1529), .C(g1088), .D(g2068), .Z(g5864) ) ;
INV     gate3385  (.A(g5864), .Z(g5884) ) ;
NAND4   gate3386  (.A(g5649), .B(g1088), .C(g1076), .D(g2068), .Z(g5865) ) ;
INV     gate3387  (.A(g5865), .Z(g5885) ) ;
NOR2    gate3388  (.A(g1477), .B(g5688), .Z(g5753) ) ;
INV     gate3389  (.A(g5753), .Z(g5886) ) ;
INV     gate3390  (.A(g5742), .Z(g5887) ) ;
NOR2    gate3391  (.A(g952), .B(g5688), .Z(g5731) ) ;
INV     gate3392  (.A(g5731), .Z(g5888) ) ;
INV     gate3393  (.A(g5742), .Z(g5889) ) ;
INV     gate3394  (.A(g5753), .Z(g5890) ) ;
INV     gate3395  (.A(g5731), .Z(g5891) ) ;
INV     gate3396  (.A(g5742), .Z(g5892) ) ;
INV     gate3397  (.A(g5753), .Z(g5893) ) ;
INV     gate3398  (.A(g5731), .Z(g5894) ) ;
INV     gate3399  (.A(g5742), .Z(g5895) ) ;
INV     gate3400  (.A(g5753), .Z(g5896) ) ;
INV     gate3401  (.A(g5731), .Z(g5897) ) ;
INV     gate3402  (.A(g5753), .Z(g5899) ) ;
INV     gate3403  (.A(g5753), .Z(g5901) ) ;
INV     gate3404  (.A(g5753), .Z(g5903) ) ;
NAND3   gate3405  (.A(g5638), .B(g2053), .C(g1661), .Z(g5852) ) ;
INV     gate3406  (.A(g5852), .Z(g5905) ) ;
INV     gate3407  (.A(g5753), .Z(g5908) ) ;
NAND3   gate3408  (.A(g5638), .B(g2053), .C(g1076), .Z(g5853) ) ;
INV     gate3409  (.A(g5853), .Z(g5912) ) ;
INV     gate3410  (.A(g5726), .Z(II7679) ) ;
INV     gate3411  (.A(II7679), .Z(g5915) ) ;
INV     gate3412  (.A(g5702), .Z(II7683) ) ;
INV     gate3413  (.A(II7683), .Z(g5917) ) ;
INV     gate3414  (.A(g5705), .Z(II7686) ) ;
INV     gate3415  (.A(II7686), .Z(g5918) ) ;
INV     gate3416  (.A(g5708), .Z(II7689) ) ;
INV     gate3417  (.A(II7689), .Z(g5919) ) ;
INV     gate3418  (.A(g5711), .Z(II7692) ) ;
INV     gate3419  (.A(II7692), .Z(g5920) ) ;
INV     gate3420  (.A(g5714), .Z(II7695) ) ;
INV     gate3421  (.A(II7695), .Z(g5921) ) ;
INV     gate3422  (.A(g5717), .Z(II7698) ) ;
INV     gate3423  (.A(II7698), .Z(g5922) ) ;
INV     gate3424  (.A(g5720), .Z(II7701) ) ;
INV     gate3425  (.A(II7701), .Z(g5923) ) ;
INV     gate3426  (.A(g5723), .Z(II7704) ) ;
INV     gate3427  (.A(II7704), .Z(g5924) ) ;
AND2    gate3428  (.A(g5683), .B(g3813), .Z(g5701) ) ;
INV     gate3429  (.A(g5701), .Z(II7707) ) ;
INV     gate3430  (.A(II7707), .Z(g5925) ) ;
INV     gate3431  (.A(g5729), .Z(g5946) ) ;
INV     gate3432  (.A(g5730), .Z(g5950) ) ;
NAND3   gate3433  (.A(g5649), .B(g1529), .C(g2081), .Z(g5866) ) ;
INV     gate3434  (.A(g5866), .Z(g5957) ) ;
NAND4   gate3435  (.A(g5638), .B(g2056), .C(g1666), .D(g1661), .Z(g5818) ) ;
INV     gate3436  (.A(g5818), .Z(g5958) ) ;
NAND4   gate3437  (.A(g5638), .B(g2056), .C(g1076), .D(g1666), .Z(g5821) ) ;
INV     gate3438  (.A(g5821), .Z(g5975) ) ;
NAND3   gate3439  (.A(g5649), .B(g1076), .C(g2081), .Z(g5869) ) ;
INV     gate3440  (.A(g5869), .Z(g5992) ) ;
NAND4   gate3441  (.A(g5649), .B(g1557), .C(g1564), .D(g2113), .Z(g5872) ) ;
INV     gate3442  (.A(g5872), .Z(g5993) ) ;
NAND4   gate3443  (.A(g5649), .B(g1017), .C(g1564), .D(g2113), .Z(g5873) ) ;
INV     gate3444  (.A(g5873), .Z(g5994) ) ;
INV     gate3445  (.A(g5824), .Z(g5995) ) ;
INV     gate3446  (.A(g5824), .Z(g5996) ) ;
NAND4   gate3447  (.A(g5638), .B(g1683), .C(g1552), .D(g2062), .Z(g5854) ) ;
INV     gate3448  (.A(g5854), .Z(g5997) ) ;
INV     gate3449  (.A(g5824), .Z(g6014) ) ;
NAND4   gate3450  (.A(g5638), .B(g1552), .C(g1017), .D(g2062), .Z(g5857) ) ;
INV     gate3451  (.A(g5857), .Z(g6015) ) ;
INV     gate3452  (.A(g5770), .Z(g6032) ) ;
INV     gate3453  (.A(g5824), .Z(g6033) ) ;
INV     gate3454  (.A(g5824), .Z(g6034) ) ;
INV     gate3455  (.A(g5824), .Z(g6035) ) ;
INV     gate3456  (.A(g5824), .Z(g6036) ) ;
INV     gate3457  (.A(g5824), .Z(g6039) ) ;
INV     gate3458  (.A(g5824), .Z(g6040) ) ;
INV     gate3459  (.A(g5824), .Z(g6043) ) ;
INV     gate3460  (.A(g5824), .Z(g6044) ) ;
INV     gate3461  (.A(g5824), .Z(g6048) ) ;
INV     gate3462  (.A(g5824), .Z(g6051) ) ;
INV     gate3463  (.A(g5824), .Z(g6052) ) ;
INV     gate3464  (.A(g5824), .Z(g6057) ) ;
INV     gate3465  (.A(g5824), .Z(g6062) ) ;
INV     gate3466  (.A(g5784), .Z(g6065) ) ;
INV     gate3467  (.A(g5788), .Z(g6067) ) ;
INV     gate3468  (.A(g5791), .Z(g6069) ) ;
INV     gate3469  (.A(g5824), .Z(g6070) ) ;
INV     gate3470  (.A(g5794), .Z(g6074) ) ;
INV     gate3471  (.A(g5797), .Z(g6076) ) ;
INV     gate3472  (.A(g5801), .Z(g6078) ) ;
INV     gate3473  (.A(g5805), .Z(g6080) ) ;
INV     gate3474  (.A(g5809), .Z(g6083) ) ;
INV     gate3475  (.A(g5813), .Z(g6087) ) ;
INV     gate3476  (.A(g5917), .Z(II7796) ) ;
INV     gate3477  (.A(g5918), .Z(II7799) ) ;
INV     gate3478  (.A(g5920), .Z(II7802) ) ;
INV     gate3479  (.A(g5923), .Z(II7805) ) ;
INV     gate3480  (.A(g5919), .Z(II7808) ) ;
INV     gate3481  (.A(g5921), .Z(II7811) ) ;
INV     gate3482  (.A(g5922), .Z(II7814) ) ;
INV     gate3483  (.A(g5924), .Z(II7817) ) ;
INV     gate3484  (.A(g5879), .Z(g6115) ) ;
INV     gate3485  (.A(g5880), .Z(g6117) ) ;
NAND2   gate3486  (.A(g5741), .B(g639), .Z(g5926) ) ;
INV     gate3487  (.A(g5926), .Z(II7829) ) ;
INV     gate3488  (.A(II7829), .Z(g6119) ) ;
NAND2   gate3489  (.A(g5818), .B(g2940), .Z(g5943) ) ;
INV     gate3490  (.A(g5943), .Z(II7832) ) ;
INV     gate3491  (.A(II7832), .Z(g6120) ) ;
INV     gate3492  (.A(g5926), .Z(II7835) ) ;
INV     gate3493  (.A(II7835), .Z(g6121) ) ;
NAND2   gate3494  (.A(g5821), .B(g2944), .Z(g5947) ) ;
INV     gate3495  (.A(g5947), .Z(II7838) ) ;
INV     gate3496  (.A(II7838), .Z(g6122) ) ;
INV     gate3497  (.A(g5993), .Z(II7852) ) ;
INV     gate3498  (.A(II7852), .Z(g6134) ) ;
INV     gate3499  (.A(g5994), .Z(II7856) ) ;
INV     gate3500  (.A(II7856), .Z(g6136) ) ;
INV     gate3501  (.A(g6032), .Z(II7859) ) ;
INV     gate3502  (.A(II7859), .Z(g6137) ) ;
NAND2   gate3503  (.A(g2952), .B(g5854), .Z(g6095) ) ;
INV     gate3504  (.A(g6095), .Z(II7865) ) ;
INV     gate3505  (.A(II7865), .Z(g6143) ) ;
NAND2   gate3506  (.A(g2954), .B(g5857), .Z(g6097) ) ;
INV     gate3507  (.A(g6097), .Z(II7871) ) ;
INV     gate3508  (.A(II7871), .Z(g6147) ) ;
INV     gate3509  (.A(g5926), .Z(g6160) ) ;
INV     gate3510  (.A(g5926), .Z(g6161) ) ;
INV     gate3511  (.A(g5926), .Z(g6162) ) ;
INV     gate3512  (.A(g5926), .Z(g6163) ) ;
INV     gate3513  (.A(g5926), .Z(g6164) ) ;
INV     gate3514  (.A(g5926), .Z(g6165) ) ;
OR2     gate3515  (.A(g5728), .B(g3781), .Z(g5916) ) ;
INV     gate3516  (.A(g5916), .Z(II7892) ) ;
INV     gate3517  (.A(II7892), .Z(g6166) ) ;
INV     gate3518  (.A(g5950), .Z(g6188) ) ;
INV     gate3519  (.A(g5946), .Z(g6192) ) ;
INV     gate3520  (.A(g5957), .Z(g6193) ) ;
INV     gate3521  (.A(g5912), .Z(II7906) ) ;
INV     gate3522  (.A(II7906), .Z(g6194) ) ;
INV     gate3523  (.A(g5992), .Z(g6211) ) ;
INV     gate3524  (.A(g5905), .Z(II7910) ) ;
INV     gate3525  (.A(II7910), .Z(g6212) ) ;
INV     gate3526  (.A(g6036), .Z(g6229) ) ;
INV     gate3527  (.A(g6040), .Z(g6230) ) ;
INV     gate3528  (.A(g6044), .Z(g6231) ) ;
INV     gate3529  (.A(g6048), .Z(g6232) ) ;
INV     gate3530  (.A(g6052), .Z(g6233) ) ;
INV     gate3531  (.A(g6057), .Z(g6234) ) ;
INV     gate3532  (.A(g6062), .Z(g6235) ) ;
INV     gate3533  (.A(g6070), .Z(g6236) ) ;
INV     gate3534  (.A(g5925), .Z(II7960) ) ;
INV     gate3535  (.A(II7960), .Z(g6276) ) ;
INV     gate3536  (.A(g6276), .Z(II7963) ) ;
INV     gate3537  (.A(g6166), .Z(II7966) ) ;
INV     gate3538  (.A(g6137), .Z(II7996) ) ;
INV     gate3539  (.A(g6137), .Z(II7999) ) ;
INV     gate3540  (.A(II7999), .Z(g6283) ) ;
OR2     gate3541  (.A(g5883), .B(g5996), .Z(g6110) ) ;
INV     gate3542  (.A(g6110), .Z(II8002) ) ;
INV     gate3543  (.A(g6110), .Z(II8005) ) ;
INV     gate3544  (.A(II8005), .Z(g6285) ) ;
OR2     gate3545  (.A(g5912), .B(g2381), .Z(g6237) ) ;
INV     gate3546  (.A(g6237), .Z(II8027) ) ;
INV     gate3547  (.A(II8027), .Z(g6305) ) ;
OR2     gate3548  (.A(g2339), .B(g6073), .Z(g6239) ) ;
INV     gate3549  (.A(g6239), .Z(II8030) ) ;
INV     gate3550  (.A(II8030), .Z(g6306) ) ;
OR2     gate3551  (.A(g2356), .B(g6075), .Z(g6242) ) ;
INV     gate3552  (.A(g6242), .Z(II8034) ) ;
INV     gate3553  (.A(II8034), .Z(g6308) ) ;
OR2     gate3554  (.A(g5909), .B(g3806), .Z(g6142) ) ;
INV     gate3555  (.A(g6142), .Z(II8040) ) ;
INV     gate3556  (.A(II8040), .Z(g6312) ) ;
OR2     gate3557  (.A(g5905), .B(g2381), .Z(g6252) ) ;
INV     gate3558  (.A(g6252), .Z(II8044) ) ;
INV     gate3559  (.A(II8044), .Z(g6314) ) ;
OR2     gate3560  (.A(g5898), .B(g5598), .Z(g6108) ) ;
INV     gate3561  (.A(g6108), .Z(II8051) ) ;
INV     gate3562  (.A(II8051), .Z(g6319) ) ;
OR2     gate3563  (.A(g5900), .B(g5599), .Z(g6109) ) ;
INV     gate3564  (.A(g6109), .Z(II8056) ) ;
INV     gate3565  (.A(II8056), .Z(g6322) ) ;
OR2     gate3566  (.A(g5902), .B(g5601), .Z(g6113) ) ;
INV     gate3567  (.A(g6113), .Z(II8061) ) ;
INV     gate3568  (.A(II8061), .Z(g6325) ) ;
OR2     gate3569  (.A(g5904), .B(g5604), .Z(g6114) ) ;
INV     gate3570  (.A(g6114), .Z(II8066) ) ;
INV     gate3571  (.A(II8066), .Z(g6328) ) ;
OR2     gate3572  (.A(g5910), .B(g5617), .Z(g6116) ) ;
INV     gate3573  (.A(g6116), .Z(II8070) ) ;
INV     gate3574  (.A(II8070), .Z(g6330) ) ;
OR2     gate3575  (.A(g5911), .B(g5619), .Z(g6118) ) ;
INV     gate3576  (.A(g6118), .Z(II8074) ) ;
INV     gate3577  (.A(II8074), .Z(g6332) ) ;
INV     gate3578  (.A(g6120), .Z(II8089) ) ;
INV     gate3579  (.A(II8089), .Z(g6337) ) ;
INV     gate3580  (.A(g6122), .Z(II8093) ) ;
INV     gate3581  (.A(II8093), .Z(g6339) ) ;
INV     gate3582  (.A(g6134), .Z(II8103) ) ;
INV     gate3583  (.A(II8103), .Z(g6347) ) ;
INV     gate3584  (.A(g6136), .Z(II8107) ) ;
INV     gate3585  (.A(II8107), .Z(g6351) ) ;
INV     gate3586  (.A(g6143), .Z(II8110) ) ;
INV     gate3587  (.A(II8110), .Z(g6352) ) ;
INV     gate3588  (.A(g6147), .Z(II8113) ) ;
INV     gate3589  (.A(II8113), .Z(g6353) ) ;
OR2     gate3590  (.A(g6047), .B(g6034), .Z(g6182) ) ;
INV     gate3591  (.A(g6182), .Z(II8144) ) ;
INV     gate3592  (.A(g6182), .Z(II8147) ) ;
INV     gate3593  (.A(II8147), .Z(g6361) ) ;
OR2     gate3594  (.A(g6055), .B(g5995), .Z(g6185) ) ;
INV     gate3595  (.A(g6185), .Z(II8150) ) ;
INV     gate3596  (.A(g6185), .Z(II8153) ) ;
INV     gate3597  (.A(II8153), .Z(g6363) ) ;
OR2     gate3598  (.A(g6056), .B(g6039), .Z(g6167) ) ;
INV     gate3599  (.A(g6167), .Z(II8156) ) ;
INV     gate3600  (.A(g6167), .Z(II8159) ) ;
INV     gate3601  (.A(II8159), .Z(g6365) ) ;
OR2     gate3602  (.A(g6060), .B(g6035), .Z(g6189) ) ;
INV     gate3603  (.A(g6189), .Z(II8162) ) ;
INV     gate3604  (.A(g6189), .Z(II8165) ) ;
INV     gate3605  (.A(II8165), .Z(g6367) ) ;
OR2     gate3606  (.A(g6061), .B(g6014), .Z(g6170) ) ;
INV     gate3607  (.A(g6170), .Z(II8168) ) ;
INV     gate3608  (.A(g6170), .Z(II8171) ) ;
INV     gate3609  (.A(II8171), .Z(g6369) ) ;
OR2     gate3610  (.A(g6066), .B(g6043), .Z(g6173) ) ;
INV     gate3611  (.A(g6173), .Z(II8174) ) ;
INV     gate3612  (.A(g6173), .Z(II8177) ) ;
INV     gate3613  (.A(II8177), .Z(g6371) ) ;
OR2     gate3614  (.A(g6068), .B(g6033), .Z(g6176) ) ;
INV     gate3615  (.A(g6176), .Z(II8180) ) ;
INV     gate3616  (.A(g6176), .Z(II8183) ) ;
INV     gate3617  (.A(II8183), .Z(g6373) ) ;
OR2     gate3618  (.A(g6077), .B(g6051), .Z(g6179) ) ;
INV     gate3619  (.A(g6179), .Z(II8186) ) ;
INV     gate3620  (.A(g6179), .Z(II8189) ) ;
INV     gate3621  (.A(II8189), .Z(g6375) ) ;
OR2     gate3622  (.A(g2953), .B(g5884), .Z(g6267) ) ;
INV     gate3623  (.A(g6267), .Z(g6376) ) ;
OR2     gate3624  (.A(g2955), .B(g5885), .Z(g6271) ) ;
INV     gate3625  (.A(g6271), .Z(g6385) ) ;
INV     gate3626  (.A(g6319), .Z(II8217) ) ;
INV     gate3627  (.A(g6322), .Z(II8220) ) ;
INV     gate3628  (.A(g6325), .Z(II8223) ) ;
INV     gate3629  (.A(g6328), .Z(II8226) ) ;
INV     gate3630  (.A(g6330), .Z(II8229) ) ;
INV     gate3631  (.A(g6332), .Z(II8232) ) ;
INV     gate3632  (.A(g6312), .Z(II8235) ) ;
INV     gate3633  (.A(g6283), .Z(g6408) ) ;
INV     gate3634  (.A(g6285), .Z(g6409) ) ;
OR2     gate3635  (.A(g6241), .B(g6082), .Z(g6287) ) ;
INV     gate3636  (.A(g6287), .Z(II8240) ) ;
INV     gate3637  (.A(II8240), .Z(g6410) ) ;
OR2     gate3638  (.A(g6238), .B(g6079), .Z(g6286) ) ;
INV     gate3639  (.A(g6286), .Z(II8243) ) ;
INV     gate3640  (.A(II8243), .Z(g6411) ) ;
OR2     gate3641  (.A(g6245), .B(g6086), .Z(g6290) ) ;
INV     gate3642  (.A(g6290), .Z(II8246) ) ;
INV     gate3643  (.A(II8246), .Z(g6412) ) ;
OR2     gate3644  (.A(g6240), .B(g6081), .Z(g6289) ) ;
INV     gate3645  (.A(g6289), .Z(II8249) ) ;
INV     gate3646  (.A(II8249), .Z(g6413) ) ;
OR2     gate3647  (.A(g6249), .B(g6090), .Z(g6294) ) ;
INV     gate3648  (.A(g6294), .Z(II8252) ) ;
INV     gate3649  (.A(II8252), .Z(g6414) ) ;
OR2     gate3650  (.A(g6243), .B(g6084), .Z(g6292) ) ;
INV     gate3651  (.A(g6292), .Z(II8255) ) ;
INV     gate3652  (.A(II8255), .Z(g6415) ) ;
OR2     gate3653  (.A(g6244), .B(g6085), .Z(g6293) ) ;
INV     gate3654  (.A(g6293), .Z(II8258) ) ;
INV     gate3655  (.A(II8258), .Z(g6416) ) ;
OR2     gate3656  (.A(g6255), .B(g6093), .Z(g6298) ) ;
INV     gate3657  (.A(g6298), .Z(II8261) ) ;
INV     gate3658  (.A(II8261), .Z(g6417) ) ;
OR2     gate3659  (.A(g6247), .B(g6088), .Z(g6296) ) ;
INV     gate3660  (.A(g6296), .Z(II8264) ) ;
INV     gate3661  (.A(II8264), .Z(g6418) ) ;
OR2     gate3662  (.A(g6248), .B(g6089), .Z(g6297) ) ;
INV     gate3663  (.A(g6297), .Z(II8267) ) ;
INV     gate3664  (.A(II8267), .Z(g6419) ) ;
OR2     gate3665  (.A(g6253), .B(g6091), .Z(g6300) ) ;
INV     gate3666  (.A(g6300), .Z(II8270) ) ;
INV     gate3667  (.A(II8270), .Z(g6420) ) ;
OR2     gate3668  (.A(g6254), .B(g6092), .Z(g6301) ) ;
INV     gate3669  (.A(g6301), .Z(II8273) ) ;
INV     gate3670  (.A(II8273), .Z(g6421) ) ;
OR2     gate3671  (.A(g6258), .B(g6094), .Z(g6303) ) ;
INV     gate3672  (.A(g6303), .Z(II8276) ) ;
INV     gate3673  (.A(II8276), .Z(g6422) ) ;
OR2     gate3674  (.A(g6262), .B(g6096), .Z(g6307) ) ;
INV     gate3675  (.A(g6307), .Z(II8279) ) ;
INV     gate3676  (.A(II8279), .Z(g6423) ) ;
OR2     gate3677  (.A(g6265), .B(g6098), .Z(g6309) ) ;
INV     gate3678  (.A(g6309), .Z(II8282) ) ;
INV     gate3679  (.A(II8282), .Z(g6424) ) ;
OR2     gate3680  (.A(g6269), .B(g6099), .Z(g6310) ) ;
INV     gate3681  (.A(g6310), .Z(II8285) ) ;
INV     gate3682  (.A(II8285), .Z(g6425) ) ;
AND2    gate3683  (.A(g5210), .B(g6161), .Z(g6291) ) ;
INV     gate3684  (.A(g6291), .Z(II8290) ) ;
INV     gate3685  (.A(II8290), .Z(g6428) ) ;
AND2    gate3686  (.A(g5379), .B(g6162), .Z(g6295) ) ;
INV     gate3687  (.A(g6295), .Z(II8295) ) ;
INV     gate3688  (.A(II8295), .Z(g6431) ) ;
AND2    gate3689  (.A(g5530), .B(g6163), .Z(g6299) ) ;
INV     gate3690  (.A(g6299), .Z(II8300) ) ;
INV     gate3691  (.A(II8300), .Z(g6434) ) ;
AND2    gate3692  (.A(g5915), .B(g6165), .Z(g6304) ) ;
INV     gate3693  (.A(g6304), .Z(II8309) ) ;
INV     gate3694  (.A(II8309), .Z(g6441) ) ;
INV     gate3695  (.A(g6305), .Z(II8329) ) ;
INV     gate3696  (.A(II8329), .Z(g6465) ) ;
INV     gate3697  (.A(g6306), .Z(II8332) ) ;
INV     gate3698  (.A(II8332), .Z(g6466) ) ;
INV     gate3699  (.A(g6308), .Z(II8335) ) ;
INV     gate3700  (.A(II8335), .Z(g6467) ) ;
INV     gate3701  (.A(g6314), .Z(II8342) ) ;
INV     gate3702  (.A(II8342), .Z(g6478) ) ;
INV     gate3703  (.A(g6361), .Z(g6484) ) ;
INV     gate3704  (.A(g6363), .Z(g6486) ) ;
INV     gate3705  (.A(g6365), .Z(g6487) ) ;
INV     gate3706  (.A(g6367), .Z(g6488) ) ;
INV     gate3707  (.A(g6369), .Z(g6489) ) ;
INV     gate3708  (.A(g6371), .Z(g6490) ) ;
INV     gate3709  (.A(g6373), .Z(g6491) ) ;
INV     gate3710  (.A(g6375), .Z(g6493) ) ;
INV     gate3711  (.A(g6415), .Z(II8411) ) ;
INV     gate3712  (.A(g6418), .Z(II8414) ) ;
INV     gate3713  (.A(g6420), .Z(II8417) ) ;
INV     gate3714  (.A(g6422), .Z(II8420) ) ;
INV     gate3715  (.A(g6423), .Z(II8423) ) ;
INV     gate3716  (.A(g6424), .Z(II8426) ) ;
INV     gate3717  (.A(g6425), .Z(II8429) ) ;
INV     gate3718  (.A(g6411), .Z(II8432) ) ;
INV     gate3719  (.A(g6413), .Z(II8435) ) ;
INV     gate3720  (.A(g6416), .Z(II8438) ) ;
INV     gate3721  (.A(g6419), .Z(II8441) ) ;
INV     gate3722  (.A(g6421), .Z(II8444) ) ;
INV     gate3723  (.A(g6410), .Z(II8447) ) ;
INV     gate3724  (.A(g6412), .Z(II8450) ) ;
INV     gate3725  (.A(g6414), .Z(II8453) ) ;
INV     gate3726  (.A(g6417), .Z(II8456) ) ;
NOR4    gate3727  (.A(g6376), .B(g4086), .C(g4074), .D(g4068), .Z(g6427) ) ;
INV     gate3728  (.A(g6427), .Z(II8459) ) ;
INV     gate3729  (.A(II8459), .Z(g6513) ) ;
NOR4    gate3730  (.A(g6385), .B(g3733), .C(g4092), .D(g4080), .Z(g6430) ) ;
INV     gate3731  (.A(g6430), .Z(II8462) ) ;
INV     gate3732  (.A(II8462), .Z(g6514) ) ;
INV     gate3733  (.A(g6408), .Z(g6515) ) ;
INV     gate3734  (.A(g6409), .Z(g6516) ) ;
OR2     gate3735  (.A(g6352), .B(g6347), .Z(g6457) ) ;
INV     gate3736  (.A(g6457), .Z(II8467) ) ;
INV     gate3737  (.A(II8467), .Z(g6517) ) ;
OR2     gate3738  (.A(g6353), .B(g6351), .Z(g6461) ) ;
INV     gate3739  (.A(g6461), .Z(II8470) ) ;
INV     gate3740  (.A(II8470), .Z(g6518) ) ;
OR3     gate3741  (.A(II8393), .B(II8394), .C(II8395), .Z(g6485) ) ;
INV     gate3742  (.A(g6485), .Z(II8473) ) ;
INV     gate3743  (.A(II8473), .Z(g6519) ) ;
INV     gate3744  (.A(g6457), .Z(II8476) ) ;
INV     gate3745  (.A(II8476), .Z(g6520) ) ;
OR4     gate3746  (.A(II8376), .B(II8377), .C(II8378), .D(II8379), .Z(g6482) ) ;
INV     gate3747  (.A(g6482), .Z(II8479) ) ;
INV     gate3748  (.A(II8479), .Z(g6521) ) ;
INV     gate3749  (.A(g6461), .Z(II8482) ) ;
INV     gate3750  (.A(II8482), .Z(g6522) ) ;
OR2     gate3751  (.A(II8349), .B(g6335), .Z(g6479) ) ;
INV     gate3752  (.A(g6479), .Z(II8485) ) ;
INV     gate3753  (.A(II8485), .Z(g6523) ) ;
OR2     gate3754  (.A(g6288), .B(g6119), .Z(g6426) ) ;
INV     gate3755  (.A(g6426), .Z(II8488) ) ;
INV     gate3756  (.A(II8488), .Z(g6524) ) ;
OR2     gate3757  (.A(II8360), .B(g6359), .Z(g6480) ) ;
INV     gate3758  (.A(g6480), .Z(II8491) ) ;
INV     gate3759  (.A(II8491), .Z(g6525) ) ;
INV     gate3760  (.A(g6428), .Z(II8494) ) ;
INV     gate3761  (.A(II8494), .Z(g6526) ) ;
OR4     gate3762  (.A(II8367), .B(II8368), .C(II8369), .D(II8370), .Z(g6481) ) ;
INV     gate3763  (.A(g6481), .Z(II8497) ) ;
INV     gate3764  (.A(II8497), .Z(g6527) ) ;
INV     gate3765  (.A(g6431), .Z(II8500) ) ;
INV     gate3766  (.A(II8500), .Z(g6528) ) ;
INV     gate3767  (.A(g6434), .Z(II8503) ) ;
INV     gate3768  (.A(II8503), .Z(g6529) ) ;
OR3     gate3769  (.A(II8385), .B(II8386), .C(II8387), .Z(g6483) ) ;
INV     gate3770  (.A(g6483), .Z(II8506) ) ;
INV     gate3771  (.A(II8506), .Z(g6530) ) ;
OR2     gate3772  (.A(g6302), .B(g6121), .Z(g6437) ) ;
INV     gate3773  (.A(g6437), .Z(II8509) ) ;
INV     gate3774  (.A(II8509), .Z(g6531) ) ;
INV     gate3775  (.A(g6441), .Z(II8512) ) ;
INV     gate3776  (.A(II8512), .Z(g6532) ) ;
NOR2    gate3777  (.A(g6348), .B(g1734), .Z(g6492) ) ;
INV     gate3778  (.A(g6492), .Z(II8515) ) ;
INV     gate3779  (.A(II8515), .Z(g6533) ) ;
NOR2    gate3780  (.A(g952), .B(g6348), .Z(g6494) ) ;
INV     gate3781  (.A(g6494), .Z(II8518) ) ;
INV     gate3782  (.A(II8518), .Z(g6534) ) ;
NOR2    gate3783  (.A(g6354), .B(g1775), .Z(g6495) ) ;
INV     gate3784  (.A(g6495), .Z(II8521) ) ;
INV     gate3785  (.A(II8521), .Z(g6535) ) ;
NOR2    gate3786  (.A(g952), .B(g6354), .Z(g6496) ) ;
INV     gate3787  (.A(g6496), .Z(II8524) ) ;
INV     gate3788  (.A(II8524), .Z(g6536) ) ;
OR2     gate3789  (.A(g6336), .B(g5935), .Z(g6440) ) ;
INV     gate3790  (.A(g6440), .Z(II8527) ) ;
INV     gate3791  (.A(II8527), .Z(g6537) ) ;
AND3    gate3792  (.A(g2121), .B(g2032), .C(g6394), .Z(g6469) ) ;
INV     gate3793  (.A(g6469), .Z(g6538) ) ;
OR2     gate3794  (.A(g6338), .B(g5936), .Z(g6444) ) ;
INV     gate3795  (.A(g6444), .Z(II8531) ) ;
INV     gate3796  (.A(II8531), .Z(g6539) ) ;
AND3    gate3797  (.A(g2138), .B(g2036), .C(g6397), .Z(g6474) ) ;
INV     gate3798  (.A(g6474), .Z(g6540) ) ;
OR2     gate3799  (.A(g6340), .B(g5938), .Z(g6447) ) ;
INV     gate3800  (.A(g6447), .Z(II8535) ) ;
INV     gate3801  (.A(II8535), .Z(g6541) ) ;
OR2     gate3802  (.A(g6341), .B(g5940), .Z(g6450) ) ;
INV     gate3803  (.A(g6450), .Z(II8538) ) ;
INV     gate3804  (.A(II8538), .Z(g6542) ) ;
OR2     gate3805  (.A(g6342), .B(g5942), .Z(g6452) ) ;
INV     gate3806  (.A(g6452), .Z(II8541) ) ;
INV     gate3807  (.A(II8541), .Z(g6543) ) ;
OR2     gate3808  (.A(g6343), .B(g5945), .Z(g6453) ) ;
INV     gate3809  (.A(g6453), .Z(II8544) ) ;
INV     gate3810  (.A(II8544), .Z(g6544) ) ;
OR2     gate3811  (.A(g6344), .B(g5949), .Z(g6454) ) ;
INV     gate3812  (.A(g6454), .Z(II8548) ) ;
INV     gate3813  (.A(II8548), .Z(g6548) ) ;
OR2     gate3814  (.A(g6345), .B(g5952), .Z(g6455) ) ;
INV     gate3815  (.A(g6455), .Z(II8552) ) ;
INV     gate3816  (.A(II8552), .Z(g6552) ) ;
OR2     gate3817  (.A(g6346), .B(g5954), .Z(g6456) ) ;
INV     gate3818  (.A(g6456), .Z(II8555) ) ;
INV     gate3819  (.A(II8555), .Z(g6553) ) ;
NOR4    gate3820  (.A(g6376), .B(g4086), .C(g4074), .D(g4302), .Z(g6429) ) ;
INV     gate3821  (.A(g6429), .Z(II8564) ) ;
INV     gate3822  (.A(II8564), .Z(g6560) ) ;
NOR4    gate3823  (.A(g6376), .B(g4086), .C(g4309), .D(g4068), .Z(g6432) ) ;
INV     gate3824  (.A(g6432), .Z(II8567) ) ;
INV     gate3825  (.A(II8567), .Z(g6561) ) ;
NOR4    gate3826  (.A(g6385), .B(g3733), .C(g4092), .D(g4314), .Z(g6433) ) ;
INV     gate3827  (.A(g6433), .Z(II8570) ) ;
INV     gate3828  (.A(II8570), .Z(g6562) ) ;
NOR4    gate3829  (.A(g6376), .B(g4086), .C(g4309), .D(g4302), .Z(g6435) ) ;
INV     gate3830  (.A(g6435), .Z(II8573) ) ;
INV     gate3831  (.A(II8573), .Z(g6563) ) ;
NOR4    gate3832  (.A(g6385), .B(g3733), .C(g4328), .D(g4080), .Z(g6436) ) ;
INV     gate3833  (.A(g6436), .Z(II8576) ) ;
INV     gate3834  (.A(II8576), .Z(g6564) ) ;
NOR4    gate3835  (.A(g6376), .B(g4323), .C(g4074), .D(g4068), .Z(g6438) ) ;
INV     gate3836  (.A(g6438), .Z(II8579) ) ;
INV     gate3837  (.A(II8579), .Z(g6565) ) ;
NOR4    gate3838  (.A(g6385), .B(g3733), .C(g4328), .D(g4314), .Z(g6439) ) ;
INV     gate3839  (.A(g6439), .Z(II8582) ) ;
INV     gate3840  (.A(II8582), .Z(g6566) ) ;
NOR4    gate3841  (.A(g6376), .B(g4323), .C(g4074), .D(g4302), .Z(g6442) ) ;
INV     gate3842  (.A(g6442), .Z(II8585) ) ;
INV     gate3843  (.A(II8585), .Z(g6567) ) ;
NOR4    gate3844  (.A(g6385), .B(g4334), .C(g4092), .D(g4080), .Z(g6443) ) ;
INV     gate3845  (.A(g6443), .Z(II8588) ) ;
INV     gate3846  (.A(II8588), .Z(g6568) ) ;
NOR4    gate3847  (.A(g6376), .B(g4323), .C(g4309), .D(g4302), .Z(g6448) ) ;
INV     gate3848  (.A(g6448), .Z(II8591) ) ;
INV     gate3849  (.A(II8591), .Z(g6569) ) ;
NOR4    gate3850  (.A(g6385), .B(g4334), .C(g4092), .D(g4314), .Z(g6446) ) ;
INV     gate3851  (.A(g6446), .Z(II8594) ) ;
INV     gate3852  (.A(II8594), .Z(g6570) ) ;
NOR4    gate3853  (.A(g6376), .B(g4323), .C(g4309), .D(g4068), .Z(g6445) ) ;
INV     gate3854  (.A(g6445), .Z(II8597) ) ;
INV     gate3855  (.A(II8597), .Z(g6571) ) ;
NOR4    gate3856  (.A(g6385), .B(g4334), .C(g4328), .D(g4314), .Z(g6451) ) ;
INV     gate3857  (.A(g6451), .Z(II8600) ) ;
INV     gate3858  (.A(II8600), .Z(g6572) ) ;
NOR4    gate3859  (.A(g6385), .B(g4334), .C(g4328), .D(g4080), .Z(g6449) ) ;
INV     gate3860  (.A(g6449), .Z(II8603) ) ;
INV     gate3861  (.A(II8603), .Z(g6573) ) ;
INV     gate3862  (.A(g6484), .Z(g6574) ) ;
INV     gate3863  (.A(g6486), .Z(g6575) ) ;
INV     gate3864  (.A(g6487), .Z(g6576) ) ;
INV     gate3865  (.A(g6488), .Z(g6577) ) ;
INV     gate3866  (.A(g6489), .Z(g6578) ) ;
INV     gate3867  (.A(g6490), .Z(g6579) ) ;
INV     gate3868  (.A(g6491), .Z(g6580) ) ;
INV     gate3869  (.A(g6493), .Z(g6581) ) ;
INV     gate3870  (.A(g6537), .Z(II8614) ) ;
INV     gate3871  (.A(g6539), .Z(II8617) ) ;
INV     gate3872  (.A(g6541), .Z(II8620) ) ;
INV     gate3873  (.A(g6542), .Z(II8623) ) ;
INV     gate3874  (.A(g6543), .Z(II8626) ) ;
INV     gate3875  (.A(g6544), .Z(II8629) ) ;
INV     gate3876  (.A(g6548), .Z(II8632) ) ;
INV     gate3877  (.A(g6552), .Z(II8635) ) ;
INV     gate3878  (.A(g6553), .Z(II8638) ) ;
INV     gate3879  (.A(g6524), .Z(II8641) ) ;
INV     gate3880  (.A(g6526), .Z(II8644) ) ;
INV     gate3881  (.A(g6528), .Z(II8647) ) ;
INV     gate3882  (.A(g6529), .Z(II8650) ) ;
INV     gate3883  (.A(g6531), .Z(II8653) ) ;
INV     gate3884  (.A(g6532), .Z(II8656) ) ;
INV     gate3885  (.A(g6523), .Z(II8659) ) ;
INV     gate3886  (.A(g6525), .Z(II8662) ) ;
INV     gate3887  (.A(g6527), .Z(II8665) ) ;
INV     gate3888  (.A(g6530), .Z(II8668) ) ;
INV     gate3889  (.A(g6519), .Z(II8671) ) ;
INV     gate3890  (.A(g6521), .Z(II8674) ) ;
INV     gate3891  (.A(g6565), .Z(II8678) ) ;
INV     gate3892  (.A(II8678), .Z(g6604) ) ;
INV     gate3893  (.A(g6566), .Z(II8681) ) ;
INV     gate3894  (.A(II8681), .Z(g6605) ) ;
INV     gate3895  (.A(g6567), .Z(II8684) ) ;
INV     gate3896  (.A(II8684), .Z(g6606) ) ;
INV     gate3897  (.A(g6568), .Z(II8687) ) ;
INV     gate3898  (.A(II8687), .Z(g6607) ) ;
INV     gate3899  (.A(g6571), .Z(II8690) ) ;
INV     gate3900  (.A(II8690), .Z(g6608) ) ;
INV     gate3901  (.A(g6570), .Z(II8693) ) ;
INV     gate3902  (.A(II8693), .Z(g6609) ) ;
INV     gate3903  (.A(g6569), .Z(II8696) ) ;
INV     gate3904  (.A(II8696), .Z(g6610) ) ;
INV     gate3905  (.A(g6573), .Z(II8699) ) ;
INV     gate3906  (.A(II8699), .Z(g6611) ) ;
INV     gate3907  (.A(g6572), .Z(II8702) ) ;
INV     gate3908  (.A(II8702), .Z(g6612) ) ;
INV     gate3909  (.A(g6520), .Z(II8707) ) ;
INV     gate3910  (.A(II8707), .Z(g6615) ) ;
INV     gate3911  (.A(g6517), .Z(II8710) ) ;
INV     gate3912  (.A(II8710), .Z(g6616) ) ;
INV     gate3913  (.A(g6522), .Z(II8713) ) ;
INV     gate3914  (.A(II8713), .Z(g6617) ) ;
INV     gate3915  (.A(g6518), .Z(II8716) ) ;
INV     gate3916  (.A(II8716), .Z(g6618) ) ;
INV     gate3917  (.A(g6534), .Z(II8721) ) ;
INV     gate3918  (.A(II8721), .Z(g6621) ) ;
INV     gate3919  (.A(g6533), .Z(II8724) ) ;
INV     gate3920  (.A(II8724), .Z(g6622) ) ;
INV     gate3921  (.A(g6536), .Z(II8727) ) ;
INV     gate3922  (.A(II8727), .Z(g6623) ) ;
INV     gate3923  (.A(g6535), .Z(II8730) ) ;
INV     gate3924  (.A(II8730), .Z(g6624) ) ;
INV     gate3925  (.A(g6513), .Z(II8745) ) ;
INV     gate3926  (.A(II8745), .Z(g6649) ) ;
INV     gate3927  (.A(g6560), .Z(II8749) ) ;
INV     gate3928  (.A(II8749), .Z(g6651) ) ;
INV     gate3929  (.A(g6514), .Z(II8752) ) ;
INV     gate3930  (.A(II8752), .Z(g6652) ) ;
INV     gate3931  (.A(g6561), .Z(II8755) ) ;
INV     gate3932  (.A(II8755), .Z(g6653) ) ;
INV     gate3933  (.A(g6562), .Z(II8758) ) ;
INV     gate3934  (.A(II8758), .Z(g6654) ) ;
INV     gate3935  (.A(g6563), .Z(II8761) ) ;
INV     gate3936  (.A(II8761), .Z(g6655) ) ;
INV     gate3937  (.A(g6564), .Z(II8764) ) ;
INV     gate3938  (.A(II8764), .Z(g6656) ) ;
AND2    gate3939  (.A(g6515), .B(g6115), .Z(g6619) ) ;
INV     gate3940  (.A(g6619), .Z(II8767) ) ;
INV     gate3941  (.A(II8767), .Z(g6657) ) ;
OR2     gate3942  (.A(g6250), .B(g6643), .Z(g6684) ) ;
INV     gate3943  (.A(g6684), .Z(II8800) ) ;
INV     gate3944  (.A(II8800), .Z(g6694) ) ;
OR2     gate3945  (.A(g6256), .B(g6644), .Z(g6685) ) ;
INV     gate3946  (.A(g6685), .Z(II8803) ) ;
INV     gate3947  (.A(II8803), .Z(g6695) ) ;
OR2     gate3948  (.A(g6259), .B(g6645), .Z(g6686) ) ;
INV     gate3949  (.A(g6686), .Z(II8806) ) ;
INV     gate3950  (.A(II8806), .Z(g6696) ) ;
OR2     gate3951  (.A(g6260), .B(g6646), .Z(g6687) ) ;
INV     gate3952  (.A(g6687), .Z(II8809) ) ;
INV     gate3953  (.A(II8809), .Z(g6697) ) ;
OR2     gate3954  (.A(g6263), .B(g6647), .Z(g6688) ) ;
INV     gate3955  (.A(g6688), .Z(II8812) ) ;
INV     gate3956  (.A(II8812), .Z(g6698) ) ;
OR2     gate3957  (.A(g6266), .B(g6648), .Z(g6689) ) ;
INV     gate3958  (.A(g6689), .Z(II8815) ) ;
INV     gate3959  (.A(II8815), .Z(g6699) ) ;
OR2     gate3960  (.A(g6270), .B(g6650), .Z(g6690) ) ;
INV     gate3961  (.A(g6690), .Z(II8818) ) ;
INV     gate3962  (.A(II8818), .Z(g6700) ) ;
OR2     gate3963  (.A(g6275), .B(g6603), .Z(g6691) ) ;
INV     gate3964  (.A(g6691), .Z(II8821) ) ;
INV     gate3965  (.A(II8821), .Z(g6701) ) ;
OR2     gate3966  (.A(II8773), .B(II8774), .Z(g6661) ) ;
INV     gate3967  (.A(g6661), .Z(II8828) ) ;
INV     gate3968  (.A(II8828), .Z(g6706) ) ;
OR2     gate3969  (.A(II8778), .B(II8779), .Z(g6665) ) ;
INV     gate3970  (.A(g6665), .Z(II8831) ) ;
INV     gate3971  (.A(II8831), .Z(g6707) ) ;
INV     gate3972  (.A(g6661), .Z(II8834) ) ;
INV     gate3973  (.A(II8834), .Z(g6708) ) ;
INV     gate3974  (.A(g6665), .Z(II8837) ) ;
INV     gate3975  (.A(II8837), .Z(g6709) ) ;
INV     gate3976  (.A(g6657), .Z(II8840) ) ;
INV     gate3977  (.A(II8840), .Z(g6710) ) ;
OR2     gate3978  (.A(g6132), .B(g6620), .Z(g6658) ) ;
INV     gate3979  (.A(g6658), .Z(II8843) ) ;
INV     gate3980  (.A(II8843), .Z(g6711) ) ;
OR2     gate3981  (.A(g6631), .B(g6555), .Z(g6676) ) ;
INV     gate3982  (.A(g6676), .Z(g6712) ) ;
OR2     gate3983  (.A(g6637), .B(g6558), .Z(g6679) ) ;
INV     gate3984  (.A(g6679), .Z(g6713) ) ;
OR4     gate3985  (.A(g6557), .B(g6634), .C(g4410), .D(g2948), .Z(g6670) ) ;
INV     gate3986  (.A(g6670), .Z(g6714) ) ;
OR4     gate3987  (.A(g6559), .B(g6640), .C(g4416), .D(g2950), .Z(g6673) ) ;
INV     gate3988  (.A(g6673), .Z(g6715) ) ;
INV     gate3989  (.A(g6696), .Z(II8854) ) ;
INV     gate3990  (.A(g6698), .Z(II8857) ) ;
INV     gate3991  (.A(g6699), .Z(II8860) ) ;
INV     gate3992  (.A(g6700), .Z(II8863) ) ;
INV     gate3993  (.A(g6701), .Z(II8866) ) ;
INV     gate3994  (.A(g6694), .Z(II8869) ) ;
INV     gate3995  (.A(g6695), .Z(II8872) ) ;
INV     gate3996  (.A(g6697), .Z(II8875) ) ;
INV     gate3997  (.A(g6710), .Z(II8878) ) ;
INV     gate3998  (.A(g6711), .Z(II8881) ) ;
OR2     gate3999  (.A(g6660), .B(g492), .Z(g6704) ) ;
INV     gate4000  (.A(g6704), .Z(II8884) ) ;
INV     gate4001  (.A(II8884), .Z(g6730) ) ;
INV     gate4002  (.A(g6708), .Z(II8888) ) ;
INV     gate4003  (.A(II8888), .Z(g6732) ) ;
INV     gate4004  (.A(g6706), .Z(II8891) ) ;
INV     gate4005  (.A(II8891), .Z(g6733) ) ;
INV     gate4006  (.A(g6709), .Z(II8894) ) ;
INV     gate4007  (.A(II8894), .Z(g6734) ) ;
INV     gate4008  (.A(g6707), .Z(II8897) ) ;
INV     gate4009  (.A(II8897), .Z(g6735) ) ;
OR2     gate4010  (.A(g6659), .B(g496), .Z(g6702) ) ;
INV     gate4011  (.A(g6702), .Z(II8907) ) ;
INV     gate4012  (.A(II8907), .Z(g6743) ) ;
INV     gate4013  (.A(g6730), .Z(II8910) ) ;
INV     gate4014  (.A(g6743), .Z(II8913) ) ;
NAND3   gate4015  (.A(g6683), .B(g932), .C(g6716), .Z(g6742) ) ;
INV     gate4016  (.A(g6742), .Z(II8916) ) ;
INV     gate4017  (.A(II8916), .Z(g6746) ) ;
NAND3   gate4018  (.A(g6747), .B(g5068), .C(g5066), .Z(g6783) ) ;
INV     gate4019  (.A(g6783), .Z(II8940) ) ;
INV     gate4020  (.A(II8940), .Z(g6784) ) ;
NAND2   gate4021  (.A(g6754), .B(g6750), .Z(g6774) ) ;
INV     gate4022  (.A(g6774), .Z(II8943) ) ;
INV     gate4023  (.A(II8943), .Z(g6785) ) ;
NAND2   gate4024  (.A(g6762), .B(g6758), .Z(g6778) ) ;
INV     gate4025  (.A(g6778), .Z(II8946) ) ;
INV     gate4026  (.A(II8946), .Z(g6786) ) ;
INV     gate4027  (.A(g6774), .Z(II8958) ) ;
INV     gate4028  (.A(II8958), .Z(g6796) ) ;
INV     gate4029  (.A(g6778), .Z(II8961) ) ;
INV     gate4030  (.A(II8961), .Z(g6797) ) ;
INV     gate4031  (.A(g6796), .Z(II8966) ) ;
INV     gate4032  (.A(g6797), .Z(II8969) ) ;
OR2     gate4033  (.A(g4867), .B(g6772), .Z(g6795) ) ;
INV     gate4034  (.A(g6795), .Z(II8972) ) ;
INV     gate4035  (.A(II8972), .Z(g6802) ) ;
OR2     gate4036  (.A(g6768), .B(g3307), .Z(g6791) ) ;
INV     gate4037  (.A(g6791), .Z(II8975) ) ;
INV     gate4038  (.A(II8975), .Z(g6803) ) ;
OR2     gate4039  (.A(g6770), .B(g3321), .Z(g6792) ) ;
INV     gate4040  (.A(g6792), .Z(II8978) ) ;
INV     gate4041  (.A(II8978), .Z(g6806) ) ;
OR2     gate4042  (.A(g6771), .B(g3323), .Z(g6793) ) ;
INV     gate4043  (.A(g6793), .Z(II8981) ) ;
INV     gate4044  (.A(II8981), .Z(g6809) ) ;
OR2     gate4045  (.A(g6777), .B(g3333), .Z(g6794) ) ;
INV     gate4046  (.A(g6794), .Z(II8984) ) ;
INV     gate4047  (.A(II8984), .Z(g6812) ) ;
OR2     gate4048  (.A(g3758), .B(g6766), .Z(g6787) ) ;
INV     gate4049  (.A(g6787), .Z(II8988) ) ;
INV     gate4050  (.A(II8988), .Z(g6817) ) ;
OR2     gate4051  (.A(g3760), .B(g6767), .Z(g6788) ) ;
INV     gate4052  (.A(g6788), .Z(II8991) ) ;
INV     gate4053  (.A(II8991), .Z(g6818) ) ;
OR2     gate4054  (.A(g3764), .B(g6769), .Z(g6789) ) ;
INV     gate4055  (.A(g6789), .Z(II8994) ) ;
INV     gate4056  (.A(II8994), .Z(g6819) ) ;
OR2     gate4057  (.A(g3765), .B(g6773), .Z(g6790) ) ;
INV     gate4058  (.A(g6790), .Z(II8997) ) ;
INV     gate4059  (.A(II8997), .Z(g6820) ) ;
INV     gate4060  (.A(g6785), .Z(g6821) ) ;
INV     gate4061  (.A(g6786), .Z(g6822) ) ;
INV     gate4062  (.A(g6802), .Z(II9002) ) ;
INV     gate4063  (.A(g6817), .Z(II9005) ) ;
INV     gate4064  (.A(g6818), .Z(II9008) ) ;
INV     gate4065  (.A(g6819), .Z(II9011) ) ;
INV     gate4066  (.A(g6820), .Z(II9014) ) ;
INV     gate4067  (.A(g6812), .Z(II9021) ) ;
INV     gate4068  (.A(II9021), .Z(g6832) ) ;
INV     gate4069  (.A(g6803), .Z(II9024) ) ;
INV     gate4070  (.A(II9024), .Z(g6833) ) ;
INV     gate4071  (.A(g6821), .Z(g6834) ) ;
INV     gate4072  (.A(g6806), .Z(II9028) ) ;
INV     gate4073  (.A(II9028), .Z(g6835) ) ;
INV     gate4074  (.A(g6809), .Z(II9031) ) ;
INV     gate4075  (.A(II9031), .Z(g6836) ) ;
INV     gate4076  (.A(g6822), .Z(g6837) ) ;
INV     gate4077  (.A(g6812), .Z(II9035) ) ;
INV     gate4078  (.A(II9035), .Z(g6838) ) ;
INV     gate4079  (.A(g6833), .Z(II9038) ) ;
INV     gate4080  (.A(g6835), .Z(II9041) ) ;
INV     gate4081  (.A(g6836), .Z(II9044) ) ;
INV     gate4082  (.A(g6838), .Z(II9047) ) ;
OR3     gate4083  (.A(II9057), .B(II9058), .C(II9059), .Z(g6844) ) ;
INV     gate4084  (.A(g6844), .Z(II9074) ) ;
INV     gate4085  (.A(II9074), .Z(g6849) ) ;
OR3     gate4086  (.A(II9064), .B(II9065), .C(II9066), .Z(g6845) ) ;
INV     gate4087  (.A(g6845), .Z(II9077) ) ;
INV     gate4088  (.A(II9077), .Z(g6850) ) ;
INV     gate4089  (.A(g6849), .Z(II9082) ) ;
INV     gate4090  (.A(g6850), .Z(II9085) ) ;
OR2     gate4091  (.A(g6851), .B(g2085), .Z(g6855) ) ;
INV     gate4092  (.A(g6855), .Z(II9092) ) ;
INV     gate4093  (.A(II9092), .Z(g6875) ) ;
INV     gate4094  (.A(g6855), .Z(II9095) ) ;
INV     gate4095  (.A(II9095), .Z(g6876) ) ;
OR2     gate4096  (.A(g6852), .B(g2089), .Z(g6864) ) ;
INV     gate4097  (.A(g6864), .Z(II9098) ) ;
INV     gate4098  (.A(II9098), .Z(g6877) ) ;
INV     gate4099  (.A(g6855), .Z(II9101) ) ;
INV     gate4100  (.A(II9101), .Z(g6878) ) ;
INV     gate4101  (.A(g6864), .Z(II9104) ) ;
INV     gate4102  (.A(II9104), .Z(g6879) ) ;
INV     gate4103  (.A(g6855), .Z(II9107) ) ;
INV     gate4104  (.A(II9107), .Z(g6880) ) ;
INV     gate4105  (.A(g6864), .Z(II9110) ) ;
INV     gate4106  (.A(II9110), .Z(g6881) ) ;
INV     gate4107  (.A(g6855), .Z(II9113) ) ;
INV     gate4108  (.A(II9113), .Z(g6882) ) ;
INV     gate4109  (.A(g6864), .Z(II9116) ) ;
INV     gate4110  (.A(II9116), .Z(g6883) ) ;
INV     gate4111  (.A(g6855), .Z(II9119) ) ;
INV     gate4112  (.A(II9119), .Z(g6884) ) ;
INV     gate4113  (.A(g6864), .Z(II9122) ) ;
INV     gate4114  (.A(II9122), .Z(g6885) ) ;
INV     gate4115  (.A(g6855), .Z(II9125) ) ;
INV     gate4116  (.A(II9125), .Z(g6886) ) ;
INV     gate4117  (.A(g6864), .Z(II9128) ) ;
INV     gate4118  (.A(II9128), .Z(g6887) ) ;
INV     gate4119  (.A(g6855), .Z(II9131) ) ;
INV     gate4120  (.A(II9131), .Z(g6888) ) ;
INV     gate4121  (.A(g6864), .Z(II9134) ) ;
INV     gate4122  (.A(II9134), .Z(g6889) ) ;
INV     gate4123  (.A(g6864), .Z(II9137) ) ;
INV     gate4124  (.A(II9137), .Z(g6890) ) ;
INV     gate4125  (.A(g6888), .Z(II9140) ) ;
INV     gate4126  (.A(II9140), .Z(g6891) ) ;
INV     gate4127  (.A(g6886), .Z(II9143) ) ;
INV     gate4128  (.A(II9143), .Z(g6892) ) ;
INV     gate4129  (.A(g6890), .Z(II9146) ) ;
INV     gate4130  (.A(II9146), .Z(g6893) ) ;
INV     gate4131  (.A(g6884), .Z(II9149) ) ;
INV     gate4132  (.A(II9149), .Z(g6894) ) ;
INV     gate4133  (.A(g6889), .Z(II9152) ) ;
INV     gate4134  (.A(II9152), .Z(g6895) ) ;
INV     gate4135  (.A(g6882), .Z(II9155) ) ;
INV     gate4136  (.A(II9155), .Z(g6896) ) ;
INV     gate4137  (.A(g6887), .Z(II9158) ) ;
INV     gate4138  (.A(II9158), .Z(g6897) ) ;
INV     gate4139  (.A(g6880), .Z(II9161) ) ;
INV     gate4140  (.A(II9161), .Z(g6898) ) ;
INV     gate4141  (.A(g6885), .Z(II9164) ) ;
INV     gate4142  (.A(II9164), .Z(g6899) ) ;
INV     gate4143  (.A(g6878), .Z(II9167) ) ;
INV     gate4144  (.A(II9167), .Z(g6900) ) ;
INV     gate4145  (.A(g6883), .Z(II9170) ) ;
INV     gate4146  (.A(II9170), .Z(g6901) ) ;
INV     gate4147  (.A(g6876), .Z(II9173) ) ;
INV     gate4148  (.A(II9173), .Z(g6902) ) ;
INV     gate4149  (.A(g6881), .Z(II9176) ) ;
INV     gate4150  (.A(II9176), .Z(g6903) ) ;
INV     gate4151  (.A(g6875), .Z(II9179) ) ;
INV     gate4152  (.A(II9179), .Z(g6904) ) ;
INV     gate4153  (.A(g6879), .Z(II9182) ) ;
INV     gate4154  (.A(II9182), .Z(g6905) ) ;
INV     gate4155  (.A(g6877), .Z(II9185) ) ;
INV     gate4156  (.A(II9185), .Z(g6906) ) ;
OR2     gate4157  (.A(g6908), .B(g6816), .Z(g6921) ) ;
INV     gate4158  (.A(g6921), .Z(II9203) ) ;
INV     gate4159  (.A(II9203), .Z(g6922) ) ;
INV     gate4160  (.A(g6922), .Z(II9208) ) ;
OR2     gate4161  (.A(g6741), .B(g6929), .Z(g6931) ) ;
INV     gate4162  (.A(g6931), .Z(II9217) ) ;
INV     gate4163  (.A(II9217), .Z(g6932) ) ;
OR2     gate4164  (.A(g6740), .B(g6928), .Z(g6930) ) ;
INV     gate4165  (.A(g6930), .Z(II9220) ) ;
INV     gate4166  (.A(II9220), .Z(g6933) ) ;
OR2     gate4167  (.A(g4616), .B(g6934), .Z(g6937) ) ;
INV     gate4168  (.A(g6937), .Z(II9227) ) ;
INV     gate4169  (.A(II9227), .Z(g6938) ) ;
OR2     gate4170  (.A(g5438), .B(g6935), .Z(g6936) ) ;
INV     gate4171  (.A(g6936), .Z(II9230) ) ;
INV     gate4172  (.A(II9230), .Z(g6939) ) ;
INV     gate4173  (.A(g6938), .Z(II9233) ) ;
INV     gate4174  (.A(g6939), .Z(II9236) ) ;
AND2    gate4175  (.A(g610), .B(g602), .Z(g918) ) ;
AND2    gate4176  (.A(g598), .B(g567), .Z(g1027) ) ;
AND2    gate4177  (.A(g913), .B(g266), .Z(g1416) ) ;
AND2    gate4178  (.A(g613), .B(g918), .Z(g1419) ) ;
AND2    gate4179  (.A(g834), .B(g830), .Z(g1436) ) ;
AND2    gate4180  (.A(g1101), .B(g1094), .Z(g1499) ) ;
AND2    gate4181  (.A(g1017), .B(g1011), .Z(g1514) ) ;
AND2    gate4182  (.A(g634), .B(g1027), .Z(g1570) ) ;
AND2    gate4183  (.A(g980), .B(g965), .Z(g1575) ) ;
AND2    gate4184  (.A(g1101), .B(g1094), .Z(g1576) ) ;
AND2    gate4185  (.A(g1017), .B(g1011), .Z(g1585) ) ;
AND3    gate4186  (.A(g749), .B(g743), .C(g736), .Z(II2566) ) ;
AND2    gate4187  (.A(g760), .B(g754), .Z(g1609) ) ;
AND3    gate4188  (.A(g804), .B(g798), .C(g791), .Z(II2574) ) ;
AND2    gate4189  (.A(g1056), .B(g1084), .Z(g1620) ) ;
AND2    gate4190  (.A(g815), .B(g809), .Z(g1628) ) ;
AND2    gate4191  (.A(g716), .B(g152), .Z(g1633) ) ;
AND2    gate4192  (.A(g766), .B(g719), .Z(g1689) ) ;
AND2    gate4193  (.A(g821), .B(g774), .Z(g1691) ) ;
AND3    gate4194  (.A(g766), .B(g719), .C(g729), .Z(g1706) ) ;
AND3    gate4195  (.A(g821), .B(g774), .C(g784), .Z(g1716) ) ;
AND2    gate4196  (.A(g478), .B(g1119), .Z(g1763) ) ;
AND2    gate4197  (.A(g858), .B(g889), .Z(g1784) ) ;
AND2    gate4198  (.A(g706), .B(g49), .Z(g1808) ) ;
AND2    gate4199  (.A(g714), .B(g710), .Z(g1826) ) ;
AND2    gate4200  (.A(g616), .B(g1419), .Z(g2015) ) ;
AND2    gate4201  (.A(g1423), .B(g1254), .Z(g2018) ) ;
AND2    gate4202  (.A(g835), .B(g1436), .Z(g2021) ) ;
NAND2   gate4203  (.A(g314), .B(g310), .Z(g901) ) ;
AND2    gate4204  (.A(g1094), .B(g1675), .Z(g2053) ) ;
AND2    gate4205  (.A(g1672), .B(g1675), .Z(g2056) ) ;
AND2    gate4206  (.A(g1499), .B(g1666), .Z(g2062) ) ;
AND2    gate4207  (.A(g1541), .B(g1546), .Z(g2068) ) ;
AND2    gate4208  (.A(g1088), .B(g1499), .Z(g2073) ) ;
AND2    gate4209  (.A(g1094), .B(g1546), .Z(g2081) ) ;
AND2    gate4210  (.A(g1577), .B(g1563), .Z(g2084) ) ;
AND2    gate4211  (.A(g1123), .B(g1567), .Z(g2085) ) ;
AND2    gate4212  (.A(g1123), .B(g1578), .Z(g2089) ) ;
AND2    gate4213  (.A(g642), .B(g1570), .Z(g2092) ) ;
AND2    gate4214  (.A(g1001), .B(g1543), .Z(g2101) ) ;
AND2    gate4215  (.A(g1583), .B(g1543), .Z(g2107) ) ;
AND2    gate4216  (.A(g1576), .B(g1535), .Z(g2113) ) ;
AND2    gate4217  (.A(g1632), .B(g754), .Z(g2121) ) ;
AND2    gate4218  (.A(g760), .B(g1638), .Z(g2137) ) ;
AND2    gate4219  (.A(g1639), .B(g809), .Z(g2138) ) ;
AND2    gate4220  (.A(g1793), .B(g1777), .Z(g2142) ) ;
AND2    gate4221  (.A(g815), .B(g1642), .Z(g2156) ) ;
AND2    gate4222  (.A(g1624), .B(g929), .Z(g2160) ) ;
AND2    gate4223  (.A(g1633), .B(g161), .Z(g2166) ) ;
AND2    gate4224  (.A(g1706), .B(g736), .Z(g2255) ) ;
AND2    gate4225  (.A(g1716), .B(g791), .Z(g2267) ) ;
AND3    gate4226  (.A(g1706), .B(g736), .C(g743), .Z(g2292) ) ;
AND3    gate4227  (.A(g1716), .B(g791), .C(g798), .Z(g2294) ) ;
AND2    gate4228  (.A(g471), .B(g1358), .Z(g2323) ) ;
AND2    gate4229  (.A(g1603), .B(g197), .Z(g2339) ) ;
AND2    gate4230  (.A(g1398), .B(g1387), .Z(g2340) ) ;
AND2    gate4231  (.A(g1603), .B(g269), .Z(g2356) ) ;
AND2    gate4232  (.A(g1808), .B(g54), .Z(g2419) ) ;
AND2    gate4233  (.A(g715), .B(g1826), .Z(g2551) ) ;
NAND2   gate4234  (.A(g102), .B(g98), .Z(g1138) ) ;
NAND2   gate4235  (.A(II2675), .B(II2676), .Z(g1686) ) ;
AND2    gate4236  (.A(g1686), .B(g2296), .Z(g2659) ) ;
NAND2   gate4237  (.A(II3399), .B(II3400), .Z(g2263) ) ;
AND2    gate4238  (.A(g2263), .B(g2296), .Z(g2671) ) ;
AND2    gate4239  (.A(g2370), .B(g1887), .Z(g2685) ) ;
AND2    gate4240  (.A(g2397), .B(g1905), .Z(g2699) ) ;
AND2    gate4241  (.A(g2370), .B(g1908), .Z(g2700) ) ;
AND2    gate4242  (.A(g2422), .B(g1919), .Z(g2720) ) ;
AND2    gate4243  (.A(g2397), .B(g1922), .Z(g2721) ) ;
AND2    gate4244  (.A(g2449), .B(g1940), .Z(g2732) ) ;
AND2    gate4245  (.A(g2422), .B(g1943), .Z(g2733) ) ;
AND2    gate4246  (.A(g2473), .B(g1954), .Z(g2746) ) ;
AND2    gate4247  (.A(g2449), .B(g1957), .Z(g2747) ) ;
AND2    gate4248  (.A(g2497), .B(g1963), .Z(g2758) ) ;
AND2    gate4249  (.A(g2473), .B(g1966), .Z(g2759) ) ;
AND2    gate4250  (.A(g2518), .B(g1972), .Z(g2770) ) ;
AND2    gate4251  (.A(g2497), .B(g1975), .Z(g2771) ) ;
AND2    gate4252  (.A(g2544), .B(g1982), .Z(g2781) ) ;
AND2    gate4253  (.A(g2518), .B(g1985), .Z(g2782) ) ;
AND2    gate4254  (.A(g2568), .B(g1991), .Z(g2793) ) ;
AND2    gate4255  (.A(g2544), .B(g1994), .Z(g2794) ) ;
AND2    gate4256  (.A(g2568), .B(g2001), .Z(g2807) ) ;
NAND3   gate4257  (.A(g901), .B(g1387), .C(g905), .Z(g2009) ) ;
AND2    gate4258  (.A(g2009), .B(g1581), .Z(g2808) ) ;
AND2    gate4259  (.A(g1890), .B(g910), .Z(g2821) ) ;
AND3    gate4260  (.A(g1279), .B(g2025), .C(g1267), .Z(II4040) ) ;
AND2    gate4261  (.A(g619), .B(g2015), .Z(g2846) ) ;
AND2    gate4262  (.A(g2018), .B(g1255), .Z(g2850) ) ;
AND2    gate4263  (.A(g836), .B(g2021), .Z(g2853) ) ;
AND2    gate4264  (.A(g710), .B(g2296), .Z(g2860) ) ;
NAND2   gate4265  (.A(II2300), .B(II2301), .Z(g1316) ) ;
AND2    gate4266  (.A(g1316), .B(g1861), .Z(g2868) ) ;
NAND2   gate4267  (.A(II2934), .B(II2935), .Z(g1845) ) ;
AND2    gate4268  (.A(g1845), .B(g1861), .Z(g2873) ) ;
AND2    gate4269  (.A(g1030), .B(g2062), .Z(g2897) ) ;
AND2    gate4270  (.A(g606), .B(g2092), .Z(g2909) ) ;
AND2    gate4271  (.A(g1030), .B(g2113), .Z(g2916) ) ;
AND2    gate4272  (.A(g2291), .B(g1788), .Z(g2935) ) ;
AND2    gate4273  (.A(g2160), .B(g931), .Z(g2937) ) ;
AND2    gate4274  (.A(g2166), .B(g170), .Z(g2941) ) ;
AND2    gate4275  (.A(g2137), .B(g1595), .Z(g2948) ) ;
AND2    gate4276  (.A(g830), .B(g1861), .Z(g2949) ) ;
AND2    gate4277  (.A(g2156), .B(g1612), .Z(g2950) ) ;
AND2    gate4278  (.A(g2381), .B(g293), .Z(g2953) ) ;
AND2    gate4279  (.A(g2381), .B(g297), .Z(g2955) ) ;
AND2    gate4280  (.A(g212), .B(g2336), .Z(g3089) ) ;
AND2    gate4281  (.A(g218), .B(g2350), .Z(g3099) ) ;
AND2    gate4282  (.A(g212), .B(g2353), .Z(g3103) ) ;
AND2    gate4283  (.A(g224), .B(g2364), .Z(g3113) ) ;
AND2    gate4284  (.A(g218), .B(g2367), .Z(g3117) ) ;
NAND3   gate4285  (.A(g1138), .B(g1777), .C(g1157), .Z(g2435) ) ;
AND2    gate4286  (.A(g2435), .B(g1394), .Z(g3122) ) ;
AND2    gate4287  (.A(g230), .B(g2391), .Z(g3123) ) ;
AND2    gate4288  (.A(g224), .B(g2394), .Z(g3127) ) ;
AND2    gate4289  (.A(g2306), .B(g1206), .Z(g3132) ) ;
AND2    gate4290  (.A(g236), .B(g2410), .Z(g3133) ) ;
AND2    gate4291  (.A(g230), .B(g2413), .Z(g3134) ) ;
AND2    gate4292  (.A(g2370), .B(g2416), .Z(g3135) ) ;
AND2    gate4293  (.A(g242), .B(g2437), .Z(g3143) ) ;
AND2    gate4294  (.A(g236), .B(g2440), .Z(g3144) ) ;
AND2    gate4295  (.A(g2397), .B(g2443), .Z(g3145) ) ;
AND2    gate4296  (.A(g2370), .B(g2446), .Z(g3146) ) ;
AND2    gate4297  (.A(g2419), .B(g59), .Z(g3147) ) ;
AND2    gate4298  (.A(g2039), .B(g1410), .Z(g3154) ) ;
AND2    gate4299  (.A(g248), .B(g2461), .Z(g3155) ) ;
AND2    gate4300  (.A(g242), .B(g2464), .Z(g3156) ) ;
AND2    gate4301  (.A(g2422), .B(g2467), .Z(g3157) ) ;
AND2    gate4302  (.A(g2397), .B(g2470), .Z(g3161) ) ;
AND2    gate4303  (.A(g2042), .B(g1233), .Z(g3166) ) ;
AND2    gate4304  (.A(g1883), .B(g921), .Z(g3167) ) ;
AND2    gate4305  (.A(g254), .B(g2485), .Z(g3170) ) ;
AND2    gate4306  (.A(g248), .B(g2488), .Z(g3171) ) ;
AND2    gate4307  (.A(g2449), .B(g2491), .Z(g3172) ) ;
AND2    gate4308  (.A(g2422), .B(g2494), .Z(g3176) ) ;
AND2    gate4309  (.A(g260), .B(g2506), .Z(g3180) ) ;
AND2    gate4310  (.A(g254), .B(g2509), .Z(g3181) ) ;
AND2    gate4311  (.A(g2473), .B(g2512), .Z(g3182) ) ;
AND2    gate4312  (.A(g2449), .B(g2515), .Z(g3186) ) ;
AND2    gate4313  (.A(g260), .B(g2535), .Z(g3190) ) ;
AND2    gate4314  (.A(g2497), .B(g2538), .Z(g3191) ) ;
AND2    gate4315  (.A(g2473), .B(g2541), .Z(g3195) ) ;
AND2    gate4316  (.A(g2497), .B(g2565), .Z(g3203) ) ;
AND2    gate4317  (.A(g895), .B(g2551), .Z(g3208) ) ;
AND2    gate4318  (.A(g2172), .B(g2615), .Z(g3275) ) ;
AND2    gate4319  (.A(g2174), .B(g2625), .Z(g3277) ) ;
AND2    gate4320  (.A(g2175), .B(g2628), .Z(g3278) ) ;
AND2    gate4321  (.A(g2599), .B(g2612), .Z(g3279) ) ;
AND2    gate4322  (.A(g2177), .B(g2637), .Z(g3280) ) ;
AND2    gate4323  (.A(g2178), .B(g2640), .Z(g3281) ) ;
AND2    gate4324  (.A(g131), .B(g2863), .Z(g3282) ) ;
AND2    gate4325  (.A(g2609), .B(g2622), .Z(g3283) ) ;
AND2    gate4326  (.A(g2195), .B(g2653), .Z(g3285) ) ;
AND2    gate4327  (.A(g2196), .B(g2656), .Z(g3286) ) ;
AND2    gate4328  (.A(g135), .B(g2865), .Z(g3287) ) ;
AND2    gate4329  (.A(g2631), .B(g2634), .Z(g3288) ) ;
AND2    gate4330  (.A(g2213), .B(g2664), .Z(g3290) ) ;
AND2    gate4331  (.A(g2214), .B(g2667), .Z(g3292) ) ;
AND2    gate4332  (.A(g212), .B(g2864), .Z(g3293) ) ;
AND2    gate4333  (.A(g139), .B(g2870), .Z(g3294) ) ;
AND2    gate4334  (.A(g2660), .B(g2647), .Z(g3295) ) ;
AND2    gate4335  (.A(g3054), .B(g2650), .Z(g3296) ) ;
AND2    gate4336  (.A(g2231), .B(g2679), .Z(g3298) ) ;
AND2    gate4337  (.A(g2232), .B(g2682), .Z(g3300) ) ;
AND2    gate4338  (.A(g218), .B(g2866), .Z(g3301) ) ;
AND2    gate4339  (.A(g212), .B(g2867), .Z(g3302) ) ;
AND2    gate4340  (.A(g2722), .B(g2890), .Z(g3303) ) ;
AND2    gate4341  (.A(g2857), .B(g1513), .Z(g3304) ) ;
NAND2   gate4342  (.A(II4151), .B(II4152), .Z(g2960) ) ;
AND2    gate4343  (.A(g2960), .B(g2296), .Z(g3305) ) ;
AND2    gate4344  (.A(g2242), .B(g2692), .Z(g3307) ) ;
AND2    gate4345  (.A(g2243), .B(g2695), .Z(g3309) ) ;
AND2    gate4346  (.A(g224), .B(g2871), .Z(g3310) ) ;
AND2    gate4347  (.A(g218), .B(g2872), .Z(g3311) ) ;
AND2    gate4348  (.A(g2701), .B(g1875), .Z(g3315) ) ;
AND2    gate4349  (.A(g2748), .B(g2894), .Z(g3316) ) ;
AND2    gate4350  (.A(g2722), .B(g2895), .Z(g3317) ) ;
AND2    gate4351  (.A(g2688), .B(g2675), .Z(g3319) ) ;
AND2    gate4352  (.A(g2252), .B(g2713), .Z(g3321) ) ;
AND2    gate4353  (.A(g2253), .B(g2716), .Z(g3323) ) ;
AND2    gate4354  (.A(g230), .B(g2875), .Z(g3324) ) ;
AND2    gate4355  (.A(g224), .B(g2876), .Z(g3325) ) ;
AND2    gate4356  (.A(g2734), .B(g1891), .Z(g3326) ) ;
AND2    gate4357  (.A(g2772), .B(g2906), .Z(g3327) ) ;
AND2    gate4358  (.A(g2701), .B(g1894), .Z(g3328) ) ;
AND2    gate4359  (.A(g2748), .B(g2907), .Z(g3329) ) ;
AND2    gate4360  (.A(g2264), .B(g2728), .Z(g3333) ) ;
AND2    gate4361  (.A(g236), .B(g2883), .Z(g3334) ) ;
AND2    gate4362  (.A(g230), .B(g2884), .Z(g3335) ) ;
AND2    gate4363  (.A(g2760), .B(g1911), .Z(g3336) ) ;
AND2    gate4364  (.A(g2796), .B(g2913), .Z(g3337) ) ;
AND2    gate4365  (.A(g3162), .B(g2914), .Z(g3338) ) ;
AND2    gate4366  (.A(g2734), .B(g1914), .Z(g3339) ) ;
AND2    gate4367  (.A(g2772), .B(g2915), .Z(g3340) ) ;
AND2    gate4368  (.A(g2998), .B(g2709), .Z(g3341) ) ;
AND2    gate4369  (.A(g242), .B(g2885), .Z(g3344) ) ;
AND2    gate4370  (.A(g236), .B(g2886), .Z(g3345) ) ;
AND2    gate4371  (.A(g2783), .B(g1925), .Z(g3349) ) ;
AND2    gate4372  (.A(g3150), .B(g1928), .Z(g3350) ) ;
AND2    gate4373  (.A(g2760), .B(g1931), .Z(g3351) ) ;
AND2    gate4374  (.A(g2796), .B(g2920), .Z(g3352) ) ;
AND2    gate4375  (.A(g3162), .B(g2921), .Z(g3353) ) ;
AND2    gate4376  (.A(g248), .B(g2888), .Z(g3356) ) ;
AND2    gate4377  (.A(g242), .B(g2889), .Z(g3357) ) ;
AND2    gate4378  (.A(g2842), .B(g1369), .Z(g3358) ) ;
AND2    gate4379  (.A(g2822), .B(g2922), .Z(g3359) ) ;
AND2    gate4380  (.A(g2783), .B(g1947), .Z(g3360) ) ;
AND2    gate4381  (.A(g3150), .B(g1950), .Z(g3361) ) ;
AND2    gate4382  (.A(g3031), .B(g2740), .Z(g3362) ) ;
AND2    gate4383  (.A(g254), .B(g2892), .Z(g3365) ) ;
AND2    gate4384  (.A(g248), .B(g2893), .Z(g3366) ) ;
AND2    gate4385  (.A(g2809), .B(g1960), .Z(g3367) ) ;
AND2    gate4386  (.A(g2822), .B(g2923), .Z(g3368) ) ;
AND2    gate4387  (.A(g260), .B(g2904), .Z(g3371) ) ;
AND2    gate4388  (.A(g254), .B(g2905), .Z(g3372) ) ;
AND2    gate4389  (.A(g3118), .B(g2927), .Z(g3373) ) ;
AND2    gate4390  (.A(g2809), .B(g1969), .Z(g3374) ) ;
AND2    gate4391  (.A(g260), .B(g2912), .Z(g3375) ) ;
AND2    gate4392  (.A(g3104), .B(g1979), .Z(g3376) ) ;
AND2    gate4393  (.A(g3118), .B(g2931), .Z(g3377) ) ;
AND2    gate4394  (.A(g3136), .B(g2932), .Z(g3378) ) ;
AND2    gate4395  (.A(g3104), .B(g1988), .Z(g3379) ) ;
AND2    gate4396  (.A(g3128), .B(g1998), .Z(g3381) ) ;
AND2    gate4397  (.A(g3136), .B(g2934), .Z(g3382) ) ;
AND2    gate4398  (.A(g3128), .B(g2004), .Z(g3383) ) ;
AND2    gate4399  (.A(g622), .B(g2846), .Z(g3421) ) ;
AND2    gate4400  (.A(g2296), .B(g3208), .Z(g3425) ) ;
NAND2   gate4401  (.A(g301), .B(g319), .Z(g905) ) ;
AND3    gate4402  (.A(g1359), .B(g2831), .C(g905), .Z(g3433) ) ;
AND2    gate4403  (.A(g2850), .B(g857), .Z(g3434) ) ;
AND2    gate4404  (.A(g837), .B(g2853), .Z(g3437) ) ;
AND2    gate4405  (.A(g128), .B(g2946), .Z(g3449) ) ;
AND2    gate4406  (.A(g341), .B(g2956), .Z(g3464) ) ;
AND2    gate4407  (.A(g345), .B(g2957), .Z(g3479) ) ;
AND2    gate4408  (.A(g349), .B(g2958), .Z(g3484) ) ;
NAND2   gate4409  (.A(II3740), .B(II3741), .Z(g2607) ) ;
AND2    gate4410  (.A(g2607), .B(g1861), .Z(g3489) ) ;
AND2    gate4411  (.A(g353), .B(g2959), .Z(g3490) ) ;
AND2    gate4412  (.A(g357), .B(g2961), .Z(g3499) ) ;
AND2    gate4413  (.A(g646), .B(g2909), .Z(g3522) ) ;
AND2    gate4414  (.A(g2937), .B(g938), .Z(g3551) ) ;
AND2    gate4415  (.A(g2941), .B(g179), .Z(g3554) ) ;
AND2    gate4416  (.A(g338), .B(g3199), .Z(g3558) ) ;
AND2    gate4417  (.A(g2688), .B(g2663), .Z(g3602) ) ;
AND2    gate4418  (.A(g2370), .B(g3019), .Z(g3603) ) ;
AND2    gate4419  (.A(g2599), .B(g2308), .Z(g3608) ) ;
AND2    gate4420  (.A(g2706), .B(g2678), .Z(g3609) ) ;
AND2    gate4421  (.A(g2397), .B(g3034), .Z(g3610) ) ;
AND2    gate4422  (.A(g2370), .B(g3037), .Z(g3611) ) ;
AND2    gate4423  (.A(g2604), .B(g2312), .Z(g3613) ) ;
AND2    gate4424  (.A(g2998), .B(g2691), .Z(g3614) ) ;
AND2    gate4425  (.A(g2422), .B(g3046), .Z(g3615) ) ;
AND2    gate4426  (.A(g2397), .B(g3049), .Z(g3616) ) ;
AND2    gate4427  (.A(g2609), .B(g2317), .Z(g3617) ) ;
AND2    gate4428  (.A(g3016), .B(g2712), .Z(g3618) ) ;
AND2    gate4429  (.A(g2449), .B(g3057), .Z(g3619) ) ;
AND2    gate4430  (.A(g2422), .B(g3060), .Z(g3620) ) ;
AND2    gate4431  (.A(g2619), .B(g2320), .Z(g3625) ) ;
AND2    gate4432  (.A(g3031), .B(g2727), .Z(g3626) ) ;
AND2    gate4433  (.A(g2473), .B(g3067), .Z(g3627) ) ;
AND2    gate4434  (.A(g2449), .B(g3070), .Z(g3628) ) ;
AND2    gate4435  (.A(g2809), .B(g2738), .Z(g3629) ) ;
AND2    gate4436  (.A(g3167), .B(g1756), .Z(g3630) ) ;
AND2    gate4437  (.A(g2631), .B(g2324), .Z(g3631) ) ;
AND2    gate4438  (.A(g3043), .B(g2743), .Z(g3632) ) ;
AND2    gate4439  (.A(g2497), .B(g3076), .Z(g3633) ) ;
AND2    gate4440  (.A(g2179), .B(g2744), .Z(g3634) ) ;
AND2    gate4441  (.A(g2473), .B(g3079), .Z(g3635) ) ;
AND2    gate4442  (.A(g2701), .B(g2327), .Z(g3636) ) ;
AND2    gate4443  (.A(g2822), .B(g2752), .Z(g3637) ) ;
AND2    gate4444  (.A(g2644), .B(g2333), .Z(g3641) ) ;
AND2    gate4445  (.A(g3054), .B(g2754), .Z(g3642) ) ;
AND2    gate4446  (.A(g2518), .B(g3086), .Z(g3643) ) ;
AND2    gate4447  (.A(g2197), .B(g2755), .Z(g3644) ) ;
AND2    gate4448  (.A(g2497), .B(g3090), .Z(g3645) ) ;
AND2    gate4449  (.A(g2179), .B(g2756), .Z(g3646) ) ;
AND2    gate4450  (.A(g2722), .B(g2343), .Z(g3648) ) ;
AND2    gate4451  (.A(g3104), .B(g2764), .Z(g3649) ) ;
AND2    gate4452  (.A(g2660), .B(g2347), .Z(g3650) ) ;
AND2    gate4453  (.A(g3064), .B(g2766), .Z(g3651) ) ;
AND2    gate4454  (.A(g2544), .B(g3096), .Z(g3652) ) ;
AND2    gate4455  (.A(g2215), .B(g2767), .Z(g3653) ) ;
AND2    gate4456  (.A(g2518), .B(g3100), .Z(g3654) ) ;
AND2    gate4457  (.A(g2197), .B(g2768), .Z(g3655) ) ;
AND2    gate4458  (.A(g2734), .B(g2357), .Z(g3657) ) ;
AND2    gate4459  (.A(g3118), .B(g2776), .Z(g3658) ) ;
AND2    gate4460  (.A(g2672), .B(g2361), .Z(g3659) ) ;
AND2    gate4461  (.A(g2568), .B(g3110), .Z(g3660) ) ;
AND2    gate4462  (.A(g2234), .B(g2778), .Z(g3661) ) ;
AND2    gate4463  (.A(g2544), .B(g3114), .Z(g3662) ) ;
AND2    gate4464  (.A(g2215), .B(g2779), .Z(g3663) ) ;
AND2    gate4465  (.A(g2748), .B(g2378), .Z(g3665) ) ;
AND2    gate4466  (.A(g3128), .B(g2787), .Z(g3666) ) ;
AND2    gate4467  (.A(g2245), .B(g2789), .Z(g3667) ) ;
AND2    gate4468  (.A(g2568), .B(g3124), .Z(g3668) ) ;
AND2    gate4469  (.A(g2234), .B(g2790), .Z(g3669) ) ;
AND2    gate4470  (.A(g2234), .B(g2792), .Z(g3670) ) ;
AND2    gate4471  (.A(g2760), .B(g2405), .Z(g3671) ) ;
AND2    gate4472  (.A(g3136), .B(g2800), .Z(g3672) ) ;
AND2    gate4473  (.A(g2256), .B(g2802), .Z(g3678) ) ;
AND2    gate4474  (.A(g2245), .B(g2803), .Z(g3679) ) ;
AND2    gate4475  (.A(g2245), .B(g2805), .Z(g3680) ) ;
AND2    gate4476  (.A(g2234), .B(g2806), .Z(g3681) ) ;
AND2    gate4477  (.A(g2772), .B(g2430), .Z(g3682) ) ;
AND2    gate4478  (.A(g3150), .B(g2813), .Z(g3683) ) ;
AND2    gate4479  (.A(g2268), .B(g2817), .Z(g3684) ) ;
AND2    gate4480  (.A(g2256), .B(g2818), .Z(g3685) ) ;
AND2    gate4481  (.A(g2256), .B(g2819), .Z(g3686) ) ;
AND2    gate4482  (.A(g2245), .B(g2820), .Z(g3687) ) ;
AND2    gate4483  (.A(g2783), .B(g2457), .Z(g3688) ) ;
AND2    gate4484  (.A(g3162), .B(g2826), .Z(g3689) ) ;
AND2    gate4485  (.A(g2276), .B(g2827), .Z(g3690) ) ;
AND2    gate4486  (.A(g2268), .B(g2828), .Z(g3691) ) ;
AND2    gate4487  (.A(g2268), .B(g2829), .Z(g3692) ) ;
AND2    gate4488  (.A(g2256), .B(g2830), .Z(g3693) ) ;
AND2    gate4489  (.A(g3147), .B(g64), .Z(g3694) ) ;
AND2    gate4490  (.A(g2796), .B(g2481), .Z(g3697) ) ;
AND2    gate4491  (.A(g2284), .B(g2835), .Z(g3698) ) ;
AND2    gate4492  (.A(g2276), .B(g2836), .Z(g3699) ) ;
AND2    gate4493  (.A(g2276), .B(g2837), .Z(g3700) ) ;
AND2    gate4494  (.A(g2268), .B(g2838), .Z(g3701) ) ;
AND2    gate4495  (.A(g2284), .B(g2839), .Z(g3702) ) ;
AND2    gate4496  (.A(g2284), .B(g2840), .Z(g3703) ) ;
AND2    gate4497  (.A(g2276), .B(g2841), .Z(g3704) ) ;
AND2    gate4498  (.A(g2284), .B(g2845), .Z(g3709) ) ;
NAND2   gate4499  (.A(g89), .B(g107), .Z(g1157) ) ;
AND3    gate4500  (.A(g1743), .B(g3140), .C(g1157), .Z(g3718) ) ;
AND2    gate4501  (.A(g2604), .B(g3481), .Z(g3755) ) ;
AND2    gate4502  (.A(g2619), .B(g3487), .Z(g3757) ) ;
AND2    gate4503  (.A(g545), .B(g3461), .Z(g3758) ) ;
AND2    gate4504  (.A(g2644), .B(g3498), .Z(g3759) ) ;
AND2    gate4505  (.A(g548), .B(g3465), .Z(g3760) ) ;
AND2    gate4506  (.A(g2672), .B(g3500), .Z(g3762) ) ;
AND2    gate4507  (.A(g3064), .B(g3501), .Z(g3763) ) ;
AND2    gate4508  (.A(g551), .B(g3480), .Z(g3764) ) ;
AND2    gate4509  (.A(g554), .B(g3485), .Z(g3765) ) ;
AND2    gate4510  (.A(g2706), .B(g3504), .Z(g3767) ) ;
AND2    gate4511  (.A(g3016), .B(g3510), .Z(g3774) ) ;
AND2    gate4512  (.A(g3043), .B(g3519), .Z(g3780) ) ;
AND2    gate4513  (.A(g114), .B(g3251), .Z(g3784) ) ;
NAND2   gate4514  (.A(II3126), .B(II3127), .Z(g2024) ) ;
AND2    gate4515  (.A(g3384), .B(g2024), .Z(g3806) ) ;
AND2    gate4516  (.A(g625), .B(g3421), .Z(g3810) ) ;
AND2    gate4517  (.A(g3434), .B(g861), .Z(g3816) ) ;
AND2    gate4518  (.A(g964), .B(g3437), .Z(g3819) ) ;
AND2    gate4519  (.A(g2330), .B(g3425), .Z(g3831) ) ;
OR2     gate4520  (.A(g3154), .B(g3166), .Z(g3533) ) ;
AND3    gate4521  (.A(g2856), .B(g945), .C(g3533), .Z(g3843) ) ;
NAND2   gate4522  (.A(II4546), .B(II4547), .Z(g3276) ) ;
AND2    gate4523  (.A(g3276), .B(g1861), .Z(g3887) ) ;
AND2    gate4524  (.A(g323), .B(g3441), .Z(g3899) ) ;
AND2    gate4525  (.A(g650), .B(g3522), .Z(g3907) ) ;
AND2    gate4526  (.A(g3505), .B(g471), .Z(g3924) ) ;
AND2    gate4527  (.A(g3512), .B(g478), .Z(g3928) ) ;
AND2    gate4528  (.A(g3551), .B(g940), .Z(g3936) ) ;
AND2    gate4529  (.A(g3554), .B(g188), .Z(g3953) ) ;
AND3    gate4530  (.A(g1250), .B(g3425), .C(g2849), .Z(g3997) ) ;
AND2    gate4531  (.A(g445), .B(g3388), .Z(g4015) ) ;
AND2    gate4532  (.A(g441), .B(g3388), .Z(g4032) ) ;
AND2    gate4533  (.A(g426), .B(g3388), .Z(g4033) ) ;
AND2    gate4534  (.A(g437), .B(g3388), .Z(g4035) ) ;
OR2     gate4535  (.A(g2323), .B(g1763), .Z(g2896) ) ;
AND2    gate4536  (.A(g2896), .B(g3388), .Z(g4037) ) ;
AND2    gate4537  (.A(g430), .B(g3388), .Z(g4038) ) ;
AND2    gate4538  (.A(g402), .B(g3388), .Z(g4039) ) ;
AND2    gate4539  (.A(g461), .B(g3388), .Z(g4041) ) ;
AND2    gate4540  (.A(g406), .B(g3388), .Z(g4042) ) ;
AND2    gate4541  (.A(g457), .B(g3388), .Z(g4043) ) ;
AND2    gate4542  (.A(g410), .B(g3388), .Z(g4044) ) ;
AND2    gate4543  (.A(g3425), .B(g123), .Z(g4045) ) ;
NAND4   gate4544  (.A(g3158), .B(g3002), .C(g2976), .D(g2968), .Z(g3511) ) ;
NAND4   gate4545  (.A(g3173), .B(g3002), .C(g2976), .D(g2179), .Z(g3517) ) ;
NAND4   gate4546  (.A(g3183), .B(g3002), .C(g2197), .D(g2968), .Z(g3520) ) ;
NAND4   gate4547  (.A(g3192), .B(g3002), .C(g2197), .D(g2179), .Z(g3525) ) ;
AND4    gate4548  (.A(g3511), .B(g3517), .C(g3520), .D(g3525), .Z(II5351) ) ;
NAND4   gate4549  (.A(g3200), .B(g2215), .C(g2976), .D(g2968), .Z(g3529) ) ;
NAND4   gate4550  (.A(g3209), .B(g2215), .C(g2976), .D(g2179), .Z(g3531) ) ;
NAND4   gate4551  (.A(g3216), .B(g2215), .C(g2197), .D(g2968), .Z(g3535) ) ;
NAND4   gate4552  (.A(g2588), .B(g2215), .C(g2197), .D(g2179), .Z(g3538) ) ;
AND4    gate4553  (.A(g3529), .B(g3531), .C(g3535), .D(g3538), .Z(II5352) ) ;
AND2    gate4554  (.A(g453), .B(g3388), .Z(g4047) ) ;
AND2    gate4555  (.A(g414), .B(g3388), .Z(g4048) ) ;
NAND4   gate4556  (.A(g3177), .B(g3023), .C(g3007), .D(g2981), .Z(g3518) ) ;
NAND4   gate4557  (.A(g3187), .B(g3023), .C(g3007), .D(g2179), .Z(g3521) ) ;
NAND4   gate4558  (.A(g3196), .B(g3023), .C(g2197), .D(g2981), .Z(g3526) ) ;
NAND4   gate4559  (.A(g3204), .B(g3023), .C(g2197), .D(g2179), .Z(g3530) ) ;
AND4    gate4560  (.A(g3518), .B(g3521), .C(g3526), .D(g3530), .Z(II5359) ) ;
NAND4   gate4561  (.A(g3212), .B(g2215), .C(g3007), .D(g2981), .Z(g3532) ) ;
NAND4   gate4562  (.A(g3219), .B(g2215), .C(g3007), .D(g2179), .Z(g3536) ) ;
NAND4   gate4563  (.A(g2591), .B(g2215), .C(g2197), .D(g2981), .Z(g3539) ) ;
NAND4   gate4564  (.A(g2594), .B(g2215), .C(g2197), .D(g2179), .Z(g3544) ) ;
AND4    gate4565  (.A(g3532), .B(g3536), .C(g3539), .D(g3544), .Z(II5360) ) ;
AND2    gate4566  (.A(g449), .B(g3388), .Z(g4051) ) ;
AND2    gate4567  (.A(g418), .B(g3388), .Z(g4052) ) ;
AND2    gate4568  (.A(g3387), .B(g1415), .Z(g4053) ) ;
AND2    gate4569  (.A(g3694), .B(g69), .Z(g4054) ) ;
AND2    gate4570  (.A(g422), .B(g3388), .Z(g4057) ) ;
AND2    gate4571  (.A(g3424), .B(g1246), .Z(g4058) ) ;
NOR2    gate4572  (.A(g3338), .B(g3350), .Z(g3926) ) ;
AND2    gate4573  (.A(g3926), .B(g2078), .Z(g4156) ) ;
NOR2    gate4574  (.A(g3378), .B(g3381), .Z(g3923) ) ;
AND2    gate4575  (.A(g3923), .B(g1345), .Z(g4160) ) ;
NOR2    gate4576  (.A(g3353), .B(g3361), .Z(g3931) ) ;
AND2    gate4577  (.A(g3931), .B(g2087), .Z(g4161) ) ;
NOR2    gate4578  (.A(g3316), .B(g3326), .Z(g3958) ) ;
AND2    gate4579  (.A(g3958), .B(g2091), .Z(g4164) ) ;
NOR2    gate4580  (.A(g3382), .B(g3383), .Z(g3927) ) ;
AND2    gate4581  (.A(g3927), .B(g1352), .Z(g4165) ) ;
NOR2    gate4582  (.A(g3303), .B(g3315), .Z(g3925) ) ;
AND2    gate4583  (.A(g3925), .B(g1355), .Z(g4168) ) ;
NOR2    gate4584  (.A(g3329), .B(g3339), .Z(g3966) ) ;
AND2    gate4585  (.A(g3966), .B(g2099), .Z(g4169) ) ;
NOR2    gate4586  (.A(g3337), .B(g3349), .Z(g3956) ) ;
AND2    gate4587  (.A(g3956), .B(g2104), .Z(g4171) ) ;
NOR2    gate4588  (.A(g3317), .B(g3328), .Z(g3930) ) ;
AND2    gate4589  (.A(g3930), .B(g1366), .Z(g4172) ) ;
NOR2    gate4590  (.A(g3327), .B(g3336), .Z(g3933) ) ;
AND2    gate4591  (.A(g3933), .B(g1372), .Z(g4177) ) ;
NOR2    gate4592  (.A(g3352), .B(g3360), .Z(g3959) ) ;
AND2    gate4593  (.A(g3959), .B(g2110), .Z(g4178) ) ;
NOR2    gate4594  (.A(g3373), .B(g3376), .Z(g3929) ) ;
AND2    gate4595  (.A(g3929), .B(g2119), .Z(g4180) ) ;
NOR2    gate4596  (.A(g3340), .B(g3351), .Z(g3939) ) ;
AND2    gate4597  (.A(g3939), .B(g1381), .Z(g4181) ) ;
NOR2    gate4598  (.A(g3359), .B(g3367), .Z(g3965) ) ;
AND2    gate4599  (.A(g3965), .B(g1391), .Z(g4183) ) ;
NOR2    gate4600  (.A(g3377), .B(g3379), .Z(g3934) ) ;
AND2    gate4601  (.A(g3934), .B(g2136), .Z(g4184) ) ;
NOR2    gate4602  (.A(g3368), .B(g3374), .Z(g3973) ) ;
AND2    gate4603  (.A(g3973), .B(g1395), .Z(g4186) ) ;
AND2    gate4604  (.A(g628), .B(g3810), .Z(g4199) ) ;
AND2    gate4605  (.A(g3816), .B(g865), .Z(g4209) ) ;
NAND2   gate4606  (.A(g1070), .B(g1084), .Z(g1822) ) ;
AND2    gate4607  (.A(g1822), .B(g4045), .Z(g4214) ) ;
NAND2   gate4608  (.A(II4940), .B(II4941), .Z(g3756) ) ;
AND2    gate4609  (.A(g3756), .B(g1861), .Z(g4230) ) ;
AND2    gate4610  (.A(g654), .B(g3907), .Z(g4236) ) ;
NAND2   gate4611  (.A(II5301), .B(II5302), .Z(g4004) ) ;
AND3    gate4612  (.A(g1749), .B(g4004), .C(g1609), .Z(g4244) ) ;
NAND2   gate4613  (.A(II5308), .B(II5309), .Z(g4007) ) ;
AND3    gate4614  (.A(g1764), .B(g4007), .C(g1628), .Z(g4247) ) ;
AND2    gate4615  (.A(g1861), .B(g3819), .Z(g4253) ) ;
AND3    gate4616  (.A(g2121), .B(g1749), .C(g4004), .Z(g4271) ) ;
AND2    gate4617  (.A(g3936), .B(g942), .Z(g4277) ) ;
AND3    gate4618  (.A(g2138), .B(g1764), .C(g4007), .Z(g4280) ) ;
OR2     gate4619  (.A(g3634), .B(g3089), .Z(g3964) ) ;
AND2    gate4620  (.A(g3964), .B(g3284), .Z(g4333) ) ;
OR2     gate4621  (.A(g3644), .B(g3099), .Z(g3971) ) ;
AND2    gate4622  (.A(g3971), .B(g3289), .Z(g4339) ) ;
OR2     gate4623  (.A(g3646), .B(g3103), .Z(g3972) ) ;
AND2    gate4624  (.A(g3972), .B(g3291), .Z(g4340) ) ;
OR2     gate4625  (.A(g3653), .B(g3113), .Z(g3977) ) ;
AND2    gate4626  (.A(g3977), .B(g3297), .Z(g4341) ) ;
OR2     gate4627  (.A(g3655), .B(g3117), .Z(g3978) ) ;
AND2    gate4628  (.A(g3978), .B(g3299), .Z(g4342) ) ;
OR2     gate4629  (.A(g3661), .B(g3123), .Z(g3981) ) ;
AND2    gate4630  (.A(g3981), .B(g3306), .Z(g4344) ) ;
OR2     gate4631  (.A(g3663), .B(g3127), .Z(g3982) ) ;
AND2    gate4632  (.A(g3982), .B(g3308), .Z(g4345) ) ;
OR2     gate4633  (.A(g3667), .B(g3133), .Z(g3986) ) ;
AND2    gate4634  (.A(g3986), .B(g3320), .Z(g4347) ) ;
OR2     gate4635  (.A(g3669), .B(g3134), .Z(g3987) ) ;
AND2    gate4636  (.A(g3987), .B(g3322), .Z(g4348) ) ;
AND2    gate4637  (.A(g441), .B(g3775), .Z(g4349) ) ;
OR2     gate4638  (.A(g3678), .B(g3143), .Z(g3988) ) ;
AND2    gate4639  (.A(g3988), .B(g3331), .Z(g4352) ) ;
OR2     gate4640  (.A(g3679), .B(g3144), .Z(g3989) ) ;
AND2    gate4641  (.A(g3989), .B(g3332), .Z(g4353) ) ;
AND2    gate4642  (.A(g437), .B(g3777), .Z(g4354) ) ;
AND2    gate4643  (.A(g430), .B(g3778), .Z(g4355) ) ;
OR2     gate4644  (.A(g3684), .B(g3155), .Z(g3990) ) ;
AND2    gate4645  (.A(g3990), .B(g3342), .Z(g4357) ) ;
OR2     gate4646  (.A(g3685), .B(g3156), .Z(g3991) ) ;
AND2    gate4647  (.A(g3991), .B(g3343), .Z(g4358) ) ;
AND2    gate4648  (.A(g434), .B(g3782), .Z(g4359) ) ;
OR2     gate4649  (.A(g3690), .B(g3170), .Z(g3995) ) ;
AND2    gate4650  (.A(g3995), .B(g3354), .Z(g4361) ) ;
OR2     gate4651  (.A(g3691), .B(g3171), .Z(g3996) ) ;
AND2    gate4652  (.A(g3996), .B(g3355), .Z(g4362) ) ;
AND2    gate4653  (.A(g402), .B(g3786), .Z(g4363) ) ;
OR2     gate4654  (.A(g3698), .B(g3180), .Z(g3998) ) ;
AND2    gate4655  (.A(g3998), .B(g3363), .Z(g4368) ) ;
OR2     gate4656  (.A(g3699), .B(g3181), .Z(g3999) ) ;
AND2    gate4657  (.A(g3999), .B(g3364), .Z(g4369) ) ;
AND2    gate4658  (.A(g461), .B(g3789), .Z(g4371) ) ;
AND2    gate4659  (.A(g406), .B(g3790), .Z(g4372) ) ;
OR2     gate4660  (.A(g3702), .B(g3190), .Z(g4001) ) ;
AND2    gate4661  (.A(g4001), .B(g3370), .Z(g4373) ) ;
AND2    gate4662  (.A(g457), .B(g3791), .Z(g4377) ) ;
AND2    gate4663  (.A(g410), .B(g3792), .Z(g4378) ) ;
AND2    gate4664  (.A(g453), .B(g3796), .Z(g4383) ) ;
AND2    gate4665  (.A(g414), .B(g3797), .Z(g4384) ) ;
AND2    gate4666  (.A(g449), .B(g3798), .Z(g4389) ) ;
AND2    gate4667  (.A(g418), .B(g3799), .Z(g4390) ) ;
AND2    gate4668  (.A(g445), .B(g3800), .Z(g4395) ) ;
AND2    gate4669  (.A(g422), .B(g3801), .Z(g4396) ) ;
AND2    gate4670  (.A(g426), .B(g3802), .Z(g4401) ) ;
AND2    gate4671  (.A(g4054), .B(g74), .Z(g4407) ) ;
NOR2    gate4672  (.A(g3505), .B(g471), .Z(g3903) ) ;
NOR2    gate4673  (.A(g760), .B(g754), .Z(g1474) ) ;
NOR2    gate4674  (.A(g3512), .B(g478), .Z(g3905) ) ;
NOR2    gate4675  (.A(g815), .B(g809), .Z(g1481) ) ;
AND3    gate4676  (.A(g923), .B(g4253), .C(g2936), .Z(g4429) ) ;
NOR2    gate4677  (.A(g3763), .B(g3296), .Z(g4239) ) ;
AND2    gate4678  (.A(g4239), .B(g2882), .Z(g4442) ) ;
NOR2    gate4679  (.A(g3780), .B(g3362), .Z(g4235) ) ;
AND2    gate4680  (.A(g4235), .B(g1854), .Z(g4445) ) ;
OR2     gate4681  (.A(g3282), .B(g2659), .Z(g3815) ) ;
AND2    gate4682  (.A(g3815), .B(g4225), .Z(g4448) ) ;
NOR2    gate4683  (.A(g3757), .B(g3283), .Z(g4266) ) ;
AND2    gate4684  (.A(g4266), .B(g2887), .Z(g4449) ) ;
OR2     gate4685  (.A(g3287), .B(g2671), .Z(g3820) ) ;
AND2    gate4686  (.A(g3820), .B(g4227), .Z(g4452) ) ;
NOR2    gate4687  (.A(g3755), .B(g3279), .Z(g4238) ) ;
AND2    gate4688  (.A(g4238), .B(g1858), .Z(g4453) ) ;
OR2     gate4689  (.A(g3294), .B(g3305), .Z(g3829) ) ;
AND2    gate4690  (.A(g3829), .B(g4229), .Z(g4456) ) ;
NOR2    gate4691  (.A(g3762), .B(g3295), .Z(g4261) ) ;
AND2    gate4692  (.A(g4261), .B(g2902), .Z(g4457) ) ;
NOR2    gate4693  (.A(g3759), .B(g3288), .Z(g4245) ) ;
AND2    gate4694  (.A(g4245), .B(g1899), .Z(g4459) ) ;
NOR2    gate4695  (.A(g3774), .B(g3341), .Z(g4241) ) ;
AND2    gate4696  (.A(g4241), .B(g2919), .Z(g4461) ) ;
NOR2    gate4697  (.A(g3767), .B(g3319), .Z(g4272) ) ;
AND2    gate4698  (.A(g4272), .B(g1937), .Z(g4464) ) ;
AND2    gate4699  (.A(g4253), .B(g332), .Z(g4471) ) ;
AND2    gate4700  (.A(g716), .B(g4195), .Z(g4486) ) ;
AND2    gate4701  (.A(g1633), .B(g4202), .Z(g4488) ) ;
AND2    gate4702  (.A(g2166), .B(g4206), .Z(g4489) ) ;
AND2    gate4703  (.A(g2941), .B(g4210), .Z(g4490) ) ;
AND2    gate4704  (.A(g3554), .B(g4215), .Z(g4491) ) ;
OR2     gate4705  (.A(g3449), .B(g2860), .Z(g3913) ) ;
AND2    gate4706  (.A(g3913), .B(g4292), .Z(g4495) ) ;
AND2    gate4707  (.A(g631), .B(g4199), .Z(g4541) ) ;
AND2    gate4708  (.A(g706), .B(g4262), .Z(g4580) ) ;
AND2    gate4709  (.A(g1808), .B(g4267), .Z(g4583) ) ;
AND2    gate4710  (.A(g2419), .B(g4273), .Z(g4588) ) ;
AND2    gate4711  (.A(g3147), .B(g4281), .Z(g4592) ) ;
AND2    gate4712  (.A(g4277), .B(g947), .Z(g4593) ) ;
AND2    gate4713  (.A(g3694), .B(g4286), .Z(g4597) ) ;
AND2    gate4714  (.A(g1978), .B(g4253), .Z(g4598) ) ;
AND2    gate4715  (.A(g4054), .B(g4289), .Z(g4600) ) ;
AND2    gate4716  (.A(g4407), .B(g4293), .Z(g4602) ) ;
NAND3   gate4717  (.A(g1138), .B(g3718), .C(g2142), .Z(g3985) ) ;
NAND2   gate4718  (.A(II5760), .B(II5761), .Z(g4300) ) ;
AND3    gate4719  (.A(g3985), .B(g119), .C(g4300), .Z(g4611) ) ;
OR2     gate4720  (.A(g3997), .B(g4000), .Z(g4231) ) ;
AND2    gate4721  (.A(g4231), .B(g3761), .Z(g4616) ) ;
AND2    gate4722  (.A(g3953), .B(g4364), .Z(g4621) ) ;
AND2    gate4723  (.A(g4407), .B(g79), .Z(g4648) ) ;
OR2     gate4724  (.A(g4344), .B(g3619), .Z(g4637) ) ;
OR2     gate4725  (.A(g4341), .B(g3615), .Z(g4634) ) ;
AND2    gate4726  (.A(g4637), .B(g4634), .Z(g4661) ) ;
OR2     gate4727  (.A(g4339), .B(g3610), .Z(g4630) ) ;
OR2     gate4728  (.A(g4333), .B(g3603), .Z(g4627) ) ;
AND2    gate4729  (.A(g4630), .B(g4627), .Z(g4666) ) ;
OR2     gate4730  (.A(g4361), .B(g3652), .Z(g4653) ) ;
OR2     gate4731  (.A(g4357), .B(g3643), .Z(g4651) ) ;
AND2    gate4732  (.A(g4653), .B(g4651), .Z(g4667) ) ;
OR2     gate4733  (.A(g4348), .B(g3628), .Z(g4642) ) ;
OR2     gate4734  (.A(g4345), .B(g3620), .Z(g4638) ) ;
AND2    gate4735  (.A(g4642), .B(g4638), .Z(g4668) ) ;
OR2     gate4736  (.A(g4352), .B(g3633), .Z(g4645) ) ;
OR2     gate4737  (.A(g4347), .B(g3627), .Z(g4641) ) ;
AND2    gate4738  (.A(g4645), .B(g4641), .Z(g4671) ) ;
OR2     gate4739  (.A(g4342), .B(g3616), .Z(g4635) ) ;
OR2     gate4740  (.A(g4340), .B(g3611), .Z(g4631) ) ;
AND2    gate4741  (.A(g4635), .B(g4631), .Z(g4672) ) ;
OR2     gate4742  (.A(g4369), .B(g3662), .Z(g4656) ) ;
OR2     gate4743  (.A(g4362), .B(g3654), .Z(g4654) ) ;
AND2    gate4744  (.A(g4656), .B(g4654), .Z(g4673) ) ;
OR2     gate4745  (.A(g4358), .B(g3645), .Z(g4652) ) ;
OR2     gate4746  (.A(g4353), .B(g3635), .Z(g4646) ) ;
AND2    gate4747  (.A(g4652), .B(g4646), .Z(g4677) ) ;
NOR2    gate4748  (.A(g4171), .B(g4177), .Z(g4585) ) ;
AND2    gate4749  (.A(g4585), .B(g2066), .Z(g4683) ) ;
NOR2    gate4750  (.A(g4164), .B(g4168), .Z(g4584) ) ;
AND2    gate4751  (.A(g4584), .B(g1341), .Z(g4684) ) ;
NOR2    gate4752  (.A(g4178), .B(g4181), .Z(g4591) ) ;
AND2    gate4753  (.A(g4591), .B(g2079), .Z(g4685) ) ;
NOR2    gate4754  (.A(g4169), .B(g4172), .Z(g4590) ) ;
AND2    gate4755  (.A(g4590), .B(g1348), .Z(g4686) ) ;
NOR2    gate4756  (.A(g4233), .B(g3924), .Z(g4568) ) ;
AND2    gate4757  (.A(g1474), .B(g4568), .Z(g4688) ) ;
NOR2    gate4758  (.A(g4156), .B(g4160), .Z(g4581) ) ;
AND2    gate4759  (.A(g4581), .B(g2098), .Z(g4691) ) ;
NOR2    gate4760  (.A(g4234), .B(g3928), .Z(g4578) ) ;
AND2    gate4761  (.A(g1481), .B(g4578), .Z(g4694) ) ;
NOR2    gate4762  (.A(g4180), .B(g4183), .Z(g4589) ) ;
AND2    gate4763  (.A(g4589), .B(g1363), .Z(g4697) ) ;
NOR2    gate4764  (.A(g4161), .B(g4165), .Z(g4586) ) ;
AND2    gate4765  (.A(g4586), .B(g2106), .Z(g4698) ) ;
NOR2    gate4766  (.A(g4184), .B(g4186), .Z(g4596) ) ;
AND2    gate4767  (.A(g4596), .B(g1378), .Z(g4701) ) ;
AND2    gate4768  (.A(g578), .B(g4541), .Z(g4708) ) ;
AND2    gate4769  (.A(g1423), .B(g4565), .Z(g4730) ) ;
AND2    gate4770  (.A(g2018), .B(g4577), .Z(g4735) ) ;
AND2    gate4771  (.A(g2850), .B(g4579), .Z(g4739) ) ;
AND2    gate4772  (.A(g3434), .B(g4582), .Z(g4744) ) ;
AND2    gate4773  (.A(g3816), .B(g4587), .Z(g4756) ) ;
OR2     gate4774  (.A(g4243), .B(g2010), .Z(g4500) ) ;
AND2    gate4775  (.A(g536), .B(g4500), .Z(g4759) ) ;
AND2    gate4776  (.A(g1624), .B(g4623), .Z(g4782) ) ;
AND2    gate4777  (.A(g2160), .B(g4625), .Z(g4785) ) ;
AND2    gate4778  (.A(g2937), .B(g4628), .Z(g4787) ) ;
AND2    gate4779  (.A(g3551), .B(g4632), .Z(g4789) ) ;
AND2    gate4780  (.A(g3936), .B(g4636), .Z(g4791) ) ;
NAND2   gate4781  (.A(g873), .B(g889), .Z(g1417) ) ;
AND2    gate4782  (.A(g1417), .B(g4471), .Z(g4792) ) ;
AND2    gate4783  (.A(g4277), .B(g4639), .Z(g4793) ) ;
AND2    gate4784  (.A(g4593), .B(g949), .Z(g4794) ) ;
AND2    gate4785  (.A(g4593), .B(g4643), .Z(g4797) ) ;
AND2    gate4786  (.A(g4648), .B(g4296), .Z(g4800) ) ;
AND2    gate4787  (.A(g4209), .B(g4463), .Z(g4826) ) ;
AND2    gate4788  (.A(g4520), .B(g4515), .Z(g4827) ) ;
AND2    gate4789  (.A(g4510), .B(g4508), .Z(g4828) ) ;
AND2    gate4790  (.A(g4526), .B(g4522), .Z(g4829) ) ;
AND2    gate4791  (.A(g4529), .B(g4525), .Z(g4830) ) ;
AND2    gate4792  (.A(g4528), .B(g4524), .Z(g4831) ) ;
AND2    gate4793  (.A(g4517), .B(g4512), .Z(g4832) ) ;
AND2    gate4794  (.A(g4521), .B(g4516), .Z(g4833) ) ;
AND2    gate4795  (.A(g4534), .B(g4531), .Z(g4834) ) ;
AND2    gate4796  (.A(g4533), .B(g4530), .Z(g4835) ) ;
AND2    gate4797  (.A(g4527), .B(g4523), .Z(g4836) ) ;
AND2    gate4798  (.A(g4648), .B(g84), .Z(g4838) ) ;
NOR2    gate4799  (.A(g4457), .B(g4459), .Z(g4777) ) ;
AND2    gate4800  (.A(g4777), .B(g2874), .Z(g4863) ) ;
NOR2    gate4801  (.A(g4449), .B(g4453), .Z(g4776) ) ;
AND2    gate4802  (.A(g4776), .B(g1849), .Z(g4865) ) ;
OR2     gate4803  (.A(g4429), .B(g4432), .Z(g4811) ) ;
AND2    gate4804  (.A(g4811), .B(g3872), .Z(g4867) ) ;
NOR2    gate4805  (.A(g4442), .B(g4445), .Z(g4774) ) ;
AND2    gate4806  (.A(g4774), .B(g2891), .Z(g4868) ) ;
NOR2    gate4807  (.A(g4461), .B(g4464), .Z(g4779) ) ;
AND2    gate4808  (.A(g4779), .B(g1884), .Z(g4870) ) ;
AND2    gate4809  (.A(g4838), .B(g4173), .Z(g4873) ) ;
AND2    gate4810  (.A(g582), .B(g4708), .Z(g4874) ) ;
AND2    gate4811  (.A(g148), .B(g4723), .Z(g4928) ) ;
AND2    gate4812  (.A(g157), .B(g4727), .Z(g4932) ) ;
AND2    gate4813  (.A(g166), .B(g4732), .Z(g4937) ) ;
AND2    gate4814  (.A(g175), .B(g4736), .Z(g4942) ) ;
AND2    gate4815  (.A(g184), .B(g4741), .Z(g4947) ) ;
AND2    gate4816  (.A(g193), .B(g4753), .Z(g4949) ) ;
OR2     gate4817  (.A(g3464), .B(g2868), .Z(g3935) ) ;
AND2    gate4818  (.A(g3935), .B(g4804), .Z(g5023) ) ;
OR2     gate4819  (.A(g3479), .B(g2873), .Z(g3941) ) ;
AND2    gate4820  (.A(g3941), .B(g4805), .Z(g5043) ) ;
OR2     gate4821  (.A(g3484), .B(g3489), .Z(g3954) ) ;
AND2    gate4822  (.A(g3954), .B(g4806), .Z(g5047) ) ;
OR2     gate4823  (.A(g3490), .B(g3887), .Z(g4285) ) ;
OR2     gate4824  (.A(g3499), .B(g4230), .Z(g4599) ) ;
AND2    gate4825  (.A(g4599), .B(g4808), .Z(g5053) ) ;
AND2    gate4826  (.A(g4794), .B(g951), .Z(g5095) ) ;
AND2    gate4827  (.A(g4794), .B(g4647), .Z(g5096) ) ;
OR2     gate4828  (.A(g3558), .B(g2949), .Z(g4021) ) ;
AND2    gate4829  (.A(g4021), .B(g4837), .Z(g5098) ) ;
AND2    gate4830  (.A(g193), .B(g4662), .Z(g5122) ) ;
NAND2   gate4831  (.A(g4611), .B(g3528), .Z(g4670) ) ;
AND2    gate4832  (.A(g4670), .B(g1936), .Z(g5123) ) ;
AND2    gate4833  (.A(g148), .B(g5099), .Z(g5142) ) ;
AND2    gate4834  (.A(g157), .B(g5099), .Z(g5143) ) ;
AND2    gate4835  (.A(g166), .B(g5099), .Z(g5144) ) ;
AND2    gate4836  (.A(g175), .B(g5099), .Z(g5145) ) ;
AND2    gate4837  (.A(g184), .B(g5099), .Z(g5146) ) ;
NOR2    gate4838  (.A(g1472), .B(g4680), .Z(g4950) ) ;
AND2    gate4839  (.A(g430), .B(g4950), .Z(g5152) ) ;
AND2    gate4840  (.A(g492), .B(g4904), .Z(g5153) ) ;
NOR2    gate4841  (.A(g4674), .B(g1477), .Z(g4993) ) ;
AND2    gate4842  (.A(g500), .B(g4993), .Z(g5154) ) ;
NOR2    gate4843  (.A(g952), .B(g4680), .Z(g4877) ) ;
AND2    gate4844  (.A(g434), .B(g4877), .Z(g5156) ) ;
AND2    gate4845  (.A(g496), .B(g4904), .Z(g5157) ) ;
AND2    gate4846  (.A(g504), .B(g4993), .Z(g5158) ) ;
NOR2    gate4847  (.A(g4674), .B(g952), .Z(g4967) ) ;
AND2    gate4848  (.A(g536), .B(g4967), .Z(g5159) ) ;
AND2    gate4849  (.A(g5095), .B(g4535), .Z(g5161) ) ;
NOR2    gate4850  (.A(g4691), .B(g4697), .Z(g5088) ) ;
AND2    gate4851  (.A(g5088), .B(g2105), .Z(g5162) ) ;
AND2    gate4852  (.A(g402), .B(g4950), .Z(g5163) ) ;
AND2    gate4853  (.A(g437), .B(g4877), .Z(g5164) ) ;
AND2    gate4854  (.A(g508), .B(g4993), .Z(g5165) ) ;
AND2    gate4855  (.A(g541), .B(g4967), .Z(g5166) ) ;
NOR2    gate4856  (.A(g4683), .B(g4684), .Z(g5093) ) ;
AND2    gate4857  (.A(g5093), .B(g1375), .Z(g5169) ) ;
NOR2    gate4858  (.A(g4698), .B(g4701), .Z(g5091) ) ;
AND2    gate4859  (.A(g5091), .B(g2111), .Z(g5170) ) ;
AND2    gate4860  (.A(g406), .B(g4950), .Z(g5171) ) ;
AND2    gate4861  (.A(g441), .B(g4877), .Z(g5172) ) ;
AND2    gate4862  (.A(g512), .B(g4993), .Z(g5173) ) ;
NOR2    gate4863  (.A(g4685), .B(g4686), .Z(g5094) ) ;
AND2    gate4864  (.A(g5094), .B(g1384), .Z(g5175) ) ;
AND2    gate4865  (.A(g410), .B(g4950), .Z(g5176) ) ;
AND2    gate4866  (.A(g445), .B(g4877), .Z(g5177) ) ;
AND2    gate4867  (.A(g516), .B(g4993), .Z(g5178) ) ;
AND2    gate4868  (.A(g414), .B(g4950), .Z(g5180) ) ;
AND2    gate4869  (.A(g449), .B(g4877), .Z(g5181) ) ;
AND2    gate4870  (.A(g520), .B(g4993), .Z(g5182) ) ;
AND2    gate4871  (.A(g418), .B(g4950), .Z(g5183) ) ;
AND2    gate4872  (.A(g453), .B(g4877), .Z(g5184) ) ;
AND2    gate4873  (.A(g524), .B(g4993), .Z(g5185) ) ;
AND2    gate4874  (.A(g422), .B(g4950), .Z(g5186) ) ;
AND2    gate4875  (.A(g457), .B(g4877), .Z(g5187) ) ;
AND2    gate4876  (.A(g1043), .B(g4894), .Z(g5188) ) ;
AND2    gate4877  (.A(g528), .B(g4993), .Z(g5189) ) ;
AND2    gate4878  (.A(g426), .B(g4950), .Z(g5190) ) ;
AND2    gate4879  (.A(g461), .B(g4877), .Z(g5191) ) ;
AND2    gate4880  (.A(g1046), .B(g4894), .Z(g5192) ) ;
AND2    gate4881  (.A(g532), .B(g4967), .Z(g5193) ) ;
AND2    gate4882  (.A(g586), .B(g4874), .Z(g5194) ) ;
AND2    gate4883  (.A(g465), .B(g4967), .Z(g5197) ) ;
AND2    gate4884  (.A(g558), .B(g5025), .Z(g5198) ) ;
AND2    gate4885  (.A(g559), .B(g5025), .Z(g5200) ) ;
OR2     gate4886  (.A(g4730), .B(g4486), .Z(g4859) ) ;
AND2    gate4887  (.A(g4859), .B(g5084), .Z(g5201) ) ;
AND2    gate4888  (.A(g560), .B(g5025), .Z(g5209) ) ;
OR2     gate4889  (.A(g4735), .B(g4488), .Z(g4860) ) ;
AND2    gate4890  (.A(g4860), .B(g5086), .Z(g5211) ) ;
AND2    gate4891  (.A(g561), .B(g5025), .Z(g5212) ) ;
OR2     gate4892  (.A(g4739), .B(g4489), .Z(g4862) ) ;
AND2    gate4893  (.A(g4862), .B(g5087), .Z(g5213) ) ;
AND2    gate4894  (.A(g562), .B(g5025), .Z(g5214) ) ;
OR2     gate4895  (.A(g4744), .B(g4490), .Z(g4864) ) ;
AND2    gate4896  (.A(g4864), .B(g5090), .Z(g5215) ) ;
AND2    gate4897  (.A(g563), .B(g5025), .Z(g5216) ) ;
OR2     gate4898  (.A(g4756), .B(g4491), .Z(g4866) ) ;
AND2    gate4899  (.A(g4866), .B(g5092), .Z(g5217) ) ;
AND2    gate4900  (.A(g564), .B(g5025), .Z(g5218) ) ;
AND2    gate4901  (.A(g669), .B(g5054), .Z(g5225) ) ;
AND2    gate4902  (.A(g672), .B(g5054), .Z(g5226) ) ;
AND2    gate4903  (.A(g545), .B(g4980), .Z(g5229) ) ;
AND2    gate4904  (.A(g548), .B(g4980), .Z(g5232) ) ;
AND2    gate4905  (.A(g551), .B(g4980), .Z(g5233) ) ;
AND2    gate4906  (.A(g197), .B(g4915), .Z(g5234) ) ;
AND2    gate4907  (.A(g554), .B(g4980), .Z(g5235) ) ;
AND2    gate4908  (.A(g269), .B(g4915), .Z(g5236) ) ;
AND2    gate4909  (.A(g293), .B(g4915), .Z(g5240) ) ;
AND2    gate4910  (.A(g297), .B(g4915), .Z(g5245) ) ;
AND2    gate4911  (.A(g557), .B(g5025), .Z(g5269) ) ;
OR2     gate4912  (.A(g4826), .B(g4621), .Z(g5013) ) ;
OR2     gate4913  (.A(g4214), .B(g3831), .Z(g4468) ) ;
AND2    gate4914  (.A(g5013), .B(g4468), .Z(g5311) ) ;
AND2    gate4915  (.A(g148), .B(g4869), .Z(g5317) ) ;
NOR3    gate4916  (.A(g5069), .B(g4410), .C(g766), .Z(g5324) ) ;
AND2    gate4917  (.A(g5324), .B(g3451), .Z(g5349) ) ;
NOR3    gate4918  (.A(g5077), .B(g4416), .C(g821), .Z(g5325) ) ;
AND2    gate4919  (.A(g5325), .B(g3453), .Z(g5350) ) ;
OR3     gate4920  (.A(g5069), .B(g4410), .C(g3012), .Z(g5326) ) ;
AND2    gate4921  (.A(g5326), .B(g3459), .Z(g5351) ) ;
OR3     gate4922  (.A(g5077), .B(g4416), .C(g3028), .Z(g5327) ) ;
AND2    gate4923  (.A(g5327), .B(g3463), .Z(g5353) ) ;
NOR2    gate4924  (.A(g4868), .B(g4870), .Z(g5249) ) ;
AND2    gate4925  (.A(g5249), .B(g2903), .Z(g5354) ) ;
NOR2    gate4926  (.A(g4863), .B(g4865), .Z(g5265) ) ;
AND2    gate4927  (.A(g5265), .B(g1902), .Z(g5356) ) ;
AND2    gate4928  (.A(g398), .B(g5220), .Z(g5357) ) ;
AND2    gate4929  (.A(g4428), .B(g5155), .Z(g5359) ) ;
AND2    gate4930  (.A(g4431), .B(g5160), .Z(g5360) ) ;
AND2    gate4931  (.A(g4435), .B(g5168), .Z(g5361) ) ;
AND2    gate4932  (.A(g4437), .B(g5174), .Z(g5362) ) ;
AND2    gate4933  (.A(g4439), .B(g5179), .Z(g5363) ) ;
AND2    gate4934  (.A(g574), .B(g5194), .Z(g5364) ) ;
AND2    gate4935  (.A(g143), .B(g5247), .Z(g5369) ) ;
AND2    gate4936  (.A(g152), .B(g5248), .Z(g5371) ) ;
AND2    gate4937  (.A(g161), .B(g5250), .Z(g5373) ) ;
AND2    gate4938  (.A(g170), .B(g5255), .Z(g5376) ) ;
AND2    gate4939  (.A(g179), .B(g5260), .Z(g5378) ) ;
AND2    gate4940  (.A(g188), .B(g5264), .Z(g5380) ) ;
AND2    gate4941  (.A(g366), .B(g5261), .Z(g5398) ) ;
AND2    gate4942  (.A(g370), .B(g5266), .Z(g5402) ) ;
AND2    gate4943  (.A(g374), .B(g5270), .Z(g5406) ) ;
AND2    gate4944  (.A(g378), .B(g5274), .Z(g5410) ) ;
AND2    gate4945  (.A(g382), .B(g5278), .Z(g5414) ) ;
AND2    gate4946  (.A(g386), .B(g5292), .Z(g5419) ) ;
AND2    gate4947  (.A(g390), .B(g5296), .Z(g5424) ) ;
AND2    gate4948  (.A(g394), .B(g5300), .Z(g5428) ) ;
AND2    gate4949  (.A(g398), .B(g5304), .Z(g5429) ) ;
OR2     gate4950  (.A(g5123), .B(g3630), .Z(g5224) ) ;
AND2    gate4951  (.A(g5224), .B(g3769), .Z(g5438) ) ;
NAND2   gate4952  (.A(II2527), .B(II2528), .Z(g1558) ) ;
AND3    gate4953  (.A(g4537), .B(g5251), .C(g1558), .Z(g5441) ) ;
NAND2   gate4954  (.A(II3446), .B(II3447), .Z(g2307) ) ;
AND3    gate4955  (.A(g4537), .B(g5251), .C(g2307), .Z(g5443) ) ;
NAND2   gate4956  (.A(II2543), .B(II2544), .Z(g1574) ) ;
AND3    gate4957  (.A(g4545), .B(g5256), .C(g1574), .Z(g5444) ) ;
OR2     gate4958  (.A(g5069), .B(g2067), .Z(g5241) ) ;
AND2    gate4959  (.A(g4537), .B(g5241), .Z(g5446) ) ;
NAND2   gate4960  (.A(II3456), .B(II3457), .Z(g2311) ) ;
AND3    gate4961  (.A(g4545), .B(g5256), .C(g2311), .Z(g5447) ) ;
OR2     gate4962  (.A(g5077), .B(g2080), .Z(g5246) ) ;
AND2    gate4963  (.A(g4545), .B(g5246), .Z(g5449) ) ;
OR2     gate4964  (.A(g4410), .B(g2995), .Z(g4544) ) ;
AND2    gate4965  (.A(g5251), .B(g4544), .Z(g5451) ) ;
OR2     gate4966  (.A(g4416), .B(g3013), .Z(g4549) ) ;
AND2    gate4967  (.A(g5256), .B(g4549), .Z(g5454) ) ;
AND2    gate4968  (.A(g366), .B(g5331), .Z(g5481) ) ;
AND2    gate4969  (.A(g370), .B(g5331), .Z(g5482) ) ;
AND2    gate4970  (.A(g374), .B(g5331), .Z(g5483) ) ;
AND2    gate4971  (.A(g378), .B(g5331), .Z(g5484) ) ;
AND2    gate4972  (.A(g382), .B(g5331), .Z(g5485) ) ;
AND2    gate4973  (.A(g386), .B(g5331), .Z(g5486) ) ;
AND2    gate4974  (.A(g390), .B(g5331), .Z(g5487) ) ;
AND2    gate4975  (.A(g394), .B(g5331), .Z(g5488) ) ;
AND2    gate4976  (.A(g5441), .B(g3452), .Z(g5492) ) ;
AND2    gate4977  (.A(g5443), .B(g3455), .Z(g5494) ) ;
AND2    gate4978  (.A(g5444), .B(g3456), .Z(g5495) ) ;
AND2    gate4979  (.A(g5446), .B(g3457), .Z(g5496) ) ;
AND2    gate4980  (.A(g5447), .B(g3458), .Z(g5497) ) ;
AND2    gate4981  (.A(g5449), .B(g3460), .Z(g5498) ) ;
AND2    gate4982  (.A(g5451), .B(g3462), .Z(g5499) ) ;
OR2     gate4983  (.A(g5161), .B(g4873), .Z(g5430) ) ;
OR2     gate4984  (.A(g4792), .B(g4598), .Z(g5074) ) ;
AND2    gate4985  (.A(g5430), .B(g5074), .Z(g5500) ) ;
AND2    gate4986  (.A(g5454), .B(g3478), .Z(g5501) ) ;
AND2    gate4987  (.A(g366), .B(g5384), .Z(g5503) ) ;
AND2    gate4988  (.A(g590), .B(g5364), .Z(g5515) ) ;
OR2     gate4989  (.A(g4782), .B(g4580), .Z(g5012) ) ;
AND2    gate4990  (.A(g5012), .B(g5440), .Z(g5553) ) ;
OR2     gate4991  (.A(g4785), .B(g4583), .Z(g5014) ) ;
AND2    gate4992  (.A(g5014), .B(g5442), .Z(g5555) ) ;
OR2     gate4993  (.A(g4787), .B(g4588), .Z(g5015) ) ;
AND2    gate4994  (.A(g5015), .B(g5445), .Z(g5556) ) ;
OR2     gate4995  (.A(g4789), .B(g4592), .Z(g5016) ) ;
AND2    gate4996  (.A(g5016), .B(g5448), .Z(g5557) ) ;
OR2     gate4997  (.A(g4791), .B(g4597), .Z(g5018) ) ;
AND2    gate4998  (.A(g5018), .B(g5450), .Z(g5558) ) ;
OR2     gate4999  (.A(g4793), .B(g4600), .Z(g5024) ) ;
AND2    gate5000  (.A(g5024), .B(g5453), .Z(g5559) ) ;
OR2     gate5001  (.A(g4797), .B(g4602), .Z(g5044) ) ;
AND2    gate5002  (.A(g5044), .B(g5456), .Z(g5560) ) ;
OR2     gate5003  (.A(g5096), .B(g4800), .Z(g5228) ) ;
AND2    gate5004  (.A(g5228), .B(g5457), .Z(g5562) ) ;
OR2     gate5005  (.A(g5317), .B(g5122), .Z(g5348) ) ;
AND2    gate5006  (.A(g5348), .B(g3772), .Z(g5569) ) ;
AND2    gate5007  (.A(g5046), .B(g5509), .Z(g5598) ) ;
AND2    gate5008  (.A(g5049), .B(g5512), .Z(g5599) ) ;
NAND2   gate5009  (.A(II7209), .B(II7210), .Z(g5502) ) ;
AND2    gate5010  (.A(g5502), .B(g4900), .Z(g5600) ) ;
AND2    gate5011  (.A(g5052), .B(g5518), .Z(g5601) ) ;
NAND2   gate5012  (.A(II7217), .B(II7218), .Z(g5504) ) ;
AND2    gate5013  (.A(g5504), .B(g4911), .Z(g5603) ) ;
AND2    gate5014  (.A(g5059), .B(g5521), .Z(g5604) ) ;
NAND2   gate5015  (.A(II7224), .B(II7225), .Z(g5505) ) ;
AND2    gate5016  (.A(g5505), .B(g4929), .Z(g5616) ) ;
AND2    gate5017  (.A(g5061), .B(g5524), .Z(g5617) ) ;
NAND2   gate5018  (.A(II7231), .B(II7232), .Z(g5506) ) ;
AND2    gate5019  (.A(g5506), .B(g4933), .Z(g5618) ) ;
AND2    gate5020  (.A(g5064), .B(g5527), .Z(g5619) ) ;
NAND2   gate5021  (.A(II7238), .B(II7239), .Z(g5507) ) ;
AND2    gate5022  (.A(g5507), .B(g4938), .Z(g5620) ) ;
NAND2   gate5023  (.A(II7245), .B(II7246), .Z(g5508) ) ;
AND2    gate5024  (.A(g5508), .B(g4943), .Z(g5621) ) ;
AND2    gate5025  (.A(g4494), .B(g5538), .Z(g5632) ) ;
AND2    gate5026  (.A(g4496), .B(g5539), .Z(g5633) ) ;
AND2    gate5027  (.A(g4498), .B(g5542), .Z(g5635) ) ;
AND2    gate5028  (.A(g4499), .B(g5543), .Z(g5637) ) ;
AND2    gate5029  (.A(g4502), .B(g5544), .Z(g5646) ) ;
AND2    gate5030  (.A(g4507), .B(g5545), .Z(g5648) ) ;
AND2    gate5031  (.A(g4509), .B(g5549), .Z(g5660) ) ;
AND2    gate5032  (.A(g4513), .B(g5550), .Z(g5663) ) ;
AND2    gate5033  (.A(g361), .B(g5570), .Z(g5665) ) ;
AND2    gate5034  (.A(g49), .B(g5571), .Z(g5668) ) ;
AND2    gate5035  (.A(g54), .B(g5572), .Z(g5671) ) ;
AND2    gate5036  (.A(g59), .B(g5573), .Z(g5673) ) ;
AND2    gate5037  (.A(g64), .B(g5574), .Z(g5675) ) ;
AND2    gate5038  (.A(g69), .B(g5575), .Z(g5677) ) ;
AND2    gate5039  (.A(g74), .B(g5576), .Z(g5679) ) ;
AND2    gate5040  (.A(g79), .B(g5577), .Z(g5681) ) ;
AND2    gate5041  (.A(g84), .B(g5578), .Z(g5682) ) ;
NAND2   gate5042  (.A(II7433), .B(II7434), .Z(g5683) ) ;
OR2     gate5043  (.A(g5503), .B(g5357), .Z(g5623) ) ;
AND2    gate5044  (.A(g5623), .B(g3889), .Z(g5728) ) ;
AND2    gate5045  (.A(g5824), .B(g3752), .Z(g5883) ) ;
OR2     gate5046  (.A(g5369), .B(g5600), .Z(g5800) ) ;
AND2    gate5047  (.A(g5800), .B(g5647), .Z(g5898) ) ;
OR2     gate5048  (.A(g5371), .B(g5603), .Z(g5804) ) ;
AND2    gate5049  (.A(g5804), .B(g5658), .Z(g5900) ) ;
OR2     gate5050  (.A(g5373), .B(g5616), .Z(g5808) ) ;
AND2    gate5051  (.A(g5808), .B(g5661), .Z(g5902) ) ;
OR2     gate5052  (.A(g5376), .B(g5618), .Z(g5812) ) ;
AND2    gate5053  (.A(g5812), .B(g5664), .Z(g5904) ) ;
AND2    gate5054  (.A(g5787), .B(g3384), .Z(g5909) ) ;
OR2     gate5055  (.A(g5378), .B(g5620), .Z(g5816) ) ;
AND2    gate5056  (.A(g5816), .B(g5667), .Z(g5910) ) ;
OR2     gate5057  (.A(g5380), .B(g5621), .Z(g5817) ) ;
AND2    gate5058  (.A(g5817), .B(g5670), .Z(g5911) ) ;
AND2    gate5059  (.A(g5112), .B(g5784), .Z(g5935) ) ;
AND2    gate5060  (.A(g5113), .B(g5788), .Z(g5936) ) ;
NAND2   gate5061  (.A(II7521), .B(II7522), .Z(g5775) ) ;
AND2    gate5062  (.A(g5775), .B(g5392), .Z(g5937) ) ;
AND2    gate5063  (.A(g5114), .B(g5791), .Z(g5938) ) ;
NAND2   gate5064  (.A(II7528), .B(II7529), .Z(g5776) ) ;
AND2    gate5065  (.A(g5776), .B(g5395), .Z(g5939) ) ;
AND2    gate5066  (.A(g5115), .B(g5794), .Z(g5940) ) ;
NAND2   gate5067  (.A(II7535), .B(II7536), .Z(g5777) ) ;
AND2    gate5068  (.A(g5777), .B(g5399), .Z(g5941) ) ;
AND2    gate5069  (.A(g5117), .B(g5797), .Z(g5942) ) ;
NAND2   gate5070  (.A(II7542), .B(II7543), .Z(g5778) ) ;
AND2    gate5071  (.A(g5778), .B(g5403), .Z(g5944) ) ;
AND2    gate5072  (.A(g5118), .B(g5801), .Z(g5945) ) ;
NAND2   gate5073  (.A(II7549), .B(II7550), .Z(g5779) ) ;
AND2    gate5074  (.A(g5779), .B(g5407), .Z(g5948) ) ;
AND2    gate5075  (.A(g5119), .B(g5805), .Z(g5949) ) ;
NAND2   gate5076  (.A(II7556), .B(II7557), .Z(g5780) ) ;
AND2    gate5077  (.A(g5780), .B(g5411), .Z(g5951) ) ;
AND2    gate5078  (.A(g5120), .B(g5809), .Z(g5952) ) ;
NAND2   gate5079  (.A(II7563), .B(II7564), .Z(g5781) ) ;
AND2    gate5080  (.A(g5781), .B(g5415), .Z(g5953) ) ;
AND2    gate5081  (.A(g5121), .B(g5813), .Z(g5954) ) ;
NAND2   gate5082  (.A(II7570), .B(II7571), .Z(g5782) ) ;
AND2    gate5083  (.A(g5782), .B(g5420), .Z(g5955) ) ;
NAND2   gate5084  (.A(II7577), .B(II7578), .Z(g5783) ) ;
AND2    gate5085  (.A(g5783), .B(g5425), .Z(g5956) ) ;
AND2    gate5086  (.A(g5824), .B(g1692), .Z(g6047) ) ;
AND2    gate5087  (.A(g5824), .B(g1696), .Z(g6055) ) ;
AND2    gate5088  (.A(g5824), .B(g1699), .Z(g6056) ) ;
AND2    gate5089  (.A(g5824), .B(g1703), .Z(g6060) ) ;
AND2    gate5090  (.A(g5824), .B(g1711), .Z(g6061) ) ;
AND2    gate5091  (.A(g5824), .B(g1721), .Z(g6066) ) ;
AND2    gate5092  (.A(g5824), .B(g1726), .Z(g6068) ) ;
AND2    gate5093  (.A(g5824), .B(g1735), .Z(g6077) ) ;
AND2    gate5094  (.A(g1236), .B(g5753), .Z(g6079) ) ;
AND2    gate5095  (.A(g1177), .B(g5731), .Z(g6081) ) ;
AND2    gate5096  (.A(g1123), .B(g5742), .Z(g6082) ) ;
AND2    gate5097  (.A(g1123), .B(g5753), .Z(g6084) ) ;
AND2    gate5098  (.A(g1161), .B(g5731), .Z(g6085) ) ;
AND2    gate5099  (.A(g1143), .B(g5742), .Z(g6086) ) ;
AND2    gate5100  (.A(g1143), .B(g5753), .Z(g6088) ) ;
AND2    gate5101  (.A(g1143), .B(g5731), .Z(g6089) ) ;
AND2    gate5102  (.A(g1161), .B(g5742), .Z(g6090) ) ;
AND2    gate5103  (.A(g1161), .B(g5753), .Z(g6091) ) ;
AND2    gate5104  (.A(g1123), .B(g5731), .Z(g6092) ) ;
AND2    gate5105  (.A(g1177), .B(g5742), .Z(g6093) ) ;
AND2    gate5106  (.A(g1177), .B(g5753), .Z(g6094) ) ;
AND2    gate5107  (.A(g1193), .B(g5753), .Z(g6096) ) ;
AND2    gate5108  (.A(g1209), .B(g5753), .Z(g6098) ) ;
AND2    gate5109  (.A(g1222), .B(g5753), .Z(g6099) ) ;
AND2    gate5110  (.A(g5702), .B(g5958), .Z(g6123) ) ;
AND2    gate5111  (.A(g5705), .B(g5958), .Z(g6124) ) ;
AND2    gate5112  (.A(g5708), .B(g5975), .Z(g6125) ) ;
AND2    gate5113  (.A(g5711), .B(g5958), .Z(g6126) ) ;
AND2    gate5114  (.A(g5714), .B(g5975), .Z(g6127) ) ;
AND2    gate5115  (.A(g5590), .B(g5958), .Z(g6128) ) ;
AND2    gate5116  (.A(g5717), .B(g5975), .Z(g6129) ) ;
AND2    gate5117  (.A(g5720), .B(g5958), .Z(g6130) ) ;
AND2    gate5118  (.A(g5593), .B(g5975), .Z(g6131) ) ;
AND2    gate5119  (.A(g3752), .B(g5880), .Z(g6132) ) ;
AND2    gate5120  (.A(g5723), .B(g5975), .Z(g6133) ) ;
AND2    gate5121  (.A(g5584), .B(g5958), .Z(g6135) ) ;
AND2    gate5122  (.A(g5587), .B(g5975), .Z(g6140) ) ;
AND2    gate5123  (.A(g3173), .B(g5997), .Z(g6141) ) ;
AND2    gate5124  (.A(g3183), .B(g5997), .Z(g6144) ) ;
AND2    gate5125  (.A(g3187), .B(g6015), .Z(g6145) ) ;
AND2    gate5126  (.A(g3192), .B(g5997), .Z(g6146) ) ;
AND2    gate5127  (.A(g3196), .B(g6015), .Z(g6148) ) ;
AND2    gate5128  (.A(g3200), .B(g5997), .Z(g6149) ) ;
AND2    gate5129  (.A(g3204), .B(g6015), .Z(g6150) ) ;
AND2    gate5130  (.A(g3209), .B(g5997), .Z(g6151) ) ;
AND2    gate5131  (.A(g3212), .B(g6015), .Z(g6152) ) ;
AND2    gate5132  (.A(g3216), .B(g5997), .Z(g6153) ) ;
AND2    gate5133  (.A(g3219), .B(g6015), .Z(g6154) ) ;
AND2    gate5134  (.A(g2588), .B(g5997), .Z(g6155) ) ;
AND2    gate5135  (.A(g2591), .B(g6015), .Z(g6156) ) ;
AND2    gate5136  (.A(g3158), .B(g5997), .Z(g6157) ) ;
AND2    gate5137  (.A(g2594), .B(g6015), .Z(g6158) ) ;
AND2    gate5138  (.A(g3177), .B(g6015), .Z(g6159) ) ;
AND2    gate5139  (.A(g528), .B(g5886), .Z(g6238) ) ;
OR2     gate5140  (.A(g3843), .B(g541), .Z(g4205) ) ;
AND2    gate5141  (.A(g4205), .B(g5888), .Z(g6240) ) ;
AND2    gate5142  (.A(g1325), .B(g5887), .Z(g6241) ) ;
AND2    gate5143  (.A(g500), .B(g5890), .Z(g6243) ) ;
AND2    gate5144  (.A(g4759), .B(g5891), .Z(g6244) ) ;
AND2    gate5145  (.A(g1329), .B(g5889), .Z(g6245) ) ;
AND2    gate5146  (.A(g504), .B(g5893), .Z(g6247) ) ;
AND2    gate5147  (.A(g465), .B(g5894), .Z(g6248) ) ;
AND2    gate5148  (.A(g1332), .B(g5892), .Z(g6249) ) ;
AND2    gate5149  (.A(g1692), .B(g6036), .Z(g6250) ) ;
AND2    gate5150  (.A(g508), .B(g5896), .Z(g6253) ) ;
AND2    gate5151  (.A(g532), .B(g5897), .Z(g6254) ) ;
AND2    gate5152  (.A(g1335), .B(g5895), .Z(g6255) ) ;
AND2    gate5153  (.A(g1696), .B(g6040), .Z(g6256) ) ;
AND2    gate5154  (.A(g512), .B(g5899), .Z(g6258) ) ;
AND2    gate5155  (.A(g1699), .B(g6044), .Z(g6259) ) ;
AND2    gate5156  (.A(g1703), .B(g6048), .Z(g6260) ) ;
AND2    gate5157  (.A(g516), .B(g5901), .Z(g6262) ) ;
AND2    gate5158  (.A(g1711), .B(g6052), .Z(g6263) ) ;
AND2    gate5159  (.A(g520), .B(g5903), .Z(g6265) ) ;
AND2    gate5160  (.A(g1721), .B(g6057), .Z(g6266) ) ;
AND2    gate5161  (.A(g524), .B(g5908), .Z(g6269) ) ;
AND2    gate5162  (.A(g1726), .B(g6062), .Z(g6270) ) ;
AND2    gate5163  (.A(g1735), .B(g6070), .Z(g6275) ) ;
AND2    gate5164  (.A(g5615), .B(g6160), .Z(g6288) ) ;
AND2    gate5165  (.A(g5740), .B(g6164), .Z(g6302) ) ;
OR2     gate5166  (.A(g3609), .B(g3613), .Z(g3837) ) ;
AND2    gate5167  (.A(g3837), .B(g6194), .Z(g6311) ) ;
OR2     gate5168  (.A(g3614), .B(g3617), .Z(g3841) ) ;
AND2    gate5169  (.A(g3841), .B(g6194), .Z(g6313) ) ;
OR2     gate5170  (.A(g3618), .B(g3625), .Z(g3849) ) ;
AND2    gate5171  (.A(g3849), .B(g6194), .Z(g6315) ) ;
OR2     gate5172  (.A(g3626), .B(g3631), .Z(g3855) ) ;
AND2    gate5173  (.A(g3855), .B(g6194), .Z(g6316) ) ;
OR2     gate5174  (.A(g3632), .B(g3641), .Z(g3862) ) ;
AND2    gate5175  (.A(g3862), .B(g6194), .Z(g6317) ) ;
OR2     gate5176  (.A(g3637), .B(g3648), .Z(g3865) ) ;
AND2    gate5177  (.A(g3865), .B(g6212), .Z(g6318) ) ;
OR2     gate5178  (.A(g3642), .B(g3650), .Z(g3869) ) ;
AND2    gate5179  (.A(g3869), .B(g6194), .Z(g6320) ) ;
OR2     gate5180  (.A(g3649), .B(g3657), .Z(g3873) ) ;
AND2    gate5181  (.A(g3873), .B(g6212), .Z(g6321) ) ;
OR2     gate5182  (.A(g3651), .B(g3659), .Z(g3877) ) ;
AND2    gate5183  (.A(g3877), .B(g6194), .Z(g6323) ) ;
OR2     gate5184  (.A(g3658), .B(g3665), .Z(g3880) ) ;
AND2    gate5185  (.A(g3880), .B(g6212), .Z(g6324) ) ;
OR2     gate5186  (.A(g3602), .B(g3608), .Z(g3833) ) ;
AND2    gate5187  (.A(g3833), .B(g6194), .Z(g6326) ) ;
OR2     gate5188  (.A(g3666), .B(g3671), .Z(g3884) ) ;
AND2    gate5189  (.A(g3884), .B(g6212), .Z(g6327) ) ;
OR2     gate5190  (.A(g3672), .B(g3682), .Z(g3888) ) ;
AND2    gate5191  (.A(g3888), .B(g6212), .Z(g6329) ) ;
OR2     gate5192  (.A(g3683), .B(g3688), .Z(g3891) ) ;
AND2    gate5193  (.A(g3891), .B(g6212), .Z(g6331) ) ;
OR2     gate5194  (.A(g3689), .B(g3697), .Z(g3896) ) ;
AND2    gate5195  (.A(g3896), .B(g6212), .Z(g6333) ) ;
OR2     gate5196  (.A(g3629), .B(g3636), .Z(g3858) ) ;
AND2    gate5197  (.A(g3858), .B(g6212), .Z(g6334) ) ;
OR2     gate5198  (.A(g5665), .B(g5937), .Z(g6246) ) ;
AND2    gate5199  (.A(g6246), .B(g6065), .Z(g6336) ) ;
OR2     gate5200  (.A(g5668), .B(g5939), .Z(g6251) ) ;
AND2    gate5201  (.A(g6251), .B(g6067), .Z(g6338) ) ;
OR2     gate5202  (.A(g5671), .B(g5941), .Z(g6257) ) ;
AND2    gate5203  (.A(g6257), .B(g6069), .Z(g6340) ) ;
OR2     gate5204  (.A(g5673), .B(g5944), .Z(g6261) ) ;
AND2    gate5205  (.A(g6261), .B(g6074), .Z(g6341) ) ;
OR2     gate5206  (.A(g5675), .B(g5948), .Z(g6264) ) ;
AND2    gate5207  (.A(g6264), .B(g6076), .Z(g6342) ) ;
OR2     gate5208  (.A(g5677), .B(g5951), .Z(g6268) ) ;
AND2    gate5209  (.A(g6268), .B(g6078), .Z(g6343) ) ;
OR2     gate5210  (.A(g5679), .B(g5953), .Z(g6272) ) ;
AND2    gate5211  (.A(g6272), .B(g6080), .Z(g6344) ) ;
OR2     gate5212  (.A(g5681), .B(g5955), .Z(g6273) ) ;
AND2    gate5213  (.A(g6273), .B(g6083), .Z(g6345) ) ;
OR2     gate5214  (.A(g5682), .B(g5956), .Z(g6274) ) ;
AND2    gate5215  (.A(g6274), .B(g6087), .Z(g6346) ) ;
AND2    gate5216  (.A(g5869), .B(g6211), .Z(g6348) ) ;
AND2    gate5217  (.A(g5866), .B(g6193), .Z(g6354) ) ;
NAND2   gate5218  (.A(II8195), .B(II8196), .Z(g6394) ) ;
AND3    gate5219  (.A(g2032), .B(g6394), .C(g1609), .Z(g6468) ) ;
NAND2   gate5220  (.A(II8202), .B(II8203), .Z(g6397) ) ;
AND3    gate5221  (.A(g2036), .B(g6397), .C(g1628), .Z(g6473) ) ;
AND2    gate5222  (.A(g1838), .B(g6469), .Z(g6555) ) ;
AND2    gate5223  (.A(g1595), .B(g6469), .Z(g6557) ) ;
AND2    gate5224  (.A(g1842), .B(g6474), .Z(g6558) ) ;
AND2    gate5225  (.A(g1612), .B(g6474), .Z(g6559) ) ;
AND2    gate5226  (.A(g6581), .B(g6236), .Z(g6603) ) ;
OR2     gate5227  (.A(g6337), .B(g6466), .Z(g6554) ) ;
AND2    gate5228  (.A(g932), .B(g6554), .Z(g6613) ) ;
OR2     gate5229  (.A(g6339), .B(g6467), .Z(g6556) ) ;
AND2    gate5230  (.A(g932), .B(g6556), .Z(g6614) ) ;
AND2    gate5231  (.A(g6516), .B(g6117), .Z(g6620) ) ;
AND3    gate5232  (.A(g2121), .B(g1595), .C(g6538), .Z(g6625) ) ;
AND3    gate5233  (.A(g2138), .B(g1612), .C(g6540), .Z(g6628) ) ;
OR2     gate5234  (.A(g6468), .B(g4244), .Z(g6545) ) ;
AND2    gate5235  (.A(g1838), .B(g6545), .Z(g6631) ) ;
AND2    gate5236  (.A(g1595), .B(g6545), .Z(g6634) ) ;
OR2     gate5237  (.A(g6473), .B(g4247), .Z(g6549) ) ;
AND2    gate5238  (.A(g1842), .B(g6549), .Z(g6637) ) ;
AND2    gate5239  (.A(g1612), .B(g6549), .Z(g6640) ) ;
AND2    gate5240  (.A(g6574), .B(g6229), .Z(g6643) ) ;
AND2    gate5241  (.A(g6575), .B(g6230), .Z(g6644) ) ;
AND2    gate5242  (.A(g6576), .B(g6231), .Z(g6645) ) ;
AND2    gate5243  (.A(g6577), .B(g6232), .Z(g6646) ) ;
AND2    gate5244  (.A(g6578), .B(g6233), .Z(g6647) ) ;
AND2    gate5245  (.A(g6579), .B(g6234), .Z(g6648) ) ;
AND2    gate5246  (.A(g6580), .B(g6235), .Z(g6650) ) ;
AND2    gate5247  (.A(g6616), .B(g6615), .Z(g6692) ) ;
AND2    gate5248  (.A(g6618), .B(g6617), .Z(g6693) ) ;
OR3     gate5249  (.A(g6478), .B(g6624), .C(g6623), .Z(g6682) ) ;
AND2    gate5250  (.A(g6682), .B(g932), .Z(g6716) ) ;
AND2    gate5251  (.A(g4511), .B(g6661), .Z(g6718) ) ;
AND2    gate5252  (.A(g4518), .B(g6665), .Z(g6719) ) ;
NAND3   gate5253  (.A(g6669), .B(g5065), .C(g5062), .Z(g6717) ) ;
OR2     gate5254  (.A(g4373), .B(g3668), .Z(g4427) ) ;
AND2    gate5255  (.A(g6717), .B(g4427), .Z(g6731) ) ;
AND3    gate5256  (.A(g6712), .B(g754), .C(g5237), .Z(g6736) ) ;
AND3    gate5257  (.A(g6714), .B(g760), .C(g5237), .Z(g6737) ) ;
AND3    gate5258  (.A(g6713), .B(g809), .C(g5242), .Z(g6738) ) ;
AND3    gate5259  (.A(g6715), .B(g815), .C(g5242), .Z(g6739) ) ;
AND2    gate5260  (.A(g6733), .B(g6732), .Z(g6748) ) ;
AND2    gate5261  (.A(g6735), .B(g6734), .Z(g6749) ) ;
OR3     gate5262  (.A(g6670), .B(g6625), .C(g6736), .Z(g6750) ) ;
AND2    gate5263  (.A(g6750), .B(g2986), .Z(g6766) ) ;
OR3     gate5264  (.A(g6676), .B(g6625), .C(g6737), .Z(g6754) ) ;
AND2    gate5265  (.A(g6754), .B(g2986), .Z(g6767) ) ;
AND2    gate5266  (.A(g6750), .B(g3477), .Z(g6768) ) ;
OR3     gate5267  (.A(g6673), .B(g6628), .C(g6738), .Z(g6758) ) ;
AND2    gate5268  (.A(g6758), .B(g2986), .Z(g6769) ) ;
AND2    gate5269  (.A(g6754), .B(g3482), .Z(g6770) ) ;
AND2    gate5270  (.A(g6758), .B(g3483), .Z(g6771) ) ;
AND2    gate5271  (.A(g6746), .B(g3312), .Z(g6772) ) ;
OR3     gate5272  (.A(g6679), .B(g6628), .C(g6739), .Z(g6762) ) ;
AND2    gate5273  (.A(g6762), .B(g2986), .Z(g6773) ) ;
AND2    gate5274  (.A(g6762), .B(g3488), .Z(g6777) ) ;
OR2     gate5275  (.A(g4830), .B(g4833), .Z(g4946) ) ;
OR2     gate5276  (.A(g6718), .B(g6748), .Z(g6781) ) ;
AND2    gate5277  (.A(g4946), .B(g6781), .Z(g6798) ) ;
OR2     gate5278  (.A(g4834), .B(g4836), .Z(g4948) ) ;
OR2     gate5279  (.A(g6719), .B(g6749), .Z(g6782) ) ;
AND2    gate5280  (.A(g4948), .B(g6782), .Z(g6799) ) ;
AND2    gate5281  (.A(g6784), .B(g3346), .Z(g6816) ) ;
AND2    gate5282  (.A(g6803), .B(g5958), .Z(g6828) ) ;
AND2    gate5283  (.A(g6806), .B(g5958), .Z(g6829) ) ;
AND2    gate5284  (.A(g6809), .B(g5975), .Z(g6830) ) ;
AND2    gate5285  (.A(g6812), .B(g5975), .Z(g6831) ) ;
NAND3   gate5286  (.A(g901), .B(g3433), .C(g2340), .Z(g3741) ) ;
NAND2   gate5287  (.A(II9051), .B(II9052), .Z(g6843) ) ;
AND3    gate5288  (.A(g3741), .B(g328), .C(g6843), .Z(g6848) ) ;
OR2     gate5289  (.A(g5860), .B(g6834), .Z(g6846) ) ;
AND2    gate5290  (.A(g6846), .B(g2293), .Z(g6851) ) ;
OR2     gate5291  (.A(g5861), .B(g6837), .Z(g6847) ) ;
AND2    gate5292  (.A(g6847), .B(g2295), .Z(g6852) ) ;
NAND2   gate5293  (.A(g6848), .B(g3621), .Z(g6873) ) ;
AND2    gate5294  (.A(g6873), .B(g2060), .Z(g6874) ) ;
OR2     gate5295  (.A(g6874), .B(g3358), .Z(g6907) ) ;
AND2    gate5296  (.A(g6907), .B(g3886), .Z(g6908) ) ;
AND2    gate5297  (.A(g6896), .B(g6894), .Z(g6909) ) ;
AND2    gate5298  (.A(g6892), .B(g6891), .Z(g6910) ) ;
AND2    gate5299  (.A(g6904), .B(g6902), .Z(g6911) ) ;
AND2    gate5300  (.A(g6899), .B(g6897), .Z(g6912) ) ;
AND2    gate5301  (.A(g6900), .B(g6898), .Z(g6913) ) ;
AND2    gate5302  (.A(g6895), .B(g6893), .Z(g6914) ) ;
AND2    gate5303  (.A(g6906), .B(g6905), .Z(g6915) ) ;
AND2    gate5304  (.A(g6903), .B(g6901), .Z(g6916) ) ;
OR2     gate5305  (.A(g6911), .B(g6913), .Z(g6918) ) ;
OR2     gate5306  (.A(g6909), .B(g6910), .Z(g6917) ) ;
AND2    gate5307  (.A(g6918), .B(g6917), .Z(g6923) ) ;
OR2     gate5308  (.A(g6915), .B(g6916), .Z(g6920) ) ;
OR2     gate5309  (.A(g6912), .B(g6914), .Z(g6919) ) ;
AND2    gate5310  (.A(g6920), .B(g6919), .Z(g6924) ) ;
AND2    gate5311  (.A(g6932), .B(g3605), .Z(g6934) ) ;
AND2    gate5312  (.A(g6933), .B(g3622), .Z(g6935) ) ;
OR2     gate5313  (.A(g1059), .B(g1045), .Z(g1589) ) ;
NAND3   gate5314  (.A(g1584), .B(g749), .C(g736), .Z(g2095) ) ;
NAND3   gate5315  (.A(g729), .B(g719), .C(g766), .Z(g1573) ) ;
NAND3   gate5316  (.A(g1588), .B(g804), .C(g791), .Z(g2100) ) ;
NAND3   gate5317  (.A(g784), .B(g774), .C(g821), .Z(g1582) ) ;
OR2     gate5318  (.A(g3122), .B(g3132), .Z(g3503) ) ;
OR2     gate5319  (.A(g2808), .B(g2821), .Z(g3598) ) ;
NAND2   gate5320  (.A(g2142), .B(g1797), .Z(g2951) ) ;
NAND2   gate5321  (.A(g2340), .B(g1402), .Z(g3215) ) ;
OR2     gate5322  (.A(g1555), .B(g3559), .Z(g3992) ) ;
NOR2    gate5323  (.A(g1250), .B(g3425), .Z(g4000) ) ;
OR2     gate5324  (.A(g3912), .B(g471), .Z(g4233) ) ;
OR2     gate5325  (.A(g3921), .B(g478), .Z(g4234) ) ;
OR2     gate5326  (.A(g4053), .B(g4058), .Z(g4243) ) ;
NAND2   gate5327  (.A(II4183), .B(II4184), .Z(g2995) ) ;
NAND2   gate5328  (.A(II4211), .B(II4212), .Z(g3013) ) ;
NOR2    gate5329  (.A(g923), .B(g4253), .Z(g4432) ) ;
OR2     gate5330  (.A(g4827), .B(g4828), .Z(g4936) ) ;
OR2     gate5331  (.A(g4829), .B(g4832), .Z(g4941) ) ;
NAND2   gate5332  (.A(II6500), .B(II6501), .Z(g4819) ) ;
OR2     gate5333  (.A(g3491), .B(g4819), .Z(g5060) ) ;
OR2     gate5334  (.A(g4661), .B(g4666), .Z(g5062) ) ;
OR2     gate5335  (.A(g4667), .B(g4671), .Z(g5065) ) ;
OR2     gate5336  (.A(g4668), .B(g4672), .Z(g5066) ) ;
OR2     gate5337  (.A(g4673), .B(g4677), .Z(g5068) ) ;
OR3     gate5338  (.A(g4904), .B(g4914), .C(g4894), .Z(g5202) ) ;
NOR3    gate5339  (.A(g4819), .B(g3491), .C(g3559), .Z(g5048) ) ;
NAND2   gate5340  (.A(II3178), .B(II3179), .Z(g2067) ) ;
NAND2   gate5341  (.A(II3189), .B(II3190), .Z(g2080) ) ;
NAND2   gate5342  (.A(II4204), .B(II4205), .Z(g3012) ) ;
NAND2   gate5343  (.A(II4234), .B(II4235), .Z(g3028) ) ;
OR2     gate5344  (.A(g5199), .B(g4928), .Z(g5367) ) ;
OR2     gate5345  (.A(g5201), .B(g4932), .Z(g5368) ) ;
OR2     gate5346  (.A(g5211), .B(g4937), .Z(g5370) ) ;
OR2     gate5347  (.A(g5213), .B(g4942), .Z(g5372) ) ;
OR2     gate5348  (.A(g5215), .B(g4947), .Z(g5374) ) ;
OR2     gate5349  (.A(g5217), .B(g4949), .Z(g5377) ) ;
NOR2    gate5350  (.A(g5019), .B(g3559), .Z(g5227) ) ;
OR2     gate5351  (.A(g5551), .B(g5398), .Z(g5659) ) ;
OR2     gate5352  (.A(g5553), .B(g5402), .Z(g5662) ) ;
OR2     gate5353  (.A(g5555), .B(g5406), .Z(g5666) ) ;
OR2     gate5354  (.A(g5556), .B(g5410), .Z(g5669) ) ;
OR2     gate5355  (.A(g5557), .B(g5414), .Z(g5672) ) ;
OR2     gate5356  (.A(g5558), .B(g5419), .Z(g5674) ) ;
OR2     gate5357  (.A(g5559), .B(g5424), .Z(g5676) ) ;
OR2     gate5358  (.A(g5560), .B(g5428), .Z(g5678) ) ;
OR2     gate5359  (.A(g5562), .B(g5429), .Z(g5680) ) ;
NOR2    gate5360  (.A(g197), .B(g5862), .Z(g6073) ) ;
NOR2    gate5361  (.A(g269), .B(g5863), .Z(g6075) ) ;
OR4     gate5362  (.A(g6194), .B(g5958), .C(g5975), .D(g5997), .Z(II7969) ) ;
OR4     gate5363  (.A(g6015), .B(g6212), .C(g4950), .D(g4877), .Z(II7970) ) ;
OR4     gate5364  (.A(g5202), .B(g4993), .C(g4967), .D(g4980), .Z(II7971) ) ;
OR2     gate5365  (.A(g4915), .B(g5025), .Z(II7972) ) ;
OR4     gate5366  (.A(g6194), .B(g5958), .C(g5975), .D(g5997), .Z(II7978) ) ;
OR4     gate5367  (.A(g6015), .B(g6212), .C(g4950), .D(g4877), .Z(II7979) ) ;
OR4     gate5368  (.A(g5202), .B(g4993), .C(g4967), .D(g4980), .Z(II7980) ) ;
OR2     gate5369  (.A(g4915), .B(g5025), .Z(II7981) ) ;
OR4     gate5370  (.A(g6194), .B(g5958), .C(g5975), .D(g5997), .Z(II7987) ) ;
OR4     gate5371  (.A(g6015), .B(g6212), .C(g4950), .D(g4877), .Z(II7988) ) ;
OR4     gate5372  (.A(g5202), .B(g4993), .C(g4967), .D(g4980), .Z(II7989) ) ;
OR2     gate5373  (.A(g4915), .B(g5025), .Z(II7990) ) ;
OR4     gate5374  (.A(g6194), .B(g5958), .C(g5975), .D(g5997), .Z(II8079) ) ;
OR4     gate5375  (.A(g6015), .B(g6212), .C(g4950), .D(g4877), .Z(II8080) ) ;
OR4     gate5376  (.A(g4894), .B(g4904), .C(g4993), .D(g4967), .Z(II8081) ) ;
OR4     gate5377  (.A(g4980), .B(g4915), .C(g5025), .D(g5054), .Z(II8082) ) ;
OR4     gate5378  (.A(g6194), .B(g5958), .C(g5975), .D(g5997), .Z(II8117) ) ;
OR4     gate5379  (.A(g6015), .B(g6212), .C(g4950), .D(g4877), .Z(II8118) ) ;
OR4     gate5380  (.A(g5202), .B(g4993), .C(g4967), .D(g4980), .Z(II8119) ) ;
OR2     gate5381  (.A(g4915), .B(g5025), .Z(II8120) ) ;
OR4     gate5382  (.A(g6194), .B(g5958), .C(g5975), .D(g5997), .Z(II8126) ) ;
OR4     gate5383  (.A(g6015), .B(g6212), .C(g4950), .D(g4877), .Z(II8127) ) ;
OR4     gate5384  (.A(g5202), .B(g4993), .C(g4967), .D(g4980), .Z(II8128) ) ;
OR2     gate5385  (.A(g4915), .B(g5025), .Z(II8129) ) ;
OR4     gate5386  (.A(g6194), .B(g5958), .C(g5975), .D(g5997), .Z(II8135) ) ;
OR4     gate5387  (.A(g6015), .B(g6212), .C(g4950), .D(g4877), .Z(II8136) ) ;
OR4     gate5388  (.A(g4894), .B(g4904), .C(g4993), .D(g4967), .Z(II8137) ) ;
OR4     gate5389  (.A(g4980), .B(g4915), .C(g5025), .D(g5054), .Z(II8138) ) ;
OR4     gate5390  (.A(g6194), .B(g5958), .C(g5975), .D(g5997), .Z(II8208) ) ;
OR4     gate5391  (.A(g6015), .B(g6212), .C(g4950), .D(g4877), .Z(II8209) ) ;
OR4     gate5392  (.A(g5202), .B(g4993), .C(g4967), .D(g4980), .Z(II8210) ) ;
OR2     gate5393  (.A(g4915), .B(g5025), .Z(II8211) ) ;
OR4     gate5394  (.A(g6326), .B(g6135), .C(g6140), .D(g6157), .Z(II8345) ) ;
OR4     gate5395  (.A(g6159), .B(g6334), .C(g5163), .D(g5191), .Z(II8346) ) ;
OR4     gate5396  (.A(g5188), .B(g5157), .C(g5154), .D(g5193), .Z(II8347) ) ;
OR4     gate5397  (.A(g5229), .B(g5234), .C(g5218), .D(g5225), .Z(II8348) ) ;
OR4     gate5398  (.A(II8345), .B(II8346), .C(II8347), .D(II8348), .Z(II8349) ) ;
NOR4    gate5399  (.A(II8079), .B(II8080), .C(II8081), .D(II8082), .Z(g6335) ) ;
OR4     gate5400  (.A(g6311), .B(g6123), .C(g6125), .D(g6141), .Z(II8356) ) ;
OR4     gate5401  (.A(g6145), .B(g6318), .C(g5171), .D(g5187), .Z(II8357) ) ;
OR4     gate5402  (.A(g5192), .B(g5153), .C(g5158), .D(g5197), .Z(II8358) ) ;
OR4     gate5403  (.A(g5232), .B(g5236), .C(g5216), .D(g5226), .Z(II8359) ) ;
OR4     gate5404  (.A(II8356), .B(II8357), .C(II8358), .D(II8359), .Z(II8360) ) ;
NOR4    gate5405  (.A(II8135), .B(II8136), .C(II8137), .D(II8138), .Z(g6359) ) ;
OR4     gate5406  (.A(g6313), .B(g6124), .C(g6127), .D(g6144), .Z(II8367) ) ;
OR4     gate5407  (.A(g6148), .B(g6321), .C(g5176), .D(g5184), .Z(II8368) ) ;
OR4     gate5408  (.A(g5165), .B(g5159), .C(g5233), .D(g5240), .Z(II8369) ) ;
NOR4    gate5409  (.A(II8126), .B(II8127), .C(II8128), .D(II8129), .Z(g6358) ) ;
OR2     gate5410  (.A(g5214), .B(g6358), .Z(II8370) ) ;
OR4     gate5411  (.A(g6315), .B(g6126), .C(g6129), .D(g6146), .Z(II8376) ) ;
OR4     gate5412  (.A(g6150), .B(g6324), .C(g5180), .D(g5181), .Z(II8377) ) ;
OR4     gate5413  (.A(g5173), .B(g5166), .C(g5235), .D(g5245), .Z(II8378) ) ;
NOR4    gate5414  (.A(II8117), .B(II8118), .C(II8119), .D(II8120), .Z(g6357) ) ;
OR2     gate5415  (.A(g5212), .B(g6357), .Z(II8379) ) ;
OR4     gate5416  (.A(g6316), .B(g6128), .C(g6131), .D(g6149), .Z(II8385) ) ;
OR4     gate5417  (.A(g6152), .B(g6327), .C(g5183), .D(g5177), .Z(II8386) ) ;
NOR4    gate5418  (.A(II7987), .B(II7988), .C(II7989), .D(II7990), .Z(g6281) ) ;
OR3     gate5419  (.A(g5178), .B(g5209), .C(g6281), .Z(II8387) ) ;
OR4     gate5420  (.A(g6317), .B(g6130), .C(g6133), .D(g6151), .Z(II8393) ) ;
OR4     gate5421  (.A(g6154), .B(g6329), .C(g5186), .D(g5172), .Z(II8394) ) ;
NOR4    gate5422  (.A(II7978), .B(II7979), .C(II7980), .D(II7981), .Z(g6280) ) ;
OR3     gate5423  (.A(g5182), .B(g5200), .C(g6280), .Z(II8395) ) ;
OR2     gate5424  (.A(g6634), .B(g6631), .Z(g6659) ) ;
OR2     gate5425  (.A(g6640), .B(g6637), .Z(g6660) ) ;
OR4     gate5426  (.A(g6610), .B(g6608), .C(g6606), .D(g6604), .Z(II8773) ) ;
OR4     gate5427  (.A(g6655), .B(g6653), .C(g6651), .D(g6649), .Z(II8774) ) ;
OR4     gate5428  (.A(g6612), .B(g6611), .C(g6609), .D(g6607), .Z(II8778) ) ;
OR4     gate5429  (.A(g6605), .B(g6656), .C(g6654), .D(g6652), .Z(II8779) ) ;
OR2     gate5430  (.A(g6613), .B(g4679), .Z(g6669) ) ;
OR3     gate5431  (.A(g6465), .B(g6622), .C(g6621), .Z(g6683) ) ;
OR2     gate5432  (.A(g6692), .B(g4831), .Z(g6703) ) ;
OR2     gate5433  (.A(g6693), .B(g4835), .Z(g6705) ) ;
OR2     gate5434  (.A(g6614), .B(g6731), .Z(g6747) ) ;
OR4     gate5435  (.A(g6320), .B(g6828), .C(g6830), .D(g6153), .Z(II9057) ) ;
OR4     gate5436  (.A(g6156), .B(g6331), .C(g5190), .D(g5164), .Z(II9058) ) ;
NOR4    gate5437  (.A(II7969), .B(II7970), .C(II7971), .D(II7972), .Z(g6279) ) ;
OR3     gate5438  (.A(g5185), .B(g5198), .C(g6279), .Z(II9059) ) ;
OR4     gate5439  (.A(g6323), .B(g6829), .C(g6831), .D(g6155), .Z(II9064) ) ;
OR4     gate5440  (.A(g6158), .B(g6333), .C(g5152), .D(g5156), .Z(II9065) ) ;
NOR4    gate5441  (.A(II8208), .B(II8209), .C(II8210), .D(II8211), .Z(g6400) ) ;
OR3     gate5442  (.A(g5189), .B(g5269), .C(g6400), .Z(II9066) ) ;
OR2     gate5443  (.A(g6798), .B(g6923), .Z(g6926) ) ;
OR2     gate5444  (.A(g6799), .B(g6924), .Z(g6927) ) ;
NAND3   gate5445  (.A(g6703), .B(g6457), .C(g4936), .Z(g6740) ) ;
NAND2   gate5446  (.A(g4532), .B(g6926), .Z(g6928) ) ;
NAND3   gate5447  (.A(g6705), .B(g6461), .C(g4941), .Z(g6741) ) ;
NAND2   gate5448  (.A(g4536), .B(g6927), .Z(g6929) ) ;
NAND2   gate5449  (.A(g524), .B(g248), .Z(II1951) ) ;
NAND2   gate5450  (.A(g524), .B(II1951), .Z(II1952) ) ;
NAND2   gate5451  (.A(g248), .B(II1951), .Z(II1953) ) ;
NAND2   gate5452  (.A(II1952), .B(II1953), .Z(g926) ) ;
NAND2   gate5453  (.A(g520), .B(g242), .Z(II1961) ) ;
NAND2   gate5454  (.A(g520), .B(II1961), .Z(II1962) ) ;
NAND2   gate5455  (.A(g242), .B(II1961), .Z(II1963) ) ;
NAND2   gate5456  (.A(II1962), .B(II1963), .Z(g928) ) ;
NAND2   gate5457  (.A(g516), .B(g236), .Z(II1969) ) ;
NAND2   gate5458  (.A(g516), .B(II1969), .Z(II1970) ) ;
NAND2   gate5459  (.A(g236), .B(II1969), .Z(II1971) ) ;
NAND2   gate5460  (.A(II1970), .B(II1971), .Z(g930) ) ;
NAND2   gate5461  (.A(g512), .B(g230), .Z(II1978) ) ;
NAND2   gate5462  (.A(g512), .B(II1978), .Z(II1979) ) ;
NAND2   gate5463  (.A(g230), .B(II1978), .Z(II1980) ) ;
NAND2   gate5464  (.A(II1979), .B(II1980), .Z(g937) ) ;
NAND2   gate5465  (.A(g508), .B(g224), .Z(II1986) ) ;
NAND2   gate5466  (.A(g508), .B(II1986), .Z(II1987) ) ;
NAND2   gate5467  (.A(g224), .B(II1986), .Z(II1988) ) ;
NAND2   gate5468  (.A(II1987), .B(II1988), .Z(g939) ) ;
NAND2   gate5469  (.A(g504), .B(g218), .Z(II1994) ) ;
NAND2   gate5470  (.A(g504), .B(II1994), .Z(II1995) ) ;
NAND2   gate5471  (.A(g218), .B(II1994), .Z(II1996) ) ;
NAND2   gate5472  (.A(II1995), .B(II1996), .Z(g941) ) ;
NAND2   gate5473  (.A(g500), .B(g212), .Z(II2003) ) ;
NAND2   gate5474  (.A(g500), .B(II2003), .Z(II2004) ) ;
NAND2   gate5475  (.A(g212), .B(II2003), .Z(II2005) ) ;
NAND2   gate5476  (.A(II2004), .B(II2005), .Z(g944) ) ;
NAND2   gate5477  (.A(g532), .B(g260), .Z(II2013) ) ;
NAND2   gate5478  (.A(g532), .B(II2013), .Z(II2014) ) ;
NAND2   gate5479  (.A(g260), .B(II2013), .Z(II2015) ) ;
NAND2   gate5480  (.A(II2014), .B(II2015), .Z(g948) ) ;
NAND2   gate5481  (.A(g528), .B(g254), .Z(II2021) ) ;
NAND2   gate5482  (.A(g528), .B(II2021), .Z(II2022) ) ;
NAND2   gate5483  (.A(g254), .B(II2021), .Z(II2023) ) ;
NAND2   gate5484  (.A(II2022), .B(II2023), .Z(g950) ) ;
NAND2   gate5485  (.A(g7), .B(g3), .Z(II2060) ) ;
NAND2   gate5486  (.A(g7), .B(II2060), .Z(II2061) ) ;
NAND2   gate5487  (.A(g3), .B(II2060), .Z(II2062) ) ;
NAND2   gate5488  (.A(II2061), .B(II2062), .Z(g1036) ) ;
NAND2   gate5489  (.A(g15), .B(g11), .Z(II2072) ) ;
NAND2   gate5490  (.A(g15), .B(II2072), .Z(II2073) ) ;
NAND2   gate5491  (.A(g11), .B(II2072), .Z(II2074) ) ;
NAND2   gate5492  (.A(II2073), .B(II2074), .Z(g1042) ) ;
NAND2   gate5493  (.A(g25), .B(g19), .Z(II2080) ) ;
NAND2   gate5494  (.A(g25), .B(II2080), .Z(II2081) ) ;
NAND2   gate5495  (.A(g19), .B(II2080), .Z(II2082) ) ;
NAND2   gate5496  (.A(II2081), .B(II2082), .Z(g1044) ) ;
NAND2   gate5497  (.A(g33), .B(g29), .Z(II2089) ) ;
NAND2   gate5498  (.A(g33), .B(II2089), .Z(II2090) ) ;
NAND2   gate5499  (.A(g29), .B(II2089), .Z(II2091) ) ;
NAND2   gate5500  (.A(II2090), .B(II2091), .Z(g1047) ) ;
NAND2   gate5501  (.A(g602), .B(g610), .Z(II2108) ) ;
NAND2   gate5502  (.A(g602), .B(II2108), .Z(II2109) ) ;
NAND2   gate5503  (.A(g610), .B(II2108), .Z(II2110) ) ;
NAND2   gate5504  (.A(g567), .B(g598), .Z(II2244) ) ;
NAND2   gate5505  (.A(g567), .B(II2244), .Z(II2245) ) ;
NAND2   gate5506  (.A(g598), .B(II2244), .Z(II2246) ) ;
NAND2   gate5507  (.A(g830), .B(g341), .Z(II2299) ) ;
NAND2   gate5508  (.A(g830), .B(II2299), .Z(II2300) ) ;
NAND2   gate5509  (.A(g341), .B(II2299), .Z(II2301) ) ;
NAND2   gate5510  (.A(g1042), .B(g1036), .Z(II2497) ) ;
NAND2   gate5511  (.A(g1042), .B(II2497), .Z(II2498) ) ;
NAND2   gate5512  (.A(g1036), .B(II2497), .Z(II2499) ) ;
NAND2   gate5513  (.A(II2498), .B(II2499), .Z(g1534) ) ;
NAND2   gate5514  (.A(g1047), .B(g1044), .Z(II2506) ) ;
NAND2   gate5515  (.A(g1047), .B(II2506), .Z(II2507) ) ;
NAND2   gate5516  (.A(g1044), .B(II2506), .Z(II2508) ) ;
NAND2   gate5517  (.A(II2507), .B(II2508), .Z(g1540) ) ;
NAND2   gate5518  (.A(g766), .B(g719), .Z(II2526) ) ;
NAND2   gate5519  (.A(g766), .B(II2526), .Z(II2527) ) ;
NAND2   gate5520  (.A(g719), .B(II2526), .Z(II2528) ) ;
NAND2   gate5521  (.A(g821), .B(g774), .Z(II2542) ) ;
NAND2   gate5522  (.A(g821), .B(II2542), .Z(II2543) ) ;
NAND2   gate5523  (.A(g774), .B(II2542), .Z(II2544) ) ;
NAND2   gate5524  (.A(g710), .B(g131), .Z(II2674) ) ;
NAND2   gate5525  (.A(g710), .B(II2674), .Z(II2675) ) ;
NAND2   gate5526  (.A(g131), .B(II2674), .Z(II2676) ) ;
NAND2   gate5527  (.A(g918), .B(g613), .Z(II2681) ) ;
NAND2   gate5528  (.A(g918), .B(II2681), .Z(II2682) ) ;
NAND2   gate5529  (.A(g613), .B(II2681), .Z(II2683) ) ;
NAND2   gate5530  (.A(g749), .B(g743), .Z(II2766) ) ;
NAND2   gate5531  (.A(g749), .B(II2766), .Z(II2767) ) ;
NAND2   gate5532  (.A(g743), .B(II2766), .Z(II2768) ) ;
NAND2   gate5533  (.A(g804), .B(g798), .Z(II2795) ) ;
NAND2   gate5534  (.A(g804), .B(II2795), .Z(II2796) ) ;
NAND2   gate5535  (.A(g798), .B(II2795), .Z(II2797) ) ;
NAND2   gate5536  (.A(g1027), .B(g634), .Z(II2897) ) ;
NAND2   gate5537  (.A(g1027), .B(II2897), .Z(II2898) ) ;
NAND2   gate5538  (.A(g634), .B(II2897), .Z(II2899) ) ;
NAND2   gate5539  (.A(g1436), .B(g345), .Z(II2933) ) ;
NAND2   gate5540  (.A(g1436), .B(II2933), .Z(II2934) ) ;
NAND2   gate5541  (.A(g345), .B(II2933), .Z(II2935) ) ;
NOR3    gate5542  (.A(g944), .B(g941), .C(g939), .Z(g1473) ) ;
NOR3    gate5543  (.A(g937), .B(g930), .C(g928), .Z(g1470) ) ;
NOR3    gate5544  (.A(g926), .B(g950), .C(g948), .Z(g1459) ) ;
NAND2   gate5545  (.A(g1279), .B(g1276), .Z(II3125) ) ;
NAND2   gate5546  (.A(g1279), .B(II3125), .Z(II3126) ) ;
NAND2   gate5547  (.A(g1276), .B(II3125), .Z(II3127) ) ;
NAND2   gate5548  (.A(g1540), .B(g1534), .Z(II3168) ) ;
NAND2   gate5549  (.A(g1540), .B(II3168), .Z(II3169) ) ;
NAND2   gate5550  (.A(g1534), .B(II3168), .Z(II3170) ) ;
NAND2   gate5551  (.A(g1706), .B(g736), .Z(II3177) ) ;
NAND2   gate5552  (.A(g1706), .B(II3177), .Z(II3178) ) ;
NAND2   gate5553  (.A(g736), .B(II3177), .Z(II3179) ) ;
NAND2   gate5554  (.A(g1716), .B(g791), .Z(II3188) ) ;
NAND2   gate5555  (.A(g1716), .B(II3188), .Z(II3189) ) ;
NAND2   gate5556  (.A(g791), .B(II3188), .Z(II3190) ) ;
NAND2   gate5557  (.A(g1826), .B(g135), .Z(II3398) ) ;
NAND2   gate5558  (.A(g1826), .B(II3398), .Z(II3399) ) ;
NAND2   gate5559  (.A(g135), .B(II3398), .Z(II3400) ) ;
NAND2   gate5560  (.A(g1419), .B(g616), .Z(II3411) ) ;
NAND2   gate5561  (.A(g1419), .B(II3411), .Z(II3412) ) ;
NAND2   gate5562  (.A(g616), .B(II3411), .Z(II3413) ) ;
NAND2   gate5563  (.A(g1689), .B(g729), .Z(II3445) ) ;
NAND2   gate5564  (.A(g1689), .B(II3445), .Z(II3446) ) ;
NAND2   gate5565  (.A(g729), .B(II3445), .Z(II3447) ) ;
NAND2   gate5566  (.A(g1691), .B(g784), .Z(II3455) ) ;
NAND2   gate5567  (.A(g1691), .B(II3455), .Z(II3456) ) ;
NAND2   gate5568  (.A(g784), .B(II3455), .Z(II3457) ) ;
NAND2   gate5569  (.A(g1570), .B(g642), .Z(II3697) ) ;
NAND2   gate5570  (.A(g1570), .B(II3697), .Z(II3698) ) ;
NAND2   gate5571  (.A(g642), .B(II3697), .Z(II3699) ) ;
NAND2   gate5572  (.A(g2021), .B(g349), .Z(II3739) ) ;
NAND2   gate5573  (.A(g2021), .B(II3739), .Z(II3740) ) ;
NAND2   gate5574  (.A(g349), .B(II3739), .Z(II3741) ) ;
NAND2   gate5575  (.A(g284), .B(g2370), .Z(II3846) ) ;
NAND2   gate5576  (.A(g284), .B(II3846), .Z(II3847) ) ;
NAND2   gate5577  (.A(g2370), .B(II3846), .Z(II3848) ) ;
NAND2   gate5578  (.A(II3847), .B(II3848), .Z(g2698) ) ;
NAND2   gate5579  (.A(g285), .B(g2397), .Z(II3874) ) ;
NAND2   gate5580  (.A(g285), .B(II3874), .Z(II3875) ) ;
NAND2   gate5581  (.A(g2397), .B(II3874), .Z(II3876) ) ;
NAND2   gate5582  (.A(II3875), .B(II3876), .Z(g2719) ) ;
NAND2   gate5583  (.A(g286), .B(g2422), .Z(II3893) ) ;
NAND2   gate5584  (.A(g286), .B(II3893), .Z(II3894) ) ;
NAND2   gate5585  (.A(g2422), .B(II3893), .Z(II3895) ) ;
NAND2   gate5586  (.A(II3894), .B(II3895), .Z(g2731) ) ;
NAND2   gate5587  (.A(g287), .B(g2449), .Z(II3914) ) ;
NAND2   gate5588  (.A(g287), .B(II3914), .Z(II3915) ) ;
NAND2   gate5589  (.A(g2449), .B(II3914), .Z(II3916) ) ;
NAND2   gate5590  (.A(II3915), .B(II3916), .Z(g2745) ) ;
NAND2   gate5591  (.A(g288), .B(g2473), .Z(II3933) ) ;
NAND2   gate5592  (.A(g288), .B(II3933), .Z(II3934) ) ;
NAND2   gate5593  (.A(g2473), .B(II3933), .Z(II3935) ) ;
NAND2   gate5594  (.A(II3934), .B(II3935), .Z(g2757) ) ;
NAND2   gate5595  (.A(g289), .B(g2497), .Z(II3952) ) ;
NAND2   gate5596  (.A(g289), .B(II3952), .Z(II3953) ) ;
NAND2   gate5597  (.A(g2497), .B(II3952), .Z(II3954) ) ;
NAND2   gate5598  (.A(II3953), .B(II3954), .Z(g2769) ) ;
NAND2   gate5599  (.A(g290), .B(g2518), .Z(II3970) ) ;
NAND2   gate5600  (.A(g290), .B(II3970), .Z(II3971) ) ;
NAND2   gate5601  (.A(g2518), .B(II3970), .Z(II3972) ) ;
NAND2   gate5602  (.A(II3971), .B(II3972), .Z(g2780) ) ;
NAND2   gate5603  (.A(g291), .B(g2544), .Z(II3988) ) ;
NAND2   gate5604  (.A(g291), .B(II3988), .Z(II3989) ) ;
NAND2   gate5605  (.A(g2544), .B(II3988), .Z(II3990) ) ;
NAND2   gate5606  (.A(II3989), .B(II3990), .Z(g2791) ) ;
NAND2   gate5607  (.A(g1997), .B(g866), .Z(g2795) ) ;
NAND2   gate5608  (.A(g292), .B(g2568), .Z(II4008) ) ;
NAND2   gate5609  (.A(g292), .B(II4008), .Z(II4009) ) ;
NAND2   gate5610  (.A(g2568), .B(II4008), .Z(II4010) ) ;
NAND2   gate5611  (.A(II4009), .B(II4010), .Z(g2804) ) ;
NAND2   gate5612  (.A(g197), .B(g2381), .Z(g2940) ) ;
NAND2   gate5613  (.A(g269), .B(g2381), .Z(g2944) ) ;
NAND2   gate5614  (.A(g2551), .B(g139), .Z(II4150) ) ;
NAND2   gate5615  (.A(g2551), .B(II4150), .Z(II4151) ) ;
NAND2   gate5616  (.A(g139), .B(II4150), .Z(II4152) ) ;
NAND2   gate5617  (.A(g2015), .B(g619), .Z(II4159) ) ;
NAND2   gate5618  (.A(g2015), .B(II4159), .Z(II4160) ) ;
NAND2   gate5619  (.A(g619), .B(II4159), .Z(II4161) ) ;
NAND2   gate5620  (.A(g2292), .B(g749), .Z(II4182) ) ;
NAND2   gate5621  (.A(g2292), .B(II4182), .Z(II4183) ) ;
NAND2   gate5622  (.A(g749), .B(II4182), .Z(II4184) ) ;
NAND2   gate5623  (.A(g2255), .B(g743), .Z(II4203) ) ;
NAND2   gate5624  (.A(g2255), .B(II4203), .Z(II4204) ) ;
NAND2   gate5625  (.A(g743), .B(II4203), .Z(II4205) ) ;
NAND2   gate5626  (.A(g2294), .B(g804), .Z(II4210) ) ;
NAND2   gate5627  (.A(g2294), .B(II4210), .Z(II4211) ) ;
NAND2   gate5628  (.A(g804), .B(II4210), .Z(II4212) ) ;
NAND2   gate5629  (.A(g2267), .B(g798), .Z(II4233) ) ;
NAND2   gate5630  (.A(g2267), .B(II4233), .Z(II4234) ) ;
NAND2   gate5631  (.A(g798), .B(II4233), .Z(II4235) ) ;
NAND2   gate5632  (.A(g2360), .B(g1064), .Z(g3109) ) ;
NAND2   gate5633  (.A(g2092), .B(g606), .Z(II4444) ) ;
NAND2   gate5634  (.A(g2092), .B(II4444), .Z(II4445) ) ;
NAND2   gate5635  (.A(g606), .B(II4444), .Z(II4446) ) ;
NAND2   gate5636  (.A(g2909), .B(g646), .Z(II4526) ) ;
NAND2   gate5637  (.A(g2909), .B(II4526), .Z(II4527) ) ;
NAND2   gate5638  (.A(g646), .B(II4526), .Z(II4528) ) ;
NAND2   gate5639  (.A(g2853), .B(g353), .Z(II4545) ) ;
NAND2   gate5640  (.A(g2853), .B(II4545), .Z(II4546) ) ;
NAND2   gate5641  (.A(g353), .B(II4545), .Z(II4547) ) ;
NAND2   gate5642  (.A(g2846), .B(g622), .Z(II4782) ) ;
NAND2   gate5643  (.A(g2846), .B(II4782), .Z(II4783) ) ;
NAND2   gate5644  (.A(g622), .B(II4782), .Z(II4784) ) ;
NAND2   gate5645  (.A(g3522), .B(g650), .Z(II4919) ) ;
NAND2   gate5646  (.A(g3522), .B(II4919), .Z(II4920) ) ;
NAND2   gate5647  (.A(g650), .B(II4919), .Z(II4921) ) ;
NAND2   gate5648  (.A(g3437), .B(g357), .Z(II4939) ) ;
NAND2   gate5649  (.A(g3437), .B(II4939), .Z(II4940) ) ;
NAND2   gate5650  (.A(g357), .B(II4939), .Z(II4941) ) ;
NOR3    gate5651  (.A(g2804), .B(g2791), .C(g2780), .Z(g3664) ) ;
NOR3    gate5652  (.A(g2769), .B(g2757), .C(g2745), .Z(g3656) ) ;
NOR3    gate5653  (.A(g2731), .B(g2719), .C(g2698), .Z(g3647) ) ;
NAND2   gate5654  (.A(g3589), .B(g3593), .Z(II5187) ) ;
NAND2   gate5655  (.A(g3589), .B(II5187), .Z(II5188) ) ;
NAND2   gate5656  (.A(g3593), .B(II5187), .Z(II5189) ) ;
NAND2   gate5657  (.A(II5188), .B(II5189), .Z(g3955) ) ;
NAND2   gate5658  (.A(g3567), .B(g3571), .Z(II5195) ) ;
NAND2   gate5659  (.A(g3567), .B(II5195), .Z(II5196) ) ;
NAND2   gate5660  (.A(g3571), .B(II5195), .Z(II5197) ) ;
NAND2   gate5661  (.A(II5196), .B(II5197), .Z(g3957) ) ;
NAND2   gate5662  (.A(g3267), .B(g3271), .Z(II5207) ) ;
NAND2   gate5663  (.A(g3267), .B(II5207), .Z(II5208) ) ;
NAND2   gate5664  (.A(g3271), .B(II5207), .Z(II5209) ) ;
NAND2   gate5665  (.A(II5208), .B(II5209), .Z(g3961) ) ;
NAND2   gate5666  (.A(g3259), .B(g3263), .Z(II5226) ) ;
NAND2   gate5667  (.A(g3259), .B(II5226), .Z(II5227) ) ;
NAND2   gate5668  (.A(g3263), .B(II5226), .Z(II5228) ) ;
NAND2   gate5669  (.A(II5227), .B(II5228), .Z(g3968) ) ;
NAND2   gate5670  (.A(g3242), .B(g3247), .Z(II5242) ) ;
NAND2   gate5671  (.A(g3242), .B(II5242), .Z(II5243) ) ;
NAND2   gate5672  (.A(g3247), .B(II5242), .Z(II5244) ) ;
NAND2   gate5673  (.A(II5243), .B(II5244), .Z(g3974) ) ;
NAND2   gate5674  (.A(g3714), .B(g3719), .Z(II5257) ) ;
NAND2   gate5675  (.A(g3714), .B(II5257), .Z(II5258) ) ;
NAND2   gate5676  (.A(g3719), .B(II5257), .Z(II5259) ) ;
NAND2   gate5677  (.A(II5258), .B(II5259), .Z(g3979) ) ;
NAND2   gate5678  (.A(g3705), .B(g3710), .Z(II5269) ) ;
NAND2   gate5679  (.A(g3705), .B(II5269), .Z(II5270) ) ;
NAND2   gate5680  (.A(g3710), .B(II5269), .Z(II5271) ) ;
NAND2   gate5681  (.A(II5270), .B(II5271), .Z(g3983) ) ;
NAND2   gate5682  (.A(g3421), .B(g625), .Z(II5292) ) ;
NAND2   gate5683  (.A(g3421), .B(II5292), .Z(II5293) ) ;
NAND2   gate5684  (.A(g625), .B(II5292), .Z(II5294) ) ;
NAND2   gate5685  (.A(g471), .B(g3505), .Z(II5300) ) ;
NAND2   gate5686  (.A(g471), .B(II5300), .Z(II5301) ) ;
NAND2   gate5687  (.A(g3505), .B(II5300), .Z(II5302) ) ;
NAND2   gate5688  (.A(g478), .B(g3512), .Z(II5307) ) ;
NAND2   gate5689  (.A(g478), .B(II5307), .Z(II5308) ) ;
NAND2   gate5690  (.A(g3512), .B(II5307), .Z(II5309) ) ;
NAND2   gate5691  (.A(g3677), .B(g3425), .Z(g4049) ) ;
NAND2   gate5692  (.A(g3907), .B(g654), .Z(II5535) ) ;
NAND2   gate5693  (.A(g3907), .B(II5535), .Z(II5536) ) ;
NAND2   gate5694  (.A(g654), .B(II5535), .Z(II5537) ) ;
NAND2   gate5695  (.A(g3974), .B(g3968), .Z(II5647) ) ;
NAND2   gate5696  (.A(g3974), .B(II5647), .Z(II5648) ) ;
NAND2   gate5697  (.A(g3968), .B(II5647), .Z(II5649) ) ;
NAND2   gate5698  (.A(II5648), .B(II5649), .Z(g4221) ) ;
NAND2   gate5699  (.A(g3983), .B(g3979), .Z(II5657) ) ;
NAND2   gate5700  (.A(g3983), .B(II5657), .Z(II5658) ) ;
NAND2   gate5701  (.A(g3979), .B(II5657), .Z(II5659) ) ;
NAND2   gate5702  (.A(II5658), .B(II5659), .Z(g4223) ) ;
NAND2   gate5703  (.A(g3836), .B(g3503), .Z(II5759) ) ;
NAND2   gate5704  (.A(g3836), .B(II5759), .Z(II5760) ) ;
NAND2   gate5705  (.A(g3503), .B(II5759), .Z(II5761) ) ;
NAND2   gate5706  (.A(g3961), .B(g3957), .Z(II5766) ) ;
NAND2   gate5707  (.A(g3961), .B(II5766), .Z(II5767) ) ;
NAND2   gate5708  (.A(g3957), .B(II5766), .Z(II5768) ) ;
NAND2   gate5709  (.A(II5767), .B(II5768), .Z(g4301) ) ;
NAND2   gate5710  (.A(g3810), .B(g628), .Z(II5782) ) ;
NAND2   gate5711  (.A(g3810), .B(II5782), .Z(II5783) ) ;
NAND2   gate5712  (.A(g628), .B(II5782), .Z(II5784) ) ;
NAND2   gate5713  (.A(g3380), .B(g4253), .Z(g4472) ) ;
NAND2   gate5714  (.A(g4223), .B(g4221), .Z(II6026) ) ;
NAND2   gate5715  (.A(g4223), .B(II6026), .Z(II6027) ) ;
NAND2   gate5716  (.A(g4221), .B(II6026), .Z(II6028) ) ;
NAND2   gate5717  (.A(II6027), .B(II6028), .Z(g4504) ) ;
NAND2   gate5718  (.A(g4236), .B(g571), .Z(II6175) ) ;
NAND2   gate5719  (.A(g4236), .B(II6175), .Z(II6176) ) ;
NAND2   gate5720  (.A(g571), .B(II6175), .Z(II6177) ) ;
NAND2   gate5721  (.A(g4301), .B(g3955), .Z(II6185) ) ;
NAND2   gate5722  (.A(g4301), .B(II6185), .Z(II6186) ) ;
NAND2   gate5723  (.A(g3955), .B(II6185), .Z(II6187) ) ;
NAND2   gate5724  (.A(II6186), .B(II6187), .Z(g4610) ) ;
NAND2   gate5725  (.A(g4199), .B(g631), .Z(II6194) ) ;
NAND2   gate5726  (.A(g4199), .B(II6194), .Z(II6195) ) ;
NAND2   gate5727  (.A(g631), .B(II6194), .Z(II6196) ) ;
NOR2    gate5728  (.A(g1802), .B(g3167), .Z(g3528) ) ;
NAND4   gate5729  (.A(g4550), .B(g1514), .C(g2107), .D(g2897), .Z(g4674) ) ;
NAND4   gate5730  (.A(g4550), .B(g1514), .C(g1006), .D(g2897), .Z(g4680) ) ;
NAND2   gate5731  (.A(g4504), .B(g4610), .Z(II6390) ) ;
NAND2   gate5732  (.A(g4504), .B(II6390), .Z(II6391) ) ;
NAND2   gate5733  (.A(g4610), .B(II6390), .Z(II6392) ) ;
NAND2   gate5734  (.A(II6391), .B(II6392), .Z(g4762) ) ;
NAND2   gate5735  (.A(g4541), .B(g578), .Z(II6473) ) ;
NAND2   gate5736  (.A(g4541), .B(II6473), .Z(II6474) ) ;
NAND2   gate5737  (.A(g578), .B(II6473), .Z(II6475) ) ;
NOR2    gate5738  (.A(g996), .B(g980), .Z(g1560) ) ;
NOR2    gate5739  (.A(g980), .B(g965), .Z(g1518) ) ;
NAND2   gate5740  (.A(g4504), .B(g3541), .Z(II6499) ) ;
NAND2   gate5741  (.A(g4504), .B(II6499), .Z(II6500) ) ;
NAND2   gate5742  (.A(g3541), .B(II6499), .Z(II6501) ) ;
NAND2   gate5743  (.A(g4762), .B(g3541), .Z(II6659) ) ;
NAND2   gate5744  (.A(g4762), .B(II6659), .Z(II6660) ) ;
NAND2   gate5745  (.A(g3541), .B(II6659), .Z(II6661) ) ;
NAND2   gate5746  (.A(g4708), .B(g582), .Z(II6743) ) ;
NAND2   gate5747  (.A(g4708), .B(II6743), .Z(II6744) ) ;
NAND2   gate5748  (.A(g582), .B(II6743), .Z(II6745) ) ;
NAND2   gate5749  (.A(g4874), .B(g586), .Z(II6962) ) ;
NAND2   gate5750  (.A(g4874), .B(II6962), .Z(II6963) ) ;
NAND2   gate5751  (.A(g586), .B(II6962), .Z(II6964) ) ;
NAND2   gate5752  (.A(g5194), .B(g574), .Z(II7097) ) ;
NAND2   gate5753  (.A(g5194), .B(II7097), .Z(II7098) ) ;
NAND2   gate5754  (.A(g574), .B(II7097), .Z(II7099) ) ;
NAND2   gate5755  (.A(g143), .B(g5367), .Z(II7208) ) ;
NAND2   gate5756  (.A(g143), .B(II7208), .Z(II7209) ) ;
NAND2   gate5757  (.A(g5367), .B(II7208), .Z(II7210) ) ;
NAND2   gate5758  (.A(g152), .B(g5368), .Z(II7216) ) ;
NAND2   gate5759  (.A(g152), .B(II7216), .Z(II7217) ) ;
NAND2   gate5760  (.A(g5368), .B(II7216), .Z(II7218) ) ;
NAND2   gate5761  (.A(g161), .B(g5370), .Z(II7223) ) ;
NAND2   gate5762  (.A(g161), .B(II7223), .Z(II7224) ) ;
NAND2   gate5763  (.A(g5370), .B(II7223), .Z(II7225) ) ;
NAND2   gate5764  (.A(g170), .B(g5372), .Z(II7230) ) ;
NAND2   gate5765  (.A(g170), .B(II7230), .Z(II7231) ) ;
NAND2   gate5766  (.A(g5372), .B(II7230), .Z(II7232) ) ;
NAND2   gate5767  (.A(g179), .B(g5374), .Z(II7237) ) ;
NAND2   gate5768  (.A(g179), .B(II7237), .Z(II7238) ) ;
NAND2   gate5769  (.A(g5374), .B(II7237), .Z(II7239) ) ;
NAND2   gate5770  (.A(g188), .B(g5377), .Z(II7244) ) ;
NAND2   gate5771  (.A(g188), .B(II7244), .Z(II7245) ) ;
NAND2   gate5772  (.A(g5377), .B(II7244), .Z(II7246) ) ;
NAND2   gate5773  (.A(g5364), .B(g590), .Z(II7311) ) ;
NAND2   gate5774  (.A(g5364), .B(II7311), .Z(II7312) ) ;
NAND2   gate5775  (.A(g590), .B(II7311), .Z(II7313) ) ;
NAND2   gate5776  (.A(g111), .B(g5554), .Z(II7432) ) ;
NAND2   gate5777  (.A(g111), .B(II7432), .Z(II7433) ) ;
NAND2   gate5778  (.A(g5554), .B(II7432), .Z(II7434) ) ;
NAND2   gate5779  (.A(g5515), .B(g594), .Z(II7439) ) ;
NAND2   gate5780  (.A(g5515), .B(II7439), .Z(II7440) ) ;
NAND2   gate5781  (.A(g594), .B(II7439), .Z(II7441) ) ;
NAND4   gate5782  (.A(g5546), .B(g1585), .C(g2084), .D(g2916), .Z(g5688) ) ;
NAND2   gate5783  (.A(g361), .B(g5659), .Z(II7520) ) ;
NAND2   gate5784  (.A(g361), .B(II7520), .Z(II7521) ) ;
NAND2   gate5785  (.A(g5659), .B(II7520), .Z(II7522) ) ;
NAND2   gate5786  (.A(g49), .B(g5662), .Z(II7527) ) ;
NAND2   gate5787  (.A(g49), .B(II7527), .Z(II7528) ) ;
NAND2   gate5788  (.A(g5662), .B(II7527), .Z(II7529) ) ;
NAND2   gate5789  (.A(g54), .B(g5666), .Z(II7534) ) ;
NAND2   gate5790  (.A(g54), .B(II7534), .Z(II7535) ) ;
NAND2   gate5791  (.A(g5666), .B(II7534), .Z(II7536) ) ;
NAND2   gate5792  (.A(g59), .B(g5669), .Z(II7541) ) ;
NAND2   gate5793  (.A(g59), .B(II7541), .Z(II7542) ) ;
NAND2   gate5794  (.A(g5669), .B(II7541), .Z(II7543) ) ;
NAND2   gate5795  (.A(g64), .B(g5672), .Z(II7548) ) ;
NAND2   gate5796  (.A(g64), .B(II7548), .Z(II7549) ) ;
NAND2   gate5797  (.A(g5672), .B(II7548), .Z(II7550) ) ;
NAND2   gate5798  (.A(g69), .B(g5674), .Z(II7555) ) ;
NAND2   gate5799  (.A(g69), .B(II7555), .Z(II7556) ) ;
NAND2   gate5800  (.A(g5674), .B(II7555), .Z(II7557) ) ;
NAND2   gate5801  (.A(g74), .B(g5676), .Z(II7562) ) ;
NAND2   gate5802  (.A(g74), .B(II7562), .Z(II7563) ) ;
NAND2   gate5803  (.A(g5676), .B(II7562), .Z(II7564) ) ;
NAND2   gate5804  (.A(g79), .B(g5678), .Z(II7569) ) ;
NAND2   gate5805  (.A(g79), .B(II7569), .Z(II7570) ) ;
NAND2   gate5806  (.A(g5678), .B(II7569), .Z(II7571) ) ;
NAND2   gate5807  (.A(g84), .B(g5680), .Z(II7576) ) ;
NAND2   gate5808  (.A(g84), .B(II7576), .Z(II7577) ) ;
NAND2   gate5809  (.A(g5680), .B(II7576), .Z(II7578) ) ;
NAND4   gate5810  (.A(g5649), .B(g1529), .C(g1535), .D(g2068), .Z(g5862) ) ;
NAND4   gate5811  (.A(g5649), .B(g1076), .C(g1535), .D(g2068), .Z(g5863) ) ;
NAND2   gate5812  (.A(g471), .B(g6188), .Z(II8194) ) ;
NAND2   gate5813  (.A(g471), .B(II8194), .Z(II8195) ) ;
NAND2   gate5814  (.A(g6188), .B(II8194), .Z(II8196) ) ;
NAND2   gate5815  (.A(g478), .B(g6192), .Z(II8201) ) ;
NAND2   gate5816  (.A(g478), .B(II8201), .Z(II8202) ) ;
NAND2   gate5817  (.A(g6192), .B(II8201), .Z(II8203) ) ;
NAND2   gate5818  (.A(g6832), .B(g3598), .Z(II9050) ) ;
NAND2   gate5819  (.A(g6832), .B(II9050), .Z(II9051) ) ;
NAND2   gate5820  (.A(g3598), .B(II9050), .Z(II9052) ) ;
NOR2    gate5821  (.A(g1407), .B(g2842), .Z(g3621) ) ;
NOR2    gate5822  (.A(g486), .B(g943), .Z(g1418) ) ;
NOR2    gate5823  (.A(g489), .B(g1048), .Z(g1449) ) ;
NOR2    gate5824  (.A(g1603), .B(g1416), .Z(g1879) ) ;

endmodule
