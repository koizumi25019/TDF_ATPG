module s38584 (g35, g36, g6744, g6745, g6746
    , g6747, g6748, g6749, g6750, g6751
    , g6752, g6753, CLK
    , g7243, g7245, g7257, g7260, g7540
    , g7916, g7946, g8132, g8178, g8215
    , g8235, g8277, g8279, g8283, g8291
    , g8342, g8344, g8353, g8358, g8398
    , g8403, g8416, g8475, g8719, g8783
    , g8784, g8785, g8786, g8787, g8788
    , g8789, g8839, g8870, g8915, g8916
    , g8917, g8918, g8919, g8920, g9019
    , g9048, g9251, g9497, g9553, g9555
    , g9615, g9617, g9680, g9682, g9741
    , g9743, g9817, g10122, g10306, g10500
    , g10527, g11349, g11388, g11418, g11447
    , g11678, g11770, g12184, g12238, g12300
    , g12350, g12368, g12422, g12470, g12832
    , g12919, g12923, g13039, g13049, g13068
    , g13085, g13099, g13259, g13272, g13865
    , g13881, g13895, g13906, g13926, g13966
    , g14096, g14125, g14147, g14167, g14189
    , g14201, g14217, g14421, g14451, g14518
    , g14597, g14635, g14662, g14673, g14694
    , g14705, g14738, g14749, g14779, g14828
    , g16603, g16624, g16627, g16656, g16659
    , g16686, g16693, g16718, g16722, g16744
    , g16748, g16775, g16874, g16924, g16955
    , g17291, g17316, g17320, g17400, g17404
    , g17423, g17519, g17577, g17580, g17604
    , g17607, g17639, g17646, g17649, g17674
    , g17678, g17685, g17688, g17711, g17715
    , g17722, g17739, g17743, g17760, g17764
    , g17778, g17787, g17813, g17819, g17845
    , g17871, g18092, g18094, g18095, g18096
    , g18097, g18098, g18099, g18100, g18101
    , g18881, g19334, g19357, g20049, g20557
    , g20652, g20654, g20763, g20899, g20901
    , g21176, g21245, g21270, g21292, g21698
    , g21727, g23002, g23190, g23612, g23652
    , g23683, g23759, g24151, g25114, g25167
    , g25219, g25259, g25582, g25583, g25584
    , g25585, g25586, g25587, g25588, g25589
    , g25590, g26801, g26875, g26876, g26877
    , g27831, g28030, g28041, g28042, g28753
    , g29210, g29211, g29212, g29213, g29214
    , g29215, g29216, g29217, g29218, g29219
    , g29220, g29221, g30327, g30329, g30330
    , g30331, g30332, g31521, g31656, g31665
    , g31793, g31860, g31861, g31862, g31863
    , g32185, g32429, g32454, g32975, g33079
    , g33435, g33533, g33636, g33659, g33874
    , g33894, g33935, g33945, g33946, g33947
    , g33948, g33949, g33950, g33959, g34201
    , g34221, g34232, g34233, g34234, g34235
    , g34236, g34237, g34238, g34239, g34240
    , g34383, g34425, g34435, g34436, g34437
    , g34597, g34788, g34839, g34913, g34915
    , g34917, g34919, g34921, g34923, g34925
    , g34927, g34956, g34972) ;

input   g35, g36, g6744, g6745, g6746
    , g6747, g6748, g6749, g6750, g6751
    , g6752, g6753, CLK ;

output  g7243, g7245, g7257, g7260, g7540
    , g7916, g7946, g8132, g8178, g8215
    , g8235, g8277, g8279, g8283, g8291
    , g8342, g8344, g8353, g8358, g8398
    , g8403, g8416, g8475, g8719, g8783
    , g8784, g8785, g8786, g8787, g8788
    , g8789, g8839, g8870, g8915, g8916
    , g8917, g8918, g8919, g8920, g9019
    , g9048, g9251, g9497, g9553, g9555
    , g9615, g9617, g9680, g9682, g9741
    , g9743, g9817, g10122, g10306, g10500
    , g10527, g11349, g11388, g11418, g11447
    , g11678, g11770, g12184, g12238, g12300
    , g12350, g12368, g12422, g12470, g12832
    , g12919, g12923, g13039, g13049, g13068
    , g13085, g13099, g13259, g13272, g13865
    , g13881, g13895, g13906, g13926, g13966
    , g14096, g14125, g14147, g14167, g14189
    , g14201, g14217, g14421, g14451, g14518
    , g14597, g14635, g14662, g14673, g14694
    , g14705, g14738, g14749, g14779, g14828
    , g16603, g16624, g16627, g16656, g16659
    , g16686, g16693, g16718, g16722, g16744
    , g16748, g16775, g16874, g16924, g16955
    , g17291, g17316, g17320, g17400, g17404
    , g17423, g17519, g17577, g17580, g17604
    , g17607, g17639, g17646, g17649, g17674
    , g17678, g17685, g17688, g17711, g17715
    , g17722, g17739, g17743, g17760, g17764
    , g17778, g17787, g17813, g17819, g17845
    , g17871, g18092, g18094, g18095, g18096
    , g18097, g18098, g18099, g18100, g18101
    , g18881, g19334, g19357, g20049, g20557
    , g20652, g20654, g20763, g20899, g20901
    , g21176, g21245, g21270, g21292, g21698
    , g21727, g23002, g23190, g23612, g23652
    , g23683, g23759, g24151, g25114, g25167
    , g25219, g25259, g25582, g25583, g25584
    , g25585, g25586, g25587, g25588, g25589
    , g25590, g26801, g26875, g26876, g26877
    , g27831, g28030, g28041, g28042, g28753
    , g29210, g29211, g29212, g29213, g29214
    , g29215, g29216, g29217, g29218, g29219
    , g29220, g29221, g30327, g30329, g30330
    , g30331, g30332, g31521, g31656, g31665
    , g31793, g31860, g31861, g31862, g31863
    , g32185, g32429, g32454, g32975, g33079
    , g33435, g33533, g33636, g33659, g33874
    , g33894, g33935, g33945, g33946, g33947
    , g33948, g33949, g33950, g33959, g34201
    , g34221, g34232, g34233, g34234, g34235
    , g34236, g34237, g34238, g34239, g34240
    , g34383, g34425, g34435, g34436, g34437
    , g34597, g34788, g34839, g34913, g34915
    , g34917, g34919, g34921, g34923, g34925
    , g34927, g34956, g34972 ;

INV     gate0  (.A(II11892), .Z(g7243) ) ;
INV     gate1  (.A(II11896), .Z(g7245) ) ;
INV     gate2  (.A(II11903), .Z(g7257) ) ;
INV     gate3  (.A(II11908), .Z(g7260) ) ;
INV     gate4  (.A(II12026), .Z(g7540) ) ;
INV     gate5  (.A(II12300), .Z(g7916) ) ;
INV     gate6  (.A(II12314), .Z(g7946) ) ;
INV     gate7  (.A(II12411), .Z(g8132) ) ;
INV     gate8  (.A(II12437), .Z(g8178) ) ;
INV     gate9  (.A(II12451), .Z(g8215) ) ;
INV     gate10  (.A(II12463), .Z(g8235) ) ;
INV     gate11  (.A(II12483), .Z(g8277) ) ;
INV     gate12  (.A(II12487), .Z(g8279) ) ;
INV     gate13  (.A(II12493), .Z(g8283) ) ;
INV     gate14  (.A(II12503), .Z(g8291) ) ;
INV     gate15  (.A(II12519), .Z(g8342) ) ;
INV     gate16  (.A(II12523), .Z(g8344) ) ;
INV     gate17  (.A(II12530), .Z(g8353) ) ;
INV     gate18  (.A(II12541), .Z(g8358) ) ;
INV     gate19  (.A(II12563), .Z(g8398) ) ;
INV     gate20  (.A(II12568), .Z(g8403) ) ;
INV     gate21  (.A(II12580), .Z(g8416) ) ;
INV     gate22  (.A(II12608), .Z(g8475) ) ;
INV     gate23  (.A(II12719), .Z(g8719) ) ;
INV     gate24  (.A(II12761), .Z(g8783) ) ;
INV     gate25  (.A(II12764), .Z(g8784) ) ;
INV     gate26  (.A(II12767), .Z(g8785) ) ;
INV     gate27  (.A(II12770), .Z(g8786) ) ;
INV     gate28  (.A(II12773), .Z(g8787) ) ;
INV     gate29  (.A(II12776), .Z(g8788) ) ;
INV     gate30  (.A(II12779), .Z(g8789) ) ;
INV     gate31  (.A(II12819), .Z(g8839) ) ;
INV     gate32  (.A(II12837), .Z(g8870) ) ;
INV     gate33  (.A(II12884), .Z(g8915) ) ;
INV     gate34  (.A(II12887), .Z(g8916) ) ;
INV     gate35  (.A(II12890), .Z(g8917) ) ;
INV     gate36  (.A(II12893), .Z(g8918) ) ;
INV     gate37  (.A(II12896), .Z(g8919) ) ;
INV     gate38  (.A(II12899), .Z(g8920) ) ;
INV     gate39  (.A(II12950), .Z(g9019) ) ;
INV     gate40  (.A(II12963), .Z(g9048) ) ;
INV     gate41  (.A(II13037), .Z(g9251) ) ;
INV     gate42  (.A(II13166), .Z(g9497) ) ;
INV     gate43  (.A(II13202), .Z(g9553) ) ;
INV     gate44  (.A(II13206), .Z(g9555) ) ;
INV     gate45  (.A(II13236), .Z(g9615) ) ;
INV     gate46  (.A(II13240), .Z(g9617) ) ;
INV     gate47  (.A(II13276), .Z(g9680) ) ;
INV     gate48  (.A(II13280), .Z(g9682) ) ;
INV     gate49  (.A(II13317), .Z(g9741) ) ;
INV     gate50  (.A(II13321), .Z(g9743) ) ;
INV     gate51  (.A(II13374), .Z(g9817) ) ;
INV     gate52  (.A(II13623), .Z(g10122) ) ;
INV     gate53  (.A(II13726), .Z(g10306) ) ;
INV     gate54  (.A(II13875), .Z(g10500) ) ;
INV     gate55  (.A(II13892), .Z(g10527) ) ;
INV     gate56  (.A(II14365), .Z(g11349) ) ;
INV     gate57  (.A(II14395), .Z(g11388) ) ;
INV     gate58  (.A(II14424), .Z(g11418) ) ;
INV     gate59  (.A(II14450), .Z(g11447) ) ;
INV     gate60  (.A(II14563), .Z(g11678) ) ;
INV     gate61  (.A(II14619), .Z(g11770) ) ;
INV     gate62  (.A(II15036), .Z(g12184) ) ;
INV     gate63  (.A(II15102), .Z(g12238) ) ;
INV     gate64  (.A(II15144), .Z(g12300) ) ;
INV     gate65  (.A(II15190), .Z(g12350) ) ;
INV     gate66  (.A(II15208), .Z(g12368) ) ;
INV     gate67  (.A(II15238), .Z(g12422) ) ;
INV     gate68  (.A(II15284), .Z(g12470) ) ;
OR2     gate69  (.A(g10347), .B(g10348), .Z(g12832) ) ;
INV     gate70  (.A(II15536), .Z(g12919) ) ;
INV     gate71  (.A(II15542), .Z(g12923) ) ;
INV     gate72  (.A(II15663), .Z(g13039) ) ;
INV     gate73  (.A(II15677), .Z(g13049) ) ;
INV     gate74  (.A(II15697), .Z(g13068) ) ;
INV     gate75  (.A(II15717), .Z(g13085) ) ;
INV     gate76  (.A(II15732), .Z(g13099) ) ;
INV     gate77  (.A(II15824), .Z(g13259) ) ;
INV     gate78  (.A(II15837), .Z(g13272) ) ;
INV     gate79  (.A(II16168), .Z(g13865) ) ;
INV     gate80  (.A(II16181), .Z(g13881) ) ;
INV     gate81  (.A(II16193), .Z(g13895) ) ;
INV     gate82  (.A(II16201), .Z(g13906) ) ;
INV     gate83  (.A(II16217), .Z(g13926) ) ;
INV     gate84  (.A(II16246), .Z(g13966) ) ;
INV     gate85  (.A(II16328), .Z(g14096) ) ;
INV     gate86  (.A(II16345), .Z(g14125) ) ;
INV     gate87  (.A(II16357), .Z(g14147) ) ;
INV     gate88  (.A(II16371), .Z(g14167) ) ;
INV     gate89  (.A(II16391), .Z(g14189) ) ;
INV     gate90  (.A(II16401), .Z(g14201) ) ;
INV     gate91  (.A(II16417), .Z(g14217) ) ;
INV     gate92  (.A(II16575), .Z(g14421) ) ;
INV     gate93  (.A(II16606), .Z(g14451) ) ;
INV     gate94  (.A(II16639), .Z(g14518) ) ;
INV     gate95  (.A(II16713), .Z(g14597) ) ;
INV     gate96  (.A(II16741), .Z(g14635) ) ;
INV     gate97  (.A(II16762), .Z(g14662) ) ;
INV     gate98  (.A(II16770), .Z(g14673) ) ;
INV     gate99  (.A(II16795), .Z(g14694) ) ;
INV     gate100  (.A(II16803), .Z(g14705) ) ;
INV     gate101  (.A(II16821), .Z(g14738) ) ;
INV     gate102  (.A(II16829), .Z(g14749) ) ;
INV     gate103  (.A(II16847), .Z(g14779) ) ;
INV     gate104  (.A(II16875), .Z(g14828) ) ;
INV     gate105  (.A(II17787), .Z(g16603) ) ;
INV     gate106  (.A(II17814), .Z(g16624) ) ;
INV     gate107  (.A(II17819), .Z(g16627) ) ;
INV     gate108  (.A(II17852), .Z(g16656) ) ;
INV     gate109  (.A(II17857), .Z(g16659) ) ;
INV     gate110  (.A(II17892), .Z(g16686) ) ;
INV     gate111  (.A(II17901), .Z(g16693) ) ;
INV     gate112  (.A(II17932), .Z(g16718) ) ;
INV     gate113  (.A(II17938), .Z(g16722) ) ;
INV     gate114  (.A(II17964), .Z(g16744) ) ;
INV     gate115  (.A(II17970), .Z(g16748) ) ;
INV     gate116  (.A(II17999), .Z(g16775) ) ;
INV     gate117  (.A(II18066), .Z(g16874) ) ;
INV     gate118  (.A(II18092), .Z(g16924) ) ;
INV     gate119  (.A(II18107), .Z(g16955) ) ;
INV     gate120  (.A(II18276), .Z(g17291) ) ;
INV     gate121  (.A(II18293), .Z(g17316) ) ;
INV     gate122  (.A(II18297), .Z(g17320) ) ;
INV     gate123  (.A(II18333), .Z(g17400) ) ;
INV     gate124  (.A(II18337), .Z(g17404) ) ;
INV     gate125  (.A(II18360), .Z(g17423) ) ;
INV     gate126  (.A(II18460), .Z(g17519) ) ;
INV     gate127  (.A(II18504), .Z(g17577) ) ;
INV     gate128  (.A(II18509), .Z(g17580) ) ;
INV     gate129  (.A(II18555), .Z(g17604) ) ;
INV     gate130  (.A(II18560), .Z(g17607) ) ;
INV     gate131  (.A(II18600), .Z(g17639) ) ;
INV     gate132  (.A(II18609), .Z(g17646) ) ;
INV     gate133  (.A(II18614), .Z(g17649) ) ;
INV     gate134  (.A(II18647), .Z(g17674) ) ;
INV     gate135  (.A(II18653), .Z(g17678) ) ;
INV     gate136  (.A(II18662), .Z(g17685) ) ;
INV     gate137  (.A(II18667), .Z(g17688) ) ;
INV     gate138  (.A(II18694), .Z(g17711) ) ;
INV     gate139  (.A(II18700), .Z(g17715) ) ;
INV     gate140  (.A(II18709), .Z(g17722) ) ;
INV     gate141  (.A(II18728), .Z(g17739) ) ;
INV     gate142  (.A(II18734), .Z(g17743) ) ;
INV     gate143  (.A(II18752), .Z(g17760) ) ;
INV     gate144  (.A(II18758), .Z(g17764) ) ;
INV     gate145  (.A(II18778), .Z(g17778) ) ;
INV     gate146  (.A(II18795), .Z(g17787) ) ;
INV     gate147  (.A(II18813), .Z(g17813) ) ;
INV     gate148  (.A(II18825), .Z(g17819) ) ;
INV     gate149  (.A(II18835), .Z(g17845) ) ;
INV     gate150  (.A(II18845), .Z(g17871) ) ;
INV     gate151  (.A(II18882), .Z(g18092) ) ;
INV     gate152  (.A(II18888), .Z(g18094) ) ;
INV     gate153  (.A(II18891), .Z(g18095) ) ;
INV     gate154  (.A(II18894), .Z(g18096) ) ;
INV     gate155  (.A(II18897), .Z(g18097) ) ;
INV     gate156  (.A(II18900), .Z(g18098) ) ;
INV     gate157  (.A(II18903), .Z(g18099) ) ;
INV     gate158  (.A(II18906), .Z(g18100) ) ;
INV     gate159  (.A(II18909), .Z(g18101) ) ;
INV     gate160  (.A(II19671), .Z(g18881) ) ;
INV     gate161  (.A(II19818), .Z(g19334) ) ;
INV     gate162  (.A(II19837), .Z(g19357) ) ;
INV     gate163  (.A(II20318), .Z(g20049) ) ;
INV     gate164  (.A(II20647), .Z(g20557) ) ;
INV     gate165  (.A(II20744), .Z(g20652) ) ;
INV     gate166  (.A(II20750), .Z(g20654) ) ;
INV     gate167  (.A(II20816), .Z(g20763) ) ;
INV     gate168  (.A(II20861), .Z(g20899) ) ;
INV     gate169  (.A(II20867), .Z(g20901) ) ;
INV     gate170  (.A(II20954), .Z(g21176) ) ;
INV     gate171  (.A(II20982), .Z(g21245) ) ;
INV     gate172  (.A(II20999), .Z(g21270) ) ;
INV     gate173  (.A(II21033), .Z(g21292) ) ;
INV     gate174  (.A(g18562), .Z(g21698) ) ;
INV     gate175  (.A(II21300), .Z(g21727) ) ;
INV     gate176  (.A(II22177), .Z(g23002) ) ;
INV     gate177  (.A(II22286), .Z(g23190) ) ;
INV     gate178  (.A(II22745), .Z(g23612) ) ;
INV     gate179  (.A(II22785), .Z(g23652) ) ;
INV     gate180  (.A(II22816), .Z(g23683) ) ;
INV     gate181  (.A(II22886), .Z(g23759) ) ;
OR2     gate182  (.A(g18088), .B(g21661), .Z(g24151) ) ;
INV     gate183  (.A(II24278), .Z(g25114) ) ;
INV     gate184  (.A(II24331), .Z(g25167) ) ;
INV     gate185  (.A(II24393), .Z(g25219) ) ;
INV     gate186  (.A(II24445), .Z(g25259) ) ;
OR2     gate187  (.A(g21662), .B(g24152), .Z(g25582) ) ;
OR2     gate188  (.A(g21666), .B(g24153), .Z(g25583) ) ;
OR2     gate189  (.A(g21670), .B(g24154), .Z(g25584) ) ;
OR2     gate190  (.A(g21674), .B(g24155), .Z(g25585) ) ;
OR2     gate191  (.A(g21678), .B(g24156), .Z(g25586) ) ;
OR2     gate192  (.A(g21682), .B(g24157), .Z(g25587) ) ;
OR2     gate193  (.A(g21686), .B(g24158), .Z(g25588) ) ;
OR2     gate194  (.A(g21690), .B(g24159), .Z(g25589) ) ;
OR2     gate195  (.A(g21694), .B(g24160), .Z(g25590) ) ;
INV     gate196  (.A(II25511), .Z(g26801) ) ;
OR2     gate197  (.A(g21652), .B(g25575), .Z(g26875) ) ;
OR2     gate198  (.A(g21655), .B(g25576), .Z(g26876) ) ;
OR2     gate199  (.A(g21658), .B(g25577), .Z(g26877) ) ;
INV     gate200  (.A(II26406), .Z(g27831) ) ;
OR2     gate201  (.A(g24018), .B(g26874), .Z(g28030) ) ;
OR2     gate202  (.A(g24145), .B(g26878), .Z(g28041) ) ;
OR2     gate203  (.A(g24148), .B(g26879), .Z(g28042) ) ;
INV     gate204  (.A(II27235), .Z(g28753) ) ;
INV     gate205  (.A(II27546), .Z(g29210) ) ;
INV     gate206  (.A(II27549), .Z(g29211) ) ;
INV     gate207  (.A(II27552), .Z(g29212) ) ;
INV     gate208  (.A(II27555), .Z(g29213) ) ;
INV     gate209  (.A(II27558), .Z(g29214) ) ;
INV     gate210  (.A(II27561), .Z(g29215) ) ;
INV     gate211  (.A(II27564), .Z(g29216) ) ;
INV     gate212  (.A(II27567), .Z(g29217) ) ;
INV     gate213  (.A(II27570), .Z(g29218) ) ;
INV     gate214  (.A(II27573), .Z(g29219) ) ;
INV     gate215  (.A(II27576), .Z(g29220) ) ;
INV     gate216  (.A(II27579), .Z(g29221) ) ;
INV     gate217  (.A(II28582), .Z(g30327) ) ;
INV     gate218  (.A(II28588), .Z(g30329) ) ;
INV     gate219  (.A(II28591), .Z(g30330) ) ;
INV     gate220  (.A(II28594), .Z(g30331) ) ;
INV     gate221  (.A(II28597), .Z(g30332) ) ;
INV     gate222  (.A(II29182), .Z(g31521) ) ;
INV     gate223  (.A(II29236), .Z(g31656) ) ;
INV     gate224  (.A(II29245), .Z(g31665) ) ;
OR2     gate225  (.A(g28031), .B(g30317), .Z(g31793) ) ;
INV     gate226  (.A(II29438), .Z(g31860) ) ;
INV     gate227  (.A(II29441), .Z(g31861) ) ;
INV     gate228  (.A(II29444), .Z(g31862) ) ;
INV     gate229  (.A(II29447), .Z(g31863) ) ;
INV     gate230  (.A(II29717), .Z(g32185) ) ;
OR2     gate231  (.A(g30318), .B(g31794), .Z(g32429) ) ;
OR2     gate232  (.A(g30322), .B(g31795), .Z(g32454) ) ;
INV     gate233  (.A(II30537), .Z(g32975) ) ;
INV     gate234  (.A(II30641), .Z(g33079) ) ;
INV     gate235  (.A(II30959), .Z(g33435) ) ;
INV     gate236  (.A(II31361), .Z(g33533) ) ;
INV     gate237  (.A(II31463), .Z(g33636) ) ;
INV     gate238  (.A(II31491), .Z(g33659) ) ;
INV     gate239  (.A(II31724), .Z(g33874) ) ;
INV     gate240  (.A(II31748), .Z(g33894) ) ;
INV     gate241  (.A(II31817), .Z(g33935) ) ;
OR2     gate242  (.A(g32430), .B(g33455), .Z(g33945) ) ;
OR2     gate243  (.A(g32434), .B(g33456), .Z(g33946) ) ;
OR2     gate244  (.A(g32438), .B(g33457), .Z(g33947) ) ;
OR2     gate245  (.A(g32442), .B(g33458), .Z(g33948) ) ;
OR2     gate246  (.A(g32446), .B(g33459), .Z(g33949) ) ;
OR2     gate247  (.A(g32450), .B(g33460), .Z(g33950) ) ;
INV     gate248  (.A(II31878), .Z(g33959) ) ;
INV     gate249  (.A(II32158), .Z(g34201) ) ;
INV     gate250  (.A(II32192), .Z(g34221) ) ;
OR2     gate251  (.A(g33451), .B(g33944), .Z(g34232) ) ;
OR2     gate252  (.A(g32455), .B(g33951), .Z(g34233) ) ;
OR2     gate253  (.A(g32520), .B(g33952), .Z(g34234) ) ;
OR2     gate254  (.A(g32585), .B(g33953), .Z(g34235) ) ;
OR2     gate255  (.A(g32650), .B(g33954), .Z(g34236) ) ;
OR2     gate256  (.A(g32715), .B(g33955), .Z(g34237) ) ;
OR2     gate257  (.A(g32780), .B(g33956), .Z(g34238) ) ;
OR2     gate258  (.A(g32845), .B(g33957), .Z(g34239) ) ;
OR2     gate259  (.A(g32910), .B(g33958), .Z(g34240) ) ;
INV     gate260  (.A(II32388), .Z(g34383) ) ;
INV     gate261  (.A(II32446), .Z(g34425) ) ;
INV     gate262  (.A(II32476), .Z(g34435) ) ;
INV     gate263  (.A(II32479), .Z(g34436) ) ;
INV     gate264  (.A(II32482), .Z(g34437) ) ;
INV     gate265  (.A(II32699), .Z(g34597) ) ;
INV     gate266  (.A(II32994), .Z(g34788) ) ;
INV     gate267  (.A(II33053), .Z(g34839) ) ;
INV     gate268  (.A(II33131), .Z(g34913) ) ;
INV     gate269  (.A(II33137), .Z(g34915) ) ;
INV     gate270  (.A(II33143), .Z(g34917) ) ;
INV     gate271  (.A(II33149), .Z(g34919) ) ;
INV     gate272  (.A(II33155), .Z(g34921) ) ;
INV     gate273  (.A(II33161), .Z(g34923) ) ;
INV     gate274  (.A(II33167), .Z(g34925) ) ;
INV     gate275  (.A(II33173), .Z(g34927) ) ;
INV     gate276  (.A(II33214), .Z(g34956) ) ;
INV     gate277  (.A(II33232), .Z(g34972) ) ;
INV     gate278  (.A(II23342), .Z(g24166) ) ;
DFF     gate279  (.D(g24166), .CP(CLK), .Q(g72) ) ;
INV     gate280  (.A(II23345), .Z(g24167) ) ;
DFF     gate281  (.D(g24167), .CP(CLK), .Q(g73) ) ;
INV     gate282  (.A(II23348), .Z(g24168) ) ;
DFF     gate283  (.D(g24168), .CP(CLK), .Q(g84) ) ;
INV     gate284  (.A(II23351), .Z(g24169) ) ;
DFF     gate285  (.D(g24169), .CP(CLK), .Q(g90) ) ;
INV     gate286  (.A(II23354), .Z(g24170) ) ;
DFF     gate287  (.D(g24170), .CP(CLK), .Q(g91) ) ;
INV     gate288  (.A(II23357), .Z(g24171) ) ;
DFF     gate289  (.D(g24171), .CP(CLK), .Q(g92) ) ;
INV     gate290  (.A(II23360), .Z(g24172) ) ;
DFF     gate291  (.D(g24172), .CP(CLK), .Q(g99) ) ;
INV     gate292  (.A(II23363), .Z(g24173) ) ;
DFF     gate293  (.D(g24173), .CP(CLK), .Q(g100) ) ;
INV     gate294  (.A(II33070), .Z(g34848) ) ;
DFF     gate295  (.D(g34848), .CP(CLK), .Q(g110) ) ;
INV     gate296  (.A(II33109), .Z(g34879) ) ;
DFF     gate297  (.D(g34879), .CP(CLK), .Q(g112) ) ;
INV     gate298  (.A(II23366), .Z(g24174) ) ;
DFF     gate299  (.D(g24174), .CP(CLK), .Q(g113) ) ;
INV     gate300  (.A(II23369), .Z(g24175) ) ;
DFF     gate301  (.D(g24175), .CP(CLK), .Q(g114) ) ;
INV     gate302  (.A(II23372), .Z(g24176) ) ;
DFF     gate303  (.D(g24176), .CP(CLK), .Q(g115) ) ;
INV     gate304  (.A(II23375), .Z(g24177) ) ;
DFF     gate305  (.D(g24177), .CP(CLK), .Q(g116) ) ;
INV     gate306  (.A(II23378), .Z(g24178) ) ;
DFF     gate307  (.D(g24178), .CP(CLK), .Q(g120) ) ;
INV     gate308  (.A(II23381), .Z(g24179) ) ;
DFF     gate309  (.D(g24179), .CP(CLK), .Q(g124) ) ;
INV     gate310  (.A(II23384), .Z(g24180) ) ;
DFF     gate311  (.D(g24180), .CP(CLK), .Q(g125) ) ;
INV     gate312  (.A(II23387), .Z(g24181) ) ;
DFF     gate313  (.D(g24181), .CP(CLK), .Q(g126) ) ;
INV     gate314  (.A(II23390), .Z(g24182) ) ;
DFF     gate315  (.D(g24182), .CP(CLK), .Q(g127) ) ;
INV     gate316  (.A(II23393), .Z(g24183) ) ;
DFF     gate317  (.D(g24183), .CP(CLK), .Q(g134) ) ;
INV     gate318  (.A(II23396), .Z(g24184) ) ;
DFF     gate319  (.D(g24184), .CP(CLK), .Q(g135) ) ;
INV     gate320  (.A(II23399), .Z(g24185) ) ;
DFF     gate321  (.D(g24185), .CP(CLK), .Q(g44) ) ;
INV     gate322  (.A(II33270), .Z(g34990) ) ;
DFF     gate323  (.D(g34990), .CP(CLK), .Q(g45) ) ;
INV     gate324  (.A(II33273), .Z(g34991) ) ;
DFF     gate325  (.D(g34991), .CP(CLK), .Q(g46) ) ;
INV     gate326  (.A(II33276), .Z(g34992) ) ;
DFF     gate327  (.D(g34992), .CP(CLK), .Q(g47) ) ;
INV     gate328  (.A(II33279), .Z(g34993) ) ;
DFF     gate329  (.D(g34993), .CP(CLK), .Q(g48) ) ;
INV     gate330  (.A(II33282), .Z(g34994) ) ;
DFF     gate331  (.D(g34994), .CP(CLK), .Q(g49) ) ;
INV     gate332  (.A(II33285), .Z(g34995) ) ;
DFF     gate333  (.D(g34995), .CP(CLK), .Q(g50) ) ;
INV     gate334  (.A(II33288), .Z(g34996) ) ;
DFF     gate335  (.D(g34996), .CP(CLK), .Q(g51) ) ;
INV     gate336  (.A(II33291), .Z(g34997) ) ;
DFF     gate337  (.D(g34997), .CP(CLK), .Q(g52) ) ;
INV     gate338  (.A(II23327), .Z(g24161) ) ;
DFF     gate339  (.D(g24161), .CP(CLK), .Q(g53) ) ;
INV     gate340  (.A(II23330), .Z(g24162) ) ;
DFF     gate341  (.D(g24162), .CP(CLK), .Q(g54) ) ;
INV     gate342  (.A(II33300), .Z(g35002) ) ;
DFF     gate343  (.D(g35002), .CP(CLK), .Q(g55) ) ;
INV     gate344  (.A(II23333), .Z(g24163) ) ;
DFF     gate345  (.D(g24163), .CP(CLK), .Q(g56) ) ;
INV     gate346  (.A(II23336), .Z(g24164) ) ;
DFF     gate347  (.D(g24164), .CP(CLK), .Q(g57) ) ;
INV     gate348  (.A(II28585), .Z(g30328) ) ;
DFF     gate349  (.D(g30328), .CP(CLK), .Q(g58) ) ;
INV     gate350  (.A(II33067), .Z(g34847) ) ;
DFF     gate351  (.D(g34847), .CP(CLK), .Q(g63) ) ;
INV     gate352  (.A(II32988), .Z(g34786) ) ;
DFF     gate353  (.D(g34786), .CP(CLK), .Q(g71) ) ;
INV     gate354  (.A(II32881), .Z(g34717) ) ;
DFF     gate355  (.D(g34717), .CP(CLK), .Q(g85) ) ;
INV     gate356  (.A(II33106), .Z(g34878) ) ;
DFF     gate357  (.D(g34878), .CP(CLK), .Q(g93) ) ;
INV     gate358  (.A(II32991), .Z(g34787) ) ;
DFF     gate359  (.D(g34787), .CP(CLK), .Q(g101) ) ;
INV     gate360  (.A(II32884), .Z(g34718) ) ;
DFF     gate361  (.D(g34718), .CP(CLK), .Q(g111) ) ;
INV     gate362  (.A(II32997), .Z(g34789) ) ;
DFF     gate363  (.D(g34789), .CP(CLK), .Q(g43) ) ;
INV     gate364  (.A(II23339), .Z(g24165) ) ;
DFF     gate365  (.D(g24165), .CP(CLK), .Q(g64) ) ;
INV     gate366  (.A(II32985), .Z(g34785) ) ;
DFF     gate367  (.D(g34785), .CP(CLK), .Q(g65) ) ;
INV     gate368  (.A(II18885), .Z(g18093) ) ;
DFF     gate369  (.D(g18093), .CP(CLK), .Q(g70) ) ;
OR2     gate370  (.A(g30005), .B(g24330), .Z(g30458) ) ;
DFF     gate371  (.D(g30458), .CP(CLK), .Q(g4507) ) ;
OR2     gate372  (.A(g34171), .B(g24300), .Z(g34253) ) ;
DFF     gate373  (.D(g34253), .CP(CLK), .Q(g4459) ) ;
OR2     gate374  (.A(g26308), .B(g24332), .Z(g26970) ) ;
DFF     gate375  (.D(g26970), .CP(CLK), .Q(g4369) ) ;
OR2     gate376  (.A(g34173), .B(g24303), .Z(g34256) ) ;
DFF     gate377  (.D(g34256), .CP(CLK), .Q(g4473) ) ;
OR2     gate378  (.A(g34116), .B(g24301), .Z(g34254) ) ;
DFF     gate379  (.D(g34254), .CP(CLK), .Q(g4462) ) ;
OR2     gate380  (.A(g26313), .B(g24329), .Z(g26969) ) ;
DFF     gate381  (.D(g26969), .CP(CLK), .Q(g4581) ) ;
OR2     gate382  (.A(g34120), .B(g24302), .Z(g34255) ) ;
DFF     gate383  (.D(g34255), .CP(CLK), .Q(g4467) ) ;
INV     gate384  (.A(II13802), .Z(g10384) ) ;
DFF     gate385  (.D(g10384), .CP(CLK), .Q(g4474) ) ;
OR2     gate386  (.A(g26258), .B(g24304), .Z(g26960) ) ;
DFF     gate387  (.D(g26960), .CP(CLK), .Q(g4477) ) ;
OR2     gate388  (.A(g31242), .B(g24305), .Z(g31896) ) ;
DFF     gate389  (.D(g31896), .CP(CLK), .Q(g4480) ) ;
OR2     gate390  (.A(g32168), .B(g24309), .Z(g33036) ) ;
DFF     gate391  (.D(g33036), .CP(CLK), .Q(g4495) ) ;
OR2     gate392  (.A(g32177), .B(g24310), .Z(g33037) ) ;
DFF     gate393  (.D(g33037), .CP(CLK), .Q(g4498) ) ;
OR2     gate394  (.A(g32184), .B(g24311), .Z(g33038) ) ;
DFF     gate395  (.D(g33038), .CP(CLK), .Q(g4501) ) ;
OR2     gate396  (.A(g32187), .B(g24312), .Z(g33039) ) ;
DFF     gate397  (.D(g33039), .CP(CLK), .Q(g4504) ) ;
OR2     gate398  (.A(g32164), .B(g24313), .Z(g33040) ) ;
DFF     gate399  (.D(g33040), .CP(CLK), .Q(g4512) ) ;
OR2     gate400  (.A(g26325), .B(g24333), .Z(g26971) ) ;
DFF     gate401  (.D(g26971), .CP(CLK), .Q(g4521) ) ;
OR2     gate402  (.A(g27369), .B(g24315), .Z(g28082) ) ;
DFF     gate403  (.D(g28082), .CP(CLK), .Q(g4527) ) ;
OR2     gate404  (.A(g26259), .B(g24316), .Z(g26964) ) ;
DFF     gate405  (.D(g26964), .CP(CLK), .Q(g4515) ) ;
OR2     gate406  (.A(g33237), .B(g24314), .Z(g33616) ) ;
DFF     gate407  (.D(g33616), .CP(CLK), .Q(g4519) ) ;
INV     gate408  (.A(II11740), .Z(g6972) ) ;
DFF     gate409  (.D(g6972), .CP(CLK), .Q(g4520) ) ;
DFF     gate410  (.D(g4520), .CP(CLK), .Q(g4483) ) ;
OR2     gate411  (.A(g26280), .B(g24306), .Z(g26961) ) ;
DFF     gate412  (.D(g26961), .CP(CLK), .Q(g4486) ) ;
OR2     gate413  (.A(g26295), .B(g24307), .Z(g26962) ) ;
DFF     gate414  (.D(g26962), .CP(CLK), .Q(g4489) ) ;
OR2     gate415  (.A(g26306), .B(g24308), .Z(g26963) ) ;
DFF     gate416  (.D(g26963), .CP(CLK), .Q(g4492) ) ;
OR2     gate417  (.A(g33807), .B(g24331), .Z(g34024) ) ;
DFF     gate418  (.D(g34024), .CP(CLK), .Q(g4537) ) ;
DFF     gate419  (.D(g4537), .CP(CLK), .Q(g4423) ) ;
OR2     gate420  (.A(g31237), .B(g24322), .Z(g31897) ) ;
DFF     gate421  (.D(g31897), .CP(CLK), .Q(g4540) ) ;
OR2     gate422  (.A(g32193), .B(g24324), .Z(g33042) ) ;
DFF     gate423  (.D(g33042), .CP(CLK), .Q(g4543) ) ;
OR2     gate424  (.A(g32195), .B(g24325), .Z(g33043) ) ;
DFF     gate425  (.D(g33043), .CP(CLK), .Q(g4567) ) ;
OR2     gate426  (.A(g32206), .B(g24328), .Z(g33045) ) ;
DFF     gate427  (.D(g33045), .CP(CLK), .Q(g4546) ) ;
OR2     gate428  (.A(g32189), .B(g24323), .Z(g33041) ) ;
DFF     gate429  (.D(g33041), .CP(CLK), .Q(g4549) ) ;
OR2     gate430  (.A(g32199), .B(g24327), .Z(g33044) ) ;
DFF     gate431  (.D(g33044), .CP(CLK), .Q(g4552) ) ;
OR2     gate432  (.A(g33263), .B(g24326), .Z(g33617) ) ;
DFF     gate433  (.D(g33617), .CP(CLK), .Q(g4570) ) ;
INV     gate434  (.A(II11746), .Z(g6974) ) ;
DFF     gate435  (.D(g6974), .CP(CLK), .Q(g4571) ) ;
DFF     gate436  (.D(g4571), .CP(CLK), .Q(g4555) ) ;
OR2     gate437  (.A(g26345), .B(g24318), .Z(g26966) ) ;
DFF     gate438  (.D(g26966), .CP(CLK), .Q(g4558) ) ;
OR2     gate439  (.A(g26307), .B(g24321), .Z(g26968) ) ;
DFF     gate440  (.D(g26968), .CP(CLK), .Q(g4561) ) ;
OR2     gate441  (.A(g26350), .B(g24319), .Z(g26967) ) ;
DFF     gate442  (.D(g26967), .CP(CLK), .Q(g4564) ) ;
OR2     gate443  (.A(g33796), .B(g24320), .Z(g34023) ) ;
DFF     gate444  (.D(g34023), .CP(CLK), .Q(g4534) ) ;
OR2     gate445  (.A(g26336), .B(g24317), .Z(g26965) ) ;
DFF     gate446  (.D(g26965), .CP(CLK), .Q(g4420) ) ;
OR2     gate447  (.A(g26486), .B(g24291), .Z(g26953) ) ;
DFF     gate448  (.D(g26953), .CP(CLK), .Q(g4438) ) ;
OR2     gate449  (.A(g26391), .B(g24293), .Z(g26955) ) ;
DFF     gate450  (.D(g26955), .CP(CLK), .Q(g4449) ) ;
DFF     gate451  (.D(g4449), .CP(CLK), .Q(g4443) ) ;
OR2     gate452  (.A(g26380), .B(g24292), .Z(g26954) ) ;
DFF     gate453  (.D(g26954), .CP(CLK), .Q(g4446) ) ;
DFF     gate454  (.D(g4446), .CP(CLK), .Q(g4452) ) ;
OR2     gate455  (.A(g26487), .B(g24294), .Z(g26956) ) ;
DFF     gate456  (.D(g26956), .CP(CLK), .Q(g4434) ) ;
OR2     gate457  (.A(g26517), .B(g24295), .Z(g26957) ) ;
DFF     gate458  (.D(g26957), .CP(CLK), .Q(g4430) ) ;
OR2     gate459  (.A(g26360), .B(g24290), .Z(g26952) ) ;
DFF     gate460  (.D(g26952), .CP(CLK), .Q(g4427) ) ;
OR2     gate461  (.A(g26390), .B(g24289), .Z(g26951) ) ;
DFF     gate462  (.D(g26951), .CP(CLK), .Q(g4375) ) ;
OR2     gate463  (.A(g26389), .B(g24284), .Z(g26946) ) ;
DFF     gate464  (.D(g26946), .CP(CLK), .Q(g4414) ) ;
DFF     gate465  (.D(g4414), .CP(CLK), .Q(g4411) ) ;
OR2     gate466  (.A(g26379), .B(g24283), .Z(g26945) ) ;
DFF     gate467  (.D(g26945), .CP(CLK), .Q(g4408) ) ;
DFF     gate468  (.D(g4408), .CP(CLK), .Q(g4405) ) ;
OR2     gate469  (.A(g26399), .B(g24286), .Z(g26948) ) ;
DFF     gate470  (.D(g26948), .CP(CLK), .Q(g4401) ) ;
OR2     gate471  (.A(g26356), .B(g24287), .Z(g26949) ) ;
DFF     gate472  (.D(g26949), .CP(CLK), .Q(g4388) ) ;
OR2     gate473  (.A(g26394), .B(g24285), .Z(g26947) ) ;
DFF     gate474  (.D(g26947), .CP(CLK), .Q(g4382) ) ;
OR2     gate475  (.A(g31505), .B(g24296), .Z(g31895) ) ;
DFF     gate476  (.D(g31895), .CP(CLK), .Q(g4417) ) ;
OR2     gate477  (.A(g26357), .B(g24288), .Z(g26950) ) ;
DFF     gate478  (.D(g26950), .CP(CLK), .Q(g4392) ) ;
INV     gate479  (.A(II24839), .Z(g25692) ) ;
DFF     gate480  (.D(g25692), .CP(CLK), .Q(g4456) ) ;
OR2     gate481  (.A(g26381), .B(g24299), .Z(g26959) ) ;
DFF     gate482  (.D(g26959), .CP(CLK), .Q(g4455) ) ;
OR2     gate483  (.A(g26395), .B(g24297), .Z(g26958) ) ;
DFF     gate484  (.D(g26958), .CP(CLK), .Q(g1) ) ;
OR2     gate485  (.A(g23397), .B(g18656), .Z(g24281) ) ;
DFF     gate486  (.D(g24281), .CP(CLK), .Q(g4304) ) ;
DFF     gate487  (.D(g4304), .CP(CLK), .Q(g4308) ) ;
OR2     gate488  (.A(g23407), .B(g18657), .Z(g24282) ) ;
DFF     gate489  (.D(g24282), .CP(CLK), .Q(g2932) ) ;
OR2     gate490  (.A(g33927), .B(g18672), .Z(g34025) ) ;
DFF     gate491  (.D(g34025), .CP(CLK), .Q(g4639) ) ;
OR2     gate492  (.A(g34301), .B(g18677), .Z(g34460) ) ;
DFF     gate493  (.D(g34460), .CP(CLK), .Q(g4621) ) ;
OR2     gate494  (.A(g34394), .B(g18670), .Z(g34457) ) ;
DFF     gate495  (.D(g34457), .CP(CLK), .Q(g4628) ) ;
OR2     gate496  (.A(g34396), .B(g18671), .Z(g34458) ) ;
DFF     gate497  (.D(g34458), .CP(CLK), .Q(g4633) ) ;
OR2     gate498  (.A(g34066), .B(g18679), .Z(g34259) ) ;
DFF     gate499  (.D(g34259), .CP(CLK), .Q(g4643) ) ;
OR2     gate500  (.A(g34415), .B(g18673), .Z(g34459) ) ;
DFF     gate501  (.D(g34459), .CP(CLK), .Q(g4340) ) ;
OR2     gate502  (.A(g34226), .B(g18674), .Z(g34257) ) ;
DFF     gate503  (.D(g34257), .CP(CLK), .Q(g4349) ) ;
OR2     gate504  (.A(g34211), .B(g18675), .Z(g34258) ) ;
DFF     gate505  (.D(g34258), .CP(CLK), .Q(g4358) ) ;
OR2     gate506  (.A(g23991), .B(g18676), .Z(g24334) ) ;
DFF     gate507  (.D(g24334), .CP(CLK), .Q(g66) ) ;
OR2     gate508  (.A(g22165), .B(g18678), .Z(g24335) ) ;
DFF     gate509  (.D(g24335), .CP(CLK), .Q(g4531) ) ;
OR2     gate510  (.A(g34279), .B(g18662), .Z(g34449) ) ;
DFF     gate511  (.D(g34449), .CP(CLK), .Q(g4311) ) ;
OR2     gate512  (.A(g34281), .B(g18663), .Z(g34450) ) ;
DFF     gate513  (.D(g34450), .CP(CLK), .Q(g4322) ) ;
OR2     gate514  (.A(g34284), .B(g18668), .Z(g34455) ) ;
DFF     gate515  (.D(g34455), .CP(CLK), .Q(g4332) ) ;
OR2     gate516  (.A(g34393), .B(g18664), .Z(g34451) ) ;
DFF     gate517  (.D(g34451), .CP(CLK), .Q(g4584) ) ;
OR2     gate518  (.A(g34401), .B(g18665), .Z(g34452) ) ;
DFF     gate519  (.D(g34452), .CP(CLK), .Q(g4593) ) ;
OR2     gate520  (.A(g34410), .B(g18666), .Z(g34453) ) ;
DFF     gate521  (.D(g34453), .CP(CLK), .Q(g4601) ) ;
OR2     gate522  (.A(g34414), .B(g18667), .Z(g34454) ) ;
DFF     gate523  (.D(g34454), .CP(CLK), .Q(g4608) ) ;
OR2     gate524  (.A(g34395), .B(g18669), .Z(g34456) ) ;
DFF     gate525  (.D(g34456), .CP(CLK), .Q(g4616) ) ;
OR2     gate526  (.A(g26130), .B(g18658), .Z(g26944) ) ;
DFF     gate527  (.D(g26944), .CP(CLK), .Q(g4366) ) ;
OR2     gate528  (.A(g34876), .B(g18659), .Z(g34882) ) ;
DFF     gate529  (.D(g34882), .CP(CLK), .Q(g4372) ) ;
OR2     gate530  (.A(g34117), .B(g18711), .Z(g34265) ) ;
DFF     gate531  (.D(g34265), .CP(CLK), .Q(g4836) ) ;
OR2     gate532  (.A(g33719), .B(g18713), .Z(g34034) ) ;
DFF     gate533  (.D(g34034), .CP(CLK), .Q(g4864) ) ;
OR2     gate534  (.A(g33721), .B(g18714), .Z(g34035) ) ;
DFF     gate535  (.D(g34035), .CP(CLK), .Q(g4871) ) ;
OR2     gate536  (.A(g33722), .B(g18715), .Z(g34036) ) ;
DFF     gate537  (.D(g34036), .CP(CLK), .Q(g4878) ) ;
OR2     gate538  (.A(g34337), .B(g18716), .Z(g34466) ) ;
DFF     gate539  (.D(g34466), .CP(CLK), .Q(g4843) ) ;
OR2     gate540  (.A(g34295), .B(g18712), .Z(g34465) ) ;
DFF     gate541  (.D(g34465), .CP(CLK), .Q(g4849) ) ;
OR2     gate542  (.A(g34341), .B(g18717), .Z(g34467) ) ;
DFF     gate543  (.D(g34467), .CP(CLK), .Q(g4854) ) ;
OR2     gate544  (.A(g34342), .B(g18718), .Z(g34468) ) ;
DFF     gate545  (.D(g34468), .CP(CLK), .Q(g4859) ) ;
OR2     gate546  (.A(g34484), .B(g18721), .Z(g34638) ) ;
DFF     gate547  (.D(g34638), .CP(CLK), .Q(g4917) ) ;
OR2     gate548  (.A(g34486), .B(g18722), .Z(g34639) ) ;
DFF     gate549  (.D(g34639), .CP(CLK), .Q(g4922) ) ;
OR2     gate550  (.A(g34487), .B(g18723), .Z(g34640) ) ;
DFF     gate551  (.D(g34640), .CP(CLK), .Q(g4907) ) ;
OR2     gate552  (.A(g34479), .B(g18724), .Z(g34641) ) ;
DFF     gate553  (.D(g34641), .CP(CLK), .Q(g4912) ) ;
OR2     gate554  (.A(g34482), .B(g18725), .Z(g34642) ) ;
DFF     gate555  (.D(g34642), .CP(CLK), .Q(g4927) ) ;
INV     gate556  (.A(II21483), .Z(g21904) ) ;
DFF     gate557  (.D(g21904), .CP(CLK), .Q(g4931) ) ;
INV     gate558  (.A(II21486), .Z(g21905) ) ;
DFF     gate559  (.D(g21905), .CP(CLK), .Q(g4932) ) ;
OR2     gate560  (.A(g28442), .B(g18741), .Z(g29279) ) ;
DFF     gate561  (.D(g29279), .CP(CLK), .Q(g4572) ) ;
OR2     gate562  (.A(g28626), .B(g18740), .Z(g29278) ) ;
DFF     gate563  (.D(g29278), .CP(CLK), .Q(g4578) ) ;
OR2     gate564  (.A(g24638), .B(g18738), .Z(g25694) ) ;
DFF     gate565  (.D(g25694), .CP(CLK), .Q(g4999) ) ;
DFF     gate566  (.D(g4999), .CP(CLK), .Q(g5002) ) ;
DFF     gate567  (.D(g5002), .CP(CLK), .Q(g5005) ) ;
DFF     gate568  (.D(g5005), .CP(CLK), .Q(g5008) ) ;
OR2     gate569  (.A(g33829), .B(g18739), .Z(g34041) ) ;
DFF     gate570  (.D(g34041), .CP(CLK), .Q(g4983) ) ;
OR2     gate571  (.A(g33731), .B(g18735), .Z(g34038) ) ;
DFF     gate572  (.D(g34038), .CP(CLK), .Q(g4991) ) ;
OR2     gate573  (.A(g33743), .B(g18736), .Z(g34039) ) ;
DFF     gate574  (.D(g34039), .CP(CLK), .Q(g4966) ) ;
OR2     gate575  (.A(g33803), .B(g18734), .Z(g34037) ) ;
DFF     gate576  (.D(g34037), .CP(CLK), .Q(g4975) ) ;
OR2     gate577  (.A(g33818), .B(g18737), .Z(g34040) ) ;
DFF     gate578  (.D(g34040), .CP(CLK), .Q(g4899) ) ;
OR2     gate579  (.A(g27255), .B(g18720), .Z(g28087) ) ;
DFF     gate580  (.D(g28087), .CP(CLK), .Q(g4894) ) ;
OR2     gate581  (.A(g34076), .B(g18719), .Z(g34266) ) ;
DFF     gate582  (.D(g34266), .CP(CLK), .Q(g4888) ) ;
OR2     gate583  (.A(g27264), .B(g18729), .Z(g28088) ) ;
DFF     gate584  (.D(g28088), .CP(CLK), .Q(g4939) ) ;
OR2     gate585  (.A(g34079), .B(g18728), .Z(g34267) ) ;
DFF     gate586  (.D(g34267), .CP(CLK), .Q(g4933) ) ;
OR2     gate587  (.A(g27269), .B(g18731), .Z(g28089) ) ;
DFF     gate588  (.D(g28089), .CP(CLK), .Q(g4950) ) ;
OR2     gate589  (.A(g34082), .B(g18730), .Z(g34268) ) ;
DFF     gate590  (.D(g34268), .CP(CLK), .Q(g4944) ) ;
OR2     gate591  (.A(g27275), .B(g18733), .Z(g28090) ) ;
DFF     gate592  (.D(g28090), .CP(CLK), .Q(g4961) ) ;
OR2     gate593  (.A(g34083), .B(g18732), .Z(g34269) ) ;
DFF     gate594  (.D(g34269), .CP(CLK), .Q(g4955) ) ;
OR2     gate595  (.A(g34113), .B(g18680), .Z(g34260) ) ;
DFF     gate596  (.D(g34260), .CP(CLK), .Q(g4646) ) ;
OR2     gate597  (.A(g33715), .B(g18682), .Z(g34026) ) ;
DFF     gate598  (.D(g34026), .CP(CLK), .Q(g4674) ) ;
OR2     gate599  (.A(g33718), .B(g18683), .Z(g34027) ) ;
DFF     gate600  (.D(g34027), .CP(CLK), .Q(g4681) ) ;
OR2     gate601  (.A(g33720), .B(g18684), .Z(g34028) ) ;
DFF     gate602  (.D(g34028), .CP(CLK), .Q(g4688) ) ;
OR2     gate603  (.A(g34334), .B(g18685), .Z(g34462) ) ;
DFF     gate604  (.D(g34462), .CP(CLK), .Q(g4653) ) ;
OR2     gate605  (.A(g34291), .B(g18681), .Z(g34461) ) ;
DFF     gate606  (.D(g34461), .CP(CLK), .Q(g4659) ) ;
OR2     gate607  (.A(g34338), .B(g18686), .Z(g34463) ) ;
DFF     gate608  (.D(g34463), .CP(CLK), .Q(g4664) ) ;
OR2     gate609  (.A(g34340), .B(g18687), .Z(g34464) ) ;
DFF     gate610  (.D(g34464), .CP(CLK), .Q(g4669) ) ;
OR2     gate611  (.A(g34481), .B(g18690), .Z(g34633) ) ;
DFF     gate612  (.D(g34633), .CP(CLK), .Q(g4727) ) ;
OR2     gate613  (.A(g34483), .B(g18691), .Z(g34634) ) ;
DFF     gate614  (.D(g34634), .CP(CLK), .Q(g4732) ) ;
OR2     gate615  (.A(g34485), .B(g18692), .Z(g34635) ) ;
DFF     gate616  (.D(g34635), .CP(CLK), .Q(g4717) ) ;
OR2     gate617  (.A(g34476), .B(g18693), .Z(g34636) ) ;
DFF     gate618  (.D(g34636), .CP(CLK), .Q(g4722) ) ;
OR2     gate619  (.A(g34478), .B(g18694), .Z(g34637) ) ;
DFF     gate620  (.D(g34637), .CP(CLK), .Q(g4737) ) ;
INV     gate621  (.A(II21477), .Z(g21902) ) ;
DFF     gate622  (.D(g21902), .CP(CLK), .Q(g4741) ) ;
INV     gate623  (.A(II21480), .Z(g21903) ) ;
DFF     gate624  (.D(g21903), .CP(CLK), .Q(g4742) ) ;
OR2     gate625  (.A(g28440), .B(g18710), .Z(g29277) ) ;
DFF     gate626  (.D(g29277), .CP(CLK), .Q(g59) ) ;
OR2     gate627  (.A(g28616), .B(g18709), .Z(g29276) ) ;
DFF     gate628  (.D(g29276), .CP(CLK), .Q(g4575) ) ;
OR2     gate629  (.A(g24627), .B(g18707), .Z(g25693) ) ;
DFF     gate630  (.D(g25693), .CP(CLK), .Q(g4809) ) ;
DFF     gate631  (.D(g4809), .CP(CLK), .Q(g4812) ) ;
DFF     gate632  (.D(g4812), .CP(CLK), .Q(g4815) ) ;
DFF     gate633  (.D(g4815), .CP(CLK), .Q(g4818) ) ;
OR2     gate634  (.A(g33821), .B(g18708), .Z(g34033) ) ;
DFF     gate635  (.D(g34033), .CP(CLK), .Q(g4793) ) ;
OR2     gate636  (.A(g33727), .B(g18704), .Z(g34030) ) ;
DFF     gate637  (.D(g34030), .CP(CLK), .Q(g4801) ) ;
OR2     gate638  (.A(g33735), .B(g18705), .Z(g34031) ) ;
DFF     gate639  (.D(g34031), .CP(CLK), .Q(g4776) ) ;
OR2     gate640  (.A(g33798), .B(g18703), .Z(g34029) ) ;
DFF     gate641  (.D(g34029), .CP(CLK), .Q(g4785) ) ;
OR2     gate642  (.A(g33816), .B(g18706), .Z(g34032) ) ;
DFF     gate643  (.D(g34032), .CP(CLK), .Q(g4709) ) ;
OR2     gate644  (.A(g27249), .B(g18689), .Z(g28083) ) ;
DFF     gate645  (.D(g28083), .CP(CLK), .Q(g4704) ) ;
OR2     gate646  (.A(g34074), .B(g18688), .Z(g34261) ) ;
DFF     gate647  (.D(g34261), .CP(CLK), .Q(g4698) ) ;
OR2     gate648  (.A(g27254), .B(g18698), .Z(g28084) ) ;
DFF     gate649  (.D(g28084), .CP(CLK), .Q(g4749) ) ;
OR2     gate650  (.A(g34075), .B(g18697), .Z(g34262) ) ;
DFF     gate651  (.D(g34262), .CP(CLK), .Q(g4743) ) ;
OR2     gate652  (.A(g27263), .B(g18700), .Z(g28085) ) ;
DFF     gate653  (.D(g28085), .CP(CLK), .Q(g4760) ) ;
OR2     gate654  (.A(g34078), .B(g18699), .Z(g34263) ) ;
DFF     gate655  (.D(g34263), .CP(CLK), .Q(g4754) ) ;
OR2     gate656  (.A(g27268), .B(g18702), .Z(g28086) ) ;
DFF     gate657  (.D(g28086), .CP(CLK), .Q(g4771) ) ;
OR2     gate658  (.A(g34081), .B(g18701), .Z(g34264) ) ;
DFF     gate659  (.D(g34264), .CP(CLK), .Q(g4765) ) ;
OR2     gate660  (.A(g24012), .B(g18753), .Z(g24336) ) ;
DFF     gate661  (.D(g24336), .CP(CLK), .Q(g5313) ) ;
DFF     gate662  (.D(g5313), .CP(CLK), .Q(g5290) ) ;
DFF     gate663  (.D(g5290), .CP(CLK), .Q(g5320) ) ;
DFF     gate664  (.D(g5320), .CP(CLK), .Q(g5276) ) ;
DFF     gate665  (.D(g5276), .CP(CLK), .Q(g5283) ) ;
DFF     gate666  (.D(g5283), .CP(CLK), .Q(g5308) ) ;
DFF     gate667  (.D(g5308), .CP(CLK), .Q(g5327) ) ;
DFF     gate668  (.D(g5327), .CP(CLK), .Q(g5331) ) ;
DFF     gate669  (.D(g5331), .CP(CLK), .Q(g5335) ) ;
DFF     gate670  (.D(g5335), .CP(CLK), .Q(g5339) ) ;
OR2     gate671  (.A(g23540), .B(g18754), .Z(g24337) ) ;
DFF     gate672  (.D(g24337), .CP(CLK), .Q(g5343) ) ;
OR2     gate673  (.A(g23658), .B(g18755), .Z(g24338) ) ;
DFF     gate674  (.D(g24338), .CP(CLK), .Q(g5348) ) ;
OR2     gate675  (.A(g23690), .B(g18756), .Z(g24339) ) ;
DFF     gate676  (.D(g24339), .CP(CLK), .Q(g5352) ) ;
OR2     gate677  (.A(g33353), .B(g18757), .Z(g33618) ) ;
DFF     gate678  (.D(g33618), .CP(CLK), .Q(g5357) ) ;
OR2     gate679  (.A(g33359), .B(g18758), .Z(g33619) ) ;
DFF     gate680  (.D(g33619), .CP(CLK), .Q(g5297) ) ;
OR2     gate681  (.A(g25040), .B(g21919), .Z(g25700) ) ;
DFF     gate682  (.D(g25700), .CP(CLK), .Q(g5101) ) ;
DFF     gate683  (.D(g5101), .CP(CLK), .Q(g5109) ) ;
OR2     gate684  (.A(g25068), .B(g21921), .Z(g25702) ) ;
DFF     gate685  (.D(g25702), .CP(CLK), .Q(g5062) ) ;
OR2     gate686  (.A(g25054), .B(g21920), .Z(g25701) ) ;
DFF     gate687  (.D(g25701), .CP(CLK), .Q(g5105) ) ;
DFF     gate688  (.D(g5105), .CP(CLK), .Q(g5112) ) ;
OR2     gate689  (.A(g25087), .B(g21922), .Z(g25703) ) ;
DFF     gate690  (.D(g25703), .CP(CLK), .Q(g5022) ) ;
OR2     gate691  (.A(g31707), .B(g21906), .Z(g31898) ) ;
DFF     gate692  (.D(g31898), .CP(CLK), .Q(g5016) ) ;
OR2     gate693  (.A(g31744), .B(g21910), .Z(g31902) ) ;
DFF     gate694  (.D(g31902), .CP(CLK), .Q(g5029) ) ;
OR2     gate695  (.A(g31780), .B(g21923), .Z(g31904) ) ;
DFF     gate696  (.D(g31904), .CP(CLK), .Q(g5033) ) ;
OR2     gate697  (.A(g31470), .B(g21907), .Z(g31899) ) ;
DFF     gate698  (.D(g31899), .CP(CLK), .Q(g5037) ) ;
OR2     gate699  (.A(g31484), .B(g21908), .Z(g31900) ) ;
DFF     gate700  (.D(g31900), .CP(CLK), .Q(g5041) ) ;
OR2     gate701  (.A(g31516), .B(g21909), .Z(g31901) ) ;
DFF     gate702  (.D(g31901), .CP(CLK), .Q(g5046) ) ;
OR2     gate703  (.A(g31374), .B(g21911), .Z(g31903) ) ;
DFF     gate704  (.D(g31903), .CP(CLK), .Q(g5052) ) ;
OR2     gate705  (.A(g32308), .B(g21912), .Z(g33046) ) ;
DFF     gate706  (.D(g33046), .CP(CLK), .Q(g5057) ) ;
OR2     gate707  (.A(g27666), .B(g21924), .Z(g28092) ) ;
DFF     gate708  (.D(g28092), .CP(CLK), .Q(g5069) ) ;
OR2     gate709  (.A(g27665), .B(g21913), .Z(g28091) ) ;
DFF     gate710  (.D(g28091), .CP(CLK), .Q(g5073) ) ;
OR2     gate711  (.A(g25173), .B(g21925), .Z(g25704) ) ;
DFF     gate712  (.D(g25704), .CP(CLK), .Q(g5077) ) ;
OR2     gate713  (.A(g24998), .B(g21914), .Z(g25695) ) ;
DFF     gate714  (.D(g25695), .CP(CLK), .Q(g5080) ) ;
OR2     gate715  (.A(g25012), .B(g21915), .Z(g25696) ) ;
DFF     gate716  (.D(g25696), .CP(CLK), .Q(g5084) ) ;
OR2     gate717  (.A(g25086), .B(g21916), .Z(g25697) ) ;
DFF     gate718  (.D(g25697), .CP(CLK), .Q(g5092) ) ;
OR2     gate719  (.A(g25104), .B(g21917), .Z(g25698) ) ;
DFF     gate720  (.D(g25698), .CP(CLK), .Q(g5097) ) ;
OR2     gate721  (.A(g25125), .B(g21918), .Z(g25699) ) ;
DFF     gate722  (.D(g25699), .CP(CLK), .Q(g86) ) ;
OR2     gate723  (.A(g29314), .B(g21926), .Z(g30459) ) ;
DFF     gate724  (.D(g30459), .CP(CLK), .Q(g5164) ) ;
OR2     gate725  (.A(g31944), .B(g21927), .Z(g33047) ) ;
DFF     gate726  (.D(g33047), .CP(CLK), .Q(g5170) ) ;
OR2     gate727  (.A(g31960), .B(g21928), .Z(g33048) ) ;
DFF     gate728  (.D(g33048), .CP(CLK), .Q(g5176) ) ;
OR2     gate729  (.A(g31966), .B(g21929), .Z(g33049) ) ;
DFF     gate730  (.D(g33049), .CP(CLK), .Q(g5180) ) ;
OR2     gate731  (.A(g31974), .B(g21930), .Z(g33050) ) ;
DFF     gate732  (.D(g33050), .CP(CLK), .Q(g5188) ) ;
OR2     gate733  (.A(g30207), .B(g21931), .Z(g30460) ) ;
DFF     gate734  (.D(g30460), .CP(CLK), .Q(g5196) ) ;
OR2     gate735  (.A(g30152), .B(g21935), .Z(g30464) ) ;
DFF     gate736  (.D(g30464), .CP(CLK), .Q(g5224) ) ;
OR2     gate737  (.A(g30238), .B(g21939), .Z(g30468) ) ;
DFF     gate738  (.D(g30468), .CP(CLK), .Q(g5240) ) ;
OR2     gate739  (.A(g30186), .B(g21943), .Z(g30472) ) ;
DFF     gate740  (.D(g30472), .CP(CLK), .Q(g5256) ) ;
OR2     gate741  (.A(g30229), .B(g21947), .Z(g30476) ) ;
DFF     gate742  (.D(g30476), .CP(CLK), .Q(g5204) ) ;
OR2     gate743  (.A(g30219), .B(g21932), .Z(g30461) ) ;
DFF     gate744  (.D(g30461), .CP(CLK), .Q(g5200) ) ;
OR2     gate745  (.A(g30164), .B(g21936), .Z(g30465) ) ;
DFF     gate746  (.D(g30465), .CP(CLK), .Q(g5228) ) ;
OR2     gate747  (.A(g30153), .B(g21940), .Z(g30469) ) ;
DFF     gate748  (.D(g30469), .CP(CLK), .Q(g5244) ) ;
OR2     gate749  (.A(g30196), .B(g21944), .Z(g30473) ) ;
DFF     gate750  (.D(g30473), .CP(CLK), .Q(g5260) ) ;
OR2     gate751  (.A(g30239), .B(g21948), .Z(g30477) ) ;
DFF     gate752  (.D(g30477), .CP(CLK), .Q(g5212) ) ;
OR2     gate753  (.A(g30228), .B(g21933), .Z(g30462) ) ;
DFF     gate754  (.D(g30462), .CP(CLK), .Q(g5208) ) ;
OR2     gate755  (.A(g30174), .B(g21937), .Z(g30466) ) ;
DFF     gate756  (.D(g30466), .CP(CLK), .Q(g5232) ) ;
OR2     gate757  (.A(g30165), .B(g21941), .Z(g30470) ) ;
DFF     gate758  (.D(g30470), .CP(CLK), .Q(g5248) ) ;
OR2     gate759  (.A(g30208), .B(g21945), .Z(g30474) ) ;
DFF     gate760  (.D(g30474), .CP(CLK), .Q(g5264) ) ;
OR2     gate761  (.A(g30248), .B(g21949), .Z(g30478) ) ;
DFF     gate762  (.D(g30478), .CP(CLK), .Q(g5220) ) ;
OR2     gate763  (.A(g30140), .B(g21934), .Z(g30463) ) ;
DFF     gate764  (.D(g30463), .CP(CLK), .Q(g5216) ) ;
OR2     gate765  (.A(g30185), .B(g21938), .Z(g30467) ) ;
DFF     gate766  (.D(g30467), .CP(CLK), .Q(g5236) ) ;
OR2     gate767  (.A(g30175), .B(g21942), .Z(g30471) ) ;
DFF     gate768  (.D(g30471), .CP(CLK), .Q(g5252) ) ;
OR2     gate769  (.A(g30220), .B(g21946), .Z(g30475) ) ;
DFF     gate770  (.D(g30475), .CP(CLK), .Q(g5268) ) ;
OR2     gate771  (.A(g29320), .B(g21950), .Z(g30479) ) ;
DFF     gate772  (.D(g30479), .CP(CLK), .Q(g5272) ) ;
OR2     gate773  (.A(g27981), .B(g21951), .Z(g28093) ) ;
DFF     gate774  (.D(g28093), .CP(CLK), .Q(g128) ) ;
OR2     gate775  (.A(g28639), .B(g18750), .Z(g29285) ) ;
DFF     gate776  (.D(g29285), .CP(CLK), .Q(g5156) ) ;
OR2     gate777  (.A(g25526), .B(g18751), .Z(g25708) ) ;
DFF     gate778  (.D(g25708), .CP(CLK), .Q(g5120) ) ;
OR2     gate779  (.A(g28530), .B(g18742), .Z(g29280) ) ;
DFF     gate780  (.D(g29280), .CP(CLK), .Q(g5115) ) ;
OR2     gate781  (.A(g28541), .B(g18743), .Z(g29281) ) ;
DFF     gate782  (.D(g29281), .CP(CLK), .Q(g5124) ) ;
OR2     gate783  (.A(g25069), .B(g18744), .Z(g25705) ) ;
DFF     gate784  (.D(g25705), .CP(CLK), .Q(g5128) ) ;
OR2     gate785  (.A(g28617), .B(g18745), .Z(g29282) ) ;
DFF     gate786  (.D(g29282), .CP(CLK), .Q(g5134) ) ;
OR2     gate787  (.A(g28627), .B(g18746), .Z(g29283) ) ;
DFF     gate788  (.D(g29283), .CP(CLK), .Q(g5138) ) ;
OR2     gate789  (.A(g28554), .B(g18747), .Z(g29284) ) ;
DFF     gate790  (.D(g29284), .CP(CLK), .Q(g5142) ) ;
OR2     gate791  (.A(g25030), .B(g18748), .Z(g25706) ) ;
DFF     gate792  (.D(g25706), .CP(CLK), .Q(g5148) ) ;
OR2     gate793  (.A(g25041), .B(g18749), .Z(g25707) ) ;
DFF     gate794  (.D(g25707), .CP(CLK), .Q(g5152) ) ;
OR2     gate795  (.A(g34554), .B(g18752), .Z(g34643) ) ;
DFF     gate796  (.D(g34643), .CP(CLK), .Q(g5160) ) ;
OR2     gate797  (.A(g24016), .B(g18770), .Z(g24340) ) ;
DFF     gate798  (.D(g24340), .CP(CLK), .Q(g5659) ) ;
DFF     gate799  (.D(g5659), .CP(CLK), .Q(g5637) ) ;
DFF     gate800  (.D(g5637), .CP(CLK), .Q(g5666) ) ;
DFF     gate801  (.D(g5666), .CP(CLK), .Q(g5623) ) ;
DFF     gate802  (.D(g5623), .CP(CLK), .Q(g5630) ) ;
DFF     gate803  (.D(g5630), .CP(CLK), .Q(g5654) ) ;
DFF     gate804  (.D(g5654), .CP(CLK), .Q(g5673) ) ;
DFF     gate805  (.D(g5673), .CP(CLK), .Q(g5677) ) ;
DFF     gate806  (.D(g5677), .CP(CLK), .Q(g5681) ) ;
DFF     gate807  (.D(g5681), .CP(CLK), .Q(g5685) ) ;
OR2     gate808  (.A(g23564), .B(g18771), .Z(g24341) ) ;
DFF     gate809  (.D(g24341), .CP(CLK), .Q(g5689) ) ;
OR2     gate810  (.A(g23691), .B(g18772), .Z(g24342) ) ;
DFF     gate811  (.D(g24342), .CP(CLK), .Q(g5694) ) ;
OR2     gate812  (.A(g23724), .B(g18773), .Z(g24343) ) ;
DFF     gate813  (.D(g24343), .CP(CLK), .Q(g5698) ) ;
OR2     gate814  (.A(g33360), .B(g18774), .Z(g33620) ) ;
DFF     gate815  (.D(g33620), .CP(CLK), .Q(g5703) ) ;
OR2     gate816  (.A(g33365), .B(g18775), .Z(g33621) ) ;
DFF     gate817  (.D(g33621), .CP(CLK), .Q(g5644) ) ;
OR2     gate818  (.A(g25056), .B(g21965), .Z(g25714) ) ;
DFF     gate819  (.D(g25714), .CP(CLK), .Q(g5448) ) ;
DFF     gate820  (.D(g5448), .CP(CLK), .Q(g5456) ) ;
OR2     gate821  (.A(g25088), .B(g21967), .Z(g25716) ) ;
DFF     gate822  (.D(g25716), .CP(CLK), .Q(g5406) ) ;
OR2     gate823  (.A(g25071), .B(g21966), .Z(g25715) ) ;
DFF     gate824  (.D(g25715), .CP(CLK), .Q(g5452) ) ;
DFF     gate825  (.D(g5452), .CP(CLK), .Q(g5459) ) ;
OR2     gate826  (.A(g25106), .B(g21968), .Z(g25717) ) ;
DFF     gate827  (.D(g25717), .CP(CLK), .Q(g5366) ) ;
OR2     gate828  (.A(g31746), .B(g21952), .Z(g31905) ) ;
DFF     gate829  (.D(g31905), .CP(CLK), .Q(g5360) ) ;
OR2     gate830  (.A(g31750), .B(g21956), .Z(g31909) ) ;
DFF     gate831  (.D(g31909), .CP(CLK), .Q(g5373) ) ;
OR2     gate832  (.A(g31784), .B(g21969), .Z(g31911) ) ;
DFF     gate833  (.D(g31911), .CP(CLK), .Q(g5377) ) ;
OR2     gate834  (.A(g31477), .B(g21953), .Z(g31906) ) ;
DFF     gate835  (.D(g31906), .CP(CLK), .Q(g5381) ) ;
OR2     gate836  (.A(g31492), .B(g21954), .Z(g31907) ) ;
DFF     gate837  (.D(g31907), .CP(CLK), .Q(g5385) ) ;
OR2     gate838  (.A(g31519), .B(g21955), .Z(g31908) ) ;
DFF     gate839  (.D(g31908), .CP(CLK), .Q(g5390) ) ;
OR2     gate840  (.A(g31471), .B(g21957), .Z(g31910) ) ;
DFF     gate841  (.D(g31910), .CP(CLK), .Q(g5396) ) ;
OR2     gate842  (.A(g32316), .B(g21958), .Z(g33051) ) ;
DFF     gate843  (.D(g33051), .CP(CLK), .Q(g5401) ) ;
OR2     gate844  (.A(g27674), .B(g21970), .Z(g28095) ) ;
DFF     gate845  (.D(g28095), .CP(CLK), .Q(g5413) ) ;
OR2     gate846  (.A(g27673), .B(g21959), .Z(g28094) ) ;
DFF     gate847  (.D(g28094), .CP(CLK), .Q(g5417) ) ;
OR2     gate848  (.A(g25187), .B(g21971), .Z(g25718) ) ;
DFF     gate849  (.D(g25718), .CP(CLK), .Q(g5421) ) ;
OR2     gate850  (.A(g25014), .B(g21960), .Z(g25709) ) ;
DFF     gate851  (.D(g25709), .CP(CLK), .Q(g5424) ) ;
OR2     gate852  (.A(g25031), .B(g21961), .Z(g25710) ) ;
DFF     gate853  (.D(g25710), .CP(CLK), .Q(g5428) ) ;
OR2     gate854  (.A(g25105), .B(g21962), .Z(g25711) ) ;
DFF     gate855  (.D(g25711), .CP(CLK), .Q(g5436) ) ;
OR2     gate856  (.A(g25126), .B(g21963), .Z(g25712) ) ;
DFF     gate857  (.D(g25712), .CP(CLK), .Q(g5441) ) ;
OR2     gate858  (.A(g25147), .B(g21964), .Z(g25713) ) ;
DFF     gate859  (.D(g25713), .CP(CLK), .Q(g5445) ) ;
OR2     gate860  (.A(g29321), .B(g21972), .Z(g30480) ) ;
DFF     gate861  (.D(g30480), .CP(CLK), .Q(g5511) ) ;
OR2     gate862  (.A(g31961), .B(g21973), .Z(g33052) ) ;
DFF     gate863  (.D(g33052), .CP(CLK), .Q(g5517) ) ;
OR2     gate864  (.A(g31967), .B(g21974), .Z(g33053) ) ;
DFF     gate865  (.D(g33053), .CP(CLK), .Q(g5523) ) ;
OR2     gate866  (.A(g31975), .B(g21975), .Z(g33054) ) ;
DFF     gate867  (.D(g33054), .CP(CLK), .Q(g5527) ) ;
OR2     gate868  (.A(g31986), .B(g21976), .Z(g33055) ) ;
DFF     gate869  (.D(g33055), .CP(CLK), .Q(g5535) ) ;
OR2     gate870  (.A(g30221), .B(g21977), .Z(g30481) ) ;
DFF     gate871  (.D(g30481), .CP(CLK), .Q(g5543) ) ;
OR2     gate872  (.A(g30166), .B(g21981), .Z(g30485) ) ;
DFF     gate873  (.D(g30485), .CP(CLK), .Q(g5571) ) ;
OR2     gate874  (.A(g30250), .B(g21985), .Z(g30489) ) ;
DFF     gate875  (.D(g30489), .CP(CLK), .Q(g5587) ) ;
OR2     gate876  (.A(g30198), .B(g21989), .Z(g30493) ) ;
DFF     gate877  (.D(g30493), .CP(CLK), .Q(g5603) ) ;
OR2     gate878  (.A(g30242), .B(g21993), .Z(g30497) ) ;
DFF     gate879  (.D(g30497), .CP(CLK), .Q(g5551) ) ;
OR2     gate880  (.A(g30230), .B(g21978), .Z(g30482) ) ;
DFF     gate881  (.D(g30482), .CP(CLK), .Q(g5547) ) ;
OR2     gate882  (.A(g30177), .B(g21982), .Z(g30486) ) ;
DFF     gate883  (.D(g30486), .CP(CLK), .Q(g5575) ) ;
OR2     gate884  (.A(g30167), .B(g21986), .Z(g30490) ) ;
DFF     gate885  (.D(g30490), .CP(CLK), .Q(g5591) ) ;
OR2     gate886  (.A(g30209), .B(g21990), .Z(g30494) ) ;
DFF     gate887  (.D(g30494), .CP(CLK), .Q(g5607) ) ;
OR2     gate888  (.A(g30251), .B(g21994), .Z(g30498) ) ;
DFF     gate889  (.D(g30498), .CP(CLK), .Q(g5559) ) ;
OR2     gate890  (.A(g30241), .B(g21979), .Z(g30483) ) ;
DFF     gate891  (.D(g30483), .CP(CLK), .Q(g5555) ) ;
OR2     gate892  (.A(g30187), .B(g21983), .Z(g30487) ) ;
DFF     gate893  (.D(g30487), .CP(CLK), .Q(g5579) ) ;
OR2     gate894  (.A(g30178), .B(g21987), .Z(g30491) ) ;
DFF     gate895  (.D(g30491), .CP(CLK), .Q(g5595) ) ;
OR2     gate896  (.A(g30222), .B(g21991), .Z(g30495) ) ;
DFF     gate897  (.D(g30495), .CP(CLK), .Q(g5611) ) ;
OR2     gate898  (.A(g30261), .B(g21995), .Z(g30499) ) ;
DFF     gate899  (.D(g30499), .CP(CLK), .Q(g5567) ) ;
OR2     gate900  (.A(g30154), .B(g21980), .Z(g30484) ) ;
DFF     gate901  (.D(g30484), .CP(CLK), .Q(g5563) ) ;
OR2     gate902  (.A(g30197), .B(g21984), .Z(g30488) ) ;
DFF     gate903  (.D(g30488), .CP(CLK), .Q(g5583) ) ;
OR2     gate904  (.A(g30188), .B(g21988), .Z(g30492) ) ;
DFF     gate905  (.D(g30492), .CP(CLK), .Q(g5599) ) ;
OR2     gate906  (.A(g30231), .B(g21992), .Z(g30496) ) ;
DFF     gate907  (.D(g30496), .CP(CLK), .Q(g5615) ) ;
OR2     gate908  (.A(g29326), .B(g21996), .Z(g30500) ) ;
DFF     gate909  (.D(g30500), .CP(CLK), .Q(g5619) ) ;
OR2     gate910  (.A(g27988), .B(g21997), .Z(g28096) ) ;
DFF     gate911  (.D(g28096), .CP(CLK), .Q(g4821) ) ;
OR2     gate912  (.A(g28660), .B(g18767), .Z(g29291) ) ;
DFF     gate913  (.D(g29291), .CP(CLK), .Q(g5503) ) ;
OR2     gate914  (.A(g25530), .B(g18768), .Z(g25722) ) ;
DFF     gate915  (.D(g25722), .CP(CLK), .Q(g5467) ) ;
OR2     gate916  (.A(g28542), .B(g18759), .Z(g29286) ) ;
DFF     gate917  (.D(g29286), .CP(CLK), .Q(g5462) ) ;
OR2     gate918  (.A(g28555), .B(g18760), .Z(g29287) ) ;
DFF     gate919  (.D(g29287), .CP(CLK), .Q(g5471) ) ;
OR2     gate920  (.A(g25089), .B(g18761), .Z(g25719) ) ;
DFF     gate921  (.D(g25719), .CP(CLK), .Q(g5475) ) ;
OR2     gate922  (.A(g28630), .B(g18762), .Z(g29288) ) ;
DFF     gate923  (.D(g29288), .CP(CLK), .Q(g5481) ) ;
OR2     gate924  (.A(g28642), .B(g18763), .Z(g29289) ) ;
DFF     gate925  (.D(g29289), .CP(CLK), .Q(g5485) ) ;
OR2     gate926  (.A(g28569), .B(g18764), .Z(g29290) ) ;
DFF     gate927  (.D(g29290), .CP(CLK), .Q(g5489) ) ;
OR2     gate928  (.A(g25042), .B(g18765), .Z(g25720) ) ;
DFF     gate929  (.D(g25720), .CP(CLK), .Q(g5495) ) ;
OR2     gate930  (.A(g25057), .B(g18766), .Z(g25721) ) ;
DFF     gate931  (.D(g25721), .CP(CLK), .Q(g5499) ) ;
OR2     gate932  (.A(g34555), .B(g18769), .Z(g34644) ) ;
DFF     gate933  (.D(g34644), .CP(CLK), .Q(g5507) ) ;
OR2     gate934  (.A(g22145), .B(g18787), .Z(g24344) ) ;
DFF     gate935  (.D(g24344), .CP(CLK), .Q(g6005) ) ;
DFF     gate936  (.D(g6005), .CP(CLK), .Q(g5983) ) ;
DFF     gate937  (.D(g5983), .CP(CLK), .Q(g6012) ) ;
DFF     gate938  (.D(g6012), .CP(CLK), .Q(g5969) ) ;
DFF     gate939  (.D(g5969), .CP(CLK), .Q(g5976) ) ;
DFF     gate940  (.D(g5976), .CP(CLK), .Q(g6000) ) ;
DFF     gate941  (.D(g6000), .CP(CLK), .Q(g6019) ) ;
DFF     gate942  (.D(g6019), .CP(CLK), .Q(g6023) ) ;
DFF     gate943  (.D(g6023), .CP(CLK), .Q(g6027) ) ;
DFF     gate944  (.D(g6027), .CP(CLK), .Q(g6031) ) ;
OR2     gate945  (.A(g23606), .B(g18788), .Z(g24345) ) ;
DFF     gate946  (.D(g24345), .CP(CLK), .Q(g6035) ) ;
OR2     gate947  (.A(g23725), .B(g18789), .Z(g24346) ) ;
DFF     gate948  (.D(g24346), .CP(CLK), .Q(g6040) ) ;
OR2     gate949  (.A(g23754), .B(g18790), .Z(g24347) ) ;
DFF     gate950  (.D(g24347), .CP(CLK), .Q(g6044) ) ;
OR2     gate951  (.A(g33366), .B(g18791), .Z(g33622) ) ;
DFF     gate952  (.D(g33622), .CP(CLK), .Q(g6049) ) ;
OR2     gate953  (.A(g33370), .B(g18792), .Z(g33623) ) ;
DFF     gate954  (.D(g33623), .CP(CLK), .Q(g5990) ) ;
OR2     gate955  (.A(g25076), .B(g22011), .Z(g25728) ) ;
DFF     gate956  (.D(g25728), .CP(CLK), .Q(g5794) ) ;
DFF     gate957  (.D(g5794), .CP(CLK), .Q(g5802) ) ;
OR2     gate958  (.A(g25107), .B(g22013), .Z(g25730) ) ;
DFF     gate959  (.D(g25730), .CP(CLK), .Q(g5752) ) ;
OR2     gate960  (.A(g25091), .B(g22012), .Z(g25729) ) ;
DFF     gate961  (.D(g25729), .CP(CLK), .Q(g5798) ) ;
DFF     gate962  (.D(g5798), .CP(CLK), .Q(g5805) ) ;
OR2     gate963  (.A(g25128), .B(g22014), .Z(g25731) ) ;
DFF     gate964  (.D(g25731), .CP(CLK), .Q(g5712) ) ;
OR2     gate965  (.A(g31752), .B(g21998), .Z(g31912) ) ;
DFF     gate966  (.D(g31912), .CP(CLK), .Q(g5706) ) ;
OR2     gate967  (.A(g31756), .B(g22002), .Z(g31916) ) ;
DFF     gate968  (.D(g31916), .CP(CLK), .Q(g5719) ) ;
OR2     gate969  (.A(g31786), .B(g22015), .Z(g31918) ) ;
DFF     gate970  (.D(g31918), .CP(CLK), .Q(g5723) ) ;
OR2     gate971  (.A(g31485), .B(g21999), .Z(g31913) ) ;
DFF     gate972  (.D(g31913), .CP(CLK), .Q(g5727) ) ;
OR2     gate973  (.A(g31499), .B(g22000), .Z(g31914) ) ;
DFF     gate974  (.D(g31914), .CP(CLK), .Q(g5731) ) ;
OR2     gate975  (.A(g31520), .B(g22001), .Z(g31915) ) ;
DFF     gate976  (.D(g31915), .CP(CLK), .Q(g5736) ) ;
OR2     gate977  (.A(g31478), .B(g22003), .Z(g31917) ) ;
DFF     gate978  (.D(g31917), .CP(CLK), .Q(g5742) ) ;
OR2     gate979  (.A(g32327), .B(g22004), .Z(g33056) ) ;
DFF     gate980  (.D(g33056), .CP(CLK), .Q(g5747) ) ;
OR2     gate981  (.A(g27683), .B(g22016), .Z(g28098) ) ;
DFF     gate982  (.D(g28098), .CP(CLK), .Q(g5759) ) ;
OR2     gate983  (.A(g27682), .B(g22005), .Z(g28097) ) ;
DFF     gate984  (.D(g28097), .CP(CLK), .Q(g5763) ) ;
OR2     gate985  (.A(g25201), .B(g22017), .Z(g25732) ) ;
DFF     gate986  (.D(g25732), .CP(CLK), .Q(g5767) ) ;
OR2     gate987  (.A(g25033), .B(g22006), .Z(g25723) ) ;
DFF     gate988  (.D(g25723), .CP(CLK), .Q(g5770) ) ;
OR2     gate989  (.A(g25043), .B(g22007), .Z(g25724) ) ;
DFF     gate990  (.D(g25724), .CP(CLK), .Q(g5774) ) ;
OR2     gate991  (.A(g25127), .B(g22008), .Z(g25725) ) ;
DFF     gate992  (.D(g25725), .CP(CLK), .Q(g5782) ) ;
OR2     gate993  (.A(g25148), .B(g22009), .Z(g25726) ) ;
DFF     gate994  (.D(g25726), .CP(CLK), .Q(g5787) ) ;
OR2     gate995  (.A(g25163), .B(g22010), .Z(g25727) ) ;
DFF     gate996  (.D(g25727), .CP(CLK), .Q(g5791) ) ;
OR2     gate997  (.A(g29327), .B(g22018), .Z(g30501) ) ;
DFF     gate998  (.D(g30501), .CP(CLK), .Q(g5857) ) ;
OR2     gate999  (.A(g31968), .B(g22019), .Z(g33057) ) ;
DFF     gate1000  (.D(g33057), .CP(CLK), .Q(g5863) ) ;
OR2     gate1001  (.A(g31976), .B(g22020), .Z(g33058) ) ;
DFF     gate1002  (.D(g33058), .CP(CLK), .Q(g5869) ) ;
OR2     gate1003  (.A(g31987), .B(g22021), .Z(g33059) ) ;
DFF     gate1004  (.D(g33059), .CP(CLK), .Q(g5873) ) ;
OR2     gate1005  (.A(g31992), .B(g22022), .Z(g33060) ) ;
DFF     gate1006  (.D(g33060), .CP(CLK), .Q(g5881) ) ;
OR2     gate1007  (.A(g30232), .B(g22023), .Z(g30502) ) ;
DFF     gate1008  (.D(g30502), .CP(CLK), .Q(g5889) ) ;
OR2     gate1009  (.A(g30179), .B(g22027), .Z(g30506) ) ;
DFF     gate1010  (.D(g30506), .CP(CLK), .Q(g5917) ) ;
OR2     gate1011  (.A(g30263), .B(g22031), .Z(g30510) ) ;
DFF     gate1012  (.D(g30510), .CP(CLK), .Q(g5933) ) ;
OR2     gate1013  (.A(g30211), .B(g22035), .Z(g30514) ) ;
DFF     gate1014  (.D(g30514), .CP(CLK), .Q(g5949) ) ;
OR2     gate1015  (.A(g30254), .B(g22039), .Z(g30518) ) ;
DFF     gate1016  (.D(g30518), .CP(CLK), .Q(g5897) ) ;
OR2     gate1017  (.A(g30243), .B(g22024), .Z(g30503) ) ;
DFF     gate1018  (.D(g30503), .CP(CLK), .Q(g5893) ) ;
OR2     gate1019  (.A(g30190), .B(g22028), .Z(g30507) ) ;
DFF     gate1020  (.D(g30507), .CP(CLK), .Q(g5921) ) ;
OR2     gate1021  (.A(g30180), .B(g22032), .Z(g30511) ) ;
DFF     gate1022  (.D(g30511), .CP(CLK), .Q(g5937) ) ;
OR2     gate1023  (.A(g30223), .B(g22036), .Z(g30515) ) ;
DFF     gate1024  (.D(g30515), .CP(CLK), .Q(g5953) ) ;
OR2     gate1025  (.A(g30264), .B(g22040), .Z(g30519) ) ;
DFF     gate1026  (.D(g30519), .CP(CLK), .Q(g5905) ) ;
OR2     gate1027  (.A(g30253), .B(g22025), .Z(g30504) ) ;
DFF     gate1028  (.D(g30504), .CP(CLK), .Q(g5901) ) ;
OR2     gate1029  (.A(g30199), .B(g22029), .Z(g30508) ) ;
DFF     gate1030  (.D(g30508), .CP(CLK), .Q(g5925) ) ;
OR2     gate1031  (.A(g30191), .B(g22033), .Z(g30512) ) ;
DFF     gate1032  (.D(g30512), .CP(CLK), .Q(g5941) ) ;
OR2     gate1033  (.A(g30233), .B(g22037), .Z(g30516) ) ;
DFF     gate1034  (.D(g30516), .CP(CLK), .Q(g5957) ) ;
OR2     gate1035  (.A(g30272), .B(g22041), .Z(g30520) ) ;
DFF     gate1036  (.D(g30520), .CP(CLK), .Q(g5913) ) ;
OR2     gate1037  (.A(g30168), .B(g22026), .Z(g30505) ) ;
DFF     gate1038  (.D(g30505), .CP(CLK), .Q(g5909) ) ;
OR2     gate1039  (.A(g30210), .B(g22030), .Z(g30509) ) ;
DFF     gate1040  (.D(g30509), .CP(CLK), .Q(g5929) ) ;
OR2     gate1041  (.A(g30200), .B(g22034), .Z(g30513) ) ;
DFF     gate1042  (.D(g30513), .CP(CLK), .Q(g5945) ) ;
OR2     gate1043  (.A(g30244), .B(g22038), .Z(g30517) ) ;
DFF     gate1044  (.D(g30517), .CP(CLK), .Q(g5961) ) ;
OR2     gate1045  (.A(g29331), .B(g22042), .Z(g30521) ) ;
DFF     gate1046  (.D(g30521), .CP(CLK), .Q(g5965) ) ;
OR2     gate1047  (.A(g27992), .B(g22043), .Z(g28099) ) ;
DFF     gate1048  (.D(g28099), .CP(CLK), .Q(g4831) ) ;
OR2     gate1049  (.A(g28683), .B(g18784), .Z(g29297) ) ;
DFF     gate1050  (.D(g29297), .CP(CLK), .Q(g5849) ) ;
OR2     gate1051  (.A(g25536), .B(g18785), .Z(g25736) ) ;
DFF     gate1052  (.D(g25736), .CP(CLK), .Q(g5813) ) ;
OR2     gate1053  (.A(g28556), .B(g18776), .Z(g29292) ) ;
DFF     gate1054  (.D(g29292), .CP(CLK), .Q(g5808) ) ;
OR2     gate1055  (.A(g28570), .B(g18777), .Z(g29293) ) ;
DFF     gate1056  (.D(g29293), .CP(CLK), .Q(g5817) ) ;
OR2     gate1057  (.A(g25108), .B(g18778), .Z(g25733) ) ;
DFF     gate1058  (.D(g25733), .CP(CLK), .Q(g5821) ) ;
OR2     gate1059  (.A(g28645), .B(g18779), .Z(g29294) ) ;
DFF     gate1060  (.D(g29294), .CP(CLK), .Q(g5827) ) ;
OR2     gate1061  (.A(g28663), .B(g18780), .Z(g29295) ) ;
DFF     gate1062  (.D(g29295), .CP(CLK), .Q(g5831) ) ;
OR2     gate1063  (.A(g28586), .B(g18781), .Z(g29296) ) ;
DFF     gate1064  (.D(g29296), .CP(CLK), .Q(g5835) ) ;
OR2     gate1065  (.A(g25058), .B(g18782), .Z(g25734) ) ;
DFF     gate1066  (.D(g25734), .CP(CLK), .Q(g5841) ) ;
OR2     gate1067  (.A(g25077), .B(g18783), .Z(g25735) ) ;
DFF     gate1068  (.D(g25735), .CP(CLK), .Q(g5845) ) ;
OR2     gate1069  (.A(g34556), .B(g18786), .Z(g34645) ) ;
DFF     gate1070  (.D(g34645), .CP(CLK), .Q(g5853) ) ;
OR2     gate1071  (.A(g22149), .B(g18804), .Z(g24348) ) ;
DFF     gate1072  (.D(g24348), .CP(CLK), .Q(g6351) ) ;
DFF     gate1073  (.D(g6351), .CP(CLK), .Q(g6329) ) ;
DFF     gate1074  (.D(g6329), .CP(CLK), .Q(g6358) ) ;
DFF     gate1075  (.D(g6358), .CP(CLK), .Q(g6315) ) ;
DFF     gate1076  (.D(g6315), .CP(CLK), .Q(g6322) ) ;
DFF     gate1077  (.D(g6322), .CP(CLK), .Q(g6346) ) ;
DFF     gate1078  (.D(g6346), .CP(CLK), .Q(g6365) ) ;
DFF     gate1079  (.D(g6365), .CP(CLK), .Q(g6369) ) ;
DFF     gate1080  (.D(g6369), .CP(CLK), .Q(g6373) ) ;
DFF     gate1081  (.D(g6373), .CP(CLK), .Q(g6377) ) ;
OR2     gate1082  (.A(g23646), .B(g18805), .Z(g24349) ) ;
DFF     gate1083  (.D(g24349), .CP(CLK), .Q(g6381) ) ;
OR2     gate1084  (.A(g23755), .B(g18806), .Z(g24350) ) ;
DFF     gate1085  (.D(g24350), .CP(CLK), .Q(g6386) ) ;
OR2     gate1086  (.A(g23774), .B(g18807), .Z(g24351) ) ;
DFF     gate1087  (.D(g24351), .CP(CLK), .Q(g6390) ) ;
OR2     gate1088  (.A(g33371), .B(g18808), .Z(g33624) ) ;
DFF     gate1089  (.D(g33624), .CP(CLK), .Q(g6395) ) ;
OR2     gate1090  (.A(g33373), .B(g18809), .Z(g33625) ) ;
DFF     gate1091  (.D(g33625), .CP(CLK), .Q(g6336) ) ;
OR2     gate1092  (.A(g25093), .B(g22057), .Z(g25742) ) ;
DFF     gate1093  (.D(g25742), .CP(CLK), .Q(g6140) ) ;
DFF     gate1094  (.D(g6140), .CP(CLK), .Q(g6148) ) ;
OR2     gate1095  (.A(g25129), .B(g22059), .Z(g25744) ) ;
DFF     gate1096  (.D(g25744), .CP(CLK), .Q(g6098) ) ;
OR2     gate1097  (.A(g25110), .B(g22058), .Z(g25743) ) ;
DFF     gate1098  (.D(g25743), .CP(CLK), .Q(g6144) ) ;
DFF     gate1099  (.D(g6144), .CP(CLK), .Q(g6151) ) ;
OR2     gate1100  (.A(g25150), .B(g22060), .Z(g25745) ) ;
DFF     gate1101  (.D(g25745), .CP(CLK), .Q(g6058) ) ;
OR2     gate1102  (.A(g31758), .B(g22044), .Z(g31919) ) ;
DFF     gate1103  (.D(g31919), .CP(CLK), .Q(g6052) ) ;
OR2     gate1104  (.A(g31763), .B(g22048), .Z(g31923) ) ;
DFF     gate1105  (.D(g31923), .CP(CLK), .Q(g6065) ) ;
OR2     gate1106  (.A(g31789), .B(g22061), .Z(g31925) ) ;
DFF     gate1107  (.D(g31925), .CP(CLK), .Q(g6069) ) ;
OR2     gate1108  (.A(g31493), .B(g22045), .Z(g31920) ) ;
DFF     gate1109  (.D(g31920), .CP(CLK), .Q(g6073) ) ;
OR2     gate1110  (.A(g31508), .B(g22046), .Z(g31921) ) ;
DFF     gate1111  (.D(g31921), .CP(CLK), .Q(g6077) ) ;
OR2     gate1112  (.A(g31525), .B(g22047), .Z(g31922) ) ;
DFF     gate1113  (.D(g31922), .CP(CLK), .Q(g6082) ) ;
OR2     gate1114  (.A(g31486), .B(g22049), .Z(g31924) ) ;
DFF     gate1115  (.D(g31924), .CP(CLK), .Q(g6088) ) ;
OR2     gate1116  (.A(g32334), .B(g22050), .Z(g33061) ) ;
DFF     gate1117  (.D(g33061), .CP(CLK), .Q(g6093) ) ;
OR2     gate1118  (.A(g27691), .B(g22062), .Z(g28101) ) ;
DFF     gate1119  (.D(g28101), .CP(CLK), .Q(g6105) ) ;
OR2     gate1120  (.A(g27690), .B(g22051), .Z(g28100) ) ;
DFF     gate1121  (.D(g28100), .CP(CLK), .Q(g6109) ) ;
OR2     gate1122  (.A(g25217), .B(g22063), .Z(g25746) ) ;
DFF     gate1123  (.D(g25746), .CP(CLK), .Q(g6113) ) ;
OR2     gate1124  (.A(g25045), .B(g22052), .Z(g25737) ) ;
DFF     gate1125  (.D(g25737), .CP(CLK), .Q(g6116) ) ;
OR2     gate1126  (.A(g25059), .B(g22053), .Z(g25738) ) ;
DFF     gate1127  (.D(g25738), .CP(CLK), .Q(g6120) ) ;
OR2     gate1128  (.A(g25149), .B(g22054), .Z(g25739) ) ;
DFF     gate1129  (.D(g25739), .CP(CLK), .Q(g6128) ) ;
OR2     gate1130  (.A(g25164), .B(g22055), .Z(g25740) ) ;
DFF     gate1131  (.D(g25740), .CP(CLK), .Q(g6133) ) ;
OR2     gate1132  (.A(g25178), .B(g22056), .Z(g25741) ) ;
DFF     gate1133  (.D(g25741), .CP(CLK), .Q(g6137) ) ;
OR2     gate1134  (.A(g29332), .B(g22064), .Z(g30522) ) ;
DFF     gate1135  (.D(g30522), .CP(CLK), .Q(g6203) ) ;
OR2     gate1136  (.A(g31977), .B(g22065), .Z(g33062) ) ;
DFF     gate1137  (.D(g33062), .CP(CLK), .Q(g6209) ) ;
OR2     gate1138  (.A(g31988), .B(g22066), .Z(g33063) ) ;
DFF     gate1139  (.D(g33063), .CP(CLK), .Q(g6215) ) ;
OR2     gate1140  (.A(g31993), .B(g22067), .Z(g33064) ) ;
DFF     gate1141  (.D(g33064), .CP(CLK), .Q(g6219) ) ;
OR2     gate1142  (.A(g32008), .B(g22068), .Z(g33065) ) ;
DFF     gate1143  (.D(g33065), .CP(CLK), .Q(g6227) ) ;
OR2     gate1144  (.A(g30245), .B(g22069), .Z(g30523) ) ;
DFF     gate1145  (.D(g30523), .CP(CLK), .Q(g6235) ) ;
OR2     gate1146  (.A(g30192), .B(g22073), .Z(g30527) ) ;
DFF     gate1147  (.D(g30527), .CP(CLK), .Q(g6263) ) ;
OR2     gate1148  (.A(g30274), .B(g22077), .Z(g30531) ) ;
DFF     gate1149  (.D(g30531), .CP(CLK), .Q(g6279) ) ;
OR2     gate1150  (.A(g30225), .B(g22081), .Z(g30535) ) ;
DFF     gate1151  (.D(g30535), .CP(CLK), .Q(g6295) ) ;
OR2     gate1152  (.A(g30267), .B(g22085), .Z(g30539) ) ;
DFF     gate1153  (.D(g30539), .CP(CLK), .Q(g6243) ) ;
OR2     gate1154  (.A(g30255), .B(g22070), .Z(g30524) ) ;
DFF     gate1155  (.D(g30524), .CP(CLK), .Q(g6239) ) ;
OR2     gate1156  (.A(g30202), .B(g22074), .Z(g30528) ) ;
DFF     gate1157  (.D(g30528), .CP(CLK), .Q(g6267) ) ;
OR2     gate1158  (.A(g30193), .B(g22078), .Z(g30532) ) ;
DFF     gate1159  (.D(g30532), .CP(CLK), .Q(g6283) ) ;
OR2     gate1160  (.A(g30234), .B(g22082), .Z(g30536) ) ;
DFF     gate1161  (.D(g30536), .CP(CLK), .Q(g6299) ) ;
OR2     gate1162  (.A(g30275), .B(g22086), .Z(g30540) ) ;
DFF     gate1163  (.D(g30540), .CP(CLK), .Q(g6251) ) ;
OR2     gate1164  (.A(g30266), .B(g22071), .Z(g30525) ) ;
DFF     gate1165  (.D(g30525), .CP(CLK), .Q(g6247) ) ;
OR2     gate1166  (.A(g30212), .B(g22075), .Z(g30529) ) ;
DFF     gate1167  (.D(g30529), .CP(CLK), .Q(g6271) ) ;
OR2     gate1168  (.A(g30203), .B(g22079), .Z(g30533) ) ;
DFF     gate1169  (.D(g30533), .CP(CLK), .Q(g6287) ) ;
OR2     gate1170  (.A(g30246), .B(g22083), .Z(g30537) ) ;
DFF     gate1171  (.D(g30537), .CP(CLK), .Q(g6303) ) ;
OR2     gate1172  (.A(g30281), .B(g22087), .Z(g30541) ) ;
DFF     gate1173  (.D(g30541), .CP(CLK), .Q(g6259) ) ;
OR2     gate1174  (.A(g30181), .B(g22072), .Z(g30526) ) ;
DFF     gate1175  (.D(g30526), .CP(CLK), .Q(g6255) ) ;
OR2     gate1176  (.A(g30224), .B(g22076), .Z(g30530) ) ;
DFF     gate1177  (.D(g30530), .CP(CLK), .Q(g6275) ) ;
OR2     gate1178  (.A(g30213), .B(g22080), .Z(g30534) ) ;
DFF     gate1179  (.D(g30534), .CP(CLK), .Q(g6291) ) ;
OR2     gate1180  (.A(g30256), .B(g22084), .Z(g30538) ) ;
DFF     gate1181  (.D(g30538), .CP(CLK), .Q(g6307) ) ;
OR2     gate1182  (.A(g29337), .B(g22088), .Z(g30542) ) ;
DFF     gate1183  (.D(g30542), .CP(CLK), .Q(g6311) ) ;
OR2     gate1184  (.A(g27995), .B(g22089), .Z(g28102) ) ;
DFF     gate1185  (.D(g28102), .CP(CLK), .Q(g4826) ) ;
OR2     gate1186  (.A(g28703), .B(g18801), .Z(g29303) ) ;
DFF     gate1187  (.D(g29303), .CP(CLK), .Q(g6195) ) ;
OR2     gate1188  (.A(g25543), .B(g18802), .Z(g25750) ) ;
DFF     gate1189  (.D(g25750), .CP(CLK), .Q(g6159) ) ;
OR2     gate1190  (.A(g28571), .B(g18793), .Z(g29298) ) ;
DFF     gate1191  (.D(g29298), .CP(CLK), .Q(g6154) ) ;
OR2     gate1192  (.A(g28587), .B(g18794), .Z(g29299) ) ;
DFF     gate1193  (.D(g29299), .CP(CLK), .Q(g6163) ) ;
OR2     gate1194  (.A(g25130), .B(g18795), .Z(g25747) ) ;
DFF     gate1195  (.D(g25747), .CP(CLK), .Q(g6167) ) ;
OR2     gate1196  (.A(g28666), .B(g18796), .Z(g29300) ) ;
DFF     gate1197  (.D(g29300), .CP(CLK), .Q(g6173) ) ;
OR2     gate1198  (.A(g28686), .B(g18797), .Z(g29301) ) ;
DFF     gate1199  (.D(g29301), .CP(CLK), .Q(g6177) ) ;
OR2     gate1200  (.A(g28601), .B(g18798), .Z(g29302) ) ;
DFF     gate1201  (.D(g29302), .CP(CLK), .Q(g6181) ) ;
OR2     gate1202  (.A(g25078), .B(g18799), .Z(g25748) ) ;
DFF     gate1203  (.D(g25748), .CP(CLK), .Q(g6187) ) ;
OR2     gate1204  (.A(g25094), .B(g18800), .Z(g25749) ) ;
DFF     gate1205  (.D(g25749), .CP(CLK), .Q(g6191) ) ;
OR2     gate1206  (.A(g34557), .B(g18803), .Z(g34646) ) ;
DFF     gate1207  (.D(g34646), .CP(CLK), .Q(g6199) ) ;
OR2     gate1208  (.A(g22157), .B(g18821), .Z(g24352) ) ;
DFF     gate1209  (.D(g24352), .CP(CLK), .Q(g6697) ) ;
DFF     gate1210  (.D(g6697), .CP(CLK), .Q(g6675) ) ;
DFF     gate1211  (.D(g6675), .CP(CLK), .Q(g6704) ) ;
DFF     gate1212  (.D(g6704), .CP(CLK), .Q(g6661) ) ;
DFF     gate1213  (.D(g6661), .CP(CLK), .Q(g6668) ) ;
DFF     gate1214  (.D(g6668), .CP(CLK), .Q(g6692) ) ;
DFF     gate1215  (.D(g6692), .CP(CLK), .Q(g6711) ) ;
DFF     gate1216  (.D(g6711), .CP(CLK), .Q(g6715) ) ;
DFF     gate1217  (.D(g6715), .CP(CLK), .Q(g6719) ) ;
DFF     gate1218  (.D(g6719), .CP(CLK), .Q(g6723) ) ;
OR2     gate1219  (.A(g23682), .B(g18822), .Z(g24353) ) ;
DFF     gate1220  (.D(g24353), .CP(CLK), .Q(g6727) ) ;
OR2     gate1221  (.A(g23775), .B(g18823), .Z(g24354) ) ;
DFF     gate1222  (.D(g24354), .CP(CLK), .Q(g6732) ) ;
OR2     gate1223  (.A(g23799), .B(g18824), .Z(g24355) ) ;
DFF     gate1224  (.D(g24355), .CP(CLK), .Q(g6736) ) ;
OR2     gate1225  (.A(g33374), .B(g18825), .Z(g33626) ) ;
DFF     gate1226  (.D(g33626), .CP(CLK), .Q(g6741) ) ;
OR2     gate1227  (.A(g33376), .B(g18826), .Z(g33627) ) ;
DFF     gate1228  (.D(g33627), .CP(CLK), .Q(g6682) ) ;
OR2     gate1229  (.A(g25112), .B(g22103), .Z(g25756) ) ;
DFF     gate1230  (.D(g25756), .CP(CLK), .Q(g6486) ) ;
DFF     gate1231  (.D(g6486), .CP(CLK), .Q(g6494) ) ;
OR2     gate1232  (.A(g25151), .B(g22105), .Z(g25758) ) ;
DFF     gate1233  (.D(g25758), .CP(CLK), .Q(g6444) ) ;
OR2     gate1234  (.A(g25132), .B(g22104), .Z(g25757) ) ;
DFF     gate1235  (.D(g25757), .CP(CLK), .Q(g6490) ) ;
DFF     gate1236  (.D(g6490), .CP(CLK), .Q(g6497) ) ;
OR2     gate1237  (.A(g25166), .B(g22106), .Z(g25759) ) ;
DFF     gate1238  (.D(g25759), .CP(CLK), .Q(g6404) ) ;
OR2     gate1239  (.A(g31765), .B(g22090), .Z(g31926) ) ;
DFF     gate1240  (.D(g31926), .CP(CLK), .Q(g6398) ) ;
OR2     gate1241  (.A(g31769), .B(g22094), .Z(g31930) ) ;
DFF     gate1242  (.D(g31930), .CP(CLK), .Q(g6411) ) ;
OR2     gate1243  (.A(g31792), .B(g22107), .Z(g31932) ) ;
DFF     gate1244  (.D(g31932), .CP(CLK), .Q(g6415) ) ;
OR2     gate1245  (.A(g31500), .B(g22091), .Z(g31927) ) ;
DFF     gate1246  (.D(g31927), .CP(CLK), .Q(g6419) ) ;
OR2     gate1247  (.A(g31517), .B(g22092), .Z(g31928) ) ;
DFF     gate1248  (.D(g31928), .CP(CLK), .Q(g6423) ) ;
OR2     gate1249  (.A(g31540), .B(g22093), .Z(g31929) ) ;
DFF     gate1250  (.D(g31929), .CP(CLK), .Q(g6428) ) ;
OR2     gate1251  (.A(g31494), .B(g22095), .Z(g31931) ) ;
DFF     gate1252  (.D(g31931), .CP(CLK), .Q(g6434) ) ;
OR2     gate1253  (.A(g32341), .B(g22096), .Z(g33066) ) ;
DFF     gate1254  (.D(g33066), .CP(CLK), .Q(g6439) ) ;
OR2     gate1255  (.A(g27697), .B(g22108), .Z(g28104) ) ;
DFF     gate1256  (.D(g28104), .CP(CLK), .Q(g6451) ) ;
OR2     gate1257  (.A(g27696), .B(g22097), .Z(g28103) ) ;
DFF     gate1258  (.D(g28103), .CP(CLK), .Q(g6455) ) ;
OR2     gate1259  (.A(g25238), .B(g22109), .Z(g25760) ) ;
DFF     gate1260  (.D(g25760), .CP(CLK), .Q(g6459) ) ;
OR2     gate1261  (.A(g25061), .B(g22098), .Z(g25751) ) ;
DFF     gate1262  (.D(g25751), .CP(CLK), .Q(g6462) ) ;
OR2     gate1263  (.A(g25079), .B(g22099), .Z(g25752) ) ;
DFF     gate1264  (.D(g25752), .CP(CLK), .Q(g6466) ) ;
OR2     gate1265  (.A(g25165), .B(g22100), .Z(g25753) ) ;
DFF     gate1266  (.D(g25753), .CP(CLK), .Q(g6474) ) ;
OR2     gate1267  (.A(g25179), .B(g22101), .Z(g25754) ) ;
DFF     gate1268  (.D(g25754), .CP(CLK), .Q(g6479) ) ;
OR2     gate1269  (.A(g25192), .B(g22102), .Z(g25755) ) ;
DFF     gate1270  (.D(g25755), .CP(CLK), .Q(g6483) ) ;
OR2     gate1271  (.A(g29338), .B(g22110), .Z(g30543) ) ;
DFF     gate1272  (.D(g30543), .CP(CLK), .Q(g6549) ) ;
OR2     gate1273  (.A(g31989), .B(g22111), .Z(g33067) ) ;
DFF     gate1274  (.D(g33067), .CP(CLK), .Q(g6555) ) ;
OR2     gate1275  (.A(g31994), .B(g22112), .Z(g33068) ) ;
DFF     gate1276  (.D(g33068), .CP(CLK), .Q(g6561) ) ;
OR2     gate1277  (.A(g32009), .B(g22113), .Z(g33069) ) ;
DFF     gate1278  (.D(g33069), .CP(CLK), .Q(g6565) ) ;
OR2     gate1279  (.A(g32010), .B(g22114), .Z(g33070) ) ;
DFF     gate1280  (.D(g33070), .CP(CLK), .Q(g6573) ) ;
OR2     gate1281  (.A(g30257), .B(g22115), .Z(g30544) ) ;
DFF     gate1282  (.D(g30544), .CP(CLK), .Q(g6581) ) ;
OR2     gate1283  (.A(g30204), .B(g22119), .Z(g30548) ) ;
DFF     gate1284  (.D(g30548), .CP(CLK), .Q(g6609) ) ;
OR2     gate1285  (.A(g30283), .B(g22123), .Z(g30552) ) ;
DFF     gate1286  (.D(g30552), .CP(CLK), .Q(g6625) ) ;
OR2     gate1287  (.A(g30236), .B(g22127), .Z(g30556) ) ;
DFF     gate1288  (.D(g30556), .CP(CLK), .Q(g6641) ) ;
OR2     gate1289  (.A(g30278), .B(g22131), .Z(g30560) ) ;
DFF     gate1290  (.D(g30560), .CP(CLK), .Q(g6589) ) ;
OR2     gate1291  (.A(g30268), .B(g22116), .Z(g30545) ) ;
DFF     gate1292  (.D(g30545), .CP(CLK), .Q(g6585) ) ;
OR2     gate1293  (.A(g30215), .B(g22120), .Z(g30549) ) ;
DFF     gate1294  (.D(g30549), .CP(CLK), .Q(g6613) ) ;
OR2     gate1295  (.A(g30205), .B(g22124), .Z(g30553) ) ;
DFF     gate1296  (.D(g30553), .CP(CLK), .Q(g6629) ) ;
OR2     gate1297  (.A(g30247), .B(g22128), .Z(g30557) ) ;
DFF     gate1298  (.D(g30557), .CP(CLK), .Q(g6645) ) ;
OR2     gate1299  (.A(g30284), .B(g22132), .Z(g30561) ) ;
DFF     gate1300  (.D(g30561), .CP(CLK), .Q(g6597) ) ;
OR2     gate1301  (.A(g30277), .B(g22117), .Z(g30546) ) ;
DFF     gate1302  (.D(g30546), .CP(CLK), .Q(g6593) ) ;
OR2     gate1303  (.A(g30226), .B(g22121), .Z(g30550) ) ;
DFF     gate1304  (.D(g30550), .CP(CLK), .Q(g6617) ) ;
OR2     gate1305  (.A(g30216), .B(g22125), .Z(g30554) ) ;
DFF     gate1306  (.D(g30554), .CP(CLK), .Q(g6633) ) ;
OR2     gate1307  (.A(g30258), .B(g22129), .Z(g30558) ) ;
DFF     gate1308  (.D(g30558), .CP(CLK), .Q(g6649) ) ;
OR2     gate1309  (.A(g30289), .B(g22133), .Z(g30562) ) ;
DFF     gate1310  (.D(g30562), .CP(CLK), .Q(g6605) ) ;
OR2     gate1311  (.A(g30194), .B(g22118), .Z(g30547) ) ;
DFF     gate1312  (.D(g30547), .CP(CLK), .Q(g6601) ) ;
OR2     gate1313  (.A(g30235), .B(g22122), .Z(g30551) ) ;
DFF     gate1314  (.D(g30551), .CP(CLK), .Q(g6621) ) ;
OR2     gate1315  (.A(g30227), .B(g22126), .Z(g30555) ) ;
DFF     gate1316  (.D(g30555), .CP(CLK), .Q(g6637) ) ;
OR2     gate1317  (.A(g30269), .B(g22130), .Z(g30559) ) ;
DFF     gate1318  (.D(g30559), .CP(CLK), .Q(g6653) ) ;
OR2     gate1319  (.A(g29347), .B(g22134), .Z(g30563) ) ;
DFF     gate1320  (.D(g30563), .CP(CLK), .Q(g6657) ) ;
OR2     gate1321  (.A(g27997), .B(g22135), .Z(g28105) ) ;
DFF     gate1322  (.D(g28105), .CP(CLK), .Q(g5011) ) ;
OR2     gate1323  (.A(g28722), .B(g18818), .Z(g29309) ) ;
DFF     gate1324  (.D(g29309), .CP(CLK), .Q(g6541) ) ;
OR2     gate1325  (.A(g25551), .B(g18819), .Z(g25764) ) ;
DFF     gate1326  (.D(g25764), .CP(CLK), .Q(g6505) ) ;
OR2     gate1327  (.A(g28588), .B(g18810), .Z(g29304) ) ;
DFF     gate1328  (.D(g29304), .CP(CLK), .Q(g6500) ) ;
OR2     gate1329  (.A(g28602), .B(g18811), .Z(g29305) ) ;
DFF     gate1330  (.D(g29305), .CP(CLK), .Q(g6509) ) ;
OR2     gate1331  (.A(g25152), .B(g18812), .Z(g25761) ) ;
DFF     gate1332  (.D(g25761), .CP(CLK), .Q(g6513) ) ;
OR2     gate1333  (.A(g28689), .B(g18813), .Z(g29306) ) ;
DFF     gate1334  (.D(g29306), .CP(CLK), .Q(g6519) ) ;
OR2     gate1335  (.A(g28706), .B(g18814), .Z(g29307) ) ;
DFF     gate1336  (.D(g29307), .CP(CLK), .Q(g6523) ) ;
OR2     gate1337  (.A(g28612), .B(g18815), .Z(g29308) ) ;
DFF     gate1338  (.D(g29308), .CP(CLK), .Q(g6527) ) ;
OR2     gate1339  (.A(g25095), .B(g18816), .Z(g25762) ) ;
DFF     gate1340  (.D(g25762), .CP(CLK), .Q(g6533) ) ;
OR2     gate1341  (.A(g25113), .B(g18817), .Z(g25763) ) ;
DFF     gate1342  (.D(g25763), .CP(CLK), .Q(g6537) ) ;
OR2     gate1343  (.A(g34558), .B(g18820), .Z(g34647) ) ;
DFF     gate1344  (.D(g34647), .CP(CLK), .Q(g6545) ) ;
OR2     gate1345  (.A(g23439), .B(g18611), .Z(g24267) ) ;
DFF     gate1346  (.D(g24267), .CP(CLK), .Q(g3303) ) ;
DFF     gate1347  (.D(g3303), .CP(CLK), .Q(g3281) ) ;
DFF     gate1348  (.D(g3281), .CP(CLK), .Q(g3310) ) ;
DFF     gate1349  (.D(g3310), .CP(CLK), .Q(g3267) ) ;
DFF     gate1350  (.D(g3267), .CP(CLK), .Q(g3274) ) ;
DFF     gate1351  (.D(g3274), .CP(CLK), .Q(g3298) ) ;
DFF     gate1352  (.D(g3298), .CP(CLK), .Q(g3317) ) ;
DFF     gate1353  (.D(g3317), .CP(CLK), .Q(g3321) ) ;
DFF     gate1354  (.D(g3321), .CP(CLK), .Q(g3325) ) ;
DFF     gate1355  (.D(g3325), .CP(CLK), .Q(g3329) ) ;
OR2     gate1356  (.A(g23025), .B(g18612), .Z(g24268) ) ;
DFF     gate1357  (.D(g24268), .CP(CLK), .Q(g3338) ) ;
OR2     gate1358  (.A(g23131), .B(g18613), .Z(g24269) ) ;
DFF     gate1359  (.D(g24269), .CP(CLK), .Q(g3343) ) ;
OR2     gate1360  (.A(g23165), .B(g18614), .Z(g24270) ) ;
DFF     gate1361  (.D(g24270), .CP(CLK), .Q(g3347) ) ;
OR2     gate1362  (.A(g33239), .B(g18615), .Z(g33609) ) ;
DFF     gate1363  (.D(g33609), .CP(CLK), .Q(g3352) ) ;
OR2     gate1364  (.A(g33242), .B(g18616), .Z(g33610) ) ;
DFF     gate1365  (.D(g33610), .CP(CLK), .Q(g3288) ) ;
OR2     gate1366  (.A(g24644), .B(g21741), .Z(g25648) ) ;
DFF     gate1367  (.D(g25648), .CP(CLK), .Q(g3092) ) ;
DFF     gate1368  (.D(g3092), .CP(CLK), .Q(g3100) ) ;
OR2     gate1369  (.A(g24663), .B(g21743), .Z(g25650) ) ;
DFF     gate1370  (.D(g25650), .CP(CLK), .Q(g3050) ) ;
OR2     gate1371  (.A(g24654), .B(g21742), .Z(g25649) ) ;
DFF     gate1372  (.D(g25649), .CP(CLK), .Q(g3096) ) ;
DFF     gate1373  (.D(g3096), .CP(CLK), .Q(g3103) ) ;
OR2     gate1374  (.A(g24680), .B(g21744), .Z(g25651) ) ;
DFF     gate1375  (.D(g25651), .CP(CLK), .Q(g3010) ) ;
OR2     gate1376  (.A(g31270), .B(g21728), .Z(g31873) ) ;
DFF     gate1377  (.D(g31873), .CP(CLK), .Q(g3004) ) ;
OR2     gate1378  (.A(g31278), .B(g21732), .Z(g31877) ) ;
DFF     gate1379  (.D(g31877), .CP(CLK), .Q(g3017) ) ;
OR2     gate1380  (.A(g31475), .B(g21745), .Z(g31879) ) ;
DFF     gate1381  (.D(g31879), .CP(CLK), .Q(g3021) ) ;
OR2     gate1382  (.A(g31016), .B(g21729), .Z(g31874) ) ;
DFF     gate1383  (.D(g31874), .CP(CLK), .Q(g3025) ) ;
OR2     gate1384  (.A(g31066), .B(g21730), .Z(g31875) ) ;
DFF     gate1385  (.D(g31875), .CP(CLK), .Q(g3029) ) ;
OR2     gate1386  (.A(g31125), .B(g21731), .Z(g31876) ) ;
DFF     gate1387  (.D(g31876), .CP(CLK), .Q(g3034) ) ;
OR2     gate1388  (.A(g31015), .B(g21733), .Z(g31878) ) ;
DFF     gate1389  (.D(g31878), .CP(CLK), .Q(g3040) ) ;
OR2     gate1390  (.A(g32160), .B(g21734), .Z(g33020) ) ;
DFF     gate1391  (.D(g33020), .CP(CLK), .Q(g3045) ) ;
OR2     gate1392  (.A(g27288), .B(g21746), .Z(g28062) ) ;
DFF     gate1393  (.D(g28062), .CP(CLK), .Q(g3057) ) ;
OR2     gate1394  (.A(g27287), .B(g21735), .Z(g28061) ) ;
DFF     gate1395  (.D(g28061), .CP(CLK), .Q(g3061) ) ;
OR2     gate1396  (.A(g24777), .B(g21747), .Z(g25652) ) ;
DFF     gate1397  (.D(g25652), .CP(CLK), .Q(g3065) ) ;
OR2     gate1398  (.A(g24602), .B(g21736), .Z(g25643) ) ;
DFF     gate1399  (.D(g25643), .CP(CLK), .Q(g3068) ) ;
OR2     gate1400  (.A(g24622), .B(g21737), .Z(g25644) ) ;
DFF     gate1401  (.D(g25644), .CP(CLK), .Q(g3072) ) ;
OR2     gate1402  (.A(g24679), .B(g21738), .Z(g25645) ) ;
DFF     gate1403  (.D(g25645), .CP(CLK), .Q(g3080) ) ;
OR2     gate1404  (.A(g24706), .B(g21739), .Z(g25646) ) ;
DFF     gate1405  (.D(g25646), .CP(CLK), .Q(g3085) ) ;
OR2     gate1406  (.A(g24725), .B(g21740), .Z(g25647) ) ;
DFF     gate1407  (.D(g25647), .CP(CLK), .Q(g3089) ) ;
OR2     gate1408  (.A(g29986), .B(g21748), .Z(g30393) ) ;
DFF     gate1409  (.D(g30393), .CP(CLK), .Q(g3155) ) ;
OR2     gate1410  (.A(g32302), .B(g21749), .Z(g33021) ) ;
DFF     gate1411  (.D(g33021), .CP(CLK), .Q(g3161) ) ;
OR2     gate1412  (.A(g32306), .B(g21750), .Z(g33022) ) ;
DFF     gate1413  (.D(g33022), .CP(CLK), .Q(g3167) ) ;
OR2     gate1414  (.A(g32313), .B(g21751), .Z(g33023) ) ;
DFF     gate1415  (.D(g33023), .CP(CLK), .Q(g3171) ) ;
OR2     gate1416  (.A(g32324), .B(g21752), .Z(g33024) ) ;
DFF     gate1417  (.D(g33024), .CP(CLK), .Q(g3179) ) ;
OR2     gate1418  (.A(g29805), .B(g21753), .Z(g30394) ) ;
DFF     gate1419  (.D(g30394), .CP(CLK), .Q(g3187) ) ;
OR2     gate1420  (.A(g29749), .B(g21757), .Z(g30398) ) ;
DFF     gate1421  (.D(g30398), .CP(CLK), .Q(g3215) ) ;
OR2     gate1422  (.A(g29871), .B(g21761), .Z(g30402) ) ;
DFF     gate1423  (.D(g30402), .CP(CLK), .Q(g3231) ) ;
OR2     gate1424  (.A(g29783), .B(g21765), .Z(g30406) ) ;
DFF     gate1425  (.D(g30406), .CP(CLK), .Q(g3247) ) ;
OR2     gate1426  (.A(g29857), .B(g21769), .Z(g30410) ) ;
DFF     gate1427  (.D(g30410), .CP(CLK), .Q(g3195) ) ;
OR2     gate1428  (.A(g29841), .B(g21754), .Z(g30395) ) ;
DFF     gate1429  (.D(g30395), .CP(CLK), .Q(g3191) ) ;
OR2     gate1430  (.A(g29757), .B(g21758), .Z(g30399) ) ;
DFF     gate1431  (.D(g30399), .CP(CLK), .Q(g3219) ) ;
OR2     gate1432  (.A(g29750), .B(g21762), .Z(g30403) ) ;
DFF     gate1433  (.D(g30403), .CP(CLK), .Q(g3235) ) ;
OR2     gate1434  (.A(g29794), .B(g21766), .Z(g30407) ) ;
DFF     gate1435  (.D(g30407), .CP(CLK), .Q(g3251) ) ;
OR2     gate1436  (.A(g29872), .B(g21770), .Z(g30411) ) ;
DFF     gate1437  (.D(g30411), .CP(CLK), .Q(g3203) ) ;
OR2     gate1438  (.A(g29856), .B(g21755), .Z(g30396) ) ;
DFF     gate1439  (.D(g30396), .CP(CLK), .Q(g3199) ) ;
OR2     gate1440  (.A(g29766), .B(g21759), .Z(g30400) ) ;
DFF     gate1441  (.D(g30400), .CP(CLK), .Q(g3223) ) ;
OR2     gate1442  (.A(g29758), .B(g21763), .Z(g30404) ) ;
DFF     gate1443  (.D(g30404), .CP(CLK), .Q(g3239) ) ;
OR2     gate1444  (.A(g29806), .B(g21767), .Z(g30408) ) ;
DFF     gate1445  (.D(g30408), .CP(CLK), .Q(g3255) ) ;
OR2     gate1446  (.A(g29885), .B(g21771), .Z(g30412) ) ;
DFF     gate1447  (.D(g30412), .CP(CLK), .Q(g3211) ) ;
OR2     gate1448  (.A(g29747), .B(g21756), .Z(g30397) ) ;
DFF     gate1449  (.D(g30397), .CP(CLK), .Q(g3207) ) ;
OR2     gate1450  (.A(g29782), .B(g21760), .Z(g30401) ) ;
DFF     gate1451  (.D(g30401), .CP(CLK), .Q(g3227) ) ;
OR2     gate1452  (.A(g29767), .B(g21764), .Z(g30405) ) ;
DFF     gate1453  (.D(g30405), .CP(CLK), .Q(g3243) ) ;
OR2     gate1454  (.A(g29842), .B(g21768), .Z(g30409) ) ;
DFF     gate1455  (.D(g30409), .CP(CLK), .Q(g3259) ) ;
OR2     gate1456  (.A(g30001), .B(g21772), .Z(g30413) ) ;
DFF     gate1457  (.D(g30413), .CP(CLK), .Q(g3263) ) ;
OR2     gate1458  (.A(g27541), .B(g21773), .Z(g28063) ) ;
DFF     gate1459  (.D(g28063), .CP(CLK), .Q(g3333) ) ;
OR2     gate1460  (.A(g28327), .B(g18608), .Z(g29262) ) ;
DFF     gate1461  (.D(g29262), .CP(CLK), .Q(g3147) ) ;
OR2     gate1462  (.A(g24945), .B(g18609), .Z(g25656) ) ;
DFF     gate1463  (.D(g25656), .CP(CLK), .Q(g3111) ) ;
OR2     gate1464  (.A(g28228), .B(g18600), .Z(g29257) ) ;
DFF     gate1465  (.D(g29257), .CP(CLK), .Q(g3106) ) ;
OR2     gate1466  (.A(g28238), .B(g18601), .Z(g29258) ) ;
DFF     gate1467  (.D(g29258), .CP(CLK), .Q(g3115) ) ;
OR2     gate1468  (.A(g24664), .B(g18602), .Z(g25653) ) ;
DFF     gate1469  (.D(g25653), .CP(CLK), .Q(g3119) ) ;
OR2     gate1470  (.A(g28304), .B(g18603), .Z(g29259) ) ;
DFF     gate1471  (.D(g29259), .CP(CLK), .Q(g3125) ) ;
OR2     gate1472  (.A(g28315), .B(g18604), .Z(g29260) ) ;
DFF     gate1473  (.D(g29260), .CP(CLK), .Q(g3129) ) ;
OR2     gate1474  (.A(g28247), .B(g18605), .Z(g29261) ) ;
DFF     gate1475  (.D(g29261), .CP(CLK), .Q(g3133) ) ;
OR2     gate1476  (.A(g24634), .B(g18606), .Z(g25654) ) ;
DFF     gate1477  (.D(g25654), .CP(CLK), .Q(g3139) ) ;
OR2     gate1478  (.A(g24645), .B(g18607), .Z(g25655) ) ;
DFF     gate1479  (.D(g25655), .CP(CLK), .Q(g3143) ) ;
OR2     gate1480  (.A(g34532), .B(g18610), .Z(g34625) ) ;
DFF     gate1481  (.D(g34625), .CP(CLK), .Q(g3151) ) ;
OR2     gate1482  (.A(g23451), .B(g18628), .Z(g24271) ) ;
DFF     gate1483  (.D(g24271), .CP(CLK), .Q(g3654) ) ;
DFF     gate1484  (.D(g3654), .CP(CLK), .Q(g3632) ) ;
DFF     gate1485  (.D(g3632), .CP(CLK), .Q(g3661) ) ;
DFF     gate1486  (.D(g3661), .CP(CLK), .Q(g3618) ) ;
DFF     gate1487  (.D(g3618), .CP(CLK), .Q(g3625) ) ;
DFF     gate1488  (.D(g3625), .CP(CLK), .Q(g3649) ) ;
DFF     gate1489  (.D(g3649), .CP(CLK), .Q(g3668) ) ;
DFF     gate1490  (.D(g3668), .CP(CLK), .Q(g3672) ) ;
DFF     gate1491  (.D(g3672), .CP(CLK), .Q(g3676) ) ;
DFF     gate1492  (.D(g3676), .CP(CLK), .Q(g3680) ) ;
OR2     gate1493  (.A(g23056), .B(g18629), .Z(g24272) ) ;
DFF     gate1494  (.D(g24272), .CP(CLK), .Q(g3689) ) ;
OR2     gate1495  (.A(g23166), .B(g18630), .Z(g24273) ) ;
DFF     gate1496  (.D(g24273), .CP(CLK), .Q(g3694) ) ;
OR2     gate1497  (.A(g23187), .B(g18631), .Z(g24274) ) ;
DFF     gate1498  (.D(g24274), .CP(CLK), .Q(g3698) ) ;
OR2     gate1499  (.A(g33243), .B(g18632), .Z(g33611) ) ;
DFF     gate1500  (.D(g33611), .CP(CLK), .Q(g3703) ) ;
OR2     gate1501  (.A(g33247), .B(g18633), .Z(g33612) ) ;
DFF     gate1502  (.D(g33612), .CP(CLK), .Q(g3639) ) ;
OR2     gate1503  (.A(g24656), .B(g21787), .Z(g25662) ) ;
DFF     gate1504  (.D(g25662), .CP(CLK), .Q(g3443) ) ;
DFF     gate1505  (.D(g3443), .CP(CLK), .Q(g3451) ) ;
OR2     gate1506  (.A(g24681), .B(g21789), .Z(g25664) ) ;
DFF     gate1507  (.D(g25664), .CP(CLK), .Q(g3401) ) ;
OR2     gate1508  (.A(g24666), .B(g21788), .Z(g25663) ) ;
DFF     gate1509  (.D(g25663), .CP(CLK), .Q(g3447) ) ;
DFF     gate1510  (.D(g3447), .CP(CLK), .Q(g3454) ) ;
OR2     gate1511  (.A(g24708), .B(g21790), .Z(g25665) ) ;
DFF     gate1512  (.D(g25665), .CP(CLK), .Q(g3361) ) ;
OR2     gate1513  (.A(g31280), .B(g21774), .Z(g31880) ) ;
DFF     gate1514  (.D(g31880), .CP(CLK), .Q(g3355) ) ;
OR2     gate1515  (.A(g31290), .B(g21778), .Z(g31884) ) ;
DFF     gate1516  (.D(g31884), .CP(CLK), .Q(g3368) ) ;
OR2     gate1517  (.A(g31481), .B(g21791), .Z(g31886) ) ;
DFF     gate1518  (.D(g31886), .CP(CLK), .Q(g3372) ) ;
OR2     gate1519  (.A(g31018), .B(g21775), .Z(g31881) ) ;
DFF     gate1520  (.D(g31881), .CP(CLK), .Q(g3376) ) ;
OR2     gate1521  (.A(g31115), .B(g21776), .Z(g31882) ) ;
DFF     gate1522  (.D(g31882), .CP(CLK), .Q(g3380) ) ;
OR2     gate1523  (.A(g31132), .B(g21777), .Z(g31883) ) ;
DFF     gate1524  (.D(g31883), .CP(CLK), .Q(g3385) ) ;
OR2     gate1525  (.A(g31017), .B(g21779), .Z(g31885) ) ;
DFF     gate1526  (.D(g31885), .CP(CLK), .Q(g3391) ) ;
OR2     gate1527  (.A(g32162), .B(g21780), .Z(g33025) ) ;
DFF     gate1528  (.D(g33025), .CP(CLK), .Q(g3396) ) ;
OR2     gate1529  (.A(g27299), .B(g21792), .Z(g28065) ) ;
DFF     gate1530  (.D(g28065), .CP(CLK), .Q(g3408) ) ;
OR2     gate1531  (.A(g27298), .B(g21781), .Z(g28064) ) ;
DFF     gate1532  (.D(g28064), .CP(CLK), .Q(g3412) ) ;
OR2     gate1533  (.A(g24788), .B(g21793), .Z(g25666) ) ;
DFF     gate1534  (.D(g25666), .CP(CLK), .Q(g3416) ) ;
OR2     gate1535  (.A(g24624), .B(g21782), .Z(g25657) ) ;
DFF     gate1536  (.D(g25657), .CP(CLK), .Q(g3419) ) ;
OR2     gate1537  (.A(g24635), .B(g21783), .Z(g25658) ) ;
DFF     gate1538  (.D(g25658), .CP(CLK), .Q(g3423) ) ;
OR2     gate1539  (.A(g24707), .B(g21784), .Z(g25659) ) ;
DFF     gate1540  (.D(g25659), .CP(CLK), .Q(g3431) ) ;
OR2     gate1541  (.A(g24726), .B(g21785), .Z(g25660) ) ;
DFF     gate1542  (.D(g25660), .CP(CLK), .Q(g3436) ) ;
OR2     gate1543  (.A(g24754), .B(g21786), .Z(g25661) ) ;
DFF     gate1544  (.D(g25661), .CP(CLK), .Q(g3440) ) ;
OR2     gate1545  (.A(g30002), .B(g21794), .Z(g30414) ) ;
DFF     gate1546  (.D(g30414), .CP(CLK), .Q(g3506) ) ;
OR2     gate1547  (.A(g32307), .B(g21795), .Z(g33026) ) ;
DFF     gate1548  (.D(g33026), .CP(CLK), .Q(g3512) ) ;
OR2     gate1549  (.A(g32314), .B(g21796), .Z(g33027) ) ;
DFF     gate1550  (.D(g33027), .CP(CLK), .Q(g3518) ) ;
OR2     gate1551  (.A(g32325), .B(g21797), .Z(g33028) ) ;
DFF     gate1552  (.D(g33028), .CP(CLK), .Q(g3522) ) ;
OR2     gate1553  (.A(g32332), .B(g21798), .Z(g33029) ) ;
DFF     gate1554  (.D(g33029), .CP(CLK), .Q(g3530) ) ;
OR2     gate1555  (.A(g29843), .B(g21799), .Z(g30415) ) ;
DFF     gate1556  (.D(g30415), .CP(CLK), .Q(g3538) ) ;
OR2     gate1557  (.A(g29759), .B(g21803), .Z(g30419) ) ;
DFF     gate1558  (.D(g30419), .CP(CLK), .Q(g3566) ) ;
OR2     gate1559  (.A(g29887), .B(g21807), .Z(g30423) ) ;
DFF     gate1560  (.D(g30423), .CP(CLK), .Q(g3582) ) ;
OR2     gate1561  (.A(g29796), .B(g21811), .Z(g30427) ) ;
DFF     gate1562  (.D(g30427), .CP(CLK), .Q(g3598) ) ;
OR2     gate1563  (.A(g29875), .B(g21815), .Z(g30431) ) ;
DFF     gate1564  (.D(g30431), .CP(CLK), .Q(g3546) ) ;
OR2     gate1565  (.A(g29858), .B(g21800), .Z(g30416) ) ;
DFF     gate1566  (.D(g30416), .CP(CLK), .Q(g3542) ) ;
OR2     gate1567  (.A(g29769), .B(g21804), .Z(g30420) ) ;
DFF     gate1568  (.D(g30420), .CP(CLK), .Q(g3570) ) ;
OR2     gate1569  (.A(g29760), .B(g21808), .Z(g30424) ) ;
DFF     gate1570  (.D(g30424), .CP(CLK), .Q(g3586) ) ;
OR2     gate1571  (.A(g29807), .B(g21812), .Z(g30428) ) ;
DFF     gate1572  (.D(g30428), .CP(CLK), .Q(g3602) ) ;
OR2     gate1573  (.A(g29888), .B(g21816), .Z(g30432) ) ;
DFF     gate1574  (.D(g30432), .CP(CLK), .Q(g3554) ) ;
OR2     gate1575  (.A(g29874), .B(g21801), .Z(g30417) ) ;
DFF     gate1576  (.D(g30417), .CP(CLK), .Q(g3550) ) ;
OR2     gate1577  (.A(g29784), .B(g21805), .Z(g30421) ) ;
DFF     gate1578  (.D(g30421), .CP(CLK), .Q(g3574) ) ;
OR2     gate1579  (.A(g29770), .B(g21809), .Z(g30425) ) ;
DFF     gate1580  (.D(g30425), .CP(CLK), .Q(g3590) ) ;
OR2     gate1581  (.A(g29844), .B(g21813), .Z(g30429) ) ;
DFF     gate1582  (.D(g30429), .CP(CLK), .Q(g3606) ) ;
OR2     gate1583  (.A(g29899), .B(g21817), .Z(g30433) ) ;
DFF     gate1584  (.D(g30433), .CP(CLK), .Q(g3562) ) ;
OR2     gate1585  (.A(g29751), .B(g21802), .Z(g30418) ) ;
DFF     gate1586  (.D(g30418), .CP(CLK), .Q(g3558) ) ;
OR2     gate1587  (.A(g29795), .B(g21806), .Z(g30422) ) ;
DFF     gate1588  (.D(g30422), .CP(CLK), .Q(g3578) ) ;
OR2     gate1589  (.A(g29785), .B(g21810), .Z(g30426) ) ;
DFF     gate1590  (.D(g30426), .CP(CLK), .Q(g3594) ) ;
OR2     gate1591  (.A(g29859), .B(g21814), .Z(g30430) ) ;
DFF     gate1592  (.D(g30430), .CP(CLK), .Q(g3610) ) ;
OR2     gate1593  (.A(g30024), .B(g21818), .Z(g30434) ) ;
DFF     gate1594  (.D(g30434), .CP(CLK), .Q(g3614) ) ;
OR2     gate1595  (.A(g27553), .B(g21819), .Z(g28066) ) ;
DFF     gate1596  (.D(g28066), .CP(CLK), .Q(g3684) ) ;
OR2     gate1597  (.A(g28343), .B(g18625), .Z(g29268) ) ;
DFF     gate1598  (.D(g29268), .CP(CLK), .Q(g3498) ) ;
OR2     gate1599  (.A(g24967), .B(g18626), .Z(g25670) ) ;
DFF     gate1600  (.D(g25670), .CP(CLK), .Q(g3462) ) ;
OR2     gate1601  (.A(g28239), .B(g18617), .Z(g29263) ) ;
DFF     gate1602  (.D(g29263), .CP(CLK), .Q(g3457) ) ;
OR2     gate1603  (.A(g28248), .B(g18618), .Z(g29264) ) ;
DFF     gate1604  (.D(g29264), .CP(CLK), .Q(g3466) ) ;
OR2     gate1605  (.A(g24682), .B(g18619), .Z(g25667) ) ;
DFF     gate1606  (.D(g25667), .CP(CLK), .Q(g3470) ) ;
OR2     gate1607  (.A(g28318), .B(g18620), .Z(g29265) ) ;
DFF     gate1608  (.D(g29265), .CP(CLK), .Q(g3476) ) ;
OR2     gate1609  (.A(g28330), .B(g18621), .Z(g29266) ) ;
DFF     gate1610  (.D(g29266), .CP(CLK), .Q(g3480) ) ;
OR2     gate1611  (.A(g28257), .B(g18622), .Z(g29267) ) ;
DFF     gate1612  (.D(g29267), .CP(CLK), .Q(g3484) ) ;
OR2     gate1613  (.A(g24646), .B(g18623), .Z(g25668) ) ;
DFF     gate1614  (.D(g25668), .CP(CLK), .Q(g3490) ) ;
OR2     gate1615  (.A(g24657), .B(g18624), .Z(g25669) ) ;
DFF     gate1616  (.D(g25669), .CP(CLK), .Q(g3494) ) ;
OR2     gate1617  (.A(g34533), .B(g18627), .Z(g34626) ) ;
DFF     gate1618  (.D(g34626), .CP(CLK), .Q(g3502) ) ;
OR2     gate1619  (.A(g23474), .B(g18645), .Z(g24275) ) ;
DFF     gate1620  (.D(g24275), .CP(CLK), .Q(g4005) ) ;
DFF     gate1621  (.D(g4005), .CP(CLK), .Q(g3983) ) ;
DFF     gate1622  (.D(g3983), .CP(CLK), .Q(g4012) ) ;
DFF     gate1623  (.D(g4012), .CP(CLK), .Q(g3969) ) ;
DFF     gate1624  (.D(g3969), .CP(CLK), .Q(g3976) ) ;
DFF     gate1625  (.D(g3976), .CP(CLK), .Q(g4000) ) ;
DFF     gate1626  (.D(g4000), .CP(CLK), .Q(g4019) ) ;
DFF     gate1627  (.D(g4019), .CP(CLK), .Q(g4023) ) ;
DFF     gate1628  (.D(g4023), .CP(CLK), .Q(g4027) ) ;
DFF     gate1629  (.D(g4027), .CP(CLK), .Q(g4031) ) ;
OR2     gate1630  (.A(g23083), .B(g18646), .Z(g24276) ) ;
DFF     gate1631  (.D(g24276), .CP(CLK), .Q(g4040) ) ;
OR2     gate1632  (.A(g23188), .B(g18647), .Z(g24277) ) ;
DFF     gate1633  (.D(g24277), .CP(CLK), .Q(g4045) ) ;
OR2     gate1634  (.A(g23201), .B(g18648), .Z(g24278) ) ;
DFF     gate1635  (.D(g24278), .CP(CLK), .Q(g4049) ) ;
OR2     gate1636  (.A(g33248), .B(g18649), .Z(g33613) ) ;
DFF     gate1637  (.D(g33613), .CP(CLK), .Q(g4054) ) ;
OR2     gate1638  (.A(g33249), .B(g18650), .Z(g33614) ) ;
DFF     gate1639  (.D(g33614), .CP(CLK), .Q(g3990) ) ;
OR2     gate1640  (.A(g24668), .B(g21833), .Z(g25676) ) ;
DFF     gate1641  (.D(g25676), .CP(CLK), .Q(g3794) ) ;
DFF     gate1642  (.D(g3794), .CP(CLK), .Q(g3802) ) ;
OR2     gate1643  (.A(g24709), .B(g21835), .Z(g25678) ) ;
DFF     gate1644  (.D(g25678), .CP(CLK), .Q(g3752) ) ;
OR2     gate1645  (.A(g24684), .B(g21834), .Z(g25677) ) ;
DFF     gate1646  (.D(g25677), .CP(CLK), .Q(g3798) ) ;
DFF     gate1647  (.D(g3798), .CP(CLK), .Q(g3805) ) ;
OR2     gate1648  (.A(g24728), .B(g21836), .Z(g25679) ) ;
DFF     gate1649  (.D(g25679), .CP(CLK), .Q(g3712) ) ;
OR2     gate1650  (.A(g31292), .B(g21820), .Z(g31887) ) ;
DFF     gate1651  (.D(g31887), .CP(CLK), .Q(g3706) ) ;
OR2     gate1652  (.A(g31305), .B(g21824), .Z(g31891) ) ;
DFF     gate1653  (.D(g31891), .CP(CLK), .Q(g3719) ) ;
OR2     gate1654  (.A(g31490), .B(g21837), .Z(g31893) ) ;
DFF     gate1655  (.D(g31893), .CP(CLK), .Q(g3723) ) ;
OR2     gate1656  (.A(g31067), .B(g21821), .Z(g31888) ) ;
DFF     gate1657  (.D(g31888), .CP(CLK), .Q(g3727) ) ;
OR2     gate1658  (.A(g31118), .B(g21822), .Z(g31889) ) ;
DFF     gate1659  (.D(g31889), .CP(CLK), .Q(g3731) ) ;
OR2     gate1660  (.A(g31143), .B(g21823), .Z(g31890) ) ;
DFF     gate1661  (.D(g31890), .CP(CLK), .Q(g3736) ) ;
OR2     gate1662  (.A(g31019), .B(g21825), .Z(g31892) ) ;
DFF     gate1663  (.D(g31892), .CP(CLK), .Q(g3742) ) ;
OR2     gate1664  (.A(g32166), .B(g21826), .Z(g33030) ) ;
DFF     gate1665  (.D(g33030), .CP(CLK), .Q(g3747) ) ;
OR2     gate1666  (.A(g27310), .B(g21838), .Z(g28068) ) ;
DFF     gate1667  (.D(g28068), .CP(CLK), .Q(g3759) ) ;
OR2     gate1668  (.A(g27309), .B(g21827), .Z(g28067) ) ;
DFF     gate1669  (.D(g28067), .CP(CLK), .Q(g3763) ) ;
OR2     gate1670  (.A(g24794), .B(g21839), .Z(g25680) ) ;
DFF     gate1671  (.D(g25680), .CP(CLK), .Q(g3767) ) ;
OR2     gate1672  (.A(g24637), .B(g21828), .Z(g25671) ) ;
DFF     gate1673  (.D(g25671), .CP(CLK), .Q(g3770) ) ;
OR2     gate1674  (.A(g24647), .B(g21829), .Z(g25672) ) ;
DFF     gate1675  (.D(g25672), .CP(CLK), .Q(g3774) ) ;
OR2     gate1676  (.A(g24727), .B(g21830), .Z(g25673) ) ;
DFF     gate1677  (.D(g25673), .CP(CLK), .Q(g3782) ) ;
OR2     gate1678  (.A(g24755), .B(g21831), .Z(g25674) ) ;
DFF     gate1679  (.D(g25674), .CP(CLK), .Q(g3787) ) ;
OR2     gate1680  (.A(g24769), .B(g21832), .Z(g25675) ) ;
DFF     gate1681  (.D(g25675), .CP(CLK), .Q(g3791) ) ;
OR2     gate1682  (.A(g30025), .B(g21840), .Z(g30435) ) ;
DFF     gate1683  (.D(g30435), .CP(CLK), .Q(g3857) ) ;
OR2     gate1684  (.A(g32315), .B(g21841), .Z(g33031) ) ;
DFF     gate1685  (.D(g33031), .CP(CLK), .Q(g3863) ) ;
OR2     gate1686  (.A(g32326), .B(g21842), .Z(g33032) ) ;
DFF     gate1687  (.D(g33032), .CP(CLK), .Q(g3869) ) ;
OR2     gate1688  (.A(g32333), .B(g21843), .Z(g33033) ) ;
DFF     gate1689  (.D(g33033), .CP(CLK), .Q(g3873) ) ;
OR2     gate1690  (.A(g32340), .B(g21844), .Z(g33034) ) ;
DFF     gate1691  (.D(g33034), .CP(CLK), .Q(g3881) ) ;
OR2     gate1692  (.A(g29860), .B(g21845), .Z(g30436) ) ;
DFF     gate1693  (.D(g30436), .CP(CLK), .Q(g3889) ) ;
OR2     gate1694  (.A(g29771), .B(g21849), .Z(g30440) ) ;
DFF     gate1695  (.D(g30440), .CP(CLK), .Q(g3917) ) ;
OR2     gate1696  (.A(g29901), .B(g21853), .Z(g30444) ) ;
DFF     gate1697  (.D(g30444), .CP(CLK), .Q(g3933) ) ;
OR2     gate1698  (.A(g29809), .B(g21857), .Z(g30448) ) ;
DFF     gate1699  (.D(g30448), .CP(CLK), .Q(g3949) ) ;
OR2     gate1700  (.A(g29891), .B(g21861), .Z(g30452) ) ;
DFF     gate1701  (.D(g30452), .CP(CLK), .Q(g3897) ) ;
OR2     gate1702  (.A(g29876), .B(g21846), .Z(g30437) ) ;
DFF     gate1703  (.D(g30437), .CP(CLK), .Q(g3893) ) ;
OR2     gate1704  (.A(g29787), .B(g21850), .Z(g30441) ) ;
DFF     gate1705  (.D(g30441), .CP(CLK), .Q(g3921) ) ;
OR2     gate1706  (.A(g29772), .B(g21854), .Z(g30445) ) ;
DFF     gate1707  (.D(g30445), .CP(CLK), .Q(g3937) ) ;
OR2     gate1708  (.A(g29845), .B(g21858), .Z(g30449) ) ;
DFF     gate1709  (.D(g30449), .CP(CLK), .Q(g3953) ) ;
OR2     gate1710  (.A(g29902), .B(g21862), .Z(g30453) ) ;
DFF     gate1711  (.D(g30453), .CP(CLK), .Q(g3905) ) ;
OR2     gate1712  (.A(g29890), .B(g21847), .Z(g30438) ) ;
DFF     gate1713  (.D(g30438), .CP(CLK), .Q(g3901) ) ;
OR2     gate1714  (.A(g29797), .B(g21851), .Z(g30442) ) ;
DFF     gate1715  (.D(g30442), .CP(CLK), .Q(g3925) ) ;
OR2     gate1716  (.A(g29788), .B(g21855), .Z(g30446) ) ;
DFF     gate1717  (.D(g30446), .CP(CLK), .Q(g3941) ) ;
OR2     gate1718  (.A(g29861), .B(g21859), .Z(g30450) ) ;
DFF     gate1719  (.D(g30450), .CP(CLK), .Q(g3957) ) ;
OR2     gate1720  (.A(g29909), .B(g21863), .Z(g30454) ) ;
DFF     gate1721  (.D(g30454), .CP(CLK), .Q(g3913) ) ;
OR2     gate1722  (.A(g29761), .B(g21848), .Z(g30439) ) ;
DFF     gate1723  (.D(g30439), .CP(CLK), .Q(g3909) ) ;
OR2     gate1724  (.A(g29808), .B(g21852), .Z(g30443) ) ;
DFF     gate1725  (.D(g30443), .CP(CLK), .Q(g3929) ) ;
OR2     gate1726  (.A(g29798), .B(g21856), .Z(g30447) ) ;
DFF     gate1727  (.D(g30447), .CP(CLK), .Q(g3945) ) ;
OR2     gate1728  (.A(g29877), .B(g21860), .Z(g30451) ) ;
DFF     gate1729  (.D(g30451), .CP(CLK), .Q(g3961) ) ;
OR2     gate1730  (.A(g30041), .B(g21864), .Z(g30455) ) ;
DFF     gate1731  (.D(g30455), .CP(CLK), .Q(g3965) ) ;
OR2     gate1732  (.A(g27564), .B(g21865), .Z(g28069) ) ;
DFF     gate1733  (.D(g28069), .CP(CLK), .Q(g4035) ) ;
OR2     gate1734  (.A(g28360), .B(g18642), .Z(g29274) ) ;
DFF     gate1735  (.D(g29274), .CP(CLK), .Q(g3849) ) ;
OR2     gate1736  (.A(g24983), .B(g18643), .Z(g25684) ) ;
DFF     gate1737  (.D(g25684), .CP(CLK), .Q(g3813) ) ;
OR2     gate1738  (.A(g28249), .B(g18634), .Z(g29269) ) ;
DFF     gate1739  (.D(g29269), .CP(CLK), .Q(g3808) ) ;
OR2     gate1740  (.A(g28258), .B(g18635), .Z(g29270) ) ;
DFF     gate1741  (.D(g29270), .CP(CLK), .Q(g3817) ) ;
OR2     gate1742  (.A(g24710), .B(g18636), .Z(g25681) ) ;
DFF     gate1743  (.D(g25681), .CP(CLK), .Q(g3821) ) ;
OR2     gate1744  (.A(g28333), .B(g18637), .Z(g29271) ) ;
DFF     gate1745  (.D(g29271), .CP(CLK), .Q(g3827) ) ;
OR2     gate1746  (.A(g28346), .B(g18638), .Z(g29272) ) ;
DFF     gate1747  (.D(g29272), .CP(CLK), .Q(g3831) ) ;
OR2     gate1748  (.A(g28269), .B(g18639), .Z(g29273) ) ;
DFF     gate1749  (.D(g29273), .CP(CLK), .Q(g3835) ) ;
OR2     gate1750  (.A(g24658), .B(g18640), .Z(g25682) ) ;
DFF     gate1751  (.D(g25682), .CP(CLK), .Q(g3841) ) ;
OR2     gate1752  (.A(g24669), .B(g18641), .Z(g25683) ) ;
DFF     gate1753  (.D(g25683), .CP(CLK), .Q(g3845) ) ;
OR2     gate1754  (.A(g34534), .B(g18644), .Z(g34627) ) ;
DFF     gate1755  (.D(g34627), .CP(CLK), .Q(g3853) ) ;
INV     gate1756  (.A(II26578), .Z(g28079) ) ;
DFF     gate1757  (.D(g28079), .CP(CLK), .Q(g4165) ) ;
INV     gate1758  (.A(II26581), .Z(g28080) ) ;
DFF     gate1759  (.D(g28080), .CP(CLK), .Q(g4169) ) ;
INV     gate1760  (.A(II26584), .Z(g28081) ) ;
DFF     gate1761  (.D(g28081), .CP(CLK), .Q(g4125) ) ;
OR2     gate1762  (.A(g24536), .B(g21890), .Z(g25691) ) ;
DFF     gate1763  (.D(g25691), .CP(CLK), .Q(g4072) ) ;
OR2     gate1764  (.A(g24476), .B(g21866), .Z(g25685) ) ;
DFF     gate1765  (.D(g25685), .CP(CLK), .Q(g4064) ) ;
OR2     gate1766  (.A(g24712), .B(g21881), .Z(g25686) ) ;
DFF     gate1767  (.D(g25686), .CP(CLK), .Q(g4057) ) ;
OR2     gate1768  (.A(g24729), .B(g21882), .Z(g25687) ) ;
DFF     gate1769  (.D(g25687), .CP(CLK), .Q(g4141) ) ;
OR2     gate1770  (.A(g26186), .B(g21883), .Z(g26938) ) ;
DFF     gate1771  (.D(g26938), .CP(CLK), .Q(g4082) ) ;
OR2     gate1772  (.A(g27050), .B(g21867), .Z(g28070) ) ;
DFF     gate1773  (.D(g28070), .CP(CLK), .Q(g4076) ) ;
OR2     gate1774  (.A(g28165), .B(g21868), .Z(g29275) ) ;
DFF     gate1775  (.D(g29275), .CP(CLK), .Q(g4087) ) ;
OR2     gate1776  (.A(g29378), .B(g21869), .Z(g30456) ) ;
DFF     gate1777  (.D(g30456), .CP(CLK), .Q(g4093) ) ;
OR2     gate1778  (.A(g30671), .B(g21870), .Z(g31894) ) ;
DFF     gate1779  (.D(g31894), .CP(CLK), .Q(g4098) ) ;
OR2     gate1780  (.A(g32019), .B(g21872), .Z(g33035) ) ;
DFF     gate1781  (.D(g33035), .CP(CLK), .Q(g4108) ) ;
OR2     gate1782  (.A(g33113), .B(g21871), .Z(g33615) ) ;
DFF     gate1783  (.D(g33615), .CP(CLK), .Q(g4104) ) ;
OR2     gate1784  (.A(g25907), .B(g21884), .Z(g26939) ) ;
DFF     gate1785  (.D(g26939), .CP(CLK), .Q(g4145) ) ;
OR2     gate1786  (.A(g27085), .B(g21873), .Z(g28071) ) ;
DFF     gate1787  (.D(g28071), .CP(CLK), .Q(g4112) ) ;
OR2     gate1788  (.A(g27086), .B(g21874), .Z(g28072) ) ;
DFF     gate1789  (.D(g28072), .CP(CLK), .Q(g4116) ) ;
OR2     gate1790  (.A(g27097), .B(g21875), .Z(g28073) ) ;
DFF     gate1791  (.D(g28073), .CP(CLK), .Q(g4119) ) ;
OR2     gate1792  (.A(g27119), .B(g21876), .Z(g28074) ) ;
DFF     gate1793  (.D(g28074), .CP(CLK), .Q(g4122) ) ;
OR2     gate1794  (.A(g29369), .B(g21885), .Z(g30457) ) ;
DFF     gate1795  (.D(g30457), .CP(CLK), .Q(g4153) ) ;
OR2     gate1796  (.A(g25908), .B(g21886), .Z(g26940) ) ;
DFF     gate1797  (.D(g26940), .CP(CLK), .Q(g4164) ) ;
OR2     gate1798  (.A(g27083), .B(g21877), .Z(g28075) ) ;
DFF     gate1799  (.D(g28075), .CP(CLK), .Q(g4129) ) ;
OR2     gate1800  (.A(g27098), .B(g21878), .Z(g28076) ) ;
DFF     gate1801  (.D(g28076), .CP(CLK), .Q(g4132) ) ;
OR2     gate1802  (.A(g27120), .B(g21879), .Z(g28077) ) ;
DFF     gate1803  (.D(g28077), .CP(CLK), .Q(g4135) ) ;
OR2     gate1804  (.A(g27140), .B(g21880), .Z(g28078) ) ;
DFF     gate1805  (.D(g28078), .CP(CLK), .Q(g4138) ) ;
OR2     gate1806  (.A(g34678), .B(g18651), .Z(g34733) ) ;
DFF     gate1807  (.D(g34733), .CP(CLK), .Q(g4172) ) ;
OR2     gate1808  (.A(g34681), .B(g18652), .Z(g34734) ) ;
DFF     gate1809  (.D(g34734), .CP(CLK), .Q(g4176) ) ;
OR2     gate1810  (.A(g34493), .B(g18653), .Z(g34628) ) ;
DFF     gate1811  (.D(g34628), .CP(CLK), .Q(g4146) ) ;
OR2     gate1812  (.A(g34495), .B(g18654), .Z(g34629) ) ;
DFF     gate1813  (.D(g34629), .CP(CLK), .Q(g4157) ) ;
OR2     gate1814  (.A(g20094), .B(g18655), .Z(g21893) ) ;
DFF     gate1815  (.D(g21893), .CP(CLK), .Q(g4258) ) ;
OR2     gate1816  (.A(g20112), .B(g15107), .Z(g21894) ) ;
DFF     gate1817  (.D(g21894), .CP(CLK), .Q(g4264) ) ;
OR2     gate1818  (.A(g20135), .B(g15108), .Z(g21895) ) ;
DFF     gate1819  (.D(g21895), .CP(CLK), .Q(g4269) ) ;
OR2     gate1820  (.A(g23292), .B(g15109), .Z(g24280) ) ;
DFF     gate1821  (.D(g24280), .CP(CLK), .Q(g4273) ) ;
OR2     gate1822  (.A(g19788), .B(g15104), .Z(g21892) ) ;
DFF     gate1823  (.D(g21892), .CP(CLK), .Q(g4239) ) ;
OR2     gate1824  (.A(g20977), .B(g15114), .Z(g21900) ) ;
DFF     gate1825  (.D(g21900), .CP(CLK), .Q(g4294) ) ;
DFF     gate1826  (.D(g4294), .CP(CLK), .Q(g4297) ) ;
OR2     gate1827  (.A(g34709), .B(g15116), .Z(g34735) ) ;
DFF     gate1828  (.D(g34735), .CP(CLK), .Q(g4300) ) ;
OR2     gate1829  (.A(g34560), .B(g15117), .Z(g34630) ) ;
DFF     gate1830  (.D(g34630), .CP(CLK), .Q(g4253) ) ;
OR2     gate1831  (.A(g34562), .B(g15118), .Z(g34631) ) ;
DFF     gate1832  (.D(g34631), .CP(CLK), .Q(g4249) ) ;
OR2     gate1833  (.A(g34565), .B(g15119), .Z(g34632) ) ;
DFF     gate1834  (.D(g34632), .CP(CLK), .Q(g4245) ) ;
OR2     gate1835  (.A(g20084), .B(g15110), .Z(g21896) ) ;
DFF     gate1836  (.D(g21896), .CP(CLK), .Q(g4277) ) ;
DFF     gate1837  (.D(g4277), .CP(CLK), .Q(g4281) ) ;
OR2     gate1838  (.A(g20095), .B(g15111), .Z(g21897) ) ;
DFF     gate1839  (.D(g21897), .CP(CLK), .Q(g4284) ) ;
OR2     gate1840  (.A(g20152), .B(g15112), .Z(g21898) ) ;
DFF     gate1841  (.D(g21898), .CP(CLK), .Q(g4287) ) ;
DFF     gate1842  (.D(g4287), .CP(CLK), .Q(g4291) ) ;
OR2     gate1843  (.A(g20162), .B(g15113), .Z(g21899) ) ;
DFF     gate1844  (.D(g21899), .CP(CLK), .Q(g2946) ) ;
OR2     gate1845  (.A(g21251), .B(g15115), .Z(g21901) ) ;
DFF     gate1846  (.D(g21901), .CP(CLK), .Q(g4191) ) ;
DFF     gate1847  (.D(g4191), .CP(CLK), .Q(g4188) ) ;
DFF     gate1848  (.D(g4188), .CP(CLK), .Q(g4194) ) ;
DFF     gate1849  (.D(g4194), .CP(CLK), .Q(g4197) ) ;
DFF     gate1850  (.D(g4197), .CP(CLK), .Q(g4200) ) ;
DFF     gate1851  (.D(g4200), .CP(CLK), .Q(g4204) ) ;
DFF     gate1852  (.D(g4204), .CP(CLK), .Q(g4207) ) ;
DFF     gate1853  (.D(g4207), .CP(CLK), .Q(g4210) ) ;
DFF     gate1854  (.D(g4210), .CP(CLK), .Q(g4180) ) ;
OR2     gate1855  (.A(g19948), .B(g15103), .Z(g21891) ) ;
DFF     gate1856  (.D(g21891), .CP(CLK), .Q(g4185) ) ;
DFF     gate1857  (.D(g4185), .CP(CLK), .Q(g4213) ) ;
DFF     gate1858  (.D(g4213), .CP(CLK), .Q(g4216) ) ;
DFF     gate1859  (.D(g4216), .CP(CLK), .Q(g4219) ) ;
DFF     gate1860  (.D(g4219), .CP(CLK), .Q(g4222) ) ;
DFF     gate1861  (.D(g4222), .CP(CLK), .Q(g4226) ) ;
DFF     gate1862  (.D(g4226), .CP(CLK), .Q(g4229) ) ;
DFF     gate1863  (.D(g4229), .CP(CLK), .Q(g4232) ) ;
DFF     gate1864  (.D(g4232), .CP(CLK), .Q(g4235) ) ;
OR2     gate1865  (.A(g23218), .B(g15105), .Z(g24279) ) ;
DFF     gate1866  (.D(g24279), .CP(CLK), .Q(g4242) ) ;
OR2     gate1867  (.A(g26610), .B(g24186), .Z(g26880) ) ;
DFF     gate1868  (.D(g26880), .CP(CLK), .Q(g305) ) ;
OR2     gate1869  (.A(g26629), .B(g24187), .Z(g26881) ) ;
DFF     gate1870  (.D(g26881), .CP(CLK), .Q(g311) ) ;
OR2     gate1871  (.A(g26651), .B(g24192), .Z(g26886) ) ;
DFF     gate1872  (.D(g26886), .CP(CLK), .Q(g336) ) ;
OR2     gate1873  (.A(g26542), .B(g24193), .Z(g26887) ) ;
DFF     gate1874  (.D(g26887), .CP(CLK), .Q(g324) ) ;
OR2     gate1875  (.A(g26670), .B(g24189), .Z(g26883) ) ;
DFF     gate1876  (.D(g26883), .CP(CLK), .Q(g316) ) ;
OR2     gate1877  (.A(g26650), .B(g24188), .Z(g26882) ) ;
DFF     gate1878  (.D(g26882), .CP(CLK), .Q(g319) ) ;
OR2     gate1879  (.A(g26541), .B(g24191), .Z(g26885) ) ;
DFF     gate1880  (.D(g26885), .CP(CLK), .Q(g329) ) ;
OR2     gate1881  (.A(g26511), .B(g24190), .Z(g26884) ) ;
DFF     gate1882  (.D(g26884), .CP(CLK), .Q(g333) ) ;
OR2     gate1883  (.A(g26630), .B(g24196), .Z(g26890) ) ;
DFF     gate1884  (.D(g26890), .CP(CLK), .Q(g344) ) ;
DFF     gate1885  (.D(g344), .CP(CLK), .Q(g347) ) ;
OR2     gate1886  (.A(g26652), .B(g24197), .Z(g26891) ) ;
DFF     gate1887  (.D(g26891), .CP(CLK), .Q(g351) ) ;
OR2     gate1888  (.A(g26719), .B(g24198), .Z(g26892) ) ;
DFF     gate1889  (.D(g26892), .CP(CLK), .Q(g355) ) ;
OR2     gate1890  (.A(g26753), .B(g24199), .Z(g26893) ) ;
DFF     gate1891  (.D(g26893), .CP(CLK), .Q(g74) ) ;
OR2     gate1892  (.A(g26689), .B(g24195), .Z(g26889) ) ;
DFF     gate1893  (.D(g26889), .CP(CLK), .Q(g106) ) ;
OR2     gate1894  (.A(g26671), .B(g24194), .Z(g26888) ) ;
DFF     gate1895  (.D(g26888), .CP(CLK), .Q(g341) ) ;
OR2     gate1896  (.A(g23280), .B(g18155), .Z(g24212) ) ;
DFF     gate1897  (.D(g24212), .CP(CLK), .Q(g637) ) ;
DFF     gate1898  (.D(g637), .CP(CLK), .Q(g640) ) ;
DFF     gate1899  (.D(g640), .CP(CLK), .Q(g559) ) ;
OR2     gate1900  (.A(g25181), .B(g18140), .Z(g25613) ) ;
DFF     gate1901  (.D(g25613), .CP(CLK), .Q(g562) ) ;
OR2     gate1902  (.A(g26783), .B(g18148), .Z(g26895) ) ;
DFF     gate1903  (.D(g26895), .CP(CLK), .Q(g568) ) ;
OR2     gate1904  (.A(g27378), .B(g18141), .Z(g28045) ) ;
DFF     gate1905  (.D(g28045), .CP(CLK), .Q(g572) ) ;
OR2     gate1906  (.A(g28919), .B(g18156), .Z(g29224) ) ;
DFF     gate1907  (.D(g29224), .CP(CLK), .Q(g586) ) ;
OR2     gate1908  (.A(g29837), .B(g18143), .Z(g30334) ) ;
DFF     gate1909  (.D(g30334), .CP(CLK), .Q(g577) ) ;
OR2     gate1910  (.A(g31252), .B(g18142), .Z(g31866) ) ;
DFF     gate1911  (.D(g31866), .CP(CLK), .Q(g582) ) ;
OR2     gate1912  (.A(g32197), .B(g18145), .Z(g32978) ) ;
DFF     gate1913  (.D(g32978), .CP(CLK), .Q(g590) ) ;
OR2     gate1914  (.A(g33252), .B(g18144), .Z(g33538) ) ;
DFF     gate1915  (.D(g33538), .CP(CLK), .Q(g595) ) ;
OR2     gate1916  (.A(g33817), .B(g18146), .Z(g33964) ) ;
DFF     gate1917  (.D(g33964), .CP(CLK), .Q(g599) ) ;
OR2     gate1918  (.A(g34157), .B(g18147), .Z(g34251) ) ;
DFF     gate1919  (.D(g34251), .CP(CLK), .Q(g604) ) ;
OR2     gate1920  (.A(g34348), .B(g18150), .Z(g34438) ) ;
DFF     gate1921  (.D(g34438), .CP(CLK), .Q(g608) ) ;
OR2     gate1922  (.A(g34542), .B(g18149), .Z(g34599) ) ;
DFF     gate1923  (.D(g34599), .CP(CLK), .Q(g613) ) ;
OR2     gate1924  (.A(g34702), .B(g18152), .Z(g34724) ) ;
DFF     gate1925  (.D(g34724), .CP(CLK), .Q(g617) ) ;
OR2     gate1926  (.A(g34774), .B(g18151), .Z(g34790) ) ;
DFF     gate1927  (.D(g34790), .CP(CLK), .Q(g622) ) ;
OR2     gate1928  (.A(g34842), .B(g18154), .Z(g34849) ) ;
DFF     gate1929  (.D(g34849), .CP(CLK), .Q(g626) ) ;
OR2     gate1930  (.A(g34867), .B(g18153), .Z(g34880) ) ;
DFF     gate1931  (.D(g34880), .CP(CLK), .Q(g632) ) ;
OR2     gate1932  (.A(g26819), .B(g24217), .Z(g26900) ) ;
DFF     gate1933  (.D(g26900), .CP(CLK), .Q(g859) ) ;
DFF     gate1934  (.D(g859), .CP(CLK), .Q(g869) ) ;
DFF     gate1935  (.D(g869), .CP(CLK), .Q(g875) ) ;
DFF     gate1936  (.D(g875), .CP(CLK), .Q(g878) ) ;
DFF     gate1937  (.D(g878), .CP(CLK), .Q(g881) ) ;
DFF     gate1938  (.D(g881), .CP(CLK), .Q(g884) ) ;
DFF     gate1939  (.D(g884), .CP(CLK), .Q(g887) ) ;
DFF     gate1940  (.D(g887), .CP(CLK), .Q(g872) ) ;
OR2     gate1941  (.A(g26362), .B(g24218), .Z(g26901) ) ;
DFF     gate1942  (.D(g26901), .CP(CLK), .Q(g225) ) ;
OR2     gate1943  (.A(g26378), .B(g24219), .Z(g26902) ) ;
DFF     gate1944  (.D(g26902), .CP(CLK), .Q(g255) ) ;
OR2     gate1945  (.A(g26388), .B(g24220), .Z(g26903) ) ;
DFF     gate1946  (.D(g26903), .CP(CLK), .Q(g232) ) ;
OR2     gate1947  (.A(g26393), .B(g24221), .Z(g26904) ) ;
DFF     gate1948  (.D(g26904), .CP(CLK), .Q(g262) ) ;
OR2     gate1949  (.A(g26397), .B(g24222), .Z(g26905) ) ;
DFF     gate1950  (.D(g26905), .CP(CLK), .Q(g239) ) ;
OR2     gate1951  (.A(g26423), .B(g24223), .Z(g26906) ) ;
DFF     gate1952  (.D(g26906), .CP(CLK), .Q(g269) ) ;
OR2     gate1953  (.A(g26513), .B(g24224), .Z(g26907) ) ;
DFF     gate1954  (.D(g26907), .CP(CLK), .Q(g246) ) ;
OR2     gate1955  (.A(g26358), .B(g24225), .Z(g26908) ) ;
DFF     gate1956  (.D(g26908), .CP(CLK), .Q(g446) ) ;
OR2     gate1957  (.A(g34364), .B(g24226), .Z(g34440) ) ;
DFF     gate1958  (.D(g34440), .CP(CLK), .Q(g890) ) ;
OR2     gate1959  (.A(g26543), .B(g24227), .Z(g26909) ) ;
DFF     gate1960  (.D(g26909), .CP(CLK), .Q(g862) ) ;
OR2     gate1961  (.A(g26571), .B(g24228), .Z(g26910) ) ;
DFF     gate1962  (.D(g26910), .CP(CLK), .Q(g896) ) ;
INV     gate1963  (.A(II24759), .Z(g25620) ) ;
DFF     gate1964  (.D(g25620), .CP(CLK), .Q(g901) ) ;
OR2     gate1965  (.A(g26612), .B(g24230), .Z(g26911) ) ;
DFF     gate1966  (.D(g26911), .CP(CLK), .Q(g391) ) ;
OR2     gate1967  (.A(g24835), .B(g21717), .Z(g25595) ) ;
DFF     gate1968  (.D(g25595), .CP(CLK), .Q(g365) ) ;
DFF     gate1969  (.D(g365), .CP(CLK), .Q(g358) ) ;
OR2     gate1970  (.A(g24892), .B(g21719), .Z(g25597) ) ;
DFF     gate1971  (.D(g25597), .CP(CLK), .Q(g370) ) ;
OR2     gate1972  (.A(g24865), .B(g21718), .Z(g25596) ) ;
DFF     gate1973  (.D(g25596), .CP(CLK), .Q(g376) ) ;
OR2     gate1974  (.A(g24904), .B(g21720), .Z(g25598) ) ;
DFF     gate1975  (.D(g25598), .CP(CLK), .Q(g385) ) ;
OR2     gate1976  (.A(g24914), .B(g21721), .Z(g25599) ) ;
DFF     gate1977  (.D(g25599), .CP(CLK), .Q(g203) ) ;
OR2     gate1978  (.A(g32254), .B(g18198), .Z(g32980) ) ;
DFF     gate1979  (.D(g32980), .CP(CLK), .Q(g854) ) ;
OR2     gate1980  (.A(g23416), .B(g18197), .Z(g24216) ) ;
DFF     gate1981  (.D(g24216), .CP(CLK), .Q(g847) ) ;
OR2     gate1982  (.A(g23471), .B(g18195), .Z(g24214) ) ;
DFF     gate1983  (.D(g24214), .CP(CLK), .Q(g703) ) ;
OR2     gate1984  (.A(g23484), .B(g18196), .Z(g24215) ) ;
DFF     gate1985  (.D(g24215), .CP(CLK), .Q(g837) ) ;
OR2     gate1986  (.A(g24961), .B(g18193), .Z(g25619) ) ;
DFF     gate1987  (.D(g25619), .CP(CLK), .Q(g843) ) ;
OR2     gate1988  (.A(g26387), .B(g18194), .Z(g26898) ) ;
DFF     gate1989  (.D(g26898), .CP(CLK), .Q(g812) ) ;
OR2     gate1990  (.A(g25466), .B(g18189), .Z(g25617) ) ;
DFF     gate1991  (.D(g25617), .CP(CLK), .Q(g817) ) ;
OR2     gate1992  (.A(g25491), .B(g18192), .Z(g25618) ) ;
DFF     gate1993  (.D(g25618), .CP(CLK), .Q(g832) ) ;
OR2     gate1994  (.A(g26844), .B(g18199), .Z(g26899) ) ;
DFF     gate1995  (.D(g26899), .CP(CLK), .Q(g822) ) ;
OR2     gate1996  (.A(g27560), .B(g18190), .Z(g28055) ) ;
DFF     gate1997  (.D(g28055), .CP(CLK), .Q(g827) ) ;
OR2     gate1998  (.A(g28532), .B(g18191), .Z(g29229) ) ;
DFF     gate1999  (.D(g29229), .CP(CLK), .Q(g723) ) ;
OR2     gate2000  (.A(g27667), .B(g18157), .Z(g28046) ) ;
DFF     gate2001  (.D(g28046), .CP(CLK), .Q(g645) ) ;
OR2     gate2002  (.A(g27676), .B(g18160), .Z(g28047) ) ;
DFF     gate2003  (.D(g28047), .CP(CLK), .Q(g681) ) ;
OR2     gate2004  (.A(g27393), .B(g18168), .Z(g28053) ) ;
DFF     gate2005  (.D(g28053), .CP(CLK), .Q(g699) ) ;
OR2     gate2006  (.A(g27684), .B(g18164), .Z(g28049) ) ;
DFF     gate2007  (.D(g28049), .CP(CLK), .Q(g650) ) ;
OR2     gate2008  (.A(g27692), .B(g18165), .Z(g28050) ) ;
DFF     gate2009  (.D(g28050), .CP(CLK), .Q(g655) ) ;
OR2     gate2010  (.A(g27699), .B(g18166), .Z(g28051) ) ;
DFF     gate2011  (.D(g28051), .CP(CLK), .Q(g718) ) ;
OR2     gate2012  (.A(g27710), .B(g18167), .Z(g28052) ) ;
DFF     gate2013  (.D(g28052), .CP(CLK), .Q(g661) ) ;
OR2     gate2014  (.A(g27723), .B(g18170), .Z(g28054) ) ;
DFF     gate2015  (.D(g28054), .CP(CLK), .Q(g728) ) ;
OR2     gate2016  (.A(g26341), .B(g18171), .Z(g26896) ) ;
DFF     gate2017  (.D(g26896), .CP(CLK), .Q(g79) ) ;
OR2     gate2018  (.A(g27362), .B(g18163), .Z(g28048) ) ;
DFF     gate2019  (.D(g28048), .CP(CLK), .Q(g691) ) ;
OR2     gate2020  (.A(g24797), .B(g18161), .Z(g25614) ) ;
DFF     gate2021  (.D(g25614), .CP(CLK), .Q(g686) ) ;
OR2     gate2022  (.A(g24803), .B(g18162), .Z(g25615) ) ;
DFF     gate2023  (.D(g25615), .CP(CLK), .Q(g667) ) ;
OR2     gate2024  (.A(g28451), .B(g18158), .Z(g29225) ) ;
DFF     gate2025  (.D(g29225), .CP(CLK), .Q(g671) ) ;
OR2     gate2026  (.A(g28455), .B(g18159), .Z(g29226) ) ;
DFF     gate2027  (.D(g29226), .CP(CLK), .Q(g676) ) ;
OR2     gate2028  (.A(g28456), .B(g18169), .Z(g29227) ) ;
DFF     gate2029  (.D(g29227), .CP(CLK), .Q(g714) ) ;
OR2     gate2030  (.A(g24915), .B(g18126), .Z(g25609) ) ;
DFF     gate2031  (.D(g25609), .CP(CLK), .Q(g499) ) ;
OR2     gate2032  (.A(g24923), .B(g18127), .Z(g25610) ) ;
DFF     gate2033  (.D(g25610), .CP(CLK), .Q(g504) ) ;
OR2     gate2034  (.A(g24931), .B(g18128), .Z(g25611) ) ;
DFF     gate2035  (.D(g25611), .CP(CLK), .Q(g513) ) ;
OR2     gate2036  (.A(g24941), .B(g18132), .Z(g25612) ) ;
DFF     gate2037  (.D(g25612), .CP(CLK), .Q(g518) ) ;
OR2     gate2038  (.A(g25979), .B(g18129), .Z(g26894) ) ;
DFF     gate2039  (.D(g26894), .CP(CLK), .Q(g528) ) ;
OR2     gate2040  (.A(g27256), .B(g18130), .Z(g28044) ) ;
DFF     gate2041  (.D(g28044), .CP(CLK), .Q(g482) ) ;
OR2     gate2042  (.A(g28341), .B(g18131), .Z(g29223) ) ;
DFF     gate2043  (.D(g29223), .CP(CLK), .Q(g490) ) ;
OR2     gate2044  (.A(g23415), .B(g18122), .Z(g24209) ) ;
DFF     gate2045  (.D(g24209), .CP(CLK), .Q(g417) ) ;
OR2     gate2046  (.A(g28252), .B(g18105), .Z(g29222) ) ;
DFF     gate2047  (.D(g29222), .CP(CLK), .Q(g411) ) ;
OR2     gate2048  (.A(g22899), .B(g18106), .Z(g24202) ) ;
DFF     gate2049  (.D(g24202), .CP(CLK), .Q(g424) ) ;
OR2     gate2050  (.A(g23404), .B(g18121), .Z(g24208) ) ;
DFF     gate2051  (.D(g24208), .CP(CLK), .Q(g475) ) ;
OR2     gate2052  (.A(g23396), .B(g18119), .Z(g24207) ) ;
DFF     gate2053  (.D(g24207), .CP(CLK), .Q(g441) ) ;
OR2     gate2054  (.A(g23386), .B(g18110), .Z(g24206) ) ;
DFF     gate2055  (.D(g24206), .CP(CLK), .Q(g437) ) ;
OR2     gate2056  (.A(g23006), .B(g18109), .Z(g24205) ) ;
DFF     gate2057  (.D(g24205), .CP(CLK), .Q(g433) ) ;
OR2     gate2058  (.A(g22990), .B(g18108), .Z(g24204) ) ;
DFF     gate2059  (.D(g24204), .CP(CLK), .Q(g429) ) ;
OR2     gate2060  (.A(g22982), .B(g18107), .Z(g24203) ) ;
DFF     gate2061  (.D(g24203), .CP(CLK), .Q(g401) ) ;
OR2     gate2062  (.A(g22831), .B(g18103), .Z(g24200) ) ;
DFF     gate2063  (.D(g24200), .CP(CLK), .Q(g392) ) ;
OR2     gate2064  (.A(g22848), .B(g18104), .Z(g24201) ) ;
DFF     gate2065  (.D(g24201), .CP(CLK), .Q(g405) ) ;
OR2     gate2066  (.A(g24673), .B(g18113), .Z(g25602) ) ;
DFF     gate2067  (.D(g25602), .CP(CLK), .Q(g182) ) ;
OR2     gate2068  (.A(g24660), .B(g18112), .Z(g25601) ) ;
DFF     gate2069  (.D(g25601), .CP(CLK), .Q(g174) ) ;
OR2     gate2070  (.A(g24650), .B(g18111), .Z(g25600) ) ;
DFF     gate2071  (.D(g25600), .CP(CLK), .Q(g168) ) ;
OR2     gate2072  (.A(g24743), .B(g18116), .Z(g25605) ) ;
DFF     gate2073  (.D(g25605), .CP(CLK), .Q(g460) ) ;
OR2     gate2074  (.A(g24717), .B(g18115), .Z(g25604) ) ;
DFF     gate2075  (.D(g25604), .CP(CLK), .Q(g452) ) ;
OR2     gate2076  (.A(g24698), .B(g18114), .Z(g25603) ) ;
DFF     gate2077  (.D(g25603), .CP(CLK), .Q(g457) ) ;
OR2     gate2078  (.A(g24643), .B(g18120), .Z(g25608) ) ;
DFF     gate2079  (.D(g25608), .CP(CLK), .Q(g471) ) ;
OR2     gate2080  (.A(g24773), .B(g18118), .Z(g25607) ) ;
DFF     gate2081  (.D(g25607), .CP(CLK), .Q(g464) ) ;
OR2     gate2082  (.A(g24761), .B(g18117), .Z(g25606) ) ;
DFF     gate2083  (.D(g25606), .CP(CLK), .Q(g468) ) ;
OR2     gate2084  (.A(g22900), .B(g18125), .Z(g24210) ) ;
DFF     gate2085  (.D(g24210), .CP(CLK), .Q(g479) ) ;
OR2     gate2086  (.A(g33822), .B(g18123), .Z(g33962) ) ;
DFF     gate2087  (.D(g33962), .CP(CLK), .Q(g102) ) ;
OR2     gate2088  (.A(g33830), .B(g18124), .Z(g33963) ) ;
DFF     gate2089  (.D(g33963), .CP(CLK), .Q(g496) ) ;
OR2     gate2090  (.A(g25096), .B(g18172), .Z(g25616) ) ;
DFF     gate2091  (.D(g25616), .CP(CLK), .Q(g732) ) ;
OR2     gate2092  (.A(g26611), .B(g18176), .Z(g26897) ) ;
DFF     gate2093  (.D(g26897), .CP(CLK), .Q(g753) ) ;
OR2     gate2094  (.A(g23220), .B(g18186), .Z(g24213) ) ;
DFF     gate2095  (.D(g24213), .CP(CLK), .Q(g799) ) ;
DFF     gate2096  (.D(g799), .CP(CLK), .Q(g802) ) ;
DFF     gate2097  (.D(g802), .CP(CLK), .Q(g736) ) ;
OR2     gate2098  (.A(g28426), .B(g18173), .Z(g29228) ) ;
DFF     gate2099  (.D(g29228), .CP(CLK), .Q(g739) ) ;
OR2     gate2100  (.A(g29746), .B(g18174), .Z(g30335) ) ;
DFF     gate2101  (.D(g30335), .CP(CLK), .Q(g744) ) ;
OR2     gate2102  (.A(g31238), .B(g18175), .Z(g31867) ) ;
DFF     gate2103  (.D(g31867), .CP(CLK), .Q(g749) ) ;
OR2     gate2104  (.A(g32181), .B(g18177), .Z(g32979) ) ;
DFF     gate2105  (.D(g32979), .CP(CLK), .Q(g758) ) ;
OR2     gate2106  (.A(g33245), .B(g18178), .Z(g33539) ) ;
DFF     gate2107  (.D(g33539), .CP(CLK), .Q(g763) ) ;
OR2     gate2108  (.A(g33805), .B(g18179), .Z(g33965) ) ;
DFF     gate2109  (.D(g33965), .CP(CLK), .Q(g767) ) ;
OR2     gate2110  (.A(g34146), .B(g18180), .Z(g34252) ) ;
DFF     gate2111  (.D(g34252), .CP(CLK), .Q(g772) ) ;
OR2     gate2112  (.A(g34344), .B(g18181), .Z(g34439) ) ;
DFF     gate2113  (.D(g34439), .CP(CLK), .Q(g776) ) ;
OR2     gate2114  (.A(g34538), .B(g18182), .Z(g34600) ) ;
DFF     gate2115  (.D(g34600), .CP(CLK), .Q(g781) ) ;
OR2     gate2116  (.A(g34700), .B(g18183), .Z(g34725) ) ;
DFF     gate2117  (.D(g34725), .CP(CLK), .Q(g785) ) ;
OR2     gate2118  (.A(g34771), .B(g18184), .Z(g34791) ) ;
DFF     gate2119  (.D(g34791), .CP(CLK), .Q(g790) ) ;
OR2     gate2120  (.A(g34841), .B(g18185), .Z(g34850) ) ;
DFF     gate2121  (.D(g34850), .CP(CLK), .Q(g794) ) ;
OR2     gate2122  (.A(g34866), .B(g18187), .Z(g34881) ) ;
DFF     gate2123  (.D(g34881), .CP(CLK), .Q(g807) ) ;
OR2     gate2124  (.A(g34909), .B(g18188), .Z(g34911) ) ;
DFF     gate2125  (.D(g34911), .CP(CLK), .Q(g554) ) ;
OR2     gate2126  (.A(g34701), .B(g18133), .Z(g34719) ) ;
DFF     gate2127  (.D(g34719), .CP(CLK), .Q(g538) ) ;
OR2     gate2128  (.A(g34707), .B(g18137), .Z(g34722) ) ;
DFF     gate2129  (.D(g34722), .CP(CLK), .Q(g546) ) ;
OR2     gate2130  (.A(g23572), .B(g18138), .Z(g24211) ) ;
DFF     gate2131  (.D(g24211), .CP(CLK), .Q(g542) ) ;
OR2     gate2132  (.A(g34710), .B(g18139), .Z(g34723) ) ;
DFF     gate2133  (.D(g34723), .CP(CLK), .Q(g534) ) ;
OR2     gate2134  (.A(g34694), .B(g18134), .Z(g34720) ) ;
DFF     gate2135  (.D(g34720), .CP(CLK), .Q(g550) ) ;
OR2     gate2136  (.A(g34541), .B(g18136), .Z(g34598) ) ;
DFF     gate2137  (.D(g34598), .CP(CLK), .Q(g136) ) ;
OR2     gate2138  (.A(g34696), .B(g18135), .Z(g34721) ) ;
DFF     gate2139  (.D(g34721), .CP(CLK), .Q(g199) ) ;
OR2     gate2140  (.A(g24772), .B(g21708), .Z(g25594) ) ;
DFF     gate2141  (.D(g25594), .CP(CLK), .Q(g278) ) ;
OR2     gate2142  (.A(g27323), .B(g21714), .Z(g28043) ) ;
DFF     gate2143  (.D(g28043), .CP(CLK), .Q(g283) ) ;
OR2     gate2144  (.A(g31149), .B(g21709), .Z(g31865) ) ;
DFF     gate2145  (.D(g31865), .CP(CLK), .Q(g287) ) ;
OR2     gate2146  (.A(g32169), .B(g21710), .Z(g32977) ) ;
DFF     gate2147  (.D(g32977), .CP(CLK), .Q(g291) ) ;
OR2     gate2148  (.A(g33233), .B(g21711), .Z(g33535) ) ;
DFF     gate2149  (.D(g33535), .CP(CLK), .Q(g294) ) ;
OR2     gate2150  (.A(g33789), .B(g21712), .Z(g33961) ) ;
DFF     gate2151  (.D(g33961), .CP(CLK), .Q(g298) ) ;
OR2     gate2152  (.A(g34111), .B(g21713), .Z(g34250) ) ;
DFF     gate2153  (.D(g34250), .CP(CLK), .Q(g142) ) ;
OR2     gate2154  (.A(g29834), .B(g21699), .Z(g30333) ) ;
DFF     gate2155  (.D(g30333), .CP(CLK), .Q(g146) ) ;
OR2     gate2156  (.A(g31271), .B(g21703), .Z(g31864) ) ;
DFF     gate2157  (.D(g31864), .CP(CLK), .Q(g164) ) ;
OR2     gate2158  (.A(g32207), .B(g21704), .Z(g32976) ) ;
DFF     gate2159  (.D(g32976), .CP(CLK), .Q(g150) ) ;
OR2     gate2160  (.A(g33186), .B(g21700), .Z(g33534) ) ;
DFF     gate2161  (.D(g33534), .CP(CLK), .Q(g153) ) ;
OR2     gate2162  (.A(g33759), .B(g21701), .Z(g33960) ) ;
DFF     gate2163  (.D(g33960), .CP(CLK), .Q(g157) ) ;
OR2     gate2164  (.A(g34110), .B(g21702), .Z(g34249) ) ;
DFF     gate2165  (.D(g34249), .CP(CLK), .Q(g160) ) ;
OR2     gate2166  (.A(g33241), .B(g21715), .Z(g33536) ) ;
DFF     gate2167  (.D(g33536), .CP(CLK), .Q(g301) ) ;
OR2     gate2168  (.A(g33244), .B(g21716), .Z(g33537) ) ;
DFF     gate2169  (.D(g33537), .CP(CLK), .Q(g222) ) ;
OR2     gate2170  (.A(g24672), .B(g21706), .Z(g25592) ) ;
DFF     gate2171  (.D(g25592), .CP(CLK), .Q(g194) ) ;
DFF     gate2172  (.D(g194), .CP(CLK), .Q(g191) ) ;
OR2     gate2173  (.A(g24716), .B(g21707), .Z(g25593) ) ;
DFF     gate2174  (.D(g25593), .CP(CLK), .Q(g209) ) ;
OR2     gate2175  (.A(g24642), .B(g21705), .Z(g25591) ) ;
DFF     gate2176  (.D(g25591), .CP(CLK), .Q(g215) ) ;
DFF     gate2177  (.D(g215), .CP(CLK), .Q(g218) ) ;
OR2     gate2178  (.A(g22623), .B(g18259), .Z(g24247) ) ;
DFF     gate2179  (.D(g24247), .CP(CLK), .Q(g1249) ) ;
OR2     gate2180  (.A(g24532), .B(g18263), .Z(g25630) ) ;
DFF     gate2181  (.D(g25630), .CP(CLK), .Q(g1266) ) ;
OR2     gate2182  (.A(g25951), .B(g18267), .Z(g26919) ) ;
DFF     gate2183  (.D(g26919), .CP(CLK), .Q(g1280) ) ;
OR2     gate2184  (.A(g27235), .B(g18268), .Z(g28058) ) ;
DFF     gate2185  (.D(g28058), .CP(CLK), .Q(g1252) ) ;
OR2     gate2186  (.A(g28110), .B(g18260), .Z(g29235) ) ;
DFF     gate2187  (.D(g29235), .CP(CLK), .Q(g1256) ) ;
OR2     gate2188  (.A(g29330), .B(g18261), .Z(g30342) ) ;
DFF     gate2189  (.D(g30342), .CP(CLK), .Q(g1259) ) ;
OR2     gate2190  (.A(g30607), .B(g18262), .Z(g31870) ) ;
DFF     gate2191  (.D(g31870), .CP(CLK), .Q(g1263) ) ;
OR2     gate2192  (.A(g31934), .B(g18264), .Z(g32984) ) ;
DFF     gate2193  (.D(g32984), .CP(CLK), .Q(g1270) ) ;
OR2     gate2194  (.A(g33102), .B(g18265), .Z(g33542) ) ;
DFF     gate2195  (.D(g33542), .CP(CLK), .Q(g1274) ) ;
OR2     gate2196  (.A(g31963), .B(g18266), .Z(g32985) ) ;
DFF     gate2197  (.D(g32985), .CP(CLK), .Q(g1277) ) ;
OR2     gate2198  (.A(g23265), .B(g18306), .Z(g24254) ) ;
DFF     gate2199  (.D(g24254), .CP(CLK), .Q(g1418) ) ;
DFF     gate2200  (.D(g1418), .CP(CLK), .Q(g1422) ) ;
DFF     gate2201  (.D(g1422), .CP(CLK), .Q(g1426) ) ;
DFF     gate2202  (.D(g1426), .CP(CLK), .Q(g1430) ) ;
OR2     gate2203  (.A(g23373), .B(g18313), .Z(g24260) ) ;
DFF     gate2204  (.D(g24260), .CP(CLK), .Q(g1548) ) ;
OR2     gate2205  (.A(g23387), .B(g18315), .Z(g24262) ) ;
DFF     gate2206  (.D(g24262), .CP(CLK), .Q(g1564) ) ;
OR2     gate2207  (.A(g24977), .B(g18316), .Z(g25638) ) ;
DFF     gate2208  (.D(g25638), .CP(CLK), .Q(g1559) ) ;
OR2     gate2209  (.A(g24618), .B(g18307), .Z(g25637) ) ;
DFF     gate2210  (.D(g25637), .CP(CLK), .Q(g1554) ) ;
OR2     gate2211  (.A(g22851), .B(g18311), .Z(g24258) ) ;
DFF     gate2212  (.D(g24258), .CP(CLK), .Q(g1570) ) ;
DFF     gate2213  (.D(g1570), .CP(CLK), .Q(g1585) ) ;
OR2     gate2214  (.A(g22862), .B(g18314), .Z(g24261) ) ;
DFF     gate2215  (.D(g24261), .CP(CLK), .Q(g1589) ) ;
OR2     gate2216  (.A(g22835), .B(g18308), .Z(g24255) ) ;
DFF     gate2217  (.D(g24255), .CP(CLK), .Q(g1576) ) ;
DFF     gate2218  (.D(g1576), .CP(CLK), .Q(g1579) ) ;
OR2     gate2219  (.A(g23008), .B(g18312), .Z(g24259) ) ;
DFF     gate2220  (.D(g24259), .CP(CLK), .Q(g1339) ) ;
OR2     gate2221  (.A(g22873), .B(g18309), .Z(g24256) ) ;
DFF     gate2222  (.D(g24256), .CP(CLK), .Q(g1500) ) ;
DFF     gate2223  (.D(g1500), .CP(CLK), .Q(g1582) ) ;
DFF     gate2224  (.D(g1582), .CP(CLK), .Q(g1333) ) ;
OR2     gate2225  (.A(g22938), .B(g18310), .Z(g24257) ) ;
DFF     gate2226  (.D(g24257), .CP(CLK), .Q(g1399) ) ;
DFF     gate2227  (.D(g1399), .CP(CLK), .Q(g1459) ) ;
DFF     gate2228  (.D(g1459), .CP(CLK), .Q(g1322) ) ;
OR2     gate2229  (.A(g29630), .B(g18298), .Z(g30344) ) ;
DFF     gate2230  (.D(g30344), .CP(CLK), .Q(g1514) ) ;
OR2     gate2231  (.A(g29644), .B(g18302), .Z(g30345) ) ;
DFF     gate2232  (.D(g30345), .CP(CLK), .Q(g1526) ) ;
OR2     gate2233  (.A(g22518), .B(g18299), .Z(g24252) ) ;
DFF     gate2234  (.D(g24252), .CP(CLK), .Q(g1521) ) ;
OR2     gate2235  (.A(g24507), .B(g18305), .Z(g25636) ) ;
DFF     gate2236  (.D(g25636), .CP(CLK), .Q(g1306) ) ;
OR2     gate2237  (.A(g22525), .B(g18300), .Z(g24253) ) ;
DFF     gate2238  (.D(g24253), .CP(CLK), .Q(g1532) ) ;
OR2     gate2239  (.A(g25939), .B(g18301), .Z(g26925) ) ;
DFF     gate2240  (.D(g26925), .CP(CLK), .Q(g1536) ) ;
OR2     gate2241  (.A(g29381), .B(g18303), .Z(g30346) ) ;
DFF     gate2242  (.D(g30346), .CP(CLK), .Q(g1542) ) ;
OR2     gate2243  (.A(g29383), .B(g18304), .Z(g30347) ) ;
DFF     gate2244  (.D(g30347), .CP(CLK), .Q(g1413) ) ;
OR2     gate2245  (.A(g24559), .B(g18284), .Z(g25634) ) ;
DFF     gate2246  (.D(g25634), .CP(CLK), .Q(g1395) ) ;
OR2     gate2247  (.A(g25955), .B(g18285), .Z(g26921) ) ;
DFF     gate2248  (.D(g26921), .CP(CLK), .Q(g1404) ) ;
OR2     gate2249  (.A(g22710), .B(g18286), .Z(g24248) ) ;
DFF     gate2250  (.D(g24248), .CP(CLK), .Q(g1319) ) ;
OR2     gate2251  (.A(g24554), .B(g18275), .Z(g25631) ) ;
DFF     gate2252  (.D(g25631), .CP(CLK), .Q(g1312) ) ;
OR2     gate2253  (.A(g24558), .B(g18277), .Z(g25632) ) ;
DFF     gate2254  (.D(g25632), .CP(CLK), .Q(g1351) ) ;
OR2     gate2255  (.A(g27042), .B(g18276), .Z(g28059) ) ;
DFF     gate2256  (.D(g28059), .CP(CLK), .Q(g1345) ) ;
OR2     gate2257  (.A(g29344), .B(g18278), .Z(g30343) ) ;
DFF     gate2258  (.D(g30343), .CP(CLK), .Q(g1361) ) ;
OR2     gate2259  (.A(g30596), .B(g18279), .Z(g31871) ) ;
DFF     gate2260  (.D(g31871), .CP(CLK), .Q(g1367) ) ;
OR2     gate2261  (.A(g31996), .B(g18280), .Z(g32986) ) ;
DFF     gate2262  (.D(g32986), .CP(CLK), .Q(g1373) ) ;
OR2     gate2263  (.A(g33106), .B(g18281), .Z(g33543) ) ;
DFF     gate2264  (.D(g33543), .CP(CLK), .Q(g1379) ) ;
OR2     gate2265  (.A(g24420), .B(g18282), .Z(g25633) ) ;
DFF     gate2266  (.D(g25633), .CP(CLK), .Q(g1384) ) ;
OR2     gate2267  (.A(g25865), .B(g18283), .Z(g26920) ) ;
DFF     gate2268  (.D(g26920), .CP(CLK), .Q(g1389) ) ;
OR2     gate2269  (.A(g22624), .B(g18294), .Z(g24249) ) ;
DFF     gate2270  (.D(g24249), .CP(CLK), .Q(g1489) ) ;
OR2     gate2271  (.A(g22633), .B(g18295), .Z(g24250) ) ;
DFF     gate2272  (.D(g24250), .CP(CLK), .Q(g1495) ) ;
OR2     gate2273  (.A(g22637), .B(g18296), .Z(g24251) ) ;
DFF     gate2274  (.D(g24251), .CP(CLK), .Q(g1442) ) ;
OR2     gate2275  (.A(g28313), .B(g18287), .Z(g29236) ) ;
DFF     gate2276  (.D(g29236), .CP(CLK), .Q(g1437) ) ;
OR2     gate2277  (.A(g26153), .B(g18291), .Z(g26924) ) ;
DFF     gate2278  (.D(g26924), .CP(CLK), .Q(g1478) ) ;
OR2     gate2279  (.A(g28427), .B(g18297), .Z(g29239) ) ;
DFF     gate2280  (.D(g29239), .CP(CLK), .Q(g1454) ) ;
OR2     gate2281  (.A(g25902), .B(g18288), .Z(g26922) ) ;
DFF     gate2282  (.D(g26922), .CP(CLK), .Q(g1448) ) ;
OR2     gate2283  (.A(g28185), .B(g18289), .Z(g29237) ) ;
DFF     gate2284  (.D(g29237), .CP(CLK), .Q(g1467) ) ;
OR2     gate2285  (.A(g25923), .B(g18290), .Z(g26923) ) ;
DFF     gate2286  (.D(g26923), .CP(CLK), .Q(g1472) ) ;
OR2     gate2287  (.A(g28178), .B(g18292), .Z(g29238) ) ;
DFF     gate2288  (.D(g29238), .CP(CLK), .Q(g1484) ) ;
OR2     gate2289  (.A(g24504), .B(g18293), .Z(g25635) ) ;
DFF     gate2290  (.D(g25635), .CP(CLK), .Q(g1300) ) ;
OR2     gate2291  (.A(g34489), .B(g18269), .Z(g34602) ) ;
DFF     gate2292  (.D(g34602), .CP(CLK), .Q(g1291) ) ;
OR2     gate2293  (.A(g34666), .B(g18270), .Z(g34729) ) ;
DFF     gate2294  (.D(g34729), .CP(CLK), .Q(g1296) ) ;
OR2     gate2295  (.A(g34658), .B(g18271), .Z(g34730) ) ;
DFF     gate2296  (.D(g34730), .CP(CLK), .Q(g1283) ) ;
OR2     gate2297  (.A(g34662), .B(g18272), .Z(g34731) ) ;
DFF     gate2298  (.D(g34731), .CP(CLK), .Q(g1287) ) ;
INV     gate2299  (.A(II21291), .Z(g21724) ) ;
DFF     gate2300  (.D(g21724), .CP(CLK), .Q(g1311) ) ;
INV     gate2301  (.A(II21294), .Z(g21725) ) ;
DFF     gate2302  (.D(g21725), .CP(CLK), .Q(g929) ) ;
OR2     gate2303  (.A(g22589), .B(g18201), .Z(g24231) ) ;
DFF     gate2304  (.D(g24231), .CP(CLK), .Q(g904) ) ;
OR2     gate2305  (.A(g24523), .B(g18205), .Z(g25621) ) ;
DFF     gate2306  (.D(g25621), .CP(CLK), .Q(g921) ) ;
OR2     gate2307  (.A(g25946), .B(g18209), .Z(g26912) ) ;
DFF     gate2308  (.D(g26912), .CP(CLK), .Q(g936) ) ;
OR2     gate2309  (.A(g27230), .B(g18210), .Z(g28056) ) ;
DFF     gate2310  (.D(g28056), .CP(CLK), .Q(g907) ) ;
OR2     gate2311  (.A(g28107), .B(g18202), .Z(g29230) ) ;
DFF     gate2312  (.D(g29230), .CP(CLK), .Q(g911) ) ;
OR2     gate2313  (.A(g29324), .B(g18203), .Z(g30336) ) ;
DFF     gate2314  (.D(g30336), .CP(CLK), .Q(g914) ) ;
OR2     gate2315  (.A(g30600), .B(g18204), .Z(g31868) ) ;
DFF     gate2316  (.D(g31868), .CP(CLK), .Q(g918) ) ;
OR2     gate2317  (.A(g32425), .B(g18206), .Z(g32981) ) ;
DFF     gate2318  (.D(g32981), .CP(CLK), .Q(g925) ) ;
OR2     gate2319  (.A(g33099), .B(g18207), .Z(g33540) ) ;
DFF     gate2320  (.D(g33540), .CP(CLK), .Q(g930) ) ;
OR2     gate2321  (.A(g31948), .B(g18208), .Z(g32982) ) ;
DFF     gate2322  (.D(g32982), .CP(CLK), .Q(g933) ) ;
OR2     gate2323  (.A(g23254), .B(g18248), .Z(g24238) ) ;
DFF     gate2324  (.D(g24238), .CP(CLK), .Q(g1075) ) ;
DFF     gate2325  (.D(g1075), .CP(CLK), .Q(g1079) ) ;
DFF     gate2326  (.D(g1079), .CP(CLK), .Q(g1083) ) ;
DFF     gate2327  (.D(g1083), .CP(CLK), .Q(g1087) ) ;
OR2     gate2328  (.A(g23349), .B(g18255), .Z(g24244) ) ;
DFF     gate2329  (.D(g24244), .CP(CLK), .Q(g1205) ) ;
OR2     gate2330  (.A(g23372), .B(g18257), .Z(g24246) ) ;
DFF     gate2331  (.D(g24246), .CP(CLK), .Q(g1221) ) ;
OR2     gate2332  (.A(g24962), .B(g18258), .Z(g25629) ) ;
DFF     gate2333  (.D(g25629), .CP(CLK), .Q(g1216) ) ;
OR2     gate2334  (.A(g24600), .B(g18249), .Z(g25628) ) ;
DFF     gate2335  (.D(g25628), .CP(CLK), .Q(g1211) ) ;
OR2     gate2336  (.A(g22834), .B(g18253), .Z(g24242) ) ;
DFF     gate2337  (.D(g24242), .CP(CLK), .Q(g1227) ) ;
DFF     gate2338  (.D(g1227), .CP(CLK), .Q(g1242) ) ;
OR2     gate2339  (.A(g22849), .B(g18256), .Z(g24245) ) ;
DFF     gate2340  (.D(g24245), .CP(CLK), .Q(g1246) ) ;
OR2     gate2341  (.A(g22752), .B(g18250), .Z(g24239) ) ;
DFF     gate2342  (.D(g24239), .CP(CLK), .Q(g1233) ) ;
DFF     gate2343  (.D(g1233), .CP(CLK), .Q(g1236) ) ;
OR2     gate2344  (.A(g22992), .B(g18254), .Z(g24243) ) ;
DFF     gate2345  (.D(g24243), .CP(CLK), .Q(g996) ) ;
OR2     gate2346  (.A(g22861), .B(g18251), .Z(g24240) ) ;
DFF     gate2347  (.D(g24240), .CP(CLK), .Q(g1157) ) ;
DFF     gate2348  (.D(g1157), .CP(CLK), .Q(g1239) ) ;
DFF     gate2349  (.D(g1239), .CP(CLK), .Q(g990) ) ;
OR2     gate2350  (.A(g22920), .B(g18252), .Z(g24241) ) ;
DFF     gate2351  (.D(g24241), .CP(CLK), .Q(g1056) ) ;
DFF     gate2352  (.D(g1056), .CP(CLK), .Q(g1116) ) ;
DFF     gate2353  (.D(g1116), .CP(CLK), .Q(g979) ) ;
OR2     gate2354  (.A(g29613), .B(g18240), .Z(g30338) ) ;
DFF     gate2355  (.D(g30338), .CP(CLK), .Q(g1171) ) ;
OR2     gate2356  (.A(g29629), .B(g18244), .Z(g30339) ) ;
DFF     gate2357  (.D(g30339), .CP(CLK), .Q(g1183) ) ;
OR2     gate2358  (.A(g22489), .B(g18241), .Z(g24236) ) ;
DFF     gate2359  (.D(g24236), .CP(CLK), .Q(g1178) ) ;
OR2     gate2360  (.A(g24503), .B(g18247), .Z(g25627) ) ;
DFF     gate2361  (.D(g25627), .CP(CLK), .Q(g962) ) ;
OR2     gate2362  (.A(g22515), .B(g18242), .Z(g24237) ) ;
DFF     gate2363  (.D(g24237), .CP(CLK), .Q(g1189) ) ;
OR2     gate2364  (.A(g25931), .B(g18243), .Z(g26918) ) ;
DFF     gate2365  (.D(g26918), .CP(CLK), .Q(g1193) ) ;
OR2     gate2366  (.A(g29377), .B(g18245), .Z(g30340) ) ;
DFF     gate2367  (.D(g30340), .CP(CLK), .Q(g1199) ) ;
OR2     gate2368  (.A(g29380), .B(g18246), .Z(g30341) ) ;
DFF     gate2369  (.D(g30341), .CP(CLK), .Q(g1070) ) ;
OR2     gate2370  (.A(g24553), .B(g18226), .Z(g25625) ) ;
DFF     gate2371  (.D(g25625), .CP(CLK), .Q(g1052) ) ;
OR2     gate2372  (.A(g25949), .B(g18227), .Z(g26914) ) ;
DFF     gate2373  (.D(g26914), .CP(CLK), .Q(g1061) ) ;
OR2     gate2374  (.A(g22686), .B(g18228), .Z(g24232) ) ;
DFF     gate2375  (.D(g24232), .CP(CLK), .Q(g976) ) ;
OR2     gate2376  (.A(g24546), .B(g18217), .Z(g25622) ) ;
DFF     gate2377  (.D(g25622), .CP(CLK), .Q(g969) ) ;
OR2     gate2378  (.A(g24552), .B(g18219), .Z(g25623) ) ;
DFF     gate2379  (.D(g25623), .CP(CLK), .Q(g1008) ) ;
OR2     gate2380  (.A(g27033), .B(g18218), .Z(g28057) ) ;
DFF     gate2381  (.D(g28057), .CP(CLK), .Q(g1002) ) ;
OR2     gate2382  (.A(g29334), .B(g18220), .Z(g30337) ) ;
DFF     gate2383  (.D(g30337), .CP(CLK), .Q(g1018) ) ;
OR2     gate2384  (.A(g30592), .B(g18221), .Z(g31869) ) ;
DFF     gate2385  (.D(g31869), .CP(CLK), .Q(g1024) ) ;
OR2     gate2386  (.A(g31990), .B(g18222), .Z(g32983) ) ;
DFF     gate2387  (.D(g32983), .CP(CLK), .Q(g1030) ) ;
OR2     gate2388  (.A(g33101), .B(g18223), .Z(g33541) ) ;
DFF     gate2389  (.D(g33541), .CP(CLK), .Q(g1036) ) ;
OR2     gate2390  (.A(g24408), .B(g18224), .Z(g25624) ) ;
DFF     gate2391  (.D(g25624), .CP(CLK), .Q(g1041) ) ;
OR2     gate2392  (.A(g25848), .B(g18225), .Z(g26913) ) ;
DFF     gate2393  (.D(g26913), .CP(CLK), .Q(g1046) ) ;
OR2     gate2394  (.A(g22590), .B(g18236), .Z(g24233) ) ;
DFF     gate2395  (.D(g24233), .CP(CLK), .Q(g1146) ) ;
OR2     gate2396  (.A(g22622), .B(g18237), .Z(g24234) ) ;
DFF     gate2397  (.D(g24234), .CP(CLK), .Q(g1152) ) ;
OR2     gate2398  (.A(g22632), .B(g18238), .Z(g24235) ) ;
DFF     gate2399  (.D(g24235), .CP(CLK), .Q(g1099) ) ;
OR2     gate2400  (.A(g28301), .B(g18229), .Z(g29231) ) ;
DFF     gate2401  (.D(g29231), .CP(CLK), .Q(g1094) ) ;
OR2     gate2402  (.A(g26122), .B(g18233), .Z(g26917) ) ;
DFF     gate2403  (.D(g26917), .CP(CLK), .Q(g1135) ) ;
OR2     gate2404  (.A(g28415), .B(g18239), .Z(g29234) ) ;
DFF     gate2405  (.D(g29234), .CP(CLK), .Q(g1111) ) ;
OR2     gate2406  (.A(g25900), .B(g18230), .Z(g26915) ) ;
DFF     gate2407  (.D(g26915), .CP(CLK), .Q(g1105) ) ;
OR2     gate2408  (.A(g28183), .B(g18231), .Z(g29232) ) ;
DFF     gate2409  (.D(g29232), .CP(CLK), .Q(g1124) ) ;
OR2     gate2410  (.A(g25916), .B(g18232), .Z(g26916) ) ;
DFF     gate2411  (.D(g26916), .CP(CLK), .Q(g1129) ) ;
OR2     gate2412  (.A(g28171), .B(g18234), .Z(g29233) ) ;
DFF     gate2413  (.D(g29233), .CP(CLK), .Q(g1141) ) ;
OR2     gate2414  (.A(g24499), .B(g18235), .Z(g25626) ) ;
DFF     gate2415  (.D(g25626), .CP(CLK), .Q(g956) ) ;
OR2     gate2416  (.A(g34488), .B(g18211), .Z(g34601) ) ;
DFF     gate2417  (.D(g34601), .CP(CLK), .Q(g947) ) ;
OR2     gate2418  (.A(g34665), .B(g18212), .Z(g34726) ) ;
DFF     gate2419  (.D(g34726), .CP(CLK), .Q(g952) ) ;
OR2     gate2420  (.A(g34655), .B(g18213), .Z(g34727) ) ;
DFF     gate2421  (.D(g34727), .CP(CLK), .Q(g939) ) ;
OR2     gate2422  (.A(g34661), .B(g18214), .Z(g34728) ) ;
DFF     gate2423  (.D(g34728), .CP(CLK), .Q(g943) ) ;
INV     gate2424  (.A(II21285), .Z(g21722) ) ;
DFF     gate2425  (.D(g21722), .CP(CLK), .Q(g967) ) ;
INV     gate2426  (.A(II21288), .Z(g21723) ) ;
DFF     gate2427  (.D(g21723), .CP(CLK), .Q(g968) ) ;
OR2     gate2428  (.A(g33392), .B(g18317), .Z(g33544) ) ;
DFF     gate2429  (.D(g33544), .CP(CLK), .Q(g1592) ) ;
OR2     gate2430  (.A(g33446), .B(g18342), .Z(g33551) ) ;
DFF     gate2431  (.D(g33551), .CP(CLK), .Q(g1644) ) ;
OR2     gate2432  (.A(g33399), .B(g18324), .Z(g33545) ) ;
DFF     gate2433  (.D(g33545), .CP(CLK), .Q(g1636) ) ;
OR2     gate2434  (.A(g33402), .B(g18327), .Z(g33546) ) ;
DFF     gate2435  (.D(g33546), .CP(CLK), .Q(g1668) ) ;
OR2     gate2436  (.A(g33890), .B(g18330), .Z(g33971) ) ;
DFF     gate2437  (.D(g33971), .CP(CLK), .Q(g1682) ) ;
OR2     gate2438  (.A(g33349), .B(g18331), .Z(g33547) ) ;
DFF     gate2439  (.D(g33547), .CP(CLK), .Q(g1687) ) ;
OR2     gate2440  (.A(g33941), .B(g18335), .Z(g33972) ) ;
DFF     gate2441  (.D(g33972), .CP(CLK), .Q(g1604) ) ;
OR2     gate2442  (.A(g33837), .B(g18318), .Z(g33966) ) ;
DFF     gate2443  (.D(g33966), .CP(CLK), .Q(g1600) ) ;
OR2     gate2444  (.A(g33842), .B(g18319), .Z(g33967) ) ;
DFF     gate2445  (.D(g33967), .CP(CLK), .Q(g1608) ) ;
OR2     gate2446  (.A(g33868), .B(g18322), .Z(g33970) ) ;
DFF     gate2447  (.D(g33970), .CP(CLK), .Q(g1620) ) ;
OR2     gate2448  (.A(g33864), .B(g18321), .Z(g33969) ) ;
DFF     gate2449  (.D(g33969), .CP(CLK), .Q(g1616) ) ;
OR2     gate2450  (.A(g33855), .B(g18320), .Z(g33968) ) ;
DFF     gate2451  (.D(g33968), .CP(CLK), .Q(g1612) ) ;
OR2     gate2452  (.A(g30083), .B(g18329), .Z(g30348) ) ;
DFF     gate2453  (.D(g30348), .CP(CLK), .Q(g1632) ) ;
OR2     gate2454  (.A(g32311), .B(g18323), .Z(g32987) ) ;
DFF     gate2455  (.D(g32987), .CP(CLK), .Q(g1624) ) ;
OR2     gate2456  (.A(g32232), .B(g18325), .Z(g32988) ) ;
DFF     gate2457  (.D(g32988), .CP(CLK), .Q(g1648) ) ;
OR2     gate2458  (.A(g32281), .B(g18341), .Z(g32990) ) ;
DFF     gate2459  (.D(g32990), .CP(CLK), .Q(g1664) ) ;
OR2     gate2460  (.A(g32241), .B(g18326), .Z(g32989) ) ;
DFF     gate2461  (.D(g32989), .CP(CLK), .Q(g1657) ) ;
OR2     gate2462  (.A(g28655), .B(g18328), .Z(g29240) ) ;
DFF     gate2463  (.D(g29240), .CP(CLK), .Q(g1677) ) ;
OR2     gate2464  (.A(g28638), .B(g18332), .Z(g29241) ) ;
DFF     gate2465  (.D(g29241), .CP(CLK), .Q(g1691) ) ;
OR2     gate2466  (.A(g30051), .B(g18333), .Z(g30349) ) ;
DFF     gate2467  (.D(g30349), .CP(CLK), .Q(g1696) ) ;
OR2     gate2468  (.A(g30118), .B(g18334), .Z(g30350) ) ;
DFF     gate2469  (.D(g30350), .CP(CLK), .Q(g1700) ) ;
OR2     gate2470  (.A(g33327), .B(g18336), .Z(g33548) ) ;
DFF     gate2471  (.D(g33548), .CP(CLK), .Q(g1706) ) ;
OR2     gate2472  (.A(g33328), .B(g18337), .Z(g33549) ) ;
DFF     gate2473  (.D(g33549), .CP(CLK), .Q(g1710) ) ;
OR2     gate2474  (.A(g33342), .B(g18338), .Z(g33550) ) ;
DFF     gate2475  (.D(g33550), .CP(CLK), .Q(g1714) ) ;
OR2     gate2476  (.A(g30084), .B(g18339), .Z(g30351) ) ;
DFF     gate2477  (.D(g30351), .CP(CLK), .Q(g1720) ) ;
OR2     gate2478  (.A(g30094), .B(g18340), .Z(g30352) ) ;
DFF     gate2479  (.D(g30352), .CP(CLK), .Q(g1724) ) ;
OR2     gate2480  (.A(g33400), .B(g18343), .Z(g33552) ) ;
DFF     gate2481  (.D(g33552), .CP(CLK), .Q(g1728) ) ;
OR2     gate2482  (.A(g33073), .B(g18368), .Z(g33559) ) ;
DFF     gate2483  (.D(g33559), .CP(CLK), .Q(g1779) ) ;
OR2     gate2484  (.A(g33403), .B(g18350), .Z(g33553) ) ;
DFF     gate2485  (.D(g33553), .CP(CLK), .Q(g1772) ) ;
OR2     gate2486  (.A(g33407), .B(g18353), .Z(g33554) ) ;
DFF     gate2487  (.D(g33554), .CP(CLK), .Q(g1802) ) ;
OR2     gate2488  (.A(g33892), .B(g18356), .Z(g33978) ) ;
DFF     gate2489  (.D(g33978), .CP(CLK), .Q(g1816) ) ;
OR2     gate2490  (.A(g33355), .B(g18357), .Z(g33555) ) ;
DFF     gate2491  (.D(g33555), .CP(CLK), .Q(g1821) ) ;
OR2     gate2492  (.A(g33942), .B(g18361), .Z(g33979) ) ;
DFF     gate2493  (.D(g33979), .CP(CLK), .Q(g1740) ) ;
OR2     gate2494  (.A(g33840), .B(g18344), .Z(g33973) ) ;
DFF     gate2495  (.D(g33973), .CP(CLK), .Q(g1736) ) ;
OR2     gate2496  (.A(g33846), .B(g18345), .Z(g33974) ) ;
DFF     gate2497  (.D(g33974), .CP(CLK), .Q(g1744) ) ;
OR2     gate2498  (.A(g33876), .B(g18348), .Z(g33977) ) ;
DFF     gate2499  (.D(g33977), .CP(CLK), .Q(g1756) ) ;
OR2     gate2500  (.A(g33869), .B(g18347), .Z(g33976) ) ;
DFF     gate2501  (.D(g33976), .CP(CLK), .Q(g1752) ) ;
OR2     gate2502  (.A(g33860), .B(g18346), .Z(g33975) ) ;
DFF     gate2503  (.D(g33975), .CP(CLK), .Q(g1748) ) ;
OR2     gate2504  (.A(g30095), .B(g18355), .Z(g30353) ) ;
DFF     gate2505  (.D(g30353), .CP(CLK), .Q(g1768) ) ;
OR2     gate2506  (.A(g32322), .B(g18349), .Z(g32991) ) ;
DFF     gate2507  (.D(g32991), .CP(CLK), .Q(g1760) ) ;
OR2     gate2508  (.A(g32242), .B(g18351), .Z(g32992) ) ;
DFF     gate2509  (.D(g32992), .CP(CLK), .Q(g1783) ) ;
OR2     gate2510  (.A(g32290), .B(g18367), .Z(g32994) ) ;
DFF     gate2511  (.D(g32994), .CP(CLK), .Q(g1798) ) ;
OR2     gate2512  (.A(g32255), .B(g18352), .Z(g32993) ) ;
DFF     gate2513  (.D(g32993), .CP(CLK), .Q(g1792) ) ;
OR2     gate2514  (.A(g28674), .B(g18354), .Z(g29242) ) ;
DFF     gate2515  (.D(g29242), .CP(CLK), .Q(g1811) ) ;
OR2     gate2516  (.A(g28657), .B(g18358), .Z(g29243) ) ;
DFF     gate2517  (.D(g29243), .CP(CLK), .Q(g1825) ) ;
OR2     gate2518  (.A(g30064), .B(g18359), .Z(g30354) ) ;
DFF     gate2519  (.D(g30354), .CP(CLK), .Q(g1830) ) ;
OR2     gate2520  (.A(g30131), .B(g18360), .Z(g30355) ) ;
DFF     gate2521  (.D(g30355), .CP(CLK), .Q(g1834) ) ;
OR2     gate2522  (.A(g33329), .B(g18362), .Z(g33556) ) ;
DFF     gate2523  (.D(g33556), .CP(CLK), .Q(g1840) ) ;
OR2     gate2524  (.A(g33331), .B(g18363), .Z(g33557) ) ;
DFF     gate2525  (.D(g33557), .CP(CLK), .Q(g1844) ) ;
OR2     gate2526  (.A(g33350), .B(g18364), .Z(g33558) ) ;
DFF     gate2527  (.D(g33558), .CP(CLK), .Q(g1848) ) ;
OR2     gate2528  (.A(g30096), .B(g18365), .Z(g30356) ) ;
DFF     gate2529  (.D(g30356), .CP(CLK), .Q(g1854) ) ;
OR2     gate2530  (.A(g30107), .B(g18366), .Z(g30357) ) ;
DFF     gate2531  (.D(g30357), .CP(CLK), .Q(g1858) ) ;
OR2     gate2532  (.A(g33404), .B(g18369), .Z(g33560) ) ;
DFF     gate2533  (.D(g33560), .CP(CLK), .Q(g1862) ) ;
OR2     gate2534  (.A(g33081), .B(g18394), .Z(g33567) ) ;
DFF     gate2535  (.D(g33567), .CP(CLK), .Q(g1913) ) ;
OR2     gate2536  (.A(g33408), .B(g18376), .Z(g33561) ) ;
DFF     gate2537  (.D(g33561), .CP(CLK), .Q(g1906) ) ;
OR2     gate2538  (.A(g33414), .B(g18379), .Z(g33562) ) ;
DFF     gate2539  (.D(g33562), .CP(CLK), .Q(g1936) ) ;
OR2     gate2540  (.A(g33896), .B(g18382), .Z(g33985) ) ;
DFF     gate2541  (.D(g33985), .CP(CLK), .Q(g1950) ) ;
OR2     gate2542  (.A(g33361), .B(g18383), .Z(g33563) ) ;
DFF     gate2543  (.D(g33563), .CP(CLK), .Q(g1955) ) ;
OR2     gate2544  (.A(g33639), .B(g18387), .Z(g33986) ) ;
DFF     gate2545  (.D(g33986), .CP(CLK), .Q(g1874) ) ;
OR2     gate2546  (.A(g33843), .B(g18370), .Z(g33980) ) ;
DFF     gate2547  (.D(g33980), .CP(CLK), .Q(g1870) ) ;
OR2     gate2548  (.A(g33856), .B(g18371), .Z(g33981) ) ;
DFF     gate2549  (.D(g33981), .CP(CLK), .Q(g1878) ) ;
OR2     gate2550  (.A(g33881), .B(g18374), .Z(g33984) ) ;
DFF     gate2551  (.D(g33984), .CP(CLK), .Q(g1890) ) ;
OR2     gate2552  (.A(g33877), .B(g18373), .Z(g33983) ) ;
DFF     gate2553  (.D(g33983), .CP(CLK), .Q(g1886) ) ;
OR2     gate2554  (.A(g33865), .B(g18372), .Z(g33982) ) ;
DFF     gate2555  (.D(g33982), .CP(CLK), .Q(g1882) ) ;
OR2     gate2556  (.A(g30108), .B(g18381), .Z(g30358) ) ;
DFF     gate2557  (.D(g30358), .CP(CLK), .Q(g1902) ) ;
OR2     gate2558  (.A(g32330), .B(g18375), .Z(g32995) ) ;
DFF     gate2559  (.D(g32995), .CP(CLK), .Q(g1894) ) ;
OR2     gate2560  (.A(g32256), .B(g18377), .Z(g32996) ) ;
DFF     gate2561  (.D(g32996), .CP(CLK), .Q(g1917) ) ;
OR2     gate2562  (.A(g32300), .B(g18393), .Z(g32998) ) ;
DFF     gate2563  (.D(g32998), .CP(CLK), .Q(g1932) ) ;
OR2     gate2564  (.A(g32269), .B(g18378), .Z(g32997) ) ;
DFF     gate2565  (.D(g32997), .CP(CLK), .Q(g1926) ) ;
OR2     gate2566  (.A(g28692), .B(g18380), .Z(g29244) ) ;
DFF     gate2567  (.D(g29244), .CP(CLK), .Q(g1945) ) ;
OR2     gate2568  (.A(g28676), .B(g18384), .Z(g29245) ) ;
DFF     gate2569  (.D(g29245), .CP(CLK), .Q(g1959) ) ;
OR2     gate2570  (.A(g30075), .B(g18385), .Z(g30359) ) ;
DFF     gate2571  (.D(g30359), .CP(CLK), .Q(g1964) ) ;
OR2     gate2572  (.A(g30145), .B(g18386), .Z(g30360) ) ;
DFF     gate2573  (.D(g30360), .CP(CLK), .Q(g1968) ) ;
OR2     gate2574  (.A(g33332), .B(g18388), .Z(g33564) ) ;
DFF     gate2575  (.D(g33564), .CP(CLK), .Q(g1974) ) ;
OR2     gate2576  (.A(g33338), .B(g18389), .Z(g33565) ) ;
DFF     gate2577  (.D(g33565), .CP(CLK), .Q(g1978) ) ;
OR2     gate2578  (.A(g33356), .B(g18390), .Z(g33566) ) ;
DFF     gate2579  (.D(g33566), .CP(CLK), .Q(g1982) ) ;
OR2     gate2580  (.A(g30109), .B(g18391), .Z(g30361) ) ;
DFF     gate2581  (.D(g30361), .CP(CLK), .Q(g1988) ) ;
OR2     gate2582  (.A(g30120), .B(g18392), .Z(g30362) ) ;
DFF     gate2583  (.D(g30362), .CP(CLK), .Q(g1992) ) ;
OR2     gate2584  (.A(g33409), .B(g18395), .Z(g33568) ) ;
DFF     gate2585  (.D(g33568), .CP(CLK), .Q(g1996) ) ;
OR2     gate2586  (.A(g33086), .B(g18420), .Z(g33575) ) ;
DFF     gate2587  (.D(g33575), .CP(CLK), .Q(g2047) ) ;
OR2     gate2588  (.A(g33415), .B(g18402), .Z(g33569) ) ;
DFF     gate2589  (.D(g33569), .CP(CLK), .Q(g2040) ) ;
OR2     gate2590  (.A(g33420), .B(g18405), .Z(g33570) ) ;
DFF     gate2591  (.D(g33570), .CP(CLK), .Q(g2070) ) ;
OR2     gate2592  (.A(g33900), .B(g18408), .Z(g33992) ) ;
DFF     gate2593  (.D(g33992), .CP(CLK), .Q(g2084) ) ;
OR2     gate2594  (.A(g33367), .B(g18409), .Z(g33571) ) ;
DFF     gate2595  (.D(g33571), .CP(CLK), .Q(g2089) ) ;
OR2     gate2596  (.A(g33646), .B(g18413), .Z(g33993) ) ;
DFF     gate2597  (.D(g33993), .CP(CLK), .Q(g2008) ) ;
OR2     gate2598  (.A(g33847), .B(g18396), .Z(g33987) ) ;
DFF     gate2599  (.D(g33987), .CP(CLK), .Q(g2004) ) ;
OR2     gate2600  (.A(g33861), .B(g18397), .Z(g33988) ) ;
DFF     gate2601  (.D(g33988), .CP(CLK), .Q(g2012) ) ;
OR2     gate2602  (.A(g33885), .B(g18400), .Z(g33991) ) ;
DFF     gate2603  (.D(g33991), .CP(CLK), .Q(g2024) ) ;
OR2     gate2604  (.A(g33882), .B(g18399), .Z(g33990) ) ;
DFF     gate2605  (.D(g33990), .CP(CLK), .Q(g2020) ) ;
OR2     gate2606  (.A(g33870), .B(g18398), .Z(g33989) ) ;
DFF     gate2607  (.D(g33989), .CP(CLK), .Q(g2016) ) ;
OR2     gate2608  (.A(g30121), .B(g18407), .Z(g30363) ) ;
DFF     gate2609  (.D(g30363), .CP(CLK), .Q(g2036) ) ;
OR2     gate2610  (.A(g32337), .B(g18401), .Z(g32999) ) ;
DFF     gate2611  (.D(g32999), .CP(CLK), .Q(g2028) ) ;
OR2     gate2612  (.A(g32270), .B(g18403), .Z(g33000) ) ;
DFF     gate2613  (.D(g33000), .CP(CLK), .Q(g2051) ) ;
OR2     gate2614  (.A(g32304), .B(g18419), .Z(g33002) ) ;
DFF     gate2615  (.D(g33002), .CP(CLK), .Q(g2066) ) ;
OR2     gate2616  (.A(g32282), .B(g18404), .Z(g33001) ) ;
DFF     gate2617  (.D(g33001), .CP(CLK), .Q(g2060) ) ;
OR2     gate2618  (.A(g28710), .B(g18406), .Z(g29246) ) ;
DFF     gate2619  (.D(g29246), .CP(CLK), .Q(g2079) ) ;
OR2     gate2620  (.A(g28694), .B(g18410), .Z(g29247) ) ;
DFF     gate2621  (.D(g29247), .CP(CLK), .Q(g2093) ) ;
OR2     gate2622  (.A(g30086), .B(g18411), .Z(g30364) ) ;
DFF     gate2623  (.D(g30364), .CP(CLK), .Q(g2098) ) ;
OR2     gate2624  (.A(g30158), .B(g18412), .Z(g30365) ) ;
DFF     gate2625  (.D(g30365), .CP(CLK), .Q(g2102) ) ;
OR2     gate2626  (.A(g33339), .B(g18414), .Z(g33572) ) ;
DFF     gate2627  (.D(g33572), .CP(CLK), .Q(g2108) ) ;
OR2     gate2628  (.A(g33343), .B(g18415), .Z(g33573) ) ;
DFF     gate2629  (.D(g33573), .CP(CLK), .Q(g2112) ) ;
OR2     gate2630  (.A(g33362), .B(g18416), .Z(g33574) ) ;
DFF     gate2631  (.D(g33574), .CP(CLK), .Q(g2116) ) ;
OR2     gate2632  (.A(g30122), .B(g18417), .Z(g30366) ) ;
DFF     gate2633  (.D(g30366), .CP(CLK), .Q(g2122) ) ;
OR2     gate2634  (.A(g30133), .B(g18418), .Z(g30367) ) ;
DFF     gate2635  (.D(g30367), .CP(CLK), .Q(g2126) ) ;
OR2     gate2636  (.A(g34561), .B(g15075), .Z(g34603) ) ;
DFF     gate2637  (.D(g34603), .CP(CLK), .Q(g2130) ) ;
OR2     gate2638  (.A(g34563), .B(g15076), .Z(g34604) ) ;
DFF     gate2639  (.D(g34604), .CP(CLK), .Q(g2138) ) ;
OR2     gate2640  (.A(g34566), .B(g15077), .Z(g34605) ) ;
DFF     gate2641  (.D(g34605), .CP(CLK), .Q(g2145) ) ;
INV     gate2642  (.A(II19235), .Z(g18421) ) ;
DFF     gate2643  (.D(g18421), .CP(CLK), .Q(g2151) ) ;
INV     gate2644  (.A(II19238), .Z(g18422) ) ;
DFF     gate2645  (.D(g18422), .CP(CLK), .Q(g2152) ) ;
OR2     gate2646  (.A(g33401), .B(g18423), .Z(g33576) ) ;
DFF     gate2647  (.D(g33576), .CP(CLK), .Q(g2153) ) ;
OR2     gate2648  (.A(g33074), .B(g18448), .Z(g33583) ) ;
DFF     gate2649  (.D(g33583), .CP(CLK), .Q(g2204) ) ;
OR2     gate2650  (.A(g33405), .B(g18430), .Z(g33577) ) ;
DFF     gate2651  (.D(g33577), .CP(CLK), .Q(g2197) ) ;
OR2     gate2652  (.A(g33410), .B(g18433), .Z(g33578) ) ;
DFF     gate2653  (.D(g33578), .CP(CLK), .Q(g2227) ) ;
OR2     gate2654  (.A(g33893), .B(g18436), .Z(g33999) ) ;
DFF     gate2655  (.D(g33999), .CP(CLK), .Q(g2241) ) ;
OR2     gate2656  (.A(g33357), .B(g18437), .Z(g33579) ) ;
DFF     gate2657  (.D(g33579), .CP(CLK), .Q(g2246) ) ;
OR2     gate2658  (.A(g33943), .B(g18441), .Z(g34000) ) ;
DFF     gate2659  (.D(g34000), .CP(CLK), .Q(g2165) ) ;
OR2     gate2660  (.A(g33841), .B(g18424), .Z(g33994) ) ;
DFF     gate2661  (.D(g33994), .CP(CLK), .Q(g2161) ) ;
OR2     gate2662  (.A(g33848), .B(g18425), .Z(g33995) ) ;
DFF     gate2663  (.D(g33995), .CP(CLK), .Q(g2169) ) ;
OR2     gate2664  (.A(g33878), .B(g18428), .Z(g33998) ) ;
DFF     gate2665  (.D(g33998), .CP(CLK), .Q(g2181) ) ;
OR2     gate2666  (.A(g33871), .B(g18427), .Z(g33997) ) ;
DFF     gate2667  (.D(g33997), .CP(CLK), .Q(g2177) ) ;
OR2     gate2668  (.A(g33862), .B(g18426), .Z(g33996) ) ;
DFF     gate2669  (.D(g33996), .CP(CLK), .Q(g2173) ) ;
OR2     gate2670  (.A(g30098), .B(g18435), .Z(g30368) ) ;
DFF     gate2671  (.D(g30368), .CP(CLK), .Q(g2193) ) ;
OR2     gate2672  (.A(g32323), .B(g18429), .Z(g33003) ) ;
DFF     gate2673  (.D(g33003), .CP(CLK), .Q(g2185) ) ;
OR2     gate2674  (.A(g32246), .B(g18431), .Z(g33004) ) ;
DFF     gate2675  (.D(g33004), .CP(CLK), .Q(g2208) ) ;
OR2     gate2676  (.A(g32291), .B(g18447), .Z(g33006) ) ;
DFF     gate2677  (.D(g33006), .CP(CLK), .Q(g2223) ) ;
OR2     gate2678  (.A(g32260), .B(g18432), .Z(g33005) ) ;
DFF     gate2679  (.D(g33005), .CP(CLK), .Q(g2217) ) ;
OR2     gate2680  (.A(g28677), .B(g18434), .Z(g29248) ) ;
DFF     gate2681  (.D(g29248), .CP(CLK), .Q(g2236) ) ;
OR2     gate2682  (.A(g28658), .B(g18438), .Z(g29249) ) ;
DFF     gate2683  (.D(g29249), .CP(CLK), .Q(g2250) ) ;
OR2     gate2684  (.A(g30066), .B(g18439), .Z(g30369) ) ;
DFF     gate2685  (.D(g30369), .CP(CLK), .Q(g2255) ) ;
OR2     gate2686  (.A(g30135), .B(g18440), .Z(g30370) ) ;
DFF     gate2687  (.D(g30370), .CP(CLK), .Q(g2259) ) ;
OR2     gate2688  (.A(g33330), .B(g18442), .Z(g33580) ) ;
DFF     gate2689  (.D(g33580), .CP(CLK), .Q(g2265) ) ;
OR2     gate2690  (.A(g33333), .B(g18443), .Z(g33581) ) ;
DFF     gate2691  (.D(g33581), .CP(CLK), .Q(g2269) ) ;
OR2     gate2692  (.A(g33351), .B(g18444), .Z(g33582) ) ;
DFF     gate2693  (.D(g33582), .CP(CLK), .Q(g2273) ) ;
OR2     gate2694  (.A(g30099), .B(g18445), .Z(g30371) ) ;
DFF     gate2695  (.D(g30371), .CP(CLK), .Q(g2279) ) ;
OR2     gate2696  (.A(g30110), .B(g18446), .Z(g30372) ) ;
DFF     gate2697  (.D(g30372), .CP(CLK), .Q(g2283) ) ;
OR2     gate2698  (.A(g33406), .B(g18449), .Z(g33584) ) ;
DFF     gate2699  (.D(g33584), .CP(CLK), .Q(g2287) ) ;
OR2     gate2700  (.A(g33082), .B(g18474), .Z(g33591) ) ;
DFF     gate2701  (.D(g33591), .CP(CLK), .Q(g2338) ) ;
OR2     gate2702  (.A(g33411), .B(g18456), .Z(g33585) ) ;
DFF     gate2703  (.D(g33585), .CP(CLK), .Q(g2331) ) ;
OR2     gate2704  (.A(g33416), .B(g18459), .Z(g33586) ) ;
DFF     gate2705  (.D(g33586), .CP(CLK), .Q(g2361) ) ;
OR2     gate2706  (.A(g33897), .B(g18462), .Z(g34006) ) ;
DFF     gate2707  (.D(g34006), .CP(CLK), .Q(g2375) ) ;
OR2     gate2708  (.A(g33363), .B(g18463), .Z(g33587) ) ;
DFF     gate2709  (.D(g33587), .CP(CLK), .Q(g2380) ) ;
OR2     gate2710  (.A(g33640), .B(g18467), .Z(g34007) ) ;
DFF     gate2711  (.D(g34007), .CP(CLK), .Q(g2299) ) ;
OR2     gate2712  (.A(g33844), .B(g18450), .Z(g34001) ) ;
DFF     gate2713  (.D(g34001), .CP(CLK), .Q(g2295) ) ;
OR2     gate2714  (.A(g33857), .B(g18451), .Z(g34002) ) ;
DFF     gate2715  (.D(g34002), .CP(CLK), .Q(g2303) ) ;
OR2     gate2716  (.A(g33883), .B(g18454), .Z(g34005) ) ;
DFF     gate2717  (.D(g34005), .CP(CLK), .Q(g2315) ) ;
OR2     gate2718  (.A(g33879), .B(g18453), .Z(g34004) ) ;
DFF     gate2719  (.D(g34004), .CP(CLK), .Q(g2311) ) ;
OR2     gate2720  (.A(g33866), .B(g18452), .Z(g34003) ) ;
DFF     gate2721  (.D(g34003), .CP(CLK), .Q(g2307) ) ;
OR2     gate2722  (.A(g30111), .B(g18461), .Z(g30373) ) ;
DFF     gate2723  (.D(g30373), .CP(CLK), .Q(g2327) ) ;
OR2     gate2724  (.A(g32331), .B(g18455), .Z(g33007) ) ;
DFF     gate2725  (.D(g33007), .CP(CLK), .Q(g2319) ) ;
OR2     gate2726  (.A(g32261), .B(g18457), .Z(g33008) ) ;
DFF     gate2727  (.D(g33008), .CP(CLK), .Q(g2342) ) ;
OR2     gate2728  (.A(g32301), .B(g18473), .Z(g33010) ) ;
DFF     gate2729  (.D(g33010), .CP(CLK), .Q(g2357) ) ;
OR2     gate2730  (.A(g32273), .B(g18458), .Z(g33009) ) ;
DFF     gate2731  (.D(g33009), .CP(CLK), .Q(g2351) ) ;
OR2     gate2732  (.A(g28695), .B(g18460), .Z(g29250) ) ;
DFF     gate2733  (.D(g29250), .CP(CLK), .Q(g2370) ) ;
OR2     gate2734  (.A(g28679), .B(g18464), .Z(g29251) ) ;
DFF     gate2735  (.D(g29251), .CP(CLK), .Q(g2384) ) ;
OR2     gate2736  (.A(g30078), .B(g18465), .Z(g30374) ) ;
DFF     gate2737  (.D(g30374), .CP(CLK), .Q(g2389) ) ;
OR2     gate2738  (.A(g30149), .B(g18466), .Z(g30375) ) ;
DFF     gate2739  (.D(g30375), .CP(CLK), .Q(g2393) ) ;
OR2     gate2740  (.A(g33334), .B(g18468), .Z(g33588) ) ;
DFF     gate2741  (.D(g33588), .CP(CLK), .Q(g2399) ) ;
OR2     gate2742  (.A(g33340), .B(g18469), .Z(g33589) ) ;
DFF     gate2743  (.D(g33589), .CP(CLK), .Q(g2403) ) ;
OR2     gate2744  (.A(g33358), .B(g18470), .Z(g33590) ) ;
DFF     gate2745  (.D(g33590), .CP(CLK), .Q(g2407) ) ;
OR2     gate2746  (.A(g30112), .B(g18471), .Z(g30376) ) ;
DFF     gate2747  (.D(g30376), .CP(CLK), .Q(g2413) ) ;
OR2     gate2748  (.A(g30124), .B(g18472), .Z(g30377) ) ;
DFF     gate2749  (.D(g30377), .CP(CLK), .Q(g2417) ) ;
OR2     gate2750  (.A(g33412), .B(g18475), .Z(g33592) ) ;
DFF     gate2751  (.D(g33592), .CP(CLK), .Q(g2421) ) ;
OR2     gate2752  (.A(g33087), .B(g18500), .Z(g33599) ) ;
DFF     gate2753  (.D(g33599), .CP(CLK), .Q(g2472) ) ;
OR2     gate2754  (.A(g33417), .B(g18482), .Z(g33593) ) ;
DFF     gate2755  (.D(g33593), .CP(CLK), .Q(g2465) ) ;
OR2     gate2756  (.A(g33421), .B(g18485), .Z(g33594) ) ;
DFF     gate2757  (.D(g33594), .CP(CLK), .Q(g2495) ) ;
OR2     gate2758  (.A(g33901), .B(g18488), .Z(g34013) ) ;
DFF     gate2759  (.D(g34013), .CP(CLK), .Q(g2509) ) ;
OR2     gate2760  (.A(g33368), .B(g18489), .Z(g33595) ) ;
DFF     gate2761  (.D(g33595), .CP(CLK), .Q(g2514) ) ;
OR2     gate2762  (.A(g33647), .B(g18493), .Z(g34014) ) ;
DFF     gate2763  (.D(g34014), .CP(CLK), .Q(g2433) ) ;
OR2     gate2764  (.A(g33849), .B(g18476), .Z(g34008) ) ;
DFF     gate2765  (.D(g34008), .CP(CLK), .Q(g2429) ) ;
OR2     gate2766  (.A(g33863), .B(g18477), .Z(g34009) ) ;
DFF     gate2767  (.D(g34009), .CP(CLK), .Q(g2437) ) ;
OR2     gate2768  (.A(g33886), .B(g18480), .Z(g34012) ) ;
DFF     gate2769  (.D(g34012), .CP(CLK), .Q(g2449) ) ;
OR2     gate2770  (.A(g33884), .B(g18479), .Z(g34011) ) ;
DFF     gate2771  (.D(g34011), .CP(CLK), .Q(g2445) ) ;
OR2     gate2772  (.A(g33872), .B(g18478), .Z(g34010) ) ;
DFF     gate2773  (.D(g34010), .CP(CLK), .Q(g2441) ) ;
OR2     gate2774  (.A(g30125), .B(g18487), .Z(g30378) ) ;
DFF     gate2775  (.D(g30378), .CP(CLK), .Q(g2461) ) ;
OR2     gate2776  (.A(g32338), .B(g18481), .Z(g33011) ) ;
DFF     gate2777  (.D(g33011), .CP(CLK), .Q(g2453) ) ;
OR2     gate2778  (.A(g32274), .B(g18483), .Z(g33012) ) ;
DFF     gate2779  (.D(g33012), .CP(CLK), .Q(g2476) ) ;
OR2     gate2780  (.A(g32305), .B(g18499), .Z(g33014) ) ;
DFF     gate2781  (.D(g33014), .CP(CLK), .Q(g2491) ) ;
OR2     gate2782  (.A(g32283), .B(g18484), .Z(g33013) ) ;
DFF     gate2783  (.D(g33013), .CP(CLK), .Q(g2485) ) ;
OR2     gate2784  (.A(g28712), .B(g18486), .Z(g29252) ) ;
DFF     gate2785  (.D(g29252), .CP(CLK), .Q(g2504) ) ;
OR2     gate2786  (.A(g28697), .B(g18490), .Z(g29253) ) ;
DFF     gate2787  (.D(g29253), .CP(CLK), .Q(g2518) ) ;
OR2     gate2788  (.A(g30089), .B(g18491), .Z(g30379) ) ;
DFF     gate2789  (.D(g30379), .CP(CLK), .Q(g2523) ) ;
OR2     gate2790  (.A(g30161), .B(g18492), .Z(g30380) ) ;
DFF     gate2791  (.D(g30380), .CP(CLK), .Q(g2527) ) ;
OR2     gate2792  (.A(g33341), .B(g18494), .Z(g33596) ) ;
DFF     gate2793  (.D(g33596), .CP(CLK), .Q(g2533) ) ;
OR2     gate2794  (.A(g33344), .B(g18495), .Z(g33597) ) ;
DFF     gate2795  (.D(g33597), .CP(CLK), .Q(g2537) ) ;
OR2     gate2796  (.A(g33364), .B(g18496), .Z(g33598) ) ;
DFF     gate2797  (.D(g33598), .CP(CLK), .Q(g2541) ) ;
OR2     gate2798  (.A(g30126), .B(g18497), .Z(g30381) ) ;
DFF     gate2799  (.D(g30381), .CP(CLK), .Q(g2547) ) ;
OR2     gate2800  (.A(g30137), .B(g18498), .Z(g30382) ) ;
DFF     gate2801  (.D(g30382), .CP(CLK), .Q(g2551) ) ;
OR2     gate2802  (.A(g33418), .B(g18501), .Z(g33600) ) ;
DFF     gate2803  (.D(g33600), .CP(CLK), .Q(g2555) ) ;
OR2     gate2804  (.A(g33091), .B(g18526), .Z(g33607) ) ;
DFF     gate2805  (.D(g33607), .CP(CLK), .Q(g2606) ) ;
OR2     gate2806  (.A(g33422), .B(g18508), .Z(g33601) ) ;
DFF     gate2807  (.D(g33601), .CP(CLK), .Q(g2599) ) ;
OR2     gate2808  (.A(g33425), .B(g18511), .Z(g33602) ) ;
DFF     gate2809  (.D(g33602), .CP(CLK), .Q(g2629) ) ;
OR2     gate2810  (.A(g33904), .B(g18514), .Z(g34020) ) ;
DFF     gate2811  (.D(g34020), .CP(CLK), .Q(g2643) ) ;
OR2     gate2812  (.A(g33372), .B(g18515), .Z(g33603) ) ;
DFF     gate2813  (.D(g33603), .CP(CLK), .Q(g2648) ) ;
OR2     gate2814  (.A(g33652), .B(g18519), .Z(g34021) ) ;
DFF     gate2815  (.D(g34021), .CP(CLK), .Q(g2567) ) ;
OR2     gate2816  (.A(g33858), .B(g18502), .Z(g34015) ) ;
DFF     gate2817  (.D(g34015), .CP(CLK), .Q(g2563) ) ;
OR2     gate2818  (.A(g33867), .B(g18503), .Z(g34016) ) ;
DFF     gate2819  (.D(g34016), .CP(CLK), .Q(g2571) ) ;
OR2     gate2820  (.A(g33889), .B(g18506), .Z(g34019) ) ;
DFF     gate2821  (.D(g34019), .CP(CLK), .Q(g2583) ) ;
OR2     gate2822  (.A(g33887), .B(g18505), .Z(g34018) ) ;
DFF     gate2823  (.D(g34018), .CP(CLK), .Q(g2579) ) ;
OR2     gate2824  (.A(g33880), .B(g18504), .Z(g34017) ) ;
DFF     gate2825  (.D(g34017), .CP(CLK), .Q(g2575) ) ;
OR2     gate2826  (.A(g30138), .B(g18513), .Z(g30383) ) ;
DFF     gate2827  (.D(g30383), .CP(CLK), .Q(g2595) ) ;
OR2     gate2828  (.A(g32343), .B(g18507), .Z(g33015) ) ;
DFF     gate2829  (.D(g33015), .CP(CLK), .Q(g2587) ) ;
OR2     gate2830  (.A(g32284), .B(g18509), .Z(g33016) ) ;
DFF     gate2831  (.D(g33016), .CP(CLK), .Q(g2610) ) ;
OR2     gate2832  (.A(g32312), .B(g18525), .Z(g33018) ) ;
DFF     gate2833  (.D(g33018), .CP(CLK), .Q(g2625) ) ;
OR2     gate2834  (.A(g32292), .B(g18510), .Z(g33017) ) ;
DFF     gate2835  (.D(g33017), .CP(CLK), .Q(g2619) ) ;
OR2     gate2836  (.A(g28725), .B(g18512), .Z(g29254) ) ;
DFF     gate2837  (.D(g29254), .CP(CLK), .Q(g2638) ) ;
OR2     gate2838  (.A(g28714), .B(g18516), .Z(g29255) ) ;
DFF     gate2839  (.D(g29255), .CP(CLK), .Q(g2652) ) ;
OR2     gate2840  (.A(g30101), .B(g18517), .Z(g30384) ) ;
DFF     gate2841  (.D(g30384), .CP(CLK), .Q(g2657) ) ;
OR2     gate2842  (.A(g30172), .B(g18518), .Z(g30385) ) ;
DFF     gate2843  (.D(g30385), .CP(CLK), .Q(g2661) ) ;
OR2     gate2844  (.A(g33345), .B(g18520), .Z(g33604) ) ;
DFF     gate2845  (.D(g33604), .CP(CLK), .Q(g2667) ) ;
OR2     gate2846  (.A(g33352), .B(g18521), .Z(g33605) ) ;
DFF     gate2847  (.D(g33605), .CP(CLK), .Q(g2671) ) ;
OR2     gate2848  (.A(g33369), .B(g18522), .Z(g33606) ) ;
DFF     gate2849  (.D(g33606), .CP(CLK), .Q(g2675) ) ;
OR2     gate2850  (.A(g30139), .B(g18523), .Z(g30386) ) ;
DFF     gate2851  (.D(g30386), .CP(CLK), .Q(g2681) ) ;
OR2     gate2852  (.A(g30151), .B(g18524), .Z(g30387) ) ;
DFF     gate2853  (.D(g30387), .CP(CLK), .Q(g2685) ) ;
OR2     gate2854  (.A(g34564), .B(g15080), .Z(g34606) ) ;
DFF     gate2855  (.D(g34606), .CP(CLK), .Q(g2689) ) ;
OR2     gate2856  (.A(g34567), .B(g15081), .Z(g34607) ) ;
DFF     gate2857  (.D(g34607), .CP(CLK), .Q(g2697) ) ;
OR2     gate2858  (.A(g34568), .B(g15082), .Z(g34608) ) ;
DFF     gate2859  (.D(g34608), .CP(CLK), .Q(g2704) ) ;
INV     gate2860  (.A(II19345), .Z(g18527) ) ;
DFF     gate2861  (.D(g18527), .CP(CLK), .Q(g2710) ) ;
INV     gate2862  (.A(II19348), .Z(g18528) ) ;
DFF     gate2863  (.D(g18528), .CP(CLK), .Q(g2711) ) ;
INV     gate2864  (.A(II25677), .Z(g26935) ) ;
DFF     gate2865  (.D(g26935), .CP(CLK), .Q(g2837) ) ;
INV     gate2866  (.A(II25680), .Z(g26936) ) ;
DFF     gate2867  (.D(g26936), .CP(CLK), .Q(g2841) ) ;
INV     gate2868  (.A(II25683), .Z(g26937) ) ;
DFF     gate2869  (.D(g26937), .CP(CLK), .Q(g2712) ) ;
OR2     gate2870  (.A(g23497), .B(g18529), .Z(g24263) ) ;
DFF     gate2871  (.D(g24263), .CP(CLK), .Q(g2715) ) ;
OR2     gate2872  (.A(g25122), .B(g18530), .Z(g25639) ) ;
DFF     gate2873  (.D(g25639), .CP(CLK), .Q(g2719) ) ;
OR2     gate2874  (.A(g26633), .B(g18531), .Z(g26926) ) ;
DFF     gate2875  (.D(g26926), .CP(CLK), .Q(g2724) ) ;
OR2     gate2876  (.A(g27616), .B(g18532), .Z(g28060) ) ;
DFF     gate2877  (.D(g28060), .CP(CLK), .Q(g2729) ) ;
OR2     gate2878  (.A(g28597), .B(g18533), .Z(g29256) ) ;
DFF     gate2879  (.D(g29256), .CP(CLK), .Q(g2735) ) ;
OR2     gate2880  (.A(g30023), .B(g18534), .Z(g30388) ) ;
DFF     gate2881  (.D(g30388), .CP(CLK), .Q(g2741) ) ;
OR2     gate2882  (.A(g31524), .B(g18535), .Z(g31872) ) ;
DFF     gate2883  (.D(g31872), .CP(CLK), .Q(g2748) ) ;
OR2     gate2884  (.A(g32339), .B(g18536), .Z(g33019) ) ;
DFF     gate2885  (.D(g33019), .CP(CLK), .Q(g2756) ) ;
OR2     gate2886  (.A(g33322), .B(g18537), .Z(g33608) ) ;
DFF     gate2887  (.D(g33608), .CP(CLK), .Q(g2759) ) ;
OR2     gate2888  (.A(g33873), .B(g18538), .Z(g34022) ) ;
DFF     gate2889  (.D(g34022), .CP(CLK), .Q(g2763) ) ;
OR2     gate2890  (.A(g26711), .B(g18539), .Z(g26927) ) ;
DFF     gate2891  (.D(g26927), .CP(CLK), .Q(g2767) ) ;
OR2     gate2892  (.A(g26713), .B(g18541), .Z(g26928) ) ;
DFF     gate2893  (.D(g26928), .CP(CLK), .Q(g2779) ) ;
OR2     gate2894  (.A(g26635), .B(g18543), .Z(g26929) ) ;
DFF     gate2895  (.D(g26929), .CP(CLK), .Q(g2791) ) ;
OR2     gate2896  (.A(g26799), .B(g18544), .Z(g26930) ) ;
DFF     gate2897  (.D(g26930), .CP(CLK), .Q(g2795) ) ;
OR2     gate2898  (.A(g34389), .B(g18546), .Z(g34444) ) ;
DFF     gate2899  (.D(g34444), .CP(CLK), .Q(g2787) ) ;
OR2     gate2900  (.A(g34380), .B(g18542), .Z(g34442) ) ;
DFF     gate2901  (.D(g34442), .CP(CLK), .Q(g2783) ) ;
OR2     gate2902  (.A(g34385), .B(g18545), .Z(g34443) ) ;
DFF     gate2903  (.D(g34443), .CP(CLK), .Q(g2775) ) ;
OR2     gate2904  (.A(g34381), .B(g18540), .Z(g34441) ) ;
DFF     gate2905  (.D(g34441), .CP(CLK), .Q(g2771) ) ;
OR2     gate2906  (.A(g30080), .B(g18557), .Z(g30391) ) ;
DFF     gate2907  (.D(g30391), .CP(CLK), .Q(g2831) ) ;
OR2     gate2908  (.A(g29969), .B(g18554), .Z(g30389) ) ;
DFF     gate2909  (.D(g30389), .CP(CLK), .Q(g121) ) ;
OR2     gate2910  (.A(g26778), .B(g18547), .Z(g26931) ) ;
DFF     gate2911  (.D(g26931), .CP(CLK), .Q(g2799) ) ;
OR2     gate2912  (.A(g26684), .B(g18549), .Z(g26932) ) ;
DFF     gate2913  (.D(g26932), .CP(CLK), .Q(g2811) ) ;
OR2     gate2914  (.A(g26808), .B(g18551), .Z(g26933) ) ;
DFF     gate2915  (.D(g26933), .CP(CLK), .Q(g2823) ) ;
OR2     gate2916  (.A(g26845), .B(g18556), .Z(g26934) ) ;
DFF     gate2917  (.D(g26934), .CP(CLK), .Q(g2827) ) ;
OR2     gate2918  (.A(g34365), .B(g18553), .Z(g34448) ) ;
DFF     gate2919  (.D(g34448), .CP(CLK), .Q(g2819) ) ;
OR2     gate2920  (.A(g34390), .B(g18550), .Z(g34446) ) ;
DFF     gate2921  (.D(g34446), .CP(CLK), .Q(g2815) ) ;
OR2     gate2922  (.A(g34363), .B(g18552), .Z(g34447) ) ;
DFF     gate2923  (.D(g34447), .CP(CLK), .Q(g2807) ) ;
OR2     gate2924  (.A(g34382), .B(g18548), .Z(g34445) ) ;
DFF     gate2925  (.D(g34445), .CP(CLK), .Q(g2803) ) ;
OR2     gate2926  (.A(g30091), .B(g18558), .Z(g30392) ) ;
DFF     gate2927  (.D(g30392), .CP(CLK), .Q(g2834) ) ;
OR2     gate2928  (.A(g29985), .B(g18555), .Z(g30390) ) ;
DFF     gate2929  (.D(g30390), .CP(CLK), .Q(g117) ) ;
OR2     gate2930  (.A(g34748), .B(g18594), .Z(g34805) ) ;
DFF     gate2931  (.D(g34805), .CP(CLK), .Q(g2999) ) ;
OR2     gate2932  (.A(g34686), .B(g18593), .Z(g34732) ) ;
DFF     gate2933  (.D(g34732), .CP(CLK), .Q(g2994) ) ;
OR2     gate2934  (.A(g34509), .B(g18592), .Z(g34624) ) ;
DFF     gate2935  (.D(g34624), .CP(CLK), .Q(g2988) ) ;
OR2     gate2936  (.A(g34519), .B(g18577), .Z(g34616) ) ;
DFF     gate2937  (.D(g34616), .CP(CLK), .Q(g2868) ) ;
OR2     gate2938  (.A(g34516), .B(g18576), .Z(g34615) ) ;
DFF     gate2939  (.D(g34615), .CP(CLK), .Q(g2873) ) ;
OR2     gate2940  (.A(g34751), .B(g18578), .Z(g34799) ) ;
DFF     gate2941  (.D(g34799), .CP(CLK), .Q(g2890) ) ;
OR2     gate2942  (.A(g34503), .B(g18563), .Z(g34609) ) ;
DFF     gate2943  (.D(g34609), .CP(CLK), .Q(g2844) ) ;
OR2     gate2944  (.A(g34507), .B(g18564), .Z(g34610) ) ;
DFF     gate2945  (.D(g34610), .CP(CLK), .Q(g2852) ) ;
OR2     gate2946  (.A(g34508), .B(g18565), .Z(g34611) ) ;
DFF     gate2947  (.D(g34611), .CP(CLK), .Q(g2860) ) ;
OR2     gate2948  (.A(g34514), .B(g18566), .Z(g34612) ) ;
DFF     gate2949  (.D(g34612), .CP(CLK), .Q(g2894) ) ;
OR2     gate2950  (.A(g34515), .B(g18567), .Z(g34613) ) ;
DFF     gate2951  (.D(g34613), .CP(CLK), .Q(g37) ) ;
OR2     gate2952  (.A(g34518), .B(g18568), .Z(g34614) ) ;
DFF     gate2953  (.D(g34614), .CP(CLK), .Q(g94) ) ;
OR2     gate2954  (.A(g34750), .B(g18569), .Z(g34792) ) ;
DFF     gate2955  (.D(g34792), .CP(CLK), .Q(g2848) ) ;
OR2     gate2956  (.A(g34744), .B(g18570), .Z(g34793) ) ;
DFF     gate2957  (.D(g34793), .CP(CLK), .Q(g2856) ) ;
OR2     gate2958  (.A(g34746), .B(g18571), .Z(g34794) ) ;
DFF     gate2959  (.D(g34794), .CP(CLK), .Q(g2864) ) ;
OR2     gate2960  (.A(g34753), .B(g18572), .Z(g34795) ) ;
DFF     gate2961  (.D(g34795), .CP(CLK), .Q(g2898) ) ;
OR2     gate2962  (.A(g34745), .B(g18573), .Z(g34796) ) ;
DFF     gate2963  (.D(g34796), .CP(CLK), .Q(g2882) ) ;
OR2     gate2964  (.A(g34747), .B(g18574), .Z(g34797) ) ;
DFF     gate2965  (.D(g34797), .CP(CLK), .Q(g2878) ) ;
OR2     gate2966  (.A(g34754), .B(g18575), .Z(g34798) ) ;
DFF     gate2967  (.D(g34798), .CP(CLK), .Q(g2886) ) ;
OR2     gate2968  (.A(g34752), .B(g18586), .Z(g34800) ) ;
DFF     gate2969  (.D(g34800), .CP(CLK), .Q(g2980) ) ;
OR2     gate2970  (.A(g34969), .B(g18587), .Z(g34980) ) ;
DFF     gate2971  (.D(g34980), .CP(CLK), .Q(g2984) ) ;
OR2     gate2972  (.A(g34526), .B(g18579), .Z(g34617) ) ;
DFF     gate2973  (.D(g34617), .CP(CLK), .Q(g2907) ) ;
OR2     gate2974  (.A(g34527), .B(g18580), .Z(g34618) ) ;
DFF     gate2975  (.D(g34618), .CP(CLK), .Q(g2912) ) ;
OR2     gate2976  (.A(g34528), .B(g18581), .Z(g34619) ) ;
DFF     gate2977  (.D(g34619), .CP(CLK), .Q(g2922) ) ;
OR2     gate2978  (.A(g34529), .B(g18582), .Z(g34620) ) ;
DFF     gate2979  (.D(g34620), .CP(CLK), .Q(g2936) ) ;
OR2     gate2980  (.A(g34517), .B(g18583), .Z(g34621) ) ;
DFF     gate2981  (.D(g34621), .CP(CLK), .Q(g2950) ) ;
OR2     gate2982  (.A(g34520), .B(g18584), .Z(g34622) ) ;
DFF     gate2983  (.D(g34622), .CP(CLK), .Q(g2960) ) ;
OR2     gate2984  (.A(g34525), .B(g18585), .Z(g34623) ) ;
DFF     gate2985  (.D(g34623), .CP(CLK), .Q(g2970) ) ;
OR2     gate2986  (.A(g34756), .B(g18588), .Z(g34801) ) ;
DFF     gate2987  (.D(g34801), .CP(CLK), .Q(g2902) ) ;
OR2     gate2988  (.A(g34757), .B(g18589), .Z(g34802) ) ;
DFF     gate2989  (.D(g34802), .CP(CLK), .Q(g2917) ) ;
OR2     gate2990  (.A(g34758), .B(g18590), .Z(g34803) ) ;
DFF     gate2991  (.D(g34803), .CP(CLK), .Q(g2927) ) ;
OR2     gate2992  (.A(g34763), .B(g18595), .Z(g34806) ) ;
DFF     gate2993  (.D(g34806), .CP(CLK), .Q(g2941) ) ;
OR2     gate2994  (.A(g34764), .B(g18596), .Z(g34807) ) ;
DFF     gate2995  (.D(g34807), .CP(CLK), .Q(g2955) ) ;
OR2     gate2996  (.A(g34765), .B(g18599), .Z(g34808) ) ;
DFF     gate2997  (.D(g34808), .CP(CLK), .Q(g2965) ) ;
OR2     gate2998  (.A(g34740), .B(g18591), .Z(g34804) ) ;
DFF     gate2999  (.D(g34804), .CP(CLK), .Q(g2975) ) ;
INV     gate3000  (.A(II21297), .Z(g21726) ) ;
DFF     gate3001  (.D(g21726), .CP(CLK), .Q(g3003) ) ;
INV     gate3002  (.A(II15448), .Z(g12833) ) ;
DFF     gate3003  (.D(g12833), .CP(CLK), .Q(g5) ) ;
INV     gate3004  (.A(II32675), .Z(g34589) ) ;
DFF     gate3005  (.D(g34589), .CP(CLK), .Q(g6) ) ;
INV     gate3006  (.A(II32678), .Z(g34590) ) ;
DFF     gate3007  (.D(g34590), .CP(CLK), .Q(g7) ) ;
INV     gate3008  (.A(II32681), .Z(g34591) ) ;
DFF     gate3009  (.D(g34591), .CP(CLK), .Q(g8) ) ;
INV     gate3010  (.A(II32684), .Z(g34592) ) ;
DFF     gate3011  (.D(g34592), .CP(CLK), .Q(g9) ) ;
INV     gate3012  (.A(II32687), .Z(g34593) ) ;
DFF     gate3013  (.D(g34593), .CP(CLK), .Q(g16) ) ;
INV     gate3014  (.A(II32690), .Z(g34594) ) ;
DFF     gate3015  (.D(g34594), .CP(CLK), .Q(g19) ) ;
INV     gate3016  (.A(II32693), .Z(g34595) ) ;
DFF     gate3017  (.D(g34595), .CP(CLK), .Q(g28) ) ;
INV     gate3018  (.A(II32696), .Z(g34596) ) ;
DFF     gate3019  (.D(g34596), .CP(CLK), .Q(g31) ) ;
INV     gate3020  (.A(II33103), .Z(g34877) ) ;
DFF     gate3021  (.D(g34877), .CP(CLK), .Q(g34) ) ;
INV     gate3022  (.A(II28579), .Z(g30326) ) ;
DFF     gate3023  (.D(g30326), .CP(CLK), .Q(g12) ) ;
INV     gate3024  (.A(II27543), .Z(g29209) ) ;
DFF     gate3025  (.D(g29209), .CP(CLK), .Q(g22) ) ;
INV     gate3026  (.A(II16969), .Z(g15048) ) ;
DFF     gate3027  (.D(g15048), .CP(CLK), .Q(g25) ) ;
INV     gate3028  (.A(g1), .Z(II11617) ) ;
INV     gate3029  (.A(II11617), .Z(g6754) ) ;
INV     gate3030  (.A(g1), .Z(II11620) ) ;
INV     gate3031  (.A(II11620), .Z(g6755) ) ;
INV     gate3032  (.A(g28), .Z(II11623) ) ;
INV     gate3033  (.A(II11623), .Z(g6756) ) ;
INV     gate3034  (.A(g31), .Z(II11626) ) ;
INV     gate3035  (.A(II11626), .Z(g6767) ) ;
INV     gate3036  (.A(g19), .Z(II11629) ) ;
INV     gate3037  (.A(II11629), .Z(g6772) ) ;
INV     gate3038  (.A(g16), .Z(II11632) ) ;
INV     gate3039  (.A(II11632), .Z(g6782) ) ;
INV     gate3040  (.A(g9), .Z(II11635) ) ;
INV     gate3041  (.A(II11635), .Z(g6789) ) ;
INV     gate3042  (.A(g199), .Z(g6799) ) ;
INV     gate3043  (.A(g203), .Z(g6800) ) ;
INV     gate3044  (.A(g391), .Z(g6801) ) ;
INV     gate3045  (.A(g468), .Z(g6802) ) ;
INV     gate3046  (.A(g496), .Z(g6803) ) ;
INV     gate3047  (.A(g490), .Z(g6804) ) ;
INV     gate3048  (.A(g554), .Z(g6808) ) ;
INV     gate3049  (.A(g341), .Z(g6809) ) ;
INV     gate3050  (.A(g723), .Z(g6810) ) ;
INV     gate3051  (.A(g714), .Z(g6811) ) ;
INV     gate3052  (.A(g632), .Z(g6814) ) ;
INV     gate3053  (.A(g929), .Z(g6815) ) ;
INV     gate3054  (.A(g933), .Z(g6816) ) ;
INV     gate3055  (.A(g956), .Z(g6817) ) ;
INV     gate3056  (.A(g976), .Z(g6818) ) ;
INV     gate3057  (.A(g1046), .Z(g6819) ) ;
INV     gate3058  (.A(g1070), .Z(g6820) ) ;
INV     gate3059  (.A(g1246), .Z(II11655) ) ;
INV     gate3060  (.A(II11655), .Z(g6821) ) ;
INV     gate3061  (.A(g979), .Z(g6825) ) ;
INV     gate3062  (.A(g218), .Z(g6826) ) ;
INV     gate3063  (.A(g1277), .Z(g6827) ) ;
INV     gate3064  (.A(g1300), .Z(g6828) ) ;
INV     gate3065  (.A(g1319), .Z(g6829) ) ;
INV     gate3066  (.A(g1389), .Z(g6830) ) ;
INV     gate3067  (.A(g1413), .Z(g6831) ) ;
INV     gate3068  (.A(g1589), .Z(II11665) ) ;
INV     gate3069  (.A(II11665), .Z(g6832) ) ;
INV     gate3070  (.A(g1322), .Z(g6836) ) ;
INV     gate3071  (.A(g968), .Z(g6837) ) ;
INV     gate3072  (.A(g1724), .Z(g6838) ) ;
INV     gate3073  (.A(g1858), .Z(g6839) ) ;
INV     gate3074  (.A(g1992), .Z(g6840) ) ;
INV     gate3075  (.A(g2145), .Z(g6841) ) ;
INV     gate3076  (.A(g2126), .Z(g6845) ) ;
INV     gate3077  (.A(g2152), .Z(g6846) ) ;
INV     gate3078  (.A(g2283), .Z(g6847) ) ;
INV     gate3079  (.A(g2417), .Z(g6848) ) ;
INV     gate3080  (.A(g2551), .Z(g6849) ) ;
INV     gate3081  (.A(g2704), .Z(g6850) ) ;
INV     gate3082  (.A(g2685), .Z(g6854) ) ;
INV     gate3083  (.A(g2711), .Z(g6855) ) ;
INV     gate3084  (.A(g2756), .Z(II11682) ) ;
INV     gate3085  (.A(II11682), .Z(g6856) ) ;
INV     gate3086  (.A(g117), .Z(II11685) ) ;
INV     gate3087  (.A(II11685), .Z(g6867) ) ;
INV     gate3088  (.A(g70), .Z(II11688) ) ;
INV     gate3089  (.A(II11688), .Z(g6868) ) ;
INV     gate3090  (.A(g36), .Z(II11691) ) ;
INV     gate3091  (.A(II11691), .Z(g6869) ) ;
INV     gate3092  (.A(g3089), .Z(g6870) ) ;
INV     gate3093  (.A(g3151), .Z(g6873) ) ;
INV     gate3094  (.A(g3143), .Z(g6874) ) ;
INV     gate3095  (.A(g3352), .Z(II11697) ) ;
INV     gate3096  (.A(II11697), .Z(g6875) ) ;
INV     gate3097  (.A(g3333), .Z(g6887) ) ;
INV     gate3098  (.A(g4164), .Z(II11701) ) ;
INV     gate3099  (.A(II11701), .Z(g6888) ) ;
INV     gate3100  (.A(g3288), .Z(g6895) ) ;
INV     gate3101  (.A(g3440), .Z(g6900) ) ;
INV     gate3102  (.A(g3502), .Z(g6903) ) ;
INV     gate3103  (.A(g3494), .Z(g6904) ) ;
INV     gate3104  (.A(g3703), .Z(II11708) ) ;
INV     gate3105  (.A(II11708), .Z(g6905) ) ;
INV     gate3106  (.A(g3684), .Z(g6917) ) ;
INV     gate3107  (.A(g3639), .Z(g6918) ) ;
INV     gate3108  (.A(g3791), .Z(g6923) ) ;
INV     gate3109  (.A(g3853), .Z(g6926) ) ;
INV     gate3110  (.A(g3845), .Z(g6927) ) ;
INV     gate3111  (.A(g4054), .Z(II11716) ) ;
INV     gate3112  (.A(II11716), .Z(g6928) ) ;
INV     gate3113  (.A(g4035), .Z(g6940) ) ;
INV     gate3114  (.A(g3990), .Z(g6941) ) ;
INV     gate3115  (.A(g4145), .Z(II11721) ) ;
INV     gate3116  (.A(II11721), .Z(g6946) ) ;
INV     gate3117  (.A(g4157), .Z(g6953) ) ;
INV     gate3118  (.A(g4138), .Z(g6954) ) ;
INV     gate3119  (.A(g4273), .Z(II11726) ) ;
INV     gate3120  (.A(II11726), .Z(g6955) ) ;
INV     gate3121  (.A(g4242), .Z(g6956) ) ;
INV     gate3122  (.A(g2932), .Z(g6957) ) ;
INV     gate3123  (.A(g4372), .Z(g6958) ) ;
INV     gate3124  (.A(g4420), .Z(g6959) ) ;
INV     gate3125  (.A(g1), .Z(g6960) ) ;
INV     gate3126  (.A(g4473), .Z(II11734) ) ;
INV     gate3127  (.A(II11734), .Z(g6961) ) ;
INV     gate3128  (.A(g4467), .Z(II11737) ) ;
INV     gate3129  (.A(II11737), .Z(g6971) ) ;
INV     gate3130  (.A(g4519), .Z(II11740) ) ;
INV     gate3131  (.A(g4564), .Z(II11743) ) ;
INV     gate3132  (.A(II11743), .Z(g6973) ) ;
INV     gate3133  (.A(g4570), .Z(II11746) ) ;
INV     gate3134  (.A(g4507), .Z(g6975) ) ;
INV     gate3135  (.A(g4474), .Z(II11750) ) ;
INV     gate3136  (.A(II11750), .Z(g6976) ) ;
INV     gate3137  (.A(g4492), .Z(II11753) ) ;
INV     gate3138  (.A(II11753), .Z(g6977) ) ;
INV     gate3139  (.A(g4616), .Z(g6978) ) ;
INV     gate3140  (.A(g4531), .Z(g6982) ) ;
INV     gate3141  (.A(g4698), .Z(g6983) ) ;
INV     gate3142  (.A(g4709), .Z(g6984) ) ;
INV     gate3143  (.A(g4669), .Z(g6985) ) ;
INV     gate3144  (.A(g4743), .Z(g6986) ) ;
INV     gate3145  (.A(g4754), .Z(g6987) ) ;
INV     gate3146  (.A(g4765), .Z(g6988) ) ;
INV     gate3147  (.A(g4575), .Z(g6989) ) ;
INV     gate3148  (.A(g4742), .Z(g6990) ) ;
INV     gate3149  (.A(g4888), .Z(g6991) ) ;
INV     gate3150  (.A(g4899), .Z(g6992) ) ;
INV     gate3151  (.A(g4859), .Z(g6993) ) ;
INV     gate3152  (.A(g4933), .Z(g6994) ) ;
INV     gate3153  (.A(g4944), .Z(g6995) ) ;
INV     gate3154  (.A(g4955), .Z(g6996) ) ;
INV     gate3155  (.A(g4578), .Z(g6997) ) ;
INV     gate3156  (.A(g4932), .Z(g6998) ) ;
INV     gate3157  (.A(g86), .Z(g6999) ) ;
INV     gate3158  (.A(g5160), .Z(g7002) ) ;
INV     gate3159  (.A(g5152), .Z(g7003) ) ;
INV     gate3160  (.A(g5357), .Z(II11777) ) ;
INV     gate3161  (.A(II11777), .Z(g7004) ) ;
INV     gate3162  (.A(g128), .Z(g7017) ) ;
INV     gate3163  (.A(g5297), .Z(g7018) ) ;
INV     gate3164  (.A(g5445), .Z(g7023) ) ;
INV     gate3165  (.A(g5507), .Z(g7026) ) ;
INV     gate3166  (.A(g5499), .Z(g7027) ) ;
INV     gate3167  (.A(g5703), .Z(II11785) ) ;
INV     gate3168  (.A(II11785), .Z(g7028) ) ;
INV     gate3169  (.A(g4821), .Z(g7040) ) ;
INV     gate3170  (.A(g5644), .Z(g7041) ) ;
INV     gate3171  (.A(g5791), .Z(g7046) ) ;
INV     gate3172  (.A(g5853), .Z(g7049) ) ;
INV     gate3173  (.A(g5845), .Z(g7050) ) ;
INV     gate3174  (.A(g6049), .Z(II11793) ) ;
INV     gate3175  (.A(II11793), .Z(g7051) ) ;
INV     gate3176  (.A(g4831), .Z(g7063) ) ;
INV     gate3177  (.A(g5990), .Z(g7064) ) ;
INV     gate3178  (.A(g6137), .Z(g7069) ) ;
INV     gate3179  (.A(g6199), .Z(g7072) ) ;
INV     gate3180  (.A(g6191), .Z(g7073) ) ;
INV     gate3181  (.A(g6395), .Z(II11801) ) ;
INV     gate3182  (.A(II11801), .Z(g7074) ) ;
INV     gate3183  (.A(g4826), .Z(g7086) ) ;
INV     gate3184  (.A(g6336), .Z(g7087) ) ;
INV     gate3185  (.A(g6483), .Z(g7092) ) ;
INV     gate3186  (.A(g6545), .Z(g7095) ) ;
INV     gate3187  (.A(g6537), .Z(g7096) ) ;
INV     gate3188  (.A(g6741), .Z(II11809) ) ;
INV     gate3189  (.A(II11809), .Z(g7097) ) ;
INV     gate3190  (.A(g5011), .Z(g7109) ) ;
INV     gate3191  (.A(g6682), .Z(g7110) ) ;
INV     gate3192  (.A(g12), .Z(g7115) ) ;
INV     gate3193  (.A(g22), .Z(g7116) ) ;
INV     gate3194  (.A(g93), .Z(II11816) ) ;
INV     gate3195  (.A(II11816), .Z(g7117) ) ;
INV     gate3196  (.A(g832), .Z(g7118) ) ;
INV     gate3197  (.A(g3869), .Z(II11820) ) ;
INV     gate3198  (.A(II11820), .Z(g7121) ) ;
INV     gate3199  (.A(g4558), .Z(g7132) ) ;
INV     gate3200  (.A(g5029), .Z(g7134) ) ;
INV     gate3201  (.A(g5360), .Z(g7138) ) ;
INV     gate3202  (.A(g101), .Z(II11835) ) ;
INV     gate3203  (.A(II11835), .Z(g7148) ) ;
INV     gate3204  (.A(g4564), .Z(g7149) ) ;
INV     gate3205  (.A(g5373), .Z(g7153) ) ;
INV     gate3206  (.A(g5706), .Z(g7157) ) ;
INV     gate3207  (.A(g111), .Z(II11843) ) ;
INV     gate3208  (.A(II11843), .Z(g7161) ) ;
INV     gate3209  (.A(g4521), .Z(g7162) ) ;
INV     gate3210  (.A(g4593), .Z(g7163) ) ;
INV     gate3211  (.A(g4311), .Z(g7166) ) ;
INV     gate3212  (.A(g5719), .Z(g7170) ) ;
INV     gate3213  (.A(g6052), .Z(g7174) ) ;
INV     gate3214  (.A(g4392), .Z(g7178) ) ;
INV     gate3215  (.A(g4608), .Z(g7183) ) ;
INV     gate3216  (.A(g6065), .Z(g7187) ) ;
INV     gate3217  (.A(g6398), .Z(g7191) ) ;
INV     gate3218  (.A(g25), .Z(g7195) ) ;
INV     gate3219  (.A(g43), .Z(II11860) ) ;
INV     gate3220  (.A(II11860), .Z(g7196) ) ;
INV     gate3221  (.A(g812), .Z(g7197) ) ;
INV     gate3222  (.A(g4639), .Z(g7202) ) ;
INV     gate3223  (.A(g6411), .Z(g7212) ) ;
INV     gate3224  (.A(g822), .Z(g7216) ) ;
INV     gate3225  (.A(g4405), .Z(g7219) ) ;
INV     gate3226  (.A(g4427), .Z(g7222) ) ;
INV     gate3227  (.A(g4601), .Z(g7224) ) ;
INV     gate3228  (.A(g5), .Z(g7231) ) ;
INV     gate3229  (.A(g4411), .Z(g7232) ) ;
INV     gate3230  (.A(g4521), .Z(g7235) ) ;
INV     gate3231  (.A(g4608), .Z(g7236) ) ;
INV     gate3232  (.A(g5033), .Z(g7239) ) ;
INV     gate3233  (.A(g4408), .Z(II11892) ) ;
INV     gate3234  (.A(g4408), .Z(g7244) ) ;
INV     gate3235  (.A(g4446), .Z(II11896) ) ;
INV     gate3236  (.A(g4446), .Z(g7246) ) ;
INV     gate3237  (.A(g5377), .Z(g7247) ) ;
INV     gate3238  (.A(g1592), .Z(g7252) ) ;
INV     gate3239  (.A(g4414), .Z(II11903) ) ;
INV     gate3240  (.A(g4414), .Z(g7258) ) ;
INV     gate3241  (.A(g4375), .Z(g7259) ) ;
INV     gate3242  (.A(g4449), .Z(II11908) ) ;
INV     gate3243  (.A(g4449), .Z(g7261) ) ;
INV     gate3244  (.A(g5723), .Z(g7262) ) ;
INV     gate3245  (.A(g35), .Z(g7266) ) ;
INV     gate3246  (.A(g1604), .Z(g7267) ) ;
INV     gate3247  (.A(g1636), .Z(g7268) ) ;
INV     gate3248  (.A(g1728), .Z(g7275) ) ;
INV     gate3249  (.A(g2153), .Z(g7280) ) ;
INV     gate3250  (.A(g4643), .Z(g7285) ) ;
INV     gate3251  (.A(g4382), .Z(g7289) ) ;
INV     gate3252  (.A(g4452), .Z(g7293) ) ;
INV     gate3253  (.A(g5313), .Z(g7296) ) ;
INV     gate3254  (.A(g6069), .Z(g7297) ) ;
INV     gate3255  (.A(g925), .Z(g7301) ) ;
INV     gate3256  (.A(g1668), .Z(g7308) ) ;
INV     gate3257  (.A(g1740), .Z(g7314) ) ;
INV     gate3258  (.A(g1772), .Z(g7315) ) ;
INV     gate3259  (.A(g1862), .Z(g7322) ) ;
INV     gate3260  (.A(g2165), .Z(g7327) ) ;
INV     gate3261  (.A(g2197), .Z(g7328) ) ;
INV     gate3262  (.A(g2287), .Z(g7335) ) ;
INV     gate3263  (.A(g4443), .Z(g7340) ) ;
INV     gate3264  (.A(g5290), .Z(g7343) ) ;
INV     gate3265  (.A(g5659), .Z(g7344) ) ;
INV     gate3266  (.A(g6415), .Z(g7345) ) ;
INV     gate3267  (.A(g1270), .Z(g7349) ) ;
INV     gate3268  (.A(g1802), .Z(g7356) ) ;
INV     gate3269  (.A(g1874), .Z(g7361) ) ;
INV     gate3270  (.A(g1906), .Z(g7362) ) ;
INV     gate3271  (.A(g1996), .Z(g7369) ) ;
INV     gate3272  (.A(g2227), .Z(g7374) ) ;
INV     gate3273  (.A(g2299), .Z(g7379) ) ;
INV     gate3274  (.A(g2331), .Z(g7380) ) ;
INV     gate3275  (.A(g2421), .Z(g7387) ) ;
INV     gate3276  (.A(g4438), .Z(g7392) ) ;
INV     gate3277  (.A(g5320), .Z(g7393) ) ;
INV     gate3278  (.A(g5637), .Z(g7394) ) ;
INV     gate3279  (.A(g6005), .Z(g7395) ) ;
INV     gate3280  (.A(g890), .Z(g7397) ) ;
INV     gate3281  (.A(g911), .Z(g7400) ) ;
INV     gate3282  (.A(g1936), .Z(g7405) ) ;
INV     gate3283  (.A(g2008), .Z(g7410) ) ;
INV     gate3284  (.A(g2040), .Z(g7411) ) ;
INV     gate3285  (.A(g2361), .Z(g7418) ) ;
INV     gate3286  (.A(g2433), .Z(g7423) ) ;
INV     gate3287  (.A(g2465), .Z(g7424) ) ;
INV     gate3288  (.A(g2555), .Z(g7431) ) ;
INV     gate3289  (.A(g5276), .Z(g7436) ) ;
INV     gate3290  (.A(g5666), .Z(g7437) ) ;
INV     gate3291  (.A(g5983), .Z(g7438) ) ;
INV     gate3292  (.A(g6351), .Z(g7439) ) ;
INV     gate3293  (.A(g329), .Z(g7440) ) ;
INV     gate3294  (.A(g862), .Z(g7441) ) ;
INV     gate3295  (.A(g914), .Z(g7443) ) ;
INV     gate3296  (.A(g1256), .Z(g7446) ) ;
INV     gate3297  (.A(g2070), .Z(g7451) ) ;
INV     gate3298  (.A(g2495), .Z(g7456) ) ;
INV     gate3299  (.A(g2567), .Z(g7461) ) ;
INV     gate3300  (.A(g2599), .Z(g7462) ) ;
INV     gate3301  (.A(g5623), .Z(g7470) ) ;
INV     gate3302  (.A(g6012), .Z(g7471) ) ;
INV     gate3303  (.A(g6329), .Z(g7472) ) ;
INV     gate3304  (.A(g6697), .Z(g7473) ) ;
INV     gate3305  (.A(g66), .Z(II11980) ) ;
INV     gate3306  (.A(II11980), .Z(g7474) ) ;
INV     gate3307  (.A(g896), .Z(g7475) ) ;
INV     gate3308  (.A(g1008), .Z(g7479) ) ;
INV     gate3309  (.A(g1259), .Z(g7487) ) ;
INV     gate3310  (.A(g2629), .Z(g7490) ) ;
INV     gate3311  (.A(g4375), .Z(g7495) ) ;
INV     gate3312  (.A(g5969), .Z(g7496) ) ;
INV     gate3313  (.A(g6358), .Z(g7497) ) ;
INV     gate3314  (.A(g6675), .Z(g7498) ) ;
INV     gate3315  (.A(g763), .Z(II11992) ) ;
INV     gate3316  (.A(II11992), .Z(g7502) ) ;
INV     gate3317  (.A(g1351), .Z(g7503) ) ;
INV     gate3318  (.A(g5283), .Z(g7512) ) ;
INV     gate3319  (.A(g6315), .Z(g7513) ) ;
INV     gate3320  (.A(g6704), .Z(g7514) ) ;
INV     gate3321  (.A(g582), .Z(II12000) ) ;
INV     gate3322  (.A(II12000), .Z(g7515) ) ;
INV     gate3323  (.A(g767), .Z(II12003) ) ;
INV     gate3324  (.A(II12003), .Z(g7516) ) ;
INV     gate3325  (.A(g962), .Z(g7517) ) ;
INV     gate3326  (.A(g1024), .Z(g7518) ) ;
INV     gate3327  (.A(g1157), .Z(g7519) ) ;
INV     gate3328  (.A(g5630), .Z(g7521) ) ;
INV     gate3329  (.A(g6661), .Z(g7522) ) ;
INV     gate3330  (.A(g305), .Z(g7523) ) ;
INV     gate3331  (.A(g590), .Z(II12013) ) ;
INV     gate3332  (.A(II12013), .Z(g7526) ) ;
INV     gate3333  (.A(g772), .Z(II12016) ) ;
INV     gate3334  (.A(II12016), .Z(g7527) ) ;
INV     gate3335  (.A(g930), .Z(g7528) ) ;
INV     gate3336  (.A(g1157), .Z(g7532) ) ;
INV     gate3337  (.A(g1306), .Z(g7533) ) ;
INV     gate3338  (.A(g1367), .Z(g7534) ) ;
INV     gate3339  (.A(g1500), .Z(g7535) ) ;
INV     gate3340  (.A(g5976), .Z(g7536) ) ;
INV     gate3341  (.A(g311), .Z(g7537) ) ;
INV     gate3342  (.A(g344), .Z(II12026) ) ;
INV     gate3343  (.A(g344), .Z(g7541) ) ;
INV     gate3344  (.A(g595), .Z(II12030) ) ;
INV     gate3345  (.A(II12030), .Z(g7542) ) ;
INV     gate3346  (.A(g776), .Z(II12033) ) ;
INV     gate3347  (.A(II12033), .Z(g7543) ) ;
INV     gate3348  (.A(g918), .Z(g7544) ) ;
INV     gate3349  (.A(g1036), .Z(g7548) ) ;
INV     gate3350  (.A(g1274), .Z(g7553) ) ;
INV     gate3351  (.A(g1500), .Z(g7557) ) ;
INV     gate3352  (.A(g2741), .Z(II12041) ) ;
INV     gate3353  (.A(II12041), .Z(g7558) ) ;
INV     gate3354  (.A(g6322), .Z(g7563) ) ;
INV     gate3355  (.A(g336), .Z(g7564) ) ;
INV     gate3356  (.A(g613), .Z(II12046) ) ;
INV     gate3357  (.A(II12046), .Z(g7565) ) ;
INV     gate3358  (.A(g781), .Z(II12049) ) ;
INV     gate3359  (.A(II12049), .Z(g7566) ) ;
INV     gate3360  (.A(g1263), .Z(g7577) ) ;
INV     gate3361  (.A(g1379), .Z(g7581) ) ;
INV     gate3362  (.A(g2748), .Z(II12056) ) ;
INV     gate3363  (.A(II12056), .Z(g7586) ) ;
INV     gate3364  (.A(g6668), .Z(g7591) ) ;
INV     gate3365  (.A(g347), .Z(g7592) ) ;
INV     gate3366  (.A(g562), .Z(II12061) ) ;
INV     gate3367  (.A(II12061), .Z(g7593) ) ;
INV     gate3368  (.A(g617), .Z(II12064) ) ;
INV     gate3369  (.A(II12064), .Z(g7594) ) ;
INV     gate3370  (.A(g739), .Z(II12067) ) ;
INV     gate3371  (.A(II12067), .Z(g7595) ) ;
INV     gate3372  (.A(g785), .Z(II12070) ) ;
INV     gate3373  (.A(II12070), .Z(g7596) ) ;
INV     gate3374  (.A(g952), .Z(g7597) ) ;
INV     gate3375  (.A(g568), .Z(II12083) ) ;
INV     gate3376  (.A(II12083), .Z(g7615) ) ;
INV     gate3377  (.A(g622), .Z(II12086) ) ;
INV     gate3378  (.A(II12086), .Z(g7616) ) ;
INV     gate3379  (.A(g744), .Z(II12089) ) ;
INV     gate3380  (.A(II12089), .Z(g7617) ) ;
INV     gate3381  (.A(g790), .Z(II12092) ) ;
INV     gate3382  (.A(II12092), .Z(g7618) ) ;
INV     gate3383  (.A(g1296), .Z(g7619) ) ;
INV     gate3384  (.A(g572), .Z(II12103) ) ;
INV     gate3385  (.A(II12103), .Z(g7623) ) ;
INV     gate3386  (.A(g626), .Z(II12106) ) ;
INV     gate3387  (.A(II12106), .Z(g7624) ) ;
INV     gate3388  (.A(g749), .Z(II12109) ) ;
INV     gate3389  (.A(II12109), .Z(g7625) ) ;
INV     gate3390  (.A(g794), .Z(II12112) ) ;
INV     gate3391  (.A(II12112), .Z(g7626) ) ;
INV     gate3392  (.A(g4311), .Z(g7627) ) ;
INV     gate3393  (.A(g74), .Z(g7631) ) ;
INV     gate3394  (.A(g586), .Z(II12117) ) ;
INV     gate3395  (.A(II12117), .Z(g7632) ) ;
INV     gate3396  (.A(g632), .Z(II12120) ) ;
INV     gate3397  (.A(II12120), .Z(g7633) ) ;
INV     gate3398  (.A(g758), .Z(II12123) ) ;
INV     gate3399  (.A(II12123), .Z(g7634) ) ;
INV     gate3400  (.A(g1002), .Z(g7635) ) ;
INV     gate3401  (.A(g4098), .Z(g7636) ) ;
INV     gate3402  (.A(g4253), .Z(II12128) ) ;
INV     gate3403  (.A(II12128), .Z(g7640) ) ;
INV     gate3404  (.A(g4322), .Z(g7643) ) ;
INV     gate3405  (.A(g577), .Z(II12132) ) ;
INV     gate3406  (.A(II12132), .Z(g7647) ) ;
INV     gate3407  (.A(g807), .Z(II12135) ) ;
INV     gate3408  (.A(II12135), .Z(g7648) ) ;
INV     gate3409  (.A(g1345), .Z(g7649) ) ;
INV     gate3410  (.A(g4064), .Z(g7650) ) ;
INV     gate3411  (.A(g4332), .Z(g7655) ) ;
INV     gate3412  (.A(g599), .Z(II12141) ) ;
INV     gate3413  (.A(II12141), .Z(g7659) ) ;
INV     gate3414  (.A(g554), .Z(II12144) ) ;
INV     gate3415  (.A(II12144), .Z(g7660) ) ;
INV     gate3416  (.A(g4076), .Z(g7666) ) ;
INV     gate3417  (.A(g4104), .Z(g7670) ) ;
INV     gate3418  (.A(g604), .Z(II12151) ) ;
INV     gate3419  (.A(II12151), .Z(g7674) ) ;
INV     gate3420  (.A(g4108), .Z(g7680) ) ;
INV     gate3421  (.A(g4659), .Z(g7686) ) ;
INV     gate3422  (.A(g608), .Z(II12159) ) ;
INV     gate3423  (.A(II12159), .Z(g7689) ) ;
INV     gate3424  (.A(g4849), .Z(g7693) ) ;
INV     gate3425  (.A(g4087), .Z(g7697) ) ;
INV     gate3426  (.A(g5176), .Z(II12167) ) ;
INV     gate3427  (.A(II12167), .Z(g7704) ) ;
INV     gate3428  (.A(g1178), .Z(g7715) ) ;
INV     gate3429  (.A(g1199), .Z(g7716) ) ;
INV     gate3430  (.A(g2715), .Z(II12172) ) ;
INV     gate3431  (.A(II12172), .Z(g7717) ) ;
INV     gate3432  (.A(g4093), .Z(g7733) ) ;
INV     gate3433  (.A(g5523), .Z(II12176) ) ;
INV     gate3434  (.A(II12176), .Z(g7738) ) ;
INV     gate3435  (.A(g996), .Z(g7749) ) ;
INV     gate3436  (.A(g1070), .Z(g7750) ) ;
INV     gate3437  (.A(g1521), .Z(g7751) ) ;
INV     gate3438  (.A(g1542), .Z(g7752) ) ;
INV     gate3439  (.A(g2719), .Z(II12183) ) ;
INV     gate3440  (.A(II12183), .Z(g7753) ) ;
INV     gate3441  (.A(g4165), .Z(g7765) ) ;
INV     gate3442  (.A(g5869), .Z(II12189) ) ;
INV     gate3443  (.A(II12189), .Z(g7766) ) ;
INV     gate3444  (.A(g1339), .Z(g7778) ) ;
INV     gate3445  (.A(g1413), .Z(g7779) ) ;
INV     gate3446  (.A(g2878), .Z(g7780) ) ;
INV     gate3447  (.A(g4621), .Z(g7785) ) ;
INV     gate3448  (.A(g4674), .Z(g7788) ) ;
INV     gate3449  (.A(g6215), .Z(II12199) ) ;
INV     gate3450  (.A(II12199), .Z(g7791) ) ;
INV     gate3451  (.A(g324), .Z(g7802) ) ;
INV     gate3452  (.A(g4366), .Z(g7805) ) ;
INV     gate3453  (.A(g4681), .Z(g7806) ) ;
INV     gate3454  (.A(g4864), .Z(g7809) ) ;
INV     gate3455  (.A(g6561), .Z(II12214) ) ;
INV     gate3456  (.A(II12214), .Z(g7812) ) ;
INV     gate3457  (.A(g4169), .Z(g7824) ) ;
INV     gate3458  (.A(g4688), .Z(g7827) ) ;
INV     gate3459  (.A(g4871), .Z(g7828) ) ;
INV     gate3460  (.A(g34), .Z(II12227) ) ;
INV     gate3461  (.A(II12227), .Z(g7831) ) ;
INV     gate3462  (.A(g4125), .Z(g7835) ) ;
INV     gate3463  (.A(g4878), .Z(g7840) ) ;
INV     gate3464  (.A(g904), .Z(g7841) ) ;
INV     gate3465  (.A(g1146), .Z(g7845) ) ;
INV     gate3466  (.A(g921), .Z(g7851) ) ;
INV     gate3467  (.A(g1152), .Z(g7854) ) ;
INV     gate3468  (.A(g947), .Z(g7858) ) ;
INV     gate3469  (.A(g1249), .Z(g7863) ) ;
INV     gate3470  (.A(g1489), .Z(g7867) ) ;
INV     gate3471  (.A(g1099), .Z(g7868) ) ;
INV     gate3472  (.A(g1193), .Z(g7870) ) ;
INV     gate3473  (.A(g1266), .Z(g7873) ) ;
INV     gate3474  (.A(g1495), .Z(g7876) ) ;
INV     gate3475  (.A(g1291), .Z(g7880) ) ;
INV     gate3476  (.A(g1442), .Z(g7886) ) ;
INV     gate3477  (.A(g1536), .Z(g7888) ) ;
INV     gate3478  (.A(g2994), .Z(g7891) ) ;
INV     gate3479  (.A(g4801), .Z(g7892) ) ;
INV     gate3480  (.A(g4991), .Z(g7898) ) ;
INV     gate3481  (.A(g969), .Z(g7903) ) ;
INV     gate3482  (.A(g3072), .Z(g7907) ) ;
INV     gate3483  (.A(g4157), .Z(g7908) ) ;
INV     gate3484  (.A(g936), .Z(g7909) ) ;
INV     gate3485  (.A(g1052), .Z(g7913) ) ;
INV     gate3486  (.A(g1157), .Z(II12300) ) ;
INV     gate3487  (.A(g1157), .Z(g7917) ) ;
INV     gate3488  (.A(g1312), .Z(g7922) ) ;
INV     gate3489  (.A(g3423), .Z(g7926) ) ;
INV     gate3490  (.A(g4064), .Z(g7927) ) ;
INV     gate3491  (.A(g4776), .Z(g7928) ) ;
INV     gate3492  (.A(g907), .Z(g7933) ) ;
INV     gate3493  (.A(g1061), .Z(g7936) ) ;
INV     gate3494  (.A(g1280), .Z(g7939) ) ;
INV     gate3495  (.A(g1395), .Z(g7943) ) ;
INV     gate3496  (.A(g1500), .Z(II12314) ) ;
INV     gate3497  (.A(g1500), .Z(g7947) ) ;
INV     gate3498  (.A(g3774), .Z(g7952) ) ;
INV     gate3499  (.A(g4966), .Z(g7953) ) ;
INV     gate3500  (.A(g1252), .Z(g7957) ) ;
INV     gate3501  (.A(g1404), .Z(g7960) ) ;
INV     gate3502  (.A(g4146), .Z(g7963) ) ;
INV     gate3503  (.A(g3155), .Z(g7964) ) ;
INV     gate3504  (.A(g4688), .Z(g7970) ) ;
INV     gate3505  (.A(g4818), .Z(g7971) ) ;
INV     gate3506  (.A(g1046), .Z(g7972) ) ;
INV     gate3507  (.A(g3040), .Z(g7975) ) ;
INV     gate3508  (.A(g3161), .Z(g7980) ) ;
INV     gate3509  (.A(g3506), .Z(g7985) ) ;
INV     gate3510  (.A(g4878), .Z(g7991) ) ;
INV     gate3511  (.A(g5008), .Z(g7992) ) ;
INV     gate3512  (.A(g45), .Z(II12333) ) ;
INV     gate3513  (.A(II12333), .Z(g7993) ) ;
INV     gate3514  (.A(g52), .Z(II12336) ) ;
INV     gate3515  (.A(II12336), .Z(g7994) ) ;
INV     gate3516  (.A(g153), .Z(g7995) ) ;
INV     gate3517  (.A(g392), .Z(g7998) ) ;
INV     gate3518  (.A(g1389), .Z(g8002) ) ;
INV     gate3519  (.A(g3025), .Z(g8005) ) ;
INV     gate3520  (.A(g3106), .Z(g8009) ) ;
INV     gate3521  (.A(g3167), .Z(g8011) ) ;
INV     gate3522  (.A(g3391), .Z(g8016) ) ;
INV     gate3523  (.A(g3512), .Z(g8021) ) ;
INV     gate3524  (.A(g3857), .Z(g8026) ) ;
INV     gate3525  (.A(g46), .Z(II12355) ) ;
INV     gate3526  (.A(II12355), .Z(g8032) ) ;
INV     gate3527  (.A(g157), .Z(g8033) ) ;
INV     gate3528  (.A(g405), .Z(g8037) ) ;
INV     gate3529  (.A(g528), .Z(II12360) ) ;
INV     gate3530  (.A(II12360), .Z(g8038) ) ;
INV     gate3531  (.A(g528), .Z(g8046) ) ;
INV     gate3532  (.A(g1211), .Z(g8052) ) ;
INV     gate3533  (.A(g1236), .Z(g8055) ) ;
INV     gate3534  (.A(g1246), .Z(g8056) ) ;
INV     gate3535  (.A(g3068), .Z(g8057) ) ;
INV     gate3536  (.A(g3115), .Z(g8058) ) ;
INV     gate3537  (.A(g3171), .Z(g8059) ) ;
INV     gate3538  (.A(g3376), .Z(g8064) ) ;
INV     gate3539  (.A(g3457), .Z(g8068) ) ;
INV     gate3540  (.A(g3518), .Z(g8070) ) ;
INV     gate3541  (.A(g3742), .Z(g8075) ) ;
INV     gate3542  (.A(g3863), .Z(g8080) ) ;
INV     gate3543  (.A(g47), .Z(II12382) ) ;
INV     gate3544  (.A(II12382), .Z(g8085) ) ;
INV     gate3545  (.A(g1157), .Z(g8087) ) ;
INV     gate3546  (.A(g1554), .Z(g8088) ) ;
INV     gate3547  (.A(g1579), .Z(g8091) ) ;
INV     gate3548  (.A(g1589), .Z(g8092) ) ;
INV     gate3549  (.A(g1624), .Z(g8093) ) ;
INV     gate3550  (.A(g3029), .Z(g8097) ) ;
INV     gate3551  (.A(g3072), .Z(g8102) ) ;
INV     gate3552  (.A(g3133), .Z(g8106) ) ;
INV     gate3553  (.A(g3179), .Z(g8107) ) ;
INV     gate3554  (.A(g3419), .Z(g8112) ) ;
INV     gate3555  (.A(g3466), .Z(g8113) ) ;
INV     gate3556  (.A(g3522), .Z(g8114) ) ;
INV     gate3557  (.A(g3727), .Z(g8119) ) ;
INV     gate3558  (.A(g3808), .Z(g8123) ) ;
INV     gate3559  (.A(g3869), .Z(g8125) ) ;
INV     gate3560  (.A(g4515), .Z(g8130) ) ;
INV     gate3561  (.A(g4809), .Z(II12411) ) ;
INV     gate3562  (.A(g4809), .Z(g8133) ) ;
INV     gate3563  (.A(g48), .Z(II12415) ) ;
INV     gate3564  (.A(II12415), .Z(g8134) ) ;
INV     gate3565  (.A(g55), .Z(II12418) ) ;
INV     gate3566  (.A(II12418), .Z(g8135) ) ;
INV     gate3567  (.A(g269), .Z(g8136) ) ;
INV     gate3568  (.A(g411), .Z(g8137) ) ;
INV     gate3569  (.A(g1500), .Z(g8138) ) ;
INV     gate3570  (.A(g1648), .Z(g8139) ) ;
INV     gate3571  (.A(g1760), .Z(g8146) ) ;
INV     gate3572  (.A(g2185), .Z(g8150) ) ;
INV     gate3573  (.A(g3139), .Z(g8154) ) ;
INV     gate3574  (.A(g3380), .Z(g8155) ) ;
INV     gate3575  (.A(g3423), .Z(g8160) ) ;
INV     gate3576  (.A(g3484), .Z(g8164) ) ;
INV     gate3577  (.A(g3530), .Z(g8165) ) ;
INV     gate3578  (.A(g3770), .Z(g8170) ) ;
INV     gate3579  (.A(g3817), .Z(g8171) ) ;
INV     gate3580  (.A(g3873), .Z(g8172) ) ;
INV     gate3581  (.A(g4999), .Z(II12437) ) ;
INV     gate3582  (.A(g4999), .Z(g8179) ) ;
INV     gate3583  (.A(g262), .Z(g8180) ) ;
INV     gate3584  (.A(g424), .Z(g8181) ) ;
INV     gate3585  (.A(g482), .Z(g8183) ) ;
INV     gate3586  (.A(g990), .Z(g8186) ) ;
INV     gate3587  (.A(g1657), .Z(g8187) ) ;
INV     gate3588  (.A(g1783), .Z(g8195) ) ;
INV     gate3589  (.A(g1894), .Z(g8201) ) ;
INV     gate3590  (.A(g2208), .Z(g8205) ) ;
INV     gate3591  (.A(g2319), .Z(g8211) ) ;
INV     gate3592  (.A(g3092), .Z(II12451) ) ;
INV     gate3593  (.A(g3092), .Z(g8216) ) ;
INV     gate3594  (.A(g3143), .Z(g8217) ) ;
INV     gate3595  (.A(g3490), .Z(g8218) ) ;
INV     gate3596  (.A(g3731), .Z(g8219) ) ;
INV     gate3597  (.A(g3774), .Z(g8224) ) ;
INV     gate3598  (.A(g3835), .Z(g8228) ) ;
INV     gate3599  (.A(g3881), .Z(g8229) ) ;
INV     gate3600  (.A(g4812), .Z(II12463) ) ;
INV     gate3601  (.A(g4812), .Z(g8236) ) ;
INV     gate3602  (.A(g255), .Z(g8237) ) ;
INV     gate3603  (.A(g1056), .Z(g8239) ) ;
INV     gate3604  (.A(g1333), .Z(g8240) ) ;
INV     gate3605  (.A(g1792), .Z(g8241) ) ;
INV     gate3606  (.A(g1917), .Z(g8249) ) ;
INV     gate3607  (.A(g2028), .Z(g8255) ) ;
INV     gate3608  (.A(g2217), .Z(g8259) ) ;
INV     gate3609  (.A(g2342), .Z(g8267) ) ;
INV     gate3610  (.A(g2453), .Z(g8273) ) ;
INV     gate3611  (.A(g3096), .Z(II12483) ) ;
INV     gate3612  (.A(g3096), .Z(g8278) ) ;
INV     gate3613  (.A(g3443), .Z(II12487) ) ;
INV     gate3614  (.A(g3443), .Z(g8280) ) ;
INV     gate3615  (.A(g3494), .Z(g8281) ) ;
INV     gate3616  (.A(g3841), .Z(g8282) ) ;
INV     gate3617  (.A(g5002), .Z(II12493) ) ;
INV     gate3618  (.A(g5002), .Z(g8284) ) ;
INV     gate3619  (.A(g49), .Z(II12497) ) ;
INV     gate3620  (.A(II12497), .Z(g8285) ) ;
INV     gate3621  (.A(g53), .Z(g8286) ) ;
INV     gate3622  (.A(g160), .Z(g8287) ) ;
INV     gate3623  (.A(g218), .Z(g8290) ) ;
INV     gate3624  (.A(g215), .Z(II12503) ) ;
INV     gate3625  (.A(g246), .Z(g8296) ) ;
INV     gate3626  (.A(g142), .Z(g8297) ) ;
INV     gate3627  (.A(g1242), .Z(g8300) ) ;
INV     gate3628  (.A(g1399), .Z(g8301) ) ;
INV     gate3629  (.A(g1926), .Z(g8302) ) ;
INV     gate3630  (.A(g2051), .Z(g8310) ) ;
INV     gate3631  (.A(g2351), .Z(g8316) ) ;
INV     gate3632  (.A(g2476), .Z(g8324) ) ;
INV     gate3633  (.A(g2587), .Z(g8330) ) ;
INV     gate3634  (.A(g3034), .Z(g8334) ) ;
INV     gate3635  (.A(g3050), .Z(g8340) ) ;
INV     gate3636  (.A(g3119), .Z(g8341) ) ;
INV     gate3637  (.A(g3447), .Z(II12519) ) ;
INV     gate3638  (.A(g3447), .Z(g8343) ) ;
INV     gate3639  (.A(g3794), .Z(II12523) ) ;
INV     gate3640  (.A(g3794), .Z(g8345) ) ;
INV     gate3641  (.A(g3845), .Z(g8346) ) ;
INV     gate3642  (.A(g4646), .Z(g8350) ) ;
INV     gate3643  (.A(g4815), .Z(II12530) ) ;
INV     gate3644  (.A(g4815), .Z(g8354) ) ;
INV     gate3645  (.A(g50), .Z(II12534) ) ;
INV     gate3646  (.A(II12534), .Z(g8355) ) ;
INV     gate3647  (.A(g54), .Z(g8356) ) ;
INV     gate3648  (.A(g58), .Z(II12538) ) ;
INV     gate3649  (.A(II12538), .Z(g8357) ) ;
INV     gate3650  (.A(g194), .Z(II12541) ) ;
INV     gate3651  (.A(g194), .Z(g8362) ) ;
INV     gate3652  (.A(g239), .Z(g8363) ) ;
INV     gate3653  (.A(g1585), .Z(g8364) ) ;
INV     gate3654  (.A(g2060), .Z(g8365) ) ;
INV     gate3655  (.A(g2485), .Z(g8373) ) ;
INV     gate3656  (.A(g2610), .Z(g8381) ) ;
INV     gate3657  (.A(g3080), .Z(g8387) ) ;
INV     gate3658  (.A(g3010), .Z(g8388) ) ;
INV     gate3659  (.A(g3125), .Z(g8389) ) ;
INV     gate3660  (.A(g3385), .Z(g8390) ) ;
INV     gate3661  (.A(g3401), .Z(g8396) ) ;
INV     gate3662  (.A(g3470), .Z(g8397) ) ;
INV     gate3663  (.A(g3798), .Z(II12563) ) ;
INV     gate3664  (.A(g3798), .Z(g8399) ) ;
INV     gate3665  (.A(g4836), .Z(g8400) ) ;
INV     gate3666  (.A(g5005), .Z(II12568) ) ;
INV     gate3667  (.A(g5005), .Z(g8404) ) ;
INV     gate3668  (.A(g51), .Z(II12572) ) ;
INV     gate3669  (.A(II12572), .Z(g8405) ) ;
INV     gate3670  (.A(g232), .Z(g8406) ) ;
INV     gate3671  (.A(g1171), .Z(g8407) ) ;
INV     gate3672  (.A(g1227), .Z(II12577) ) ;
INV     gate3673  (.A(II12577), .Z(g8411) ) ;
INV     gate3674  (.A(g1239), .Z(II12580) ) ;
INV     gate3675  (.A(g2619), .Z(g8418) ) ;
INV     gate3676  (.A(g3045), .Z(g8426) ) ;
INV     gate3677  (.A(g3085), .Z(g8431) ) ;
INV     gate3678  (.A(g3100), .Z(g8438) ) ;
INV     gate3679  (.A(g3129), .Z(g8439) ) ;
INV     gate3680  (.A(g3431), .Z(g8440) ) ;
INV     gate3681  (.A(g3361), .Z(g8441) ) ;
INV     gate3682  (.A(g3476), .Z(g8442) ) ;
INV     gate3683  (.A(g3736), .Z(g8443) ) ;
INV     gate3684  (.A(g3752), .Z(g8449) ) ;
INV     gate3685  (.A(g3821), .Z(g8450) ) ;
INV     gate3686  (.A(g4057), .Z(g8451) ) ;
INV     gate3687  (.A(g56), .Z(g8456) ) ;
INV     gate3688  (.A(g225), .Z(g8457) ) ;
INV     gate3689  (.A(g294), .Z(g8458) ) ;
INV     gate3690  (.A(g1183), .Z(g8462) ) ;
INV     gate3691  (.A(g1514), .Z(g8466) ) ;
INV     gate3692  (.A(g1570), .Z(II12605) ) ;
INV     gate3693  (.A(II12605), .Z(g8470) ) ;
INV     gate3694  (.A(g1582), .Z(II12608) ) ;
INV     gate3695  (.A(g3061), .Z(g8477) ) ;
INV     gate3696  (.A(g3103), .Z(g8478) ) ;
INV     gate3697  (.A(g3057), .Z(g8479) ) ;
INV     gate3698  (.A(g3147), .Z(g8480) ) ;
INV     gate3699  (.A(g3338), .Z(II12618) ) ;
INV     gate3700  (.A(II12618), .Z(g8481) ) ;
INV     gate3701  (.A(g3396), .Z(g8492) ) ;
INV     gate3702  (.A(g3436), .Z(g8497) ) ;
INV     gate3703  (.A(g3451), .Z(g8504) ) ;
INV     gate3704  (.A(g3480), .Z(g8505) ) ;
INV     gate3705  (.A(g3782), .Z(g8506) ) ;
INV     gate3706  (.A(g3712), .Z(g8507) ) ;
INV     gate3707  (.A(g3827), .Z(g8508) ) ;
INV     gate3708  (.A(g4141), .Z(g8509) ) ;
INV     gate3709  (.A(g4258), .Z(g8514) ) ;
INV     gate3710  (.A(g1242), .Z(II12631) ) ;
INV     gate3711  (.A(II12631), .Z(g8515) ) ;
INV     gate3712  (.A(g287), .Z(g8519) ) ;
INV     gate3713  (.A(g298), .Z(g8522) ) ;
INV     gate3714  (.A(g1526), .Z(g8526) ) ;
INV     gate3715  (.A(g3288), .Z(g8531) ) ;
INV     gate3716  (.A(g3338), .Z(g8534) ) ;
INV     gate3717  (.A(g3412), .Z(g8538) ) ;
INV     gate3718  (.A(g3454), .Z(g8539) ) ;
INV     gate3719  (.A(g3408), .Z(g8540) ) ;
INV     gate3720  (.A(g3498), .Z(g8541) ) ;
INV     gate3721  (.A(g3689), .Z(II12644) ) ;
INV     gate3722  (.A(II12644), .Z(g8542) ) ;
INV     gate3723  (.A(g3747), .Z(g8553) ) ;
INV     gate3724  (.A(g3787), .Z(g8558) ) ;
INV     gate3725  (.A(g3802), .Z(g8565) ) ;
INV     gate3726  (.A(g3831), .Z(g8566) ) ;
INV     gate3727  (.A(g4082), .Z(g8567) ) ;
INV     gate3728  (.A(g57), .Z(g8571) ) ;
INV     gate3729  (.A(g1585), .Z(II12654) ) ;
INV     gate3730  (.A(II12654), .Z(g8572) ) ;
INV     gate3731  (.A(g291), .Z(g8575) ) ;
INV     gate3732  (.A(g2771), .Z(g8579) ) ;
INV     gate3733  (.A(g3639), .Z(g8584) ) ;
INV     gate3734  (.A(g3689), .Z(g8587) ) ;
INV     gate3735  (.A(g3763), .Z(g8591) ) ;
INV     gate3736  (.A(g3805), .Z(g8592) ) ;
INV     gate3737  (.A(g3759), .Z(g8593) ) ;
INV     gate3738  (.A(g3849), .Z(g8594) ) ;
INV     gate3739  (.A(g4040), .Z(II12666) ) ;
INV     gate3740  (.A(II12666), .Z(g8595) ) ;
INV     gate3741  (.A(g4653), .Z(g8606) ) ;
INV     gate3742  (.A(g37), .Z(g8607) ) ;
INV     gate3743  (.A(g278), .Z(g8608) ) ;
INV     gate3744  (.A(g2775), .Z(g8612) ) ;
INV     gate3745  (.A(g2803), .Z(g8616) ) ;
INV     gate3746  (.A(g3065), .Z(g8620) ) ;
INV     gate3747  (.A(g3990), .Z(g8623) ) ;
INV     gate3748  (.A(g4040), .Z(g8626) ) ;
INV     gate3749  (.A(g4843), .Z(g8630) ) ;
INV     gate3750  (.A(g283), .Z(g8631) ) ;
INV     gate3751  (.A(g2783), .Z(g8635) ) ;
INV     gate3752  (.A(g2807), .Z(g8639) ) ;
INV     gate3753  (.A(g3352), .Z(g8644) ) ;
INV     gate3754  (.A(g3416), .Z(g8647) ) ;
INV     gate3755  (.A(g4664), .Z(g8650) ) ;
INV     gate3756  (.A(g758), .Z(g8651) ) ;
INV     gate3757  (.A(g1087), .Z(g8654) ) ;
INV     gate3758  (.A(g2787), .Z(g8655) ) ;
INV     gate3759  (.A(g2815), .Z(g8659) ) ;
INV     gate3760  (.A(g3343), .Z(g8663) ) ;
INV     gate3761  (.A(g3703), .Z(g8666) ) ;
INV     gate3762  (.A(g3767), .Z(g8669) ) ;
INV     gate3763  (.A(g4669), .Z(g8672) ) ;
INV     gate3764  (.A(g4737), .Z(g8673) ) ;
INV     gate3765  (.A(g4821), .Z(g8676) ) ;
INV     gate3766  (.A(g4854), .Z(g8677) ) ;
INV     gate3767  (.A(g686), .Z(g8680) ) ;
INV     gate3768  (.A(g763), .Z(g8681) ) ;
INV     gate3769  (.A(g1430), .Z(g8685) ) ;
INV     gate3770  (.A(g2819), .Z(g8686) ) ;
INV     gate3771  (.A(g3347), .Z(g8696) ) ;
INV     gate3772  (.A(g3694), .Z(g8697) ) ;
INV     gate3773  (.A(g4054), .Z(g8700) ) ;
INV     gate3774  (.A(g4284), .Z(II12709) ) ;
INV     gate3775  (.A(II12709), .Z(g8703) ) ;
INV     gate3776  (.A(g59), .Z(II12712) ) ;
INV     gate3777  (.A(II12712), .Z(g8712) ) ;
INV     gate3778  (.A(g4826), .Z(g8713) ) ;
INV     gate3779  (.A(g4859), .Z(g8714) ) ;
INV     gate3780  (.A(g4927), .Z(g8715) ) ;
INV     gate3781  (.A(g3333), .Z(g8718) ) ;
INV     gate3782  (.A(g365), .Z(II12719) ) ;
INV     gate3783  (.A(g739), .Z(g8725) ) ;
INV     gate3784  (.A(g3698), .Z(g8733) ) ;
INV     gate3785  (.A(g4045), .Z(g8734) ) ;
INV     gate3786  (.A(g4572), .Z(II12735) ) ;
INV     gate3787  (.A(II12735), .Z(g8740) ) ;
INV     gate3788  (.A(g4821), .Z(g8741) ) ;
INV     gate3789  (.A(g4035), .Z(g8742) ) ;
INV     gate3790  (.A(g550), .Z(g8743) ) ;
INV     gate3791  (.A(g691), .Z(g8744) ) ;
INV     gate3792  (.A(g744), .Z(g8745) ) ;
INV     gate3793  (.A(g776), .Z(g8748) ) ;
INV     gate3794  (.A(g4049), .Z(g8756) ) ;
INV     gate3795  (.A(g4087), .Z(II12746) ) ;
INV     gate3796  (.A(II12746), .Z(g8757) ) ;
INV     gate3797  (.A(g4575), .Z(II12749) ) ;
INV     gate3798  (.A(II12749), .Z(g8763) ) ;
INV     gate3799  (.A(g4826), .Z(g8764) ) ;
INV     gate3800  (.A(g3333), .Z(g8765) ) ;
INV     gate3801  (.A(g572), .Z(g8766) ) ;
INV     gate3802  (.A(g749), .Z(g8770) ) ;
INV     gate3803  (.A(g781), .Z(g8774) ) ;
INV     gate3804  (.A(g4093), .Z(II12758) ) ;
INV     gate3805  (.A(II12758), .Z(g8778) ) ;
INV     gate3806  (.A(g4188), .Z(II12761) ) ;
INV     gate3807  (.A(g4194), .Z(II12764) ) ;
INV     gate3808  (.A(g4197), .Z(II12767) ) ;
INV     gate3809  (.A(g4200), .Z(II12770) ) ;
INV     gate3810  (.A(g4204), .Z(II12773) ) ;
INV     gate3811  (.A(g4207), .Z(II12776) ) ;
INV     gate3812  (.A(g4210), .Z(II12779) ) ;
INV     gate3813  (.A(g4311), .Z(II12787) ) ;
INV     gate3814  (.A(II12787), .Z(g8791) ) ;
INV     gate3815  (.A(g4340), .Z(II12790) ) ;
INV     gate3816  (.A(II12790), .Z(g8792) ) ;
INV     gate3817  (.A(g4578), .Z(II12793) ) ;
INV     gate3818  (.A(II12793), .Z(g8795) ) ;
INV     gate3819  (.A(g4785), .Z(g8796) ) ;
INV     gate3820  (.A(g4035), .Z(g8804) ) ;
INV     gate3821  (.A(g59), .Z(II12799) ) ;
INV     gate3822  (.A(II12799), .Z(g8805) ) ;
INV     gate3823  (.A(g79), .Z(g8807) ) ;
INV     gate3824  (.A(g595), .Z(g8808) ) ;
INV     gate3825  (.A(g4098), .Z(II12805) ) ;
INV     gate3826  (.A(II12805), .Z(g8812) ) ;
INV     gate3827  (.A(g4322), .Z(II12808) ) ;
INV     gate3828  (.A(II12808), .Z(g8818) ) ;
INV     gate3829  (.A(g4340), .Z(II12811) ) ;
INV     gate3830  (.A(II12811), .Z(g8821) ) ;
INV     gate3831  (.A(g4975), .Z(g8822) ) ;
INV     gate3832  (.A(g767), .Z(g8830) ) ;
INV     gate3833  (.A(g794), .Z(g8833) ) ;
INV     gate3834  (.A(g736), .Z(g8836) ) ;
INV     gate3835  (.A(g4277), .Z(II12819) ) ;
INV     gate3836  (.A(g4277), .Z(g8840) ) ;
INV     gate3837  (.A(g4311), .Z(II12823) ) ;
INV     gate3838  (.A(II12823), .Z(g8841) ) ;
INV     gate3839  (.A(g4349), .Z(II12826) ) ;
INV     gate3840  (.A(II12826), .Z(g8844) ) ;
INV     gate3841  (.A(g358), .Z(g8848) ) ;
INV     gate3842  (.A(g590), .Z(g8851) ) ;
INV     gate3843  (.A(g613), .Z(g8854) ) ;
INV     gate3844  (.A(g671), .Z(g8858) ) ;
INV     gate3845  (.A(g772), .Z(g8859) ) ;
INV     gate3846  (.A(g4222), .Z(II12837) ) ;
INV     gate3847  (.A(g4258), .Z(g8872) ) ;
INV     gate3848  (.A(g4311), .Z(II12855) ) ;
INV     gate3849  (.A(II12855), .Z(g8876) ) ;
INV     gate3850  (.A(g4340), .Z(II12858) ) ;
INV     gate3851  (.A(II12858), .Z(g8879) ) ;
INV     gate3852  (.A(g4372), .Z(II12861) ) ;
INV     gate3853  (.A(II12861), .Z(g8880) ) ;
INV     gate3854  (.A(g4709), .Z(g8883) ) ;
INV     gate3855  (.A(g376), .Z(g8890) ) ;
INV     gate3856  (.A(g582), .Z(g8891) ) ;
INV     gate3857  (.A(g599), .Z(g8895) ) ;
INV     gate3858  (.A(g676), .Z(g8898) ) ;
INV     gate3859  (.A(g807), .Z(g8899) ) ;
INV     gate3860  (.A(g1075), .Z(g8903) ) ;
INV     gate3861  (.A(g4180), .Z(g8912) ) ;
INV     gate3862  (.A(g4264), .Z(g8914) ) ;
INV     gate3863  (.A(g4213), .Z(II12884) ) ;
INV     gate3864  (.A(g4216), .Z(II12887) ) ;
INV     gate3865  (.A(g4219), .Z(II12890) ) ;
INV     gate3866  (.A(g4226), .Z(II12893) ) ;
INV     gate3867  (.A(g4229), .Z(II12896) ) ;
INV     gate3868  (.A(g4232), .Z(II12899) ) ;
INV     gate3869  (.A(g4322), .Z(II12907) ) ;
INV     gate3870  (.A(II12907), .Z(g8922) ) ;
INV     gate3871  (.A(g4340), .Z(II12910) ) ;
INV     gate3872  (.A(II12910), .Z(g8925) ) ;
INV     gate3873  (.A(g4340), .Z(g8928) ) ;
INV     gate3874  (.A(g4899), .Z(g8938) ) ;
INV     gate3875  (.A(g370), .Z(g8944) ) ;
INV     gate3876  (.A(g608), .Z(g8945) ) ;
INV     gate3877  (.A(g785), .Z(g8948) ) ;
INV     gate3878  (.A(g554), .Z(g8951) ) ;
INV     gate3879  (.A(g1079), .Z(g8954) ) ;
INV     gate3880  (.A(g1418), .Z(g8955) ) ;
INV     gate3881  (.A(g4269), .Z(g8964) ) ;
INV     gate3882  (.A(g4332), .Z(II12927) ) ;
INV     gate3883  (.A(II12927), .Z(g8971) ) ;
INV     gate3884  (.A(g4349), .Z(II12930) ) ;
INV     gate3885  (.A(II12930), .Z(g8974) ) ;
INV     gate3886  (.A(g4349), .Z(g8977) ) ;
INV     gate3887  (.A(g6753), .Z(II12935) ) ;
INV     gate3888  (.A(II12935), .Z(g8989) ) ;
INV     gate3889  (.A(g146), .Z(g8990) ) ;
INV     gate3890  (.A(g385), .Z(g8993) ) ;
INV     gate3891  (.A(g577), .Z(g8997) ) ;
INV     gate3892  (.A(g632), .Z(g9000) ) ;
INV     gate3893  (.A(g790), .Z(g9003) ) ;
INV     gate3894  (.A(g1083), .Z(g9007) ) ;
INV     gate3895  (.A(g1422), .Z(g9011) ) ;
INV     gate3896  (.A(g3004), .Z(g9014) ) ;
INV     gate3897  (.A(g4273), .Z(g9018) ) ;
INV     gate3898  (.A(g4287), .Z(II12950) ) ;
INV     gate3899  (.A(g4287), .Z(g9020) ) ;
INV     gate3900  (.A(g4358), .Z(II12954) ) ;
INV     gate3901  (.A(II12954), .Z(g9021) ) ;
INV     gate3902  (.A(g4358), .Z(g9024) ) ;
INV     gate3903  (.A(g4793), .Z(g9030) ) ;
INV     gate3904  (.A(g5084), .Z(g9036) ) ;
INV     gate3905  (.A(g164), .Z(g9037) ) ;
INV     gate3906  (.A(g499), .Z(g9040) ) ;
INV     gate3907  (.A(g604), .Z(g9044) ) ;
INV     gate3908  (.A(g640), .Z(II12963) ) ;
INV     gate3909  (.A(g640), .Z(g9049) ) ;
INV     gate3910  (.A(g1087), .Z(g9050) ) ;
INV     gate3911  (.A(g1426), .Z(g9051) ) ;
INV     gate3912  (.A(g3017), .Z(g9056) ) ;
INV     gate3913  (.A(g3355), .Z(g9060) ) ;
INV     gate3914  (.A(g4983), .Z(g9064) ) ;
INV     gate3915  (.A(g5428), .Z(g9070) ) ;
INV     gate3916  (.A(g2831), .Z(g9071) ) ;
INV     gate3917  (.A(g2994), .Z(g9072) ) ;
INV     gate3918  (.A(g150), .Z(g9073) ) ;
INV     gate3919  (.A(g504), .Z(g9077) ) ;
INV     gate3920  (.A(g626), .Z(g9083) ) ;
INV     gate3921  (.A(g847), .Z(g9086) ) ;
INV     gate3922  (.A(g1430), .Z(g9091) ) ;
INV     gate3923  (.A(g3368), .Z(g9095) ) ;
INV     gate3924  (.A(g3706), .Z(g9099) ) ;
INV     gate3925  (.A(g5774), .Z(g9103) ) ;
INV     gate3926  (.A(g12), .Z(II12987) ) ;
INV     gate3927  (.A(II12987), .Z(g9104) ) ;
INV     gate3928  (.A(g2834), .Z(g9152) ) ;
INV     gate3929  (.A(g6752), .Z(II12991) ) ;
INV     gate3930  (.A(II12991), .Z(g9153) ) ;
INV     gate3931  (.A(g6748), .Z(II12994) ) ;
INV     gate3932  (.A(II12994), .Z(g9154) ) ;
INV     gate3933  (.A(g351), .Z(II12997) ) ;
INV     gate3934  (.A(II12997), .Z(g9155) ) ;
INV     gate3935  (.A(g513), .Z(g9158) ) ;
INV     gate3936  (.A(g622), .Z(g9162) ) ;
INV     gate3937  (.A(g837), .Z(g9166) ) ;
INV     gate3938  (.A(g1205), .Z(g9174) ) ;
INV     gate3939  (.A(g3719), .Z(g9180) ) ;
INV     gate3940  (.A(g6120), .Z(g9184) ) ;
INV     gate3941  (.A(g65), .Z(II13007) ) ;
INV     gate3942  (.A(II13007), .Z(g9185) ) ;
INV     gate3943  (.A(g6749), .Z(II13010) ) ;
INV     gate3944  (.A(II13010), .Z(g9186) ) ;
INV     gate3945  (.A(g518), .Z(g9187) ) ;
INV     gate3946  (.A(g827), .Z(g9194) ) ;
INV     gate3947  (.A(g1221), .Z(g9197) ) ;
INV     gate3948  (.A(g1548), .Z(g9200) ) ;
INV     gate3949  (.A(g5164), .Z(g9206) ) ;
INV     gate3950  (.A(g6466), .Z(g9212) ) ;
INV     gate3951  (.A(g6750), .Z(II13020) ) ;
INV     gate3952  (.A(II13020), .Z(g9213) ) ;
INV     gate3953  (.A(g617), .Z(g9214) ) ;
INV     gate3954  (.A(g843), .Z(g9220) ) ;
INV     gate3955  (.A(g1216), .Z(g9223) ) ;
INV     gate3956  (.A(g1564), .Z(g9226) ) ;
INV     gate3957  (.A(g5052), .Z(g9229) ) ;
INV     gate3958  (.A(g5170), .Z(g9234) ) ;
INV     gate3959  (.A(g5511), .Z(g9239) ) ;
INV     gate3960  (.A(g6747), .Z(II13031) ) ;
INV     gate3961  (.A(II13031), .Z(g9245) ) ;
INV     gate3962  (.A(g1559), .Z(g9247) ) ;
INV     gate3963  (.A(g1600), .Z(g9250) ) ;
INV     gate3964  (.A(g4304), .Z(II13037) ) ;
INV     gate3965  (.A(g4304), .Z(g9252) ) ;
INV     gate3966  (.A(g5037), .Z(g9253) ) ;
INV     gate3967  (.A(g5115), .Z(g9257) ) ;
INV     gate3968  (.A(g5176), .Z(g9259) ) ;
INV     gate3969  (.A(g5396), .Z(g9264) ) ;
INV     gate3970  (.A(g5517), .Z(g9269) ) ;
INV     gate3971  (.A(g5857), .Z(g9274) ) ;
INV     gate3972  (.A(g6744), .Z(II13054) ) ;
INV     gate3973  (.A(II13054), .Z(g9280) ) ;
INV     gate3974  (.A(g112), .Z(II13057) ) ;
INV     gate3975  (.A(II13057), .Z(g9281) ) ;
INV     gate3976  (.A(g723), .Z(g9282) ) ;
INV     gate3977  (.A(g1736), .Z(g9283) ) ;
INV     gate3978  (.A(g2161), .Z(g9284) ) ;
INV     gate3979  (.A(g2715), .Z(g9285) ) ;
INV     gate3980  (.A(g3021), .Z(g9291) ) ;
INV     gate3981  (.A(g5080), .Z(g9298) ) ;
INV     gate3982  (.A(g5124), .Z(g9299) ) ;
INV     gate3983  (.A(g5180), .Z(g9300) ) ;
INV     gate3984  (.A(g5381), .Z(g9305) ) ;
INV     gate3985  (.A(g5462), .Z(g9309) ) ;
INV     gate3986  (.A(g5523), .Z(g9311) ) ;
INV     gate3987  (.A(g5742), .Z(g9316) ) ;
INV     gate3988  (.A(g5863), .Z(g9321) ) ;
INV     gate3989  (.A(g6203), .Z(g9326) ) ;
INV     gate3990  (.A(g64), .Z(g9332) ) ;
INV     gate3991  (.A(g417), .Z(g9333) ) ;
INV     gate3992  (.A(g1608), .Z(g9337) ) ;
INV     gate3993  (.A(g1870), .Z(g9338) ) ;
INV     gate3994  (.A(g2295), .Z(g9339) ) ;
INV     gate3995  (.A(g2724), .Z(II13094) ) ;
INV     gate3996  (.A(II13094), .Z(g9340) ) ;
INV     gate3997  (.A(g2719), .Z(g9354) ) ;
INV     gate3998  (.A(g3372), .Z(g9360) ) ;
INV     gate3999  (.A(g5041), .Z(g9364) ) ;
INV     gate4000  (.A(g5084), .Z(g9369) ) ;
INV     gate4001  (.A(g5142), .Z(g9373) ) ;
INV     gate4002  (.A(g5188), .Z(g9374) ) ;
INV     gate4003  (.A(g5424), .Z(g9379) ) ;
INV     gate4004  (.A(g5471), .Z(g9380) ) ;
INV     gate4005  (.A(g5527), .Z(g9381) ) ;
INV     gate4006  (.A(g5727), .Z(g9386) ) ;
INV     gate4007  (.A(g5808), .Z(g9390) ) ;
INV     gate4008  (.A(g5869), .Z(g9392) ) ;
INV     gate4009  (.A(g6088), .Z(g9397) ) ;
INV     gate4010  (.A(g6209), .Z(g9402) ) ;
INV     gate4011  (.A(g6549), .Z(g9407) ) ;
INV     gate4012  (.A(g1744), .Z(g9413) ) ;
INV     gate4013  (.A(g2004), .Z(g9414) ) ;
INV     gate4014  (.A(g2169), .Z(g9415) ) ;
INV     gate4015  (.A(g2429), .Z(g9416) ) ;
INV     gate4016  (.A(g2729), .Z(II13124) ) ;
INV     gate4017  (.A(II13124), .Z(g9417) ) ;
INV     gate4018  (.A(g3723), .Z(g9429) ) ;
INV     gate4019  (.A(g5148), .Z(g9433) ) ;
INV     gate4020  (.A(g5385), .Z(g9434) ) ;
INV     gate4021  (.A(g5428), .Z(g9439) ) ;
INV     gate4022  (.A(g5489), .Z(g9443) ) ;
INV     gate4023  (.A(g5535), .Z(g9444) ) ;
INV     gate4024  (.A(g5770), .Z(g9449) ) ;
INV     gate4025  (.A(g5817), .Z(g9450) ) ;
INV     gate4026  (.A(g5873), .Z(g9451) ) ;
INV     gate4027  (.A(g6073), .Z(g9456) ) ;
INV     gate4028  (.A(g6154), .Z(g9460) ) ;
INV     gate4029  (.A(g6215), .Z(g9462) ) ;
INV     gate4030  (.A(g6434), .Z(g9467) ) ;
INV     gate4031  (.A(g6555), .Z(g9472) ) ;
INV     gate4032  (.A(g6745), .Z(II13149) ) ;
INV     gate4033  (.A(II13149), .Z(g9477) ) ;
INV     gate4034  (.A(g6746), .Z(II13152) ) ;
INV     gate4035  (.A(II13152), .Z(g9478) ) ;
INV     gate4036  (.A(g559), .Z(g9480) ) ;
INV     gate4037  (.A(g1612), .Z(g9484) ) ;
INV     gate4038  (.A(g1878), .Z(g9488) ) ;
INV     gate4039  (.A(g2303), .Z(g9489) ) ;
INV     gate4040  (.A(g2563), .Z(g9490) ) ;
INV     gate4041  (.A(g2729), .Z(g9491) ) ;
INV     gate4042  (.A(g2759), .Z(g9492) ) ;
INV     gate4043  (.A(g3303), .Z(g9496) ) ;
INV     gate4044  (.A(g5101), .Z(II13166) ) ;
INV     gate4045  (.A(g5101), .Z(g9498) ) ;
INV     gate4046  (.A(g5152), .Z(g9499) ) ;
INV     gate4047  (.A(g5495), .Z(g9500) ) ;
INV     gate4048  (.A(g5731), .Z(g9501) ) ;
INV     gate4049  (.A(g5774), .Z(g9506) ) ;
INV     gate4050  (.A(g5835), .Z(g9510) ) ;
INV     gate4051  (.A(g5881), .Z(g9511) ) ;
INV     gate4052  (.A(g6116), .Z(g9516) ) ;
INV     gate4053  (.A(g6163), .Z(g9517) ) ;
INV     gate4054  (.A(g6219), .Z(g9518) ) ;
INV     gate4055  (.A(g6419), .Z(g9523) ) ;
INV     gate4056  (.A(g6500), .Z(g9527) ) ;
INV     gate4057  (.A(g6561), .Z(g9529) ) ;
INV     gate4058  (.A(g90), .Z(g9534) ) ;
INV     gate4059  (.A(g1748), .Z(g9537) ) ;
INV     gate4060  (.A(g2012), .Z(g9541) ) ;
INV     gate4061  (.A(g2173), .Z(g9542) ) ;
INV     gate4062  (.A(g2437), .Z(g9546) ) ;
INV     gate4063  (.A(g2735), .Z(g9547) ) ;
INV     gate4064  (.A(g3281), .Z(g9551) ) ;
INV     gate4065  (.A(g3654), .Z(g9552) ) ;
INV     gate4066  (.A(g5105), .Z(II13202) ) ;
INV     gate4067  (.A(g5105), .Z(g9554) ) ;
INV     gate4068  (.A(g5448), .Z(II13206) ) ;
INV     gate4069  (.A(g5448), .Z(g9556) ) ;
INV     gate4070  (.A(g5499), .Z(g9557) ) ;
INV     gate4071  (.A(g5841), .Z(g9558) ) ;
INV     gate4072  (.A(g6077), .Z(g9559) ) ;
INV     gate4073  (.A(g6120), .Z(g9564) ) ;
INV     gate4074  (.A(g6181), .Z(g9568) ) ;
INV     gate4075  (.A(g6227), .Z(g9569) ) ;
INV     gate4076  (.A(g6462), .Z(g9574) ) ;
INV     gate4077  (.A(g6509), .Z(g9575) ) ;
INV     gate4078  (.A(g6565), .Z(g9576) ) ;
INV     gate4079  (.A(g91), .Z(g9581) ) ;
INV     gate4080  (.A(g703), .Z(g9582) ) ;
INV     gate4081  (.A(g1616), .Z(g9585) ) ;
INV     gate4082  (.A(g1882), .Z(g9590) ) ;
INV     gate4083  (.A(g2307), .Z(g9594) ) ;
INV     gate4084  (.A(g2571), .Z(g9598) ) ;
INV     gate4085  (.A(g3310), .Z(g9599) ) ;
INV     gate4086  (.A(g3632), .Z(g9600) ) ;
INV     gate4087  (.A(g4005), .Z(g9601) ) ;
INV     gate4088  (.A(g5046), .Z(g9607) ) ;
INV     gate4089  (.A(g5062), .Z(g9613) ) ;
INV     gate4090  (.A(g5128), .Z(g9614) ) ;
INV     gate4091  (.A(g5452), .Z(II13236) ) ;
INV     gate4092  (.A(g5452), .Z(g9616) ) ;
INV     gate4093  (.A(g5794), .Z(II13240) ) ;
INV     gate4094  (.A(g5794), .Z(g9618) ) ;
INV     gate4095  (.A(g5845), .Z(g9619) ) ;
INV     gate4096  (.A(g6187), .Z(g9620) ) ;
INV     gate4097  (.A(g6423), .Z(g9621) ) ;
INV     gate4098  (.A(g6466), .Z(g9626) ) ;
INV     gate4099  (.A(g6527), .Z(g9630) ) ;
INV     gate4100  (.A(g6573), .Z(g9631) ) ;
INV     gate4101  (.A(g72), .Z(g9636) ) ;
INV     gate4102  (.A(g6751), .Z(II13252) ) ;
INV     gate4103  (.A(II13252), .Z(g9637) ) ;
INV     gate4104  (.A(g1620), .Z(g9638) ) ;
INV     gate4105  (.A(g1752), .Z(g9639) ) ;
INV     gate4106  (.A(g2016), .Z(g9644) ) ;
INV     gate4107  (.A(g2177), .Z(g9648) ) ;
INV     gate4108  (.A(g2441), .Z(g9653) ) ;
INV     gate4109  (.A(g2763), .Z(g9657) ) ;
INV     gate4110  (.A(g3267), .Z(g9660) ) ;
INV     gate4111  (.A(g3661), .Z(g9661) ) ;
INV     gate4112  (.A(g3983), .Z(g9662) ) ;
INV     gate4113  (.A(g5092), .Z(g9669) ) ;
INV     gate4114  (.A(g5022), .Z(g9670) ) ;
INV     gate4115  (.A(g5134), .Z(g9671) ) ;
INV     gate4116  (.A(g5390), .Z(g9672) ) ;
INV     gate4117  (.A(g5406), .Z(g9678) ) ;
INV     gate4118  (.A(g5475), .Z(g9679) ) ;
INV     gate4119  (.A(g5798), .Z(II13276) ) ;
INV     gate4120  (.A(g5798), .Z(g9681) ) ;
INV     gate4121  (.A(g6140), .Z(II13280) ) ;
INV     gate4122  (.A(g6140), .Z(g9683) ) ;
INV     gate4123  (.A(g6191), .Z(g9684) ) ;
INV     gate4124  (.A(g6533), .Z(g9685) ) ;
INV     gate4125  (.A(g73), .Z(g9686) ) ;
INV     gate4126  (.A(g110), .Z(II13287) ) ;
INV     gate4127  (.A(II13287), .Z(g9687) ) ;
INV     gate4128  (.A(g113), .Z(g9688) ) ;
INV     gate4129  (.A(g124), .Z(g9689) ) ;
INV     gate4130  (.A(g732), .Z(g9690) ) ;
INV     gate4131  (.A(g1706), .Z(g9691) ) ;
INV     gate4132  (.A(g1756), .Z(g9692) ) ;
INV     gate4133  (.A(g1886), .Z(g9693) ) ;
INV     gate4134  (.A(g2181), .Z(g9698) ) ;
INV     gate4135  (.A(g2311), .Z(g9699) ) ;
INV     gate4136  (.A(g2575), .Z(g9704) ) ;
INV     gate4137  (.A(g2741), .Z(g9708) ) ;
INV     gate4138  (.A(g3618), .Z(g9713) ) ;
INV     gate4139  (.A(g4012), .Z(g9714) ) ;
INV     gate4140  (.A(g5057), .Z(g9716) ) ;
INV     gate4141  (.A(g5097), .Z(g9721) ) ;
INV     gate4142  (.A(g5109), .Z(g9728) ) ;
INV     gate4143  (.A(g5138), .Z(g9729) ) ;
INV     gate4144  (.A(g5436), .Z(g9730) ) ;
INV     gate4145  (.A(g5366), .Z(g9731) ) ;
INV     gate4146  (.A(g5481), .Z(g9732) ) ;
INV     gate4147  (.A(g5736), .Z(g9733) ) ;
INV     gate4148  (.A(g5752), .Z(g9739) ) ;
INV     gate4149  (.A(g5821), .Z(g9740) ) ;
INV     gate4150  (.A(g6144), .Z(II13317) ) ;
INV     gate4151  (.A(g6144), .Z(g9742) ) ;
INV     gate4152  (.A(g6486), .Z(II13321) ) ;
INV     gate4153  (.A(g6486), .Z(g9744) ) ;
INV     gate4154  (.A(g6537), .Z(g9745) ) ;
INV     gate4155  (.A(g66), .Z(II13326) ) ;
INV     gate4156  (.A(II13326), .Z(g9746) ) ;
INV     gate4157  (.A(g86), .Z(II13329) ) ;
INV     gate4158  (.A(II13329), .Z(g9747) ) ;
INV     gate4159  (.A(g114), .Z(g9748) ) ;
INV     gate4160  (.A(g1691), .Z(g9749) ) ;
INV     gate4161  (.A(g1710), .Z(g9751) ) ;
INV     gate4162  (.A(g1840), .Z(g9752) ) ;
INV     gate4163  (.A(g1890), .Z(g9753) ) ;
INV     gate4164  (.A(g2020), .Z(g9754) ) ;
INV     gate4165  (.A(g2265), .Z(g9759) ) ;
INV     gate4166  (.A(g2315), .Z(g9760) ) ;
INV     gate4167  (.A(g2445), .Z(g9761) ) ;
INV     gate4168  (.A(g2748), .Z(g9766) ) ;
INV     gate4169  (.A(g3969), .Z(g9771) ) ;
INV     gate4170  (.A(g4146), .Z(II13352) ) ;
INV     gate4171  (.A(II13352), .Z(g9772) ) ;
INV     gate4172  (.A(g5073), .Z(g9776) ) ;
INV     gate4173  (.A(g5112), .Z(g9777) ) ;
INV     gate4174  (.A(g5069), .Z(g9778) ) ;
INV     gate4175  (.A(g5156), .Z(g9779) ) ;
INV     gate4176  (.A(g5343), .Z(II13360) ) ;
INV     gate4177  (.A(II13360), .Z(g9780) ) ;
INV     gate4178  (.A(g5401), .Z(g9792) ) ;
INV     gate4179  (.A(g5441), .Z(g9797) ) ;
INV     gate4180  (.A(g5456), .Z(g9804) ) ;
INV     gate4181  (.A(g5485), .Z(g9805) ) ;
INV     gate4182  (.A(g5782), .Z(g9806) ) ;
INV     gate4183  (.A(g5712), .Z(g9807) ) ;
INV     gate4184  (.A(g5827), .Z(g9808) ) ;
INV     gate4185  (.A(g6082), .Z(g9809) ) ;
INV     gate4186  (.A(g6098), .Z(g9815) ) ;
INV     gate4187  (.A(g6167), .Z(g9816) ) ;
INV     gate4188  (.A(g6490), .Z(II13374) ) ;
INV     gate4189  (.A(g6490), .Z(g9818) ) ;
INV     gate4190  (.A(g92), .Z(g9819) ) ;
INV     gate4191  (.A(g99), .Z(g9820) ) ;
INV     gate4192  (.A(g115), .Z(g9821) ) ;
INV     gate4193  (.A(g125), .Z(g9822) ) ;
INV     gate4194  (.A(g1825), .Z(g9824) ) ;
INV     gate4195  (.A(g1844), .Z(g9826) ) ;
INV     gate4196  (.A(g1974), .Z(g9827) ) ;
INV     gate4197  (.A(g2024), .Z(g9828) ) ;
INV     gate4198  (.A(g2250), .Z(g9829) ) ;
INV     gate4199  (.A(g2269), .Z(g9831) ) ;
INV     gate4200  (.A(g2399), .Z(g9832) ) ;
INV     gate4201  (.A(g2449), .Z(g9833) ) ;
INV     gate4202  (.A(g2579), .Z(g9834) ) ;
INV     gate4203  (.A(g2724), .Z(g9839) ) ;
INV     gate4204  (.A(g3274), .Z(g9842) ) ;
INV     gate4205  (.A(g4311), .Z(g9843) ) ;
INV     gate4206  (.A(g4462), .Z(g9848) ) ;
INV     gate4207  (.A(g5297), .Z(g9853) ) ;
INV     gate4208  (.A(g5343), .Z(g9856) ) ;
INV     gate4209  (.A(g5417), .Z(g9860) ) ;
INV     gate4210  (.A(g5459), .Z(g9861) ) ;
INV     gate4211  (.A(g5413), .Z(g9862) ) ;
INV     gate4212  (.A(g5503), .Z(g9863) ) ;
INV     gate4213  (.A(g5689), .Z(II13424) ) ;
INV     gate4214  (.A(II13424), .Z(g9864) ) ;
INV     gate4215  (.A(g5747), .Z(g9875) ) ;
INV     gate4216  (.A(g5787), .Z(g9880) ) ;
INV     gate4217  (.A(g5802), .Z(g9887) ) ;
INV     gate4218  (.A(g5831), .Z(g9888) ) ;
INV     gate4219  (.A(g6128), .Z(g9889) ) ;
INV     gate4220  (.A(g6058), .Z(g9890) ) ;
INV     gate4221  (.A(g6173), .Z(g9891) ) ;
INV     gate4222  (.A(g6428), .Z(g9892) ) ;
INV     gate4223  (.A(g6444), .Z(g9898) ) ;
INV     gate4224  (.A(g6513), .Z(g9899) ) ;
INV     gate4225  (.A(g6), .Z(g9900) ) ;
INV     gate4226  (.A(g84), .Z(g9901) ) ;
INV     gate4227  (.A(g100), .Z(g9902) ) ;
INV     gate4228  (.A(g681), .Z(g9903) ) ;
INV     gate4229  (.A(g802), .Z(g9905) ) ;
INV     gate4230  (.A(g1959), .Z(g9907) ) ;
INV     gate4231  (.A(g1978), .Z(g9909) ) ;
INV     gate4232  (.A(g2108), .Z(g9910) ) ;
INV     gate4233  (.A(g2384), .Z(g9911) ) ;
INV     gate4234  (.A(g2403), .Z(g9913) ) ;
INV     gate4235  (.A(g2533), .Z(g9914) ) ;
INV     gate4236  (.A(g2583), .Z(g9915) ) ;
INV     gate4237  (.A(g3625), .Z(g9916) ) ;
INV     gate4238  (.A(g4157), .Z(II13473) ) ;
INV     gate4239  (.A(II13473), .Z(g9917) ) ;
INV     gate4240  (.A(g4322), .Z(g9920) ) ;
INV     gate4241  (.A(g5644), .Z(g9924) ) ;
INV     gate4242  (.A(g5689), .Z(g9927) ) ;
INV     gate4243  (.A(g5763), .Z(g9931) ) ;
INV     gate4244  (.A(g5805), .Z(g9932) ) ;
INV     gate4245  (.A(g5759), .Z(g9933) ) ;
INV     gate4246  (.A(g5849), .Z(g9934) ) ;
INV     gate4247  (.A(g6035), .Z(II13483) ) ;
INV     gate4248  (.A(II13483), .Z(g9935) ) ;
INV     gate4249  (.A(g6093), .Z(g9946) ) ;
INV     gate4250  (.A(g6133), .Z(g9951) ) ;
INV     gate4251  (.A(g6148), .Z(g9958) ) ;
INV     gate4252  (.A(g6177), .Z(g9959) ) ;
INV     gate4253  (.A(g6474), .Z(g9960) ) ;
INV     gate4254  (.A(g6404), .Z(g9961) ) ;
INV     gate4255  (.A(g6519), .Z(g9962) ) ;
INV     gate4256  (.A(g7), .Z(g9963) ) ;
INV     gate4257  (.A(g126), .Z(g9964) ) ;
INV     gate4258  (.A(g127), .Z(g9965) ) ;
INV     gate4259  (.A(g1682), .Z(g9969) ) ;
INV     gate4260  (.A(g1714), .Z(g9970) ) ;
INV     gate4261  (.A(g2093), .Z(g9971) ) ;
INV     gate4262  (.A(g2112), .Z(g9973) ) ;
INV     gate4263  (.A(g2518), .Z(g9974) ) ;
INV     gate4264  (.A(g2537), .Z(g9976) ) ;
INV     gate4265  (.A(g2667), .Z(g9977) ) ;
INV     gate4266  (.A(g2756), .Z(g9978) ) ;
INV     gate4267  (.A(g3976), .Z(g9982) ) ;
INV     gate4268  (.A(g4239), .Z(g9983) ) ;
INV     gate4269  (.A(g4332), .Z(g9985) ) ;
INV     gate4270  (.A(g5077), .Z(g9989) ) ;
INV     gate4271  (.A(g5990), .Z(g9992) ) ;
INV     gate4272  (.A(g6035), .Z(g9995) ) ;
INV     gate4273  (.A(g6109), .Z(g9999) ) ;
INV     gate4274  (.A(g6151), .Z(g10000) ) ;
INV     gate4275  (.A(g6105), .Z(g10001) ) ;
INV     gate4276  (.A(g6195), .Z(g10002) ) ;
INV     gate4277  (.A(g6381), .Z(II13539) ) ;
INV     gate4278  (.A(II13539), .Z(g10003) ) ;
INV     gate4279  (.A(g6439), .Z(g10014) ) ;
INV     gate4280  (.A(g6479), .Z(g10019) ) ;
INV     gate4281  (.A(g6494), .Z(g10026) ) ;
INV     gate4282  (.A(g6523), .Z(g10027) ) ;
INV     gate4283  (.A(g8), .Z(g10028) ) ;
INV     gate4284  (.A(g94), .Z(II13548) ) ;
INV     gate4285  (.A(II13548), .Z(g10029) ) ;
INV     gate4286  (.A(g116), .Z(g10030) ) ;
INV     gate4287  (.A(g121), .Z(II13552) ) ;
INV     gate4288  (.A(II13552), .Z(g10031) ) ;
INV     gate4289  (.A(g562), .Z(g10032) ) ;
INV     gate4290  (.A(g655), .Z(g10033) ) ;
INV     gate4291  (.A(g1720), .Z(g10035) ) ;
INV     gate4292  (.A(g1816), .Z(g10036) ) ;
INV     gate4293  (.A(g1848), .Z(g10037) ) ;
INV     gate4294  (.A(g2241), .Z(g10038) ) ;
INV     gate4295  (.A(g2273), .Z(g10039) ) ;
INV     gate4296  (.A(g2652), .Z(g10040) ) ;
INV     gate4297  (.A(g2671), .Z(g10042) ) ;
INV     gate4298  (.A(g1632), .Z(g10043) ) ;
INV     gate4299  (.A(g5357), .Z(g10044) ) ;
INV     gate4300  (.A(g5421), .Z(g10047) ) ;
INV     gate4301  (.A(g6336), .Z(g10050) ) ;
INV     gate4302  (.A(g6381), .Z(g10053) ) ;
INV     gate4303  (.A(g6455), .Z(g10057) ) ;
INV     gate4304  (.A(g6497), .Z(g10058) ) ;
INV     gate4305  (.A(g6451), .Z(g10059) ) ;
INV     gate4306  (.A(g6541), .Z(g10060) ) ;
INV     gate4307  (.A(g6727), .Z(II13581) ) ;
INV     gate4308  (.A(II13581), .Z(g10061) ) ;
INV     gate4309  (.A(g9), .Z(g10072) ) ;
INV     gate4310  (.A(g134), .Z(g10073) ) ;
INV     gate4311  (.A(g718), .Z(g10074) ) ;
INV     gate4312  (.A(g1724), .Z(g10077) ) ;
INV     gate4313  (.A(g1854), .Z(g10078) ) ;
INV     gate4314  (.A(g1950), .Z(g10079) ) ;
INV     gate4315  (.A(g1982), .Z(g10080) ) ;
INV     gate4316  (.A(g2279), .Z(g10081) ) ;
INV     gate4317  (.A(g2375), .Z(g10082) ) ;
INV     gate4318  (.A(g2407), .Z(g10083) ) ;
INV     gate4319  (.A(g2837), .Z(g10084) ) ;
INV     gate4320  (.A(g1768), .Z(g10085) ) ;
INV     gate4321  (.A(g2193), .Z(g10086) ) ;
INV     gate4322  (.A(g4417), .Z(II13597) ) ;
INV     gate4323  (.A(II13597), .Z(g10087) ) ;
INV     gate4324  (.A(g5348), .Z(g10090) ) ;
INV     gate4325  (.A(g5703), .Z(g10093) ) ;
INV     gate4326  (.A(g5767), .Z(g10096) ) ;
INV     gate4327  (.A(g6682), .Z(g10099) ) ;
INV     gate4328  (.A(g6727), .Z(g10102) ) ;
INV     gate4329  (.A(g16), .Z(g10106) ) ;
INV     gate4330  (.A(g74), .Z(II13606) ) ;
INV     gate4331  (.A(II13606), .Z(g10107) ) ;
INV     gate4332  (.A(g120), .Z(g10108) ) ;
INV     gate4333  (.A(g135), .Z(g10109) ) ;
INV     gate4334  (.A(g661), .Z(g10110) ) ;
INV     gate4335  (.A(g1858), .Z(g10111) ) ;
INV     gate4336  (.A(g1988), .Z(g10112) ) ;
INV     gate4337  (.A(g2084), .Z(g10113) ) ;
INV     gate4338  (.A(g2116), .Z(g10114) ) ;
INV     gate4339  (.A(g2283), .Z(g10115) ) ;
INV     gate4340  (.A(g2413), .Z(g10116) ) ;
INV     gate4341  (.A(g2509), .Z(g10117) ) ;
INV     gate4342  (.A(g2541), .Z(g10118) ) ;
INV     gate4343  (.A(g2841), .Z(g10119) ) ;
INV     gate4344  (.A(g1902), .Z(g10120) ) ;
INV     gate4345  (.A(g2327), .Z(g10121) ) ;
INV     gate4346  (.A(g4294), .Z(II13623) ) ;
INV     gate4347  (.A(g5352), .Z(g10129) ) ;
INV     gate4348  (.A(g5694), .Z(g10130) ) ;
INV     gate4349  (.A(g6049), .Z(g10133) ) ;
INV     gate4350  (.A(g6113), .Z(g10136) ) ;
INV     gate4351  (.A(g136), .Z(g10139) ) ;
INV     gate4352  (.A(g19), .Z(g10140) ) ;
INV     gate4353  (.A(g79), .Z(II13634) ) ;
INV     gate4354  (.A(II13634), .Z(g10141) ) ;
INV     gate4355  (.A(g102), .Z(II13637) ) ;
INV     gate4356  (.A(II13637), .Z(g10142) ) ;
INV     gate4357  (.A(g568), .Z(g10143) ) ;
INV     gate4358  (.A(g728), .Z(g10147) ) ;
INV     gate4359  (.A(g1700), .Z(g10150) ) ;
INV     gate4360  (.A(g1992), .Z(g10151) ) ;
INV     gate4361  (.A(g2122), .Z(g10152) ) ;
INV     gate4362  (.A(g2417), .Z(g10153) ) ;
INV     gate4363  (.A(g2547), .Z(g10154) ) ;
INV     gate4364  (.A(g2643), .Z(g10155) ) ;
INV     gate4365  (.A(g2675), .Z(g10156) ) ;
INV     gate4366  (.A(g2036), .Z(g10157) ) ;
INV     gate4367  (.A(g2461), .Z(g10158) ) ;
INV     gate4368  (.A(g4477), .Z(g10159) ) ;
INV     gate4369  (.A(g5698), .Z(g10165) ) ;
INV     gate4370  (.A(g6040), .Z(g10166) ) ;
INV     gate4371  (.A(g6395), .Z(g10169) ) ;
INV     gate4372  (.A(g6459), .Z(g10172) ) ;
INV     gate4373  (.A(g28), .Z(g10175) ) ;
INV     gate4374  (.A(g44), .Z(g10176) ) ;
INV     gate4375  (.A(g1834), .Z(g10177) ) ;
INV     gate4376  (.A(g2126), .Z(g10178) ) ;
INV     gate4377  (.A(g2259), .Z(g10180) ) ;
INV     gate4378  (.A(g2551), .Z(g10181) ) ;
INV     gate4379  (.A(g2681), .Z(g10182) ) ;
INV     gate4380  (.A(g2595), .Z(g10183) ) ;
INV     gate4381  (.A(g4486), .Z(g10184) ) ;
INV     gate4382  (.A(g6044), .Z(g10190) ) ;
INV     gate4383  (.A(g6386), .Z(g10191) ) ;
INV     gate4384  (.A(g6741), .Z(g10194) ) ;
INV     gate4385  (.A(g31), .Z(g10197) ) ;
INV     gate4386  (.A(g106), .Z(II13672) ) ;
INV     gate4387  (.A(II13672), .Z(g10198) ) ;
INV     gate4388  (.A(g1968), .Z(g10199) ) ;
INV     gate4389  (.A(g2138), .Z(g10200) ) ;
INV     gate4390  (.A(g2393), .Z(g10203) ) ;
INV     gate4391  (.A(g2685), .Z(g10204) ) ;
INV     gate4392  (.A(g4489), .Z(g10206) ) ;
INV     gate4393  (.A(g6390), .Z(g10212) ) ;
INV     gate4394  (.A(g6732), .Z(g10213) ) ;
INV     gate4395  (.A(g128), .Z(II13684) ) ;
INV     gate4396  (.A(II13684), .Z(g10216) ) ;
INV     gate4397  (.A(g2102), .Z(g10217) ) ;
INV     gate4398  (.A(g2527), .Z(g10218) ) ;
INV     gate4399  (.A(g2697), .Z(g10219) ) ;
INV     gate4400  (.A(g4492), .Z(g10222) ) ;
INV     gate4401  (.A(g4561), .Z(g10223) ) ;
INV     gate4402  (.A(g6736), .Z(g10229) ) ;
INV     gate4403  (.A(g117), .Z(II13694) ) ;
INV     gate4404  (.A(II13694), .Z(g10230) ) ;
INV     gate4405  (.A(g2661), .Z(g10231) ) ;
INV     gate4406  (.A(g4527), .Z(g10232) ) ;
INV     gate4407  (.A(g4581), .Z(II13699) ) ;
INV     gate4408  (.A(II13699), .Z(g10233) ) ;
INV     gate4409  (.A(g4555), .Z(g10261) ) ;
INV     gate4410  (.A(g586), .Z(g10262) ) ;
INV     gate4411  (.A(g63), .Z(II13705) ) ;
INV     gate4412  (.A(II13705), .Z(g10272) ) ;
INV     gate4413  (.A(g136), .Z(II13708) ) ;
INV     gate4414  (.A(II13708), .Z(g10273) ) ;
INV     gate4415  (.A(g976), .Z(g10274) ) ;
INV     gate4416  (.A(g4584), .Z(g10275) ) ;
INV     gate4417  (.A(g4628), .Z(g10278) ) ;
INV     gate4418  (.A(g71), .Z(II13715) ) ;
INV     gate4419  (.A(II13715), .Z(g10287) ) ;
INV     gate4420  (.A(g890), .Z(II13718) ) ;
INV     gate4421  (.A(II13718), .Z(g10288) ) ;
INV     gate4422  (.A(g1319), .Z(g10289) ) ;
INV     gate4423  (.A(g3167), .Z(II13723) ) ;
INV     gate4424  (.A(II13723), .Z(g10295) ) ;
INV     gate4425  (.A(g4537), .Z(II13726) ) ;
INV     gate4426  (.A(g4459), .Z(g10308) ) ;
INV     gate4427  (.A(g4633), .Z(g10311) ) ;
INV     gate4428  (.A(g85), .Z(II13740) ) ;
INV     gate4429  (.A(II13740), .Z(g10319) ) ;
INV     gate4430  (.A(g817), .Z(g10320) ) ;
INV     gate4431  (.A(g3518), .Z(II13744) ) ;
INV     gate4432  (.A(II13744), .Z(g10323) ) ;
INV     gate4433  (.A(g4420), .Z(g10334) ) ;
INV     gate4434  (.A(g4483), .Z(g10335) ) ;
INV     gate4435  (.A(g5016), .Z(g10337) ) ;
INV     gate4436  (.A(g6754), .Z(II13759) ) ;
INV     gate4437  (.A(II13759), .Z(g10347) ) ;
INV     gate4438  (.A(g6755), .Z(II13762) ) ;
INV     gate4439  (.A(II13762), .Z(g10348) ) ;
INV     gate4440  (.A(g6956), .Z(g10349) ) ;
INV     gate4441  (.A(g6800), .Z(g10350) ) ;
INV     gate4442  (.A(g6802), .Z(g10351) ) ;
INV     gate4443  (.A(g6804), .Z(g10352) ) ;
INV     gate4444  (.A(g6803), .Z(g10353) ) ;
INV     gate4445  (.A(g6811), .Z(g10354) ) ;
INV     gate4446  (.A(g6816), .Z(g10355) ) ;
INV     gate4447  (.A(g6819), .Z(g10356) ) ;
INV     gate4448  (.A(g6825), .Z(g10357) ) ;
INV     gate4449  (.A(g6827), .Z(g10358) ) ;
INV     gate4450  (.A(g6830), .Z(g10359) ) ;
INV     gate4451  (.A(g6836), .Z(g10360) ) ;
INV     gate4452  (.A(g6841), .Z(g10361) ) ;
INV     gate4453  (.A(g6850), .Z(g10362) ) ;
INV     gate4454  (.A(g6868), .Z(II13779) ) ;
INV     gate4455  (.A(II13779), .Z(g10363) ) ;
INV     gate4456  (.A(g6869), .Z(g10364) ) ;
INV     gate4457  (.A(g6867), .Z(g10365) ) ;
INV     gate4458  (.A(g6895), .Z(g10366) ) ;
INV     gate4459  (.A(g6870), .Z(g10367) ) ;
INV     gate4460  (.A(g6887), .Z(g10368) ) ;
INV     gate4461  (.A(g6873), .Z(g10369) ) ;
INV     gate4462  (.A(g7095), .Z(g10370) ) ;
INV     gate4463  (.A(g6918), .Z(g10371) ) ;
INV     gate4464  (.A(g6900), .Z(g10372) ) ;
INV     gate4465  (.A(g6917), .Z(g10373) ) ;
INV     gate4466  (.A(g6903), .Z(g10374) ) ;
INV     gate4467  (.A(g6941), .Z(g10375) ) ;
INV     gate4468  (.A(g6923), .Z(g10376) ) ;
INV     gate4469  (.A(g6940), .Z(g10377) ) ;
INV     gate4470  (.A(g6926), .Z(g10378) ) ;
INV     gate4471  (.A(g6953), .Z(g10379) ) ;
INV     gate4472  (.A(g6960), .Z(g10380) ) ;
INV     gate4473  (.A(g6957), .Z(g10381) ) ;
INV     gate4474  (.A(g6958), .Z(g10382) ) ;
INV     gate4475  (.A(g6978), .Z(g10383) ) ;
INV     gate4476  (.A(g6971), .Z(II13802) ) ;
INV     gate4477  (.A(g6976), .Z(II13805) ) ;
INV     gate4478  (.A(II13805), .Z(g10385) ) ;
INV     gate4479  (.A(g6982), .Z(g10386) ) ;
INV     gate4480  (.A(g6996), .Z(g10387) ) ;
INV     gate4481  (.A(g6983), .Z(g10388) ) ;
INV     gate4482  (.A(g6986), .Z(g10389) ) ;
INV     gate4483  (.A(g6987), .Z(g10390) ) ;
INV     gate4484  (.A(g6988), .Z(g10391) ) ;
INV     gate4485  (.A(g6989), .Z(g10392) ) ;
INV     gate4486  (.A(g6991), .Z(g10393) ) ;
INV     gate4487  (.A(g6994), .Z(g10394) ) ;
INV     gate4488  (.A(g6995), .Z(g10395) ) ;
INV     gate4489  (.A(g6997), .Z(g10396) ) ;
INV     gate4490  (.A(g7018), .Z(g10397) ) ;
INV     gate4491  (.A(g6999), .Z(g10398) ) ;
INV     gate4492  (.A(g7017), .Z(g10399) ) ;
INV     gate4493  (.A(g7002), .Z(g10400) ) ;
INV     gate4494  (.A(g7041), .Z(g10401) ) ;
INV     gate4495  (.A(g7023), .Z(g10402) ) ;
INV     gate4496  (.A(g7040), .Z(g10403) ) ;
INV     gate4497  (.A(g7026), .Z(g10404) ) ;
INV     gate4498  (.A(g7064), .Z(g10405) ) ;
INV     gate4499  (.A(g7046), .Z(g10406) ) ;
INV     gate4500  (.A(g7063), .Z(g10407) ) ;
INV     gate4501  (.A(g7049), .Z(g10408) ) ;
INV     gate4502  (.A(g7087), .Z(g10409) ) ;
INV     gate4503  (.A(g7069), .Z(g10410) ) ;
INV     gate4504  (.A(g7086), .Z(g10411) ) ;
INV     gate4505  (.A(g7072), .Z(g10412) ) ;
INV     gate4506  (.A(g7110), .Z(g10413) ) ;
INV     gate4507  (.A(g7092), .Z(g10414) ) ;
INV     gate4508  (.A(g7109), .Z(g10415) ) ;
NOR2    gate4509  (.A(g25), .B(g22), .Z(g10318) ) ;
INV     gate4510  (.A(g10318), .Z(g10416) ) ;
INV     gate4511  (.A(g7117), .Z(g10417) ) ;
INV     gate4512  (.A(g8818), .Z(g10418) ) ;
INV     gate4513  (.A(g8821), .Z(g10419) ) ;
INV     gate4514  (.A(g9239), .Z(g10420) ) ;
INV     gate4515  (.A(g10053), .Z(g10427) ) ;
INV     gate4516  (.A(g9631), .Z(g10428) ) ;
INV     gate4517  (.A(g7148), .Z(g10429) ) ;
INV     gate4518  (.A(g7266), .Z(II13847) ) ;
INV     gate4519  (.A(II13847), .Z(g10430) ) ;
INV     gate4520  (.A(g9780), .Z(II13857) ) ;
INV     gate4521  (.A(II13857), .Z(g10473) ) ;
INV     gate4522  (.A(g8841), .Z(g10474) ) ;
INV     gate4523  (.A(g8844), .Z(g10475) ) ;
INV     gate4524  (.A(g10233), .Z(g10487) ) ;
INV     gate4525  (.A(g9259), .Z(g10489) ) ;
INV     gate4526  (.A(g9274), .Z(g10490) ) ;
INV     gate4527  (.A(g10102), .Z(g10497) ) ;
INV     gate4528  (.A(g7161), .Z(g10498) ) ;
INV     gate4529  (.A(g7474), .Z(II13872) ) ;
INV     gate4530  (.A(II13872), .Z(g10499) ) ;
INV     gate4531  (.A(g1233), .Z(II13875) ) ;
INV     gate4532  (.A(g8876), .Z(g10502) ) ;
INV     gate4533  (.A(g8879), .Z(g10503) ) ;
INV     gate4534  (.A(g8763), .Z(g10504) ) ;
INV     gate4535  (.A(g10233), .Z(g10509) ) ;
INV     gate4536  (.A(g9311), .Z(g10518) ) ;
INV     gate4537  (.A(g9326), .Z(g10519) ) ;
NAND2   gate4538  (.A(II12075), .B(II12076), .Z(g7598) ) ;
INV     gate4539  (.A(g7598), .Z(II13889) ) ;
INV     gate4540  (.A(II13889), .Z(g10521) ) ;
INV     gate4541  (.A(g1576), .Z(II13892) ) ;
INV     gate4542  (.A(g8922), .Z(g10530) ) ;
INV     gate4543  (.A(g8925), .Z(g10531) ) ;
INV     gate4544  (.A(g10233), .Z(g10532) ) ;
INV     gate4545  (.A(g8795), .Z(g10533) ) ;
INV     gate4546  (.A(g9392), .Z(g10540) ) ;
INV     gate4547  (.A(g9407), .Z(g10541) ) ;
INV     gate4548  (.A(g7196), .Z(g10542) ) ;
NAND2   gate4549  (.A(II12097), .B(II12098), .Z(g7620) ) ;
INV     gate4550  (.A(g7620), .Z(II13906) ) ;
INV     gate4551  (.A(II13906), .Z(g10544) ) ;
INV     gate4552  (.A(g8971), .Z(g10553) ) ;
INV     gate4553  (.A(g8974), .Z(g10554) ) ;
INV     gate4554  (.A(g9462), .Z(g10564) ) ;
INV     gate4555  (.A(g9021), .Z(g10570) ) ;
INV     gate4556  (.A(g10233), .Z(g10571) ) ;
INV     gate4557  (.A(g10233), .Z(g10572) ) ;
INV     gate4558  (.A(g9529), .Z(g10581) ) ;
INV     gate4559  (.A(g7116), .Z(g10582) ) ;
INV     gate4560  (.A(g10233), .Z(g10597) ) ;
INV     gate4561  (.A(g10233), .Z(g10606) ) ;
INV     gate4562  (.A(g10233), .Z(g10607) ) ;
INV     gate4563  (.A(g9155), .Z(g10608) ) ;
INV     gate4564  (.A(g10233), .Z(g10612) ) ;
INV     gate4565  (.A(g10233), .Z(g10613) ) ;
INV     gate4566  (.A(g10233), .Z(g10620) ) ;
NOR2    gate4567  (.A(g979), .B(g990), .Z(g7567) ) ;
INV     gate4568  (.A(g7567), .Z(g10621) ) ;
INV     gate4569  (.A(g7697), .Z(II13968) ) ;
INV     gate4570  (.A(II13968), .Z(g10627) ) ;
NOR2    gate4571  (.A(g1322), .B(g1333), .Z(g7601) ) ;
INV     gate4572  (.A(g7601), .Z(g10652) ) ;
INV     gate4573  (.A(g7733), .Z(II13979) ) ;
INV     gate4574  (.A(II13979), .Z(g10658) ) ;
INV     gate4575  (.A(g8928), .Z(g10664) ) ;
INV     gate4576  (.A(g7636), .Z(II13990) ) ;
INV     gate4577  (.A(II13990), .Z(g10678) ) ;
INV     gate4578  (.A(g8744), .Z(II13995) ) ;
INV     gate4579  (.A(II13995), .Z(g10685) ) ;
NAND2   gate4580  (.A(g4653), .B(g4688), .Z(g7836) ) ;
INV     gate4581  (.A(g7836), .Z(g10708) ) ;
INV     gate4582  (.A(g9104), .Z(II14006) ) ;
INV     gate4583  (.A(II14006), .Z(g10710) ) ;
NAND2   gate4584  (.A(g4843), .B(g4878), .Z(g7846) ) ;
INV     gate4585  (.A(g7846), .Z(g10725) ) ;
INV     gate4586  (.A(g9104), .Z(II14016) ) ;
INV     gate4587  (.A(II14016), .Z(g10727) ) ;
INV     gate4588  (.A(g8411), .Z(g10741) ) ;
INV     gate4589  (.A(g8411), .Z(g10761) ) ;
INV     gate4590  (.A(g8470), .Z(g10762) ) ;
INV     gate4591  (.A(g8912), .Z(II14033) ) ;
INV     gate4592  (.A(II14033), .Z(g10776) ) ;
INV     gate4593  (.A(g8470), .Z(g10794) ) ;
INV     gate4594  (.A(g7202), .Z(g10795) ) ;
INV     gate4595  (.A(g9772), .Z(g10804) ) ;
INV     gate4596  (.A(g9900), .Z(II14046) ) ;
INV     gate4597  (.A(II14046), .Z(g10805) ) ;
INV     gate4598  (.A(g9963), .Z(II14050) ) ;
INV     gate4599  (.A(II14050), .Z(g10812) ) ;
INV     gate4600  (.A(g9917), .Z(g10815) ) ;
INV     gate4601  (.A(g10028), .Z(II14054) ) ;
INV     gate4602  (.A(II14054), .Z(g10816) ) ;
INV     gate4603  (.A(g10087), .Z(g10830) ) ;
INV     gate4604  (.A(g9104), .Z(II14069) ) ;
INV     gate4605  (.A(II14069), .Z(g10851) ) ;
INV     gate4606  (.A(g8712), .Z(g10857) ) ;
INV     gate4607  (.A(g7567), .Z(g10872) ) ;
INV     gate4608  (.A(g7231), .Z(II14079) ) ;
INV     gate4609  (.A(II14079), .Z(g10877) ) ;
INV     gate4610  (.A(g7567), .Z(g10881) ) ;
INV     gate4611  (.A(g7601), .Z(g10882) ) ;
INV     gate4612  (.A(g7601), .Z(g10897) ) ;
INV     gate4613  (.A(g9007), .Z(g10960) ) ;
INV     gate4614  (.A(g9051), .Z(g10980) ) ;
INV     gate4615  (.A(g7824), .Z(II14119) ) ;
INV     gate4616  (.A(II14119), .Z(g10981) ) ;
INV     gate4617  (.A(g10274), .Z(g11011) ) ;
INV     gate4618  (.A(g10289), .Z(g11017) ) ;
NAND2   gate4619  (.A(g3080), .B(g3072), .Z(g8434) ) ;
INV     gate4620  (.A(g8434), .Z(g11026) ) ;
NAND2   gate4621  (.A(g218), .B(g215), .Z(g8292) ) ;
INV     gate4622  (.A(g8292), .Z(g11030) ) ;
NAND2   gate4623  (.A(g1171), .B(g1157), .Z(g8609) ) ;
INV     gate4624  (.A(g8609), .Z(g11031) ) ;
NAND2   gate4625  (.A(g3431), .B(g3423), .Z(g8500) ) ;
INV     gate4626  (.A(g8500), .Z(g11033) ) ;
NAND2   gate4627  (.A(g4057), .B(g4064), .Z(g7611) ) ;
INV     gate4628  (.A(g7611), .Z(g11034) ) ;
NAND2   gate4629  (.A(g1514), .B(g1500), .Z(g8632) ) ;
INV     gate4630  (.A(g8632), .Z(g11038) ) ;
NAND4   gate4631  (.A(g3267), .B(g3310), .C(g3281), .D(g3303), .Z(g8691) ) ;
INV     gate4632  (.A(g8691), .Z(g11042) ) ;
NAND2   gate4633  (.A(g3782), .B(g3774), .Z(g8561) ) ;
INV     gate4634  (.A(g8561), .Z(g11043) ) ;
NAND4   gate4635  (.A(g358), .B(g370), .C(g376), .D(g385), .Z(g8806) ) ;
INV     gate4636  (.A(g8806), .Z(II14158) ) ;
INV     gate4637  (.A(II14158), .Z(g11048) ) ;
NAND4   gate4638  (.A(g3618), .B(g3661), .C(g3632), .D(g3654), .Z(g8728) ) ;
INV     gate4639  (.A(g8728), .Z(g11110) ) ;
NAND4   gate4640  (.A(g3969), .B(g4012), .C(g3983), .D(g4005), .Z(g8751) ) ;
INV     gate4641  (.A(g8751), .Z(g11122) ) ;
INV     gate4642  (.A(g7993), .Z(g11128) ) ;
INV     gate4643  (.A(g7994), .Z(g11129) ) ;
INV     gate4644  (.A(g10233), .Z(II14192) ) ;
INV     gate4645  (.A(II14192), .Z(g11136) ) ;
INV     gate4646  (.A(g8032), .Z(g11143) ) ;
OR3     gate4647  (.A(g1056), .B(g1116), .C(II12583), .Z(g8417) ) ;
INV     gate4648  (.A(g8417), .Z(g11147) ) ;
INV     gate4649  (.A(g8085), .Z(g11164) ) ;
INV     gate4650  (.A(g8286), .Z(II14222) ) ;
INV     gate4651  (.A(II14222), .Z(g11165) ) ;
OR3     gate4652  (.A(g1399), .B(g1459), .C(II12611), .Z(g8476) ) ;
INV     gate4653  (.A(g8476), .Z(g11170) ) ;
INV     gate4654  (.A(g8134), .Z(g11181) ) ;
INV     gate4655  (.A(g8356), .Z(II14241) ) ;
INV     gate4656  (.A(II14241), .Z(g11182) ) ;
INV     gate4657  (.A(g8135), .Z(g11183) ) ;
INV     gate4658  (.A(g8038), .Z(g11192) ) ;
INV     gate4659  (.A(g7835), .Z(II14267) ) ;
INV     gate4660  (.A(II14267), .Z(g11202) ) ;
INV     gate4661  (.A(g8456), .Z(II14271) ) ;
INV     gate4662  (.A(II14271), .Z(g11204) ) ;
NOR4    gate4663  (.A(g4688), .B(g4681), .C(g4674), .D(g4646), .Z(g9602) ) ;
INV     gate4664  (.A(g9602), .Z(g11214) ) ;
INV     gate4665  (.A(g8285), .Z(g11215) ) ;
NOR4    gate4666  (.A(g4878), .B(g4871), .C(g4864), .D(g4836), .Z(g9664) ) ;
INV     gate4667  (.A(g9664), .Z(g11233) ) ;
INV     gate4668  (.A(g8355), .Z(g11234) ) ;
INV     gate4669  (.A(g8571), .Z(II14301) ) ;
INV     gate4670  (.A(II14301), .Z(g11235) ) ;
INV     gate4671  (.A(g8357), .Z(g11236) ) ;
INV     gate4672  (.A(g8805), .Z(II14305) ) ;
INV     gate4673  (.A(II14305), .Z(g11237) ) ;
INV     gate4674  (.A(g8405), .Z(g11249) ) ;
INV     gate4675  (.A(g7502), .Z(g11250) ) ;
INV     gate4676  (.A(g7515), .Z(g11268) ) ;
INV     gate4677  (.A(g7516), .Z(g11269) ) ;
INV     gate4678  (.A(g8607), .Z(II14326) ) ;
INV     gate4679  (.A(II14326), .Z(g11290) ) ;
INV     gate4680  (.A(g7526), .Z(g11291) ) ;
INV     gate4681  (.A(g7527), .Z(g11293) ) ;
INV     gate4682  (.A(g7598), .Z(g11294) ) ;
NAND2   gate4683  (.A(g4264), .B(g4258), .Z(g8967) ) ;
INV     gate4684  (.A(g8967), .Z(g11316) ) ;
INV     gate4685  (.A(g10233), .Z(II14346) ) ;
INV     gate4686  (.A(II14346), .Z(g11317) ) ;
INV     gate4687  (.A(g7542), .Z(g11324) ) ;
INV     gate4688  (.A(g7543), .Z(g11325) ) ;
INV     gate4689  (.A(g7620), .Z(g11336) ) ;
NOR2    gate4690  (.A(g3050), .B(g3010), .Z(g9015) ) ;
INV     gate4691  (.A(g9015), .Z(g11344) ) ;
INV     gate4692  (.A(g3303), .Z(II14365) ) ;
INV     gate4693  (.A(g8300), .Z(II14381) ) ;
INV     gate4694  (.A(II14381), .Z(g11367) ) ;
INV     gate4695  (.A(g7565), .Z(g11371) ) ;
INV     gate4696  (.A(g7566), .Z(g11373) ) ;
NOR2    gate4697  (.A(g3401), .B(g3361), .Z(g9061) ) ;
INV     gate4698  (.A(g9061), .Z(g11383) ) ;
INV     gate4699  (.A(g3654), .Z(II14395) ) ;
INV     gate4700  (.A(g8364), .Z(II14409) ) ;
INV     gate4701  (.A(II14409), .Z(g11398) ) ;
INV     gate4702  (.A(g7593), .Z(g11401) ) ;
INV     gate4703  (.A(g7594), .Z(g11402) ) ;
INV     gate4704  (.A(g7595), .Z(g11403) ) ;
INV     gate4705  (.A(g7596), .Z(g11404) ) ;
NOR2    gate4706  (.A(g3752), .B(g3712), .Z(g9100) ) ;
INV     gate4707  (.A(g9100), .Z(g11413) ) ;
INV     gate4708  (.A(g4005), .Z(II14424) ) ;
INV     gate4709  (.A(g7640), .Z(g11425) ) ;
INV     gate4710  (.A(g7615), .Z(g11428) ) ;
INV     gate4711  (.A(g7616), .Z(g11429) ) ;
INV     gate4712  (.A(g7617), .Z(g11430) ) ;
INV     gate4713  (.A(g7618), .Z(g11431) ) ;
INV     gate4714  (.A(g4191), .Z(II14450) ) ;
INV     gate4715  (.A(g10197), .Z(II14455) ) ;
INV     gate4716  (.A(II14455), .Z(g11450) ) ;
INV     gate4717  (.A(g7623), .Z(g11467) ) ;
INV     gate4718  (.A(g7624), .Z(g11468) ) ;
INV     gate4719  (.A(g7625), .Z(g11470) ) ;
INV     gate4720  (.A(g7626), .Z(g11471) ) ;
AND2    gate4721  (.A(g1205), .B(g1087), .Z(g7918) ) ;
INV     gate4722  (.A(g7918), .Z(g11472) ) ;
INV     gate4723  (.A(g10175), .Z(II14475) ) ;
INV     gate4724  (.A(II14475), .Z(g11498) ) ;
INV     gate4725  (.A(g7632), .Z(g11509) ) ;
INV     gate4726  (.A(g7633), .Z(g11510) ) ;
INV     gate4727  (.A(g7634), .Z(g11512) ) ;
AND2    gate4728  (.A(g1548), .B(g1430), .Z(g7948) ) ;
INV     gate4729  (.A(g7948), .Z(g11513) ) ;
INV     gate4730  (.A(g8481), .Z(g11519) ) ;
INV     gate4731  (.A(g10140), .Z(II14505) ) ;
INV     gate4732  (.A(II14505), .Z(g11547) ) ;
INV     gate4733  (.A(g7647), .Z(g11560) ) ;
INV     gate4734  (.A(g7648), .Z(g11562) ) ;
INV     gate4735  (.A(g8542), .Z(g11576) ) ;
INV     gate4736  (.A(g10106), .Z(II14537) ) ;
INV     gate4737  (.A(II14537), .Z(g11592) ) ;
INV     gate4738  (.A(g7659), .Z(g11608) ) ;
INV     gate4739  (.A(g7660), .Z(g11609) ) ;
INV     gate4740  (.A(g6875), .Z(g11615) ) ;
INV     gate4741  (.A(g8595), .Z(g11631) ) ;
INV     gate4742  (.A(g10072), .Z(II14550) ) ;
INV     gate4743  (.A(II14550), .Z(g11640) ) ;
INV     gate4744  (.A(g7674), .Z(g11652) ) ;
INV     gate4745  (.A(g6905), .Z(g11663) ) ;
INV     gate4746  (.A(g7689), .Z(g11677) ) ;
INV     gate4747  (.A(g802), .Z(II14563) ) ;
INV     gate4748  (.A(g9708), .Z(II14567) ) ;
INV     gate4749  (.A(II14567), .Z(g11686) ) ;
OR2     gate4750  (.A(g4072), .B(g4153), .Z(g7932) ) ;
INV     gate4751  (.A(g7932), .Z(II14570) ) ;
INV     gate4752  (.A(II14570), .Z(g11691) ) ;
INV     gate4753  (.A(g6928), .Z(g11702) ) ;
INV     gate4754  (.A(g8791), .Z(II14576) ) ;
INV     gate4755  (.A(II14576), .Z(g11705) ) ;
INV     gate4756  (.A(g8792), .Z(II14579) ) ;
INV     gate4757  (.A(II14579), .Z(g11706) ) ;
INV     gate4758  (.A(g9766), .Z(II14584) ) ;
INV     gate4759  (.A(II14584), .Z(g11709) ) ;
INV     gate4760  (.A(g8107), .Z(g11714) ) ;
INV     gate4761  (.A(g8818), .Z(II14589) ) ;
INV     gate4762  (.A(II14589), .Z(g11720) ) ;
INV     gate4763  (.A(g10074), .Z(g11721) ) ;
INV     gate4764  (.A(g9978), .Z(II14593) ) ;
INV     gate4765  (.A(II14593), .Z(g11724) ) ;
INV     gate4766  (.A(g8534), .Z(g11735) ) ;
INV     gate4767  (.A(g8165), .Z(g11736) ) ;
INV     gate4768  (.A(g10033), .Z(g11741) ) ;
INV     gate4769  (.A(g9340), .Z(II14602) ) ;
INV     gate4770  (.A(II14602), .Z(g11744) ) ;
INV     gate4771  (.A(g8587), .Z(g11753) ) ;
INV     gate4772  (.A(g8229), .Z(g11754) ) ;
INV     gate4773  (.A(g7964), .Z(g11762) ) ;
INV     gate4774  (.A(g8626), .Z(g11769) ) ;
INV     gate4775  (.A(g4185), .Z(II14619) ) ;
INV     gate4776  (.A(g8925), .Z(II14623) ) ;
INV     gate4777  (.A(II14623), .Z(g11772) ) ;
INV     gate4778  (.A(g9602), .Z(g11779) ) ;
NAND2   gate4779  (.A(g1018), .B(g1030), .Z(g7549) ) ;
INV     gate4780  (.A(g7549), .Z(g11786) ) ;
INV     gate4781  (.A(g7717), .Z(II14630) ) ;
INV     gate4782  (.A(II14630), .Z(g11790) ) ;
INV     gate4783  (.A(g9340), .Z(II14633) ) ;
INV     gate4784  (.A(II14633), .Z(g11793) ) ;
INV     gate4785  (.A(g7985), .Z(g11796) ) ;
INV     gate4786  (.A(g9664), .Z(g11810) ) ;
NAND2   gate4787  (.A(g5092), .B(g5084), .Z(g9724) ) ;
INV     gate4788  (.A(g9724), .Z(g11811) ) ;
INV     gate4789  (.A(g7567), .Z(g11812) ) ;
NAND2   gate4790  (.A(g1361), .B(g1373), .Z(g7582) ) ;
INV     gate4791  (.A(g7582), .Z(g11815) ) ;
INV     gate4792  (.A(g7717), .Z(g11819) ) ;
INV     gate4793  (.A(g7717), .Z(II14644) ) ;
INV     gate4794  (.A(II14644), .Z(g11820) ) ;
INV     gate4795  (.A(g7717), .Z(II14647) ) ;
INV     gate4796  (.A(II14647), .Z(g11823) ) ;
INV     gate4797  (.A(g9340), .Z(II14650) ) ;
INV     gate4798  (.A(II14650), .Z(g11826) ) ;
INV     gate4799  (.A(g9417), .Z(II14653) ) ;
INV     gate4800  (.A(II14653), .Z(g11829) ) ;
INV     gate4801  (.A(g8011), .Z(g11832) ) ;
INV     gate4802  (.A(g8026), .Z(g11833) ) ;
NAND2   gate4803  (.A(g5436), .B(g5428), .Z(g9800) ) ;
INV     gate4804  (.A(g9800), .Z(g11841) ) ;
INV     gate4805  (.A(g9746), .Z(II14660) ) ;
INV     gate4806  (.A(II14660), .Z(g11842) ) ;
INV     gate4807  (.A(g9747), .Z(II14663) ) ;
INV     gate4808  (.A(II14663), .Z(g11845) ) ;
INV     gate4809  (.A(g7601), .Z(g11849) ) ;
INV     gate4810  (.A(g7753), .Z(II14668) ) ;
INV     gate4811  (.A(II14668), .Z(g11852) ) ;
INV     gate4812  (.A(g7717), .Z(II14671) ) ;
INV     gate4813  (.A(II14671), .Z(g11855) ) ;
INV     gate4814  (.A(g8070), .Z(g11861) ) ;
NAND4   gate4815  (.A(g5276), .B(g5320), .C(g5290), .D(g5313), .Z(g10124) ) ;
INV     gate4816  (.A(g10124), .Z(g11865) ) ;
NAND2   gate4817  (.A(g5782), .B(g5774), .Z(g9883) ) ;
INV     gate4818  (.A(g9883), .Z(g11866) ) ;
INV     gate4819  (.A(g9332), .Z(II14679) ) ;
INV     gate4820  (.A(II14679), .Z(g11867) ) ;
INV     gate4821  (.A(g9185), .Z(g11868) ) ;
INV     gate4822  (.A(g7717), .Z(II14684) ) ;
INV     gate4823  (.A(II14684), .Z(g11872) ) ;
INV     gate4824  (.A(g7753), .Z(II14687) ) ;
INV     gate4825  (.A(II14687), .Z(g11875) ) ;
INV     gate4826  (.A(g9340), .Z(II14690) ) ;
INV     gate4827  (.A(II14690), .Z(g11878) ) ;
INV     gate4828  (.A(g8125), .Z(g11884) ) ;
NAND4   gate4829  (.A(g5623), .B(g5666), .C(g5637), .D(g5659), .Z(g10160) ) ;
INV     gate4830  (.A(g10160), .Z(g11888) ) ;
NAND2   gate4831  (.A(g6128), .B(g6120), .Z(g9954) ) ;
INV     gate4832  (.A(g9954), .Z(g11889) ) ;
INV     gate4833  (.A(g7717), .Z(II14702) ) ;
INV     gate4834  (.A(II14702), .Z(g11894) ) ;
INV     gate4835  (.A(g7717), .Z(II14705) ) ;
INV     gate4836  (.A(II14705), .Z(g11897) ) ;
INV     gate4837  (.A(g9417), .Z(II14708) ) ;
INV     gate4838  (.A(II14708), .Z(g11900) ) ;
NAND4   gate4839  (.A(g5969), .B(g6012), .C(g5983), .D(g6005), .Z(g10185) ) ;
INV     gate4840  (.A(g10185), .Z(g11910) ) ;
NAND2   gate4841  (.A(g6474), .B(g6466), .Z(g10022) ) ;
INV     gate4842  (.A(g10022), .Z(g11911) ) ;
INV     gate4843  (.A(g8989), .Z(g11912) ) ;
INV     gate4844  (.A(g7753), .Z(II14727) ) ;
INV     gate4845  (.A(II14727), .Z(g11917) ) ;
INV     gate4846  (.A(g7717), .Z(II14730) ) ;
INV     gate4847  (.A(II14730), .Z(g11920) ) ;
NAND4   gate4848  (.A(g6315), .B(g6358), .C(g6329), .D(g6351), .Z(g10207) ) ;
INV     gate4849  (.A(g10207), .Z(g11927) ) ;
INV     gate4850  (.A(g9534), .Z(II14742) ) ;
INV     gate4851  (.A(II14742), .Z(g11928) ) ;
INV     gate4852  (.A(g10029), .Z(II14745) ) ;
INV     gate4853  (.A(II14745), .Z(g11929) ) ;
INV     gate4854  (.A(g9281), .Z(g11930) ) ;
INV     gate4855  (.A(g10031), .Z(II14749) ) ;
INV     gate4856  (.A(II14749), .Z(g11931) ) ;
INV     gate4857  (.A(g7753), .Z(II14761) ) ;
INV     gate4858  (.A(II14761), .Z(g11941) ) ;
NAND4   gate4859  (.A(g6661), .B(g6704), .C(g6675), .D(g6697), .Z(g10224) ) ;
INV     gate4860  (.A(g10224), .Z(g11948) ) ;
INV     gate4861  (.A(g9581), .Z(II14773) ) ;
INV     gate4862  (.A(II14773), .Z(g11949) ) ;
INV     gate4863  (.A(g9153), .Z(g11963) ) ;
INV     gate4864  (.A(g9154), .Z(g11964) ) ;
INV     gate4865  (.A(g9636), .Z(II14797) ) ;
INV     gate4866  (.A(II14797), .Z(g11965) ) ;
INV     gate4867  (.A(g10107), .Z(II14800) ) ;
INV     gate4868  (.A(II14800), .Z(g11966) ) ;
INV     gate4869  (.A(g8056), .Z(II14823) ) ;
INV     gate4870  (.A(II14823), .Z(g11981) ) ;
INV     gate4871  (.A(g9186), .Z(g11984) ) ;
INV     gate4872  (.A(g9686), .Z(II14827) ) ;
INV     gate4873  (.A(II14827), .Z(g11985) ) ;
INV     gate4874  (.A(g10141), .Z(II14830) ) ;
INV     gate4875  (.A(II14830), .Z(g11986) ) ;
INV     gate4876  (.A(g10142), .Z(II14833) ) ;
INV     gate4877  (.A(II14833), .Z(g11987) ) ;
INV     gate4878  (.A(g9688), .Z(II14836) ) ;
INV     gate4879  (.A(II14836), .Z(g11988) ) ;
INV     gate4880  (.A(g9689), .Z(II14839) ) ;
INV     gate4881  (.A(II14839), .Z(g11989) ) ;
NAND2   gate4882  (.A(g1657), .B(g1624), .Z(g9485) ) ;
INV     gate4883  (.A(g9485), .Z(g11991) ) ;
INV     gate4884  (.A(g8092), .Z(II14862) ) ;
INV     gate4885  (.A(II14862), .Z(g12009) ) ;
INV     gate4886  (.A(g9213), .Z(g12012) ) ;
INV     gate4887  (.A(g9748), .Z(II14866) ) ;
INV     gate4888  (.A(II14866), .Z(g12013) ) ;
NAND2   gate4889  (.A(g1792), .B(g1760), .Z(g9538) ) ;
INV     gate4890  (.A(g9538), .Z(g12018) ) ;
NAND2   gate4891  (.A(g2217), .B(g2185), .Z(g9543) ) ;
INV     gate4892  (.A(g9543), .Z(g12021) ) ;
INV     gate4893  (.A(g9245), .Z(g12036) ) ;
INV     gate4894  (.A(g9819), .Z(II14893) ) ;
INV     gate4895  (.A(II14893), .Z(g12037) ) ;
INV     gate4896  (.A(g9820), .Z(II14896) ) ;
INV     gate4897  (.A(II14896), .Z(g12038) ) ;
INV     gate4898  (.A(g10198), .Z(II14899) ) ;
INV     gate4899  (.A(II14899), .Z(g12039) ) ;
INV     gate4900  (.A(g9821), .Z(II14902) ) ;
INV     gate4901  (.A(II14902), .Z(g12040) ) ;
INV     gate4902  (.A(g9822), .Z(II14905) ) ;
INV     gate4903  (.A(II14905), .Z(g12041) ) ;
NAND2   gate4904  (.A(g1926), .B(g1894), .Z(g9591) ) ;
INV     gate4905  (.A(g9591), .Z(g12047) ) ;
NAND2   gate4906  (.A(g2351), .B(g2319), .Z(g9595) ) ;
INV     gate4907  (.A(g9595), .Z(g12051) ) ;
NAND3   gate4908  (.A(g4669), .B(g4659), .C(g4653), .Z(g7690) ) ;
INV     gate4909  (.A(g7690), .Z(g12054) ) ;
INV     gate4910  (.A(g9901), .Z(II14932) ) ;
INV     gate4911  (.A(II14932), .Z(g12074) ) ;
INV     gate4912  (.A(g9902), .Z(II14935) ) ;
INV     gate4913  (.A(II14935), .Z(g12075) ) ;
INV     gate4914  (.A(g9280), .Z(g12076) ) ;
INV     gate4915  (.A(g10216), .Z(II14939) ) ;
INV     gate4916  (.A(II14939), .Z(g12077) ) ;
NAND2   gate4917  (.A(g2060), .B(g2028), .Z(g9645) ) ;
INV     gate4918  (.A(g9645), .Z(g12082) ) ;
NAND2   gate4919  (.A(g2485), .B(g2453), .Z(g9654) ) ;
INV     gate4920  (.A(g9654), .Z(g12086) ) ;
NAND3   gate4921  (.A(g4859), .B(g4849), .C(g4843), .Z(g7701) ) ;
INV     gate4922  (.A(g7701), .Z(g12088) ) ;
INV     gate4923  (.A(g9687), .Z(g12107) ) ;
INV     gate4924  (.A(g10230), .Z(II14964) ) ;
INV     gate4925  (.A(II14964), .Z(g12108) ) ;
INV     gate4926  (.A(g9964), .Z(II14967) ) ;
INV     gate4927  (.A(II14967), .Z(g12109) ) ;
INV     gate4928  (.A(g9965), .Z(II14970) ) ;
INV     gate4929  (.A(II14970), .Z(g12110) ) ;
NAND2   gate4930  (.A(g2619), .B(g2587), .Z(g9705) ) ;
INV     gate4931  (.A(g9705), .Z(g12122) ) ;
INV     gate4932  (.A(g10030), .Z(II14999) ) ;
INV     gate4933  (.A(II14999), .Z(g12143) ) ;
INV     gate4934  (.A(g9477), .Z(g12180) ) ;
INV     gate4935  (.A(g9478), .Z(g12181) ) ;
INV     gate4936  (.A(g10073), .Z(II15030) ) ;
INV     gate4937  (.A(II15030), .Z(g12182) ) ;
INV     gate4938  (.A(g10273), .Z(II15033) ) ;
INV     gate4939  (.A(II15033), .Z(g12183) ) ;
INV     gate4940  (.A(g799), .Z(II15036) ) ;
INV     gate4941  (.A(g10108), .Z(II15070) ) ;
INV     gate4942  (.A(II15070), .Z(g12217) ) ;
INV     gate4943  (.A(g10109), .Z(II15073) ) ;
INV     gate4944  (.A(II15073), .Z(g12218) ) ;
NOR2    gate4945  (.A(g5062), .B(g5022), .Z(g10338) ) ;
INV     gate4946  (.A(g10338), .Z(g12233) ) ;
INV     gate4947  (.A(g5313), .Z(II15102) ) ;
NOR2    gate4948  (.A(g5406), .B(g5366), .Z(g7139) ) ;
INV     gate4949  (.A(g7139), .Z(g12295) ) ;
INV     gate4950  (.A(g5659), .Z(II15144) ) ;
INV     gate4951  (.A(g9637), .Z(g12321) ) ;
INV     gate4952  (.A(g10176), .Z(II15162) ) ;
INV     gate4953  (.A(II15162), .Z(g12322) ) ;
INV     gate4954  (.A(g9340), .Z(g12337) ) ;
NOR2    gate4955  (.A(g5752), .B(g5712), .Z(g7158) ) ;
INV     gate4956  (.A(g7158), .Z(g12345) ) ;
INV     gate4957  (.A(g6005), .Z(II15190) ) ;
INV     gate4958  (.A(g10139), .Z(II15205) ) ;
INV     gate4959  (.A(II15205), .Z(g12367) ) ;
INV     gate4960  (.A(g637), .Z(II15208) ) ;
INV     gate4961  (.A(g9417), .Z(g12378) ) ;
INV     gate4962  (.A(g10119), .Z(II15223) ) ;
INV     gate4963  (.A(II15223), .Z(g12381) ) ;
INV     gate4964  (.A(g9920), .Z(g12399) ) ;
NOR2    gate4965  (.A(g6098), .B(g6058), .Z(g7175) ) ;
INV     gate4966  (.A(g7175), .Z(g12417) ) ;
INV     gate4967  (.A(g6351), .Z(II15238) ) ;
INV     gate4968  (.A(g9152), .Z(II15250) ) ;
INV     gate4969  (.A(II15250), .Z(g12430) ) ;
INV     gate4970  (.A(g9985), .Z(g12440) ) ;
NOR2    gate4971  (.A(g6444), .B(g6404), .Z(g7192) ) ;
INV     gate4972  (.A(g7192), .Z(g12465) ) ;
INV     gate4973  (.A(g6697), .Z(II15284) ) ;
INV     gate4974  (.A(g8515), .Z(II15295) ) ;
INV     gate4975  (.A(II15295), .Z(g12477) ) ;
INV     gate4976  (.A(g9340), .Z(g12487) ) ;
INV     gate4977  (.A(g10087), .Z(II15316) ) ;
INV     gate4978  (.A(II15316), .Z(g12490) ) ;
INV     gate4979  (.A(g9780), .Z(g12497) ) ;
INV     gate4980  (.A(g9417), .Z(g12543) ) ;
INV     gate4981  (.A(g8740), .Z(g12546) ) ;
INV     gate4982  (.A(g9864), .Z(g12563) ) ;
INV     gate4983  (.A(g7004), .Z(g12598) ) ;
INV     gate4984  (.A(g9935), .Z(g12614) ) ;
INV     gate4985  (.A(g9071), .Z(II15382) ) ;
INV     gate4986  (.A(II15382), .Z(g12640) ) ;
INV     gate4987  (.A(g7028), .Z(g12656) ) ;
INV     gate4988  (.A(g10003), .Z(g12672) ) ;
INV     gate4989  (.A(g7051), .Z(g12705) ) ;
INV     gate4990  (.A(g10061), .Z(g12721) ) ;
INV     gate4991  (.A(g9374), .Z(g12738) ) ;
INV     gate4992  (.A(g7074), .Z(g12749) ) ;
INV     gate4993  (.A(g10272), .Z(g12760) ) ;
INV     gate4994  (.A(g9856), .Z(g12778) ) ;
INV     gate4995  (.A(g9444), .Z(g12779) ) ;
INV     gate4996  (.A(g7097), .Z(g12790) ) ;
INV     gate4997  (.A(g10287), .Z(g12793) ) ;
INV     gate4998  (.A(g9927), .Z(g12804) ) ;
INV     gate4999  (.A(g9511), .Z(g12805) ) ;
INV     gate5000  (.A(g10319), .Z(g12811) ) ;
INV     gate5001  (.A(g8792), .Z(g12818) ) ;
INV     gate5002  (.A(g10233), .Z(g12820) ) ;
INV     gate5003  (.A(g9206), .Z(g12823) ) ;
INV     gate5004  (.A(g9995), .Z(g12830) ) ;
INV     gate5005  (.A(g9569), .Z(g12831) ) ;
INV     gate5006  (.A(g10877), .Z(II15448) ) ;
INV     gate5007  (.A(g10349), .Z(g12834) ) ;
INV     gate5008  (.A(g10352), .Z(g12835) ) ;
INV     gate5009  (.A(g10351), .Z(g12836) ) ;
INV     gate5010  (.A(g10354), .Z(g12837) ) ;
INV     gate5011  (.A(g10353), .Z(g12838) ) ;
INV     gate5012  (.A(g10350), .Z(g12839) ) ;
INV     gate5013  (.A(g10356), .Z(g12840) ) ;
INV     gate5014  (.A(g10357), .Z(g12841) ) ;
INV     gate5015  (.A(g10355), .Z(g12842) ) ;
INV     gate5016  (.A(g10359), .Z(g12843) ) ;
INV     gate5017  (.A(g10360), .Z(g12844) ) ;
INV     gate5018  (.A(g10358), .Z(g12845) ) ;
INV     gate5019  (.A(g10364), .Z(II15474) ) ;
INV     gate5020  (.A(II15474), .Z(g12857) ) ;
INV     gate5021  (.A(g10366), .Z(g12859) ) ;
INV     gate5022  (.A(g10368), .Z(g12860) ) ;
INV     gate5023  (.A(g10367), .Z(g12861) ) ;
INV     gate5024  (.A(g10370), .Z(g12862) ) ;
INV     gate5025  (.A(g10371), .Z(g12863) ) ;
INV     gate5026  (.A(g10373), .Z(g12864) ) ;
INV     gate5027  (.A(g10372), .Z(g12865) ) ;
INV     gate5028  (.A(g10369), .Z(g12866) ) ;
INV     gate5029  (.A(g10375), .Z(g12867) ) ;
INV     gate5030  (.A(g10377), .Z(g12868) ) ;
INV     gate5031  (.A(g10376), .Z(g12869) ) ;
INV     gate5032  (.A(g10374), .Z(g12870) ) ;
INV     gate5033  (.A(g10378), .Z(g12871) ) ;
INV     gate5034  (.A(g10379), .Z(g12872) ) ;
INV     gate5035  (.A(g10380), .Z(g12873) ) ;
INV     gate5036  (.A(g10383), .Z(g12874) ) ;
INV     gate5037  (.A(g10385), .Z(II15494) ) ;
INV     gate5038  (.A(II15494), .Z(g12875) ) ;
INV     gate5039  (.A(g10386), .Z(g12878) ) ;
INV     gate5040  (.A(g10381), .Z(g12879) ) ;
INV     gate5041  (.A(g10387), .Z(g12880) ) ;
INV     gate5042  (.A(g10388), .Z(g12881) ) ;
INV     gate5043  (.A(g10389), .Z(g12882) ) ;
INV     gate5044  (.A(g10390), .Z(g12883) ) ;
INV     gate5045  (.A(g10392), .Z(g12884) ) ;
INV     gate5046  (.A(g10382), .Z(g12885) ) ;
INV     gate5047  (.A(g10393), .Z(g12886) ) ;
INV     gate5048  (.A(g10394), .Z(g12887) ) ;
INV     gate5049  (.A(g10395), .Z(g12888) ) ;
INV     gate5050  (.A(g10396), .Z(g12889) ) ;
INV     gate5051  (.A(g10397), .Z(g12890) ) ;
INV     gate5052  (.A(g10399), .Z(g12891) ) ;
INV     gate5053  (.A(g10398), .Z(g12892) ) ;
INV     gate5054  (.A(g10391), .Z(g12893) ) ;
INV     gate5055  (.A(g10401), .Z(g12894) ) ;
INV     gate5056  (.A(g10403), .Z(g12895) ) ;
INV     gate5057  (.A(g10402), .Z(g12896) ) ;
INV     gate5058  (.A(g10400), .Z(g12897) ) ;
INV     gate5059  (.A(g10405), .Z(g12898) ) ;
INV     gate5060  (.A(g10407), .Z(g12899) ) ;
INV     gate5061  (.A(g10406), .Z(g12900) ) ;
INV     gate5062  (.A(g10404), .Z(g12901) ) ;
INV     gate5063  (.A(g10409), .Z(g12902) ) ;
INV     gate5064  (.A(g10411), .Z(g12903) ) ;
INV     gate5065  (.A(g10410), .Z(g12904) ) ;
INV     gate5066  (.A(g10408), .Z(g12905) ) ;
INV     gate5067  (.A(g10413), .Z(g12906) ) ;
INV     gate5068  (.A(g10415), .Z(g12907) ) ;
INV     gate5069  (.A(g10414), .Z(g12908) ) ;
INV     gate5070  (.A(g10412), .Z(g12909) ) ;
NOR2    gate5071  (.A(g9234), .B(g9206), .Z(g12235) ) ;
INV     gate5072  (.A(g12235), .Z(g12914) ) ;
INV     gate5073  (.A(g11867), .Z(II15533) ) ;
INV     gate5074  (.A(II15533), .Z(g12918) ) ;
INV     gate5075  (.A(g1227), .Z(II15536) ) ;
NOR4    gate5076  (.A(g10222), .B(g10206), .C(g10184), .D(g10335), .Z(g12228) ) ;
INV     gate5077  (.A(g12228), .Z(g12921) ) ;
NOR2    gate5078  (.A(g9269), .B(g9239), .Z(g12297) ) ;
INV     gate5079  (.A(g12297), .Z(g12922) ) ;
INV     gate5080  (.A(g1570), .Z(II15542) ) ;
NOR2    gate5081  (.A(g9300), .B(g9259), .Z(g12550) ) ;
INV     gate5082  (.A(g12550), .Z(g12929) ) ;
NOR2    gate5083  (.A(g9321), .B(g9274), .Z(g12347) ) ;
INV     gate5084  (.A(g12347), .Z(g12930) ) ;
INV     gate5085  (.A(g10430), .Z(II15550) ) ;
INV     gate5086  (.A(II15550), .Z(g12932) ) ;
NOR2    gate5087  (.A(g9381), .B(g9311), .Z(g12601) ) ;
INV     gate5088  (.A(g12601), .Z(g12936) ) ;
NOR2    gate5089  (.A(g9402), .B(g9326), .Z(g12419) ) ;
INV     gate5090  (.A(g12419), .Z(g12937) ) ;
INV     gate5091  (.A(g11928), .Z(II15556) ) ;
INV     gate5092  (.A(II15556), .Z(g12938) ) ;
INV     gate5093  (.A(g11744), .Z(g12940) ) ;
NOR2    gate5094  (.A(g9451), .B(g9392), .Z(g12659) ) ;
INV     gate5095  (.A(g12659), .Z(g12944) ) ;
NOR2    gate5096  (.A(g9472), .B(g9407), .Z(g12467) ) ;
INV     gate5097  (.A(g12467), .Z(g12945) ) ;
INV     gate5098  (.A(g11949), .Z(II15564) ) ;
INV     gate5099  (.A(II15564), .Z(g12946) ) ;
NOR2    gate5100  (.A(g9518), .B(g9462), .Z(g12708) ) ;
INV     gate5101  (.A(g12708), .Z(g12950) ) ;
INV     gate5102  (.A(g11965), .Z(II15569) ) ;
INV     gate5103  (.A(II15569), .Z(g12951) ) ;
INV     gate5104  (.A(g10499), .Z(II15572) ) ;
INV     gate5105  (.A(II15572), .Z(g12952) ) ;
INV     gate5106  (.A(g10430), .Z(II15577) ) ;
INV     gate5107  (.A(II15577), .Z(g12955) ) ;
INV     gate5108  (.A(g11790), .Z(g12967) ) ;
INV     gate5109  (.A(g11793), .Z(g12968) ) ;
NOR2    gate5110  (.A(g9576), .B(g9529), .Z(g12752) ) ;
INV     gate5111  (.A(g12752), .Z(g12975) ) ;
INV     gate5112  (.A(g11985), .Z(II15587) ) ;
INV     gate5113  (.A(II15587), .Z(g12976) ) ;
INV     gate5114  (.A(g11988), .Z(II15590) ) ;
INV     gate5115  (.A(II15590), .Z(g12977) ) ;
INV     gate5116  (.A(g11989), .Z(II15593) ) ;
INV     gate5117  (.A(II15593), .Z(g12978) ) ;
INV     gate5118  (.A(g10430), .Z(II15600) ) ;
INV     gate5119  (.A(II15600), .Z(g12983) ) ;
INV     gate5120  (.A(g11820), .Z(g12995) ) ;
INV     gate5121  (.A(g11823), .Z(g12996) ) ;
INV     gate5122  (.A(g11826), .Z(g12997) ) ;
INV     gate5123  (.A(g11829), .Z(g12998) ) ;
INV     gate5124  (.A(g12013), .Z(II15609) ) ;
INV     gate5125  (.A(II15609), .Z(g13003) ) ;
INV     gate5126  (.A(g11852), .Z(g13007) ) ;
INV     gate5127  (.A(g11855), .Z(g13008) ) ;
INV     gate5128  (.A(g12037), .Z(II15617) ) ;
INV     gate5129  (.A(II15617), .Z(g13009) ) ;
INV     gate5130  (.A(g12038), .Z(II15620) ) ;
INV     gate5131  (.A(II15620), .Z(g13010) ) ;
INV     gate5132  (.A(g12040), .Z(II15623) ) ;
INV     gate5133  (.A(II15623), .Z(g13011) ) ;
INV     gate5134  (.A(g12041), .Z(II15626) ) ;
INV     gate5135  (.A(II15626), .Z(g13012) ) ;
INV     gate5136  (.A(g11872), .Z(g13014) ) ;
INV     gate5137  (.A(g11875), .Z(g13015) ) ;
INV     gate5138  (.A(g11878), .Z(g13016) ) ;
INV     gate5139  (.A(g12074), .Z(II15633) ) ;
INV     gate5140  (.A(II15633), .Z(g13017) ) ;
INV     gate5141  (.A(g12075), .Z(II15636) ) ;
INV     gate5142  (.A(II15636), .Z(g13018) ) ;
INV     gate5143  (.A(g11894), .Z(g13022) ) ;
INV     gate5144  (.A(g11897), .Z(g13023) ) ;
INV     gate5145  (.A(g11900), .Z(g13024) ) ;
AND3    gate5146  (.A(g7655), .B(g7643), .C(g7627), .Z(g11018) ) ;
INV     gate5147  (.A(g11018), .Z(g13026) ) ;
INV     gate5148  (.A(g12109), .Z(II15647) ) ;
INV     gate5149  (.A(II15647), .Z(g13027) ) ;
INV     gate5150  (.A(g12110), .Z(II15650) ) ;
INV     gate5151  (.A(II15650), .Z(g13028) ) ;
INV     gate5152  (.A(g11917), .Z(g13033) ) ;
INV     gate5153  (.A(g11920), .Z(g13034) ) ;
INV     gate5154  (.A(g10981), .Z(g13036) ) ;
INV     gate5155  (.A(g10981), .Z(g13037) ) ;
INV     gate5156  (.A(g5308), .Z(II15663) ) ;
INV     gate5157  (.A(g12143), .Z(II15667) ) ;
INV     gate5158  (.A(II15667), .Z(g13041) ) ;
INV     gate5159  (.A(g11941), .Z(g13045) ) ;
INV     gate5160  (.A(g5654), .Z(II15677) ) ;
INV     gate5161  (.A(g11964), .Z(g13051) ) ;
INV     gate5162  (.A(g12182), .Z(II15682) ) ;
INV     gate5163  (.A(II15682), .Z(g13055) ) ;
INV     gate5164  (.A(g10981), .Z(g13061) ) ;
INV     gate5165  (.A(g10981), .Z(g13062) ) ;
INV     gate5166  (.A(g11705), .Z(g13064) ) ;
AND3    gate5167  (.A(g7244), .B(g7259), .C(II13862), .Z(g10476) ) ;
INV     gate5168  (.A(g10476), .Z(g13065) ) ;
INV     gate5169  (.A(g6000), .Z(II15697) ) ;
INV     gate5170  (.A(g11984), .Z(g13070) ) ;
INV     gate5171  (.A(g12217), .Z(II15702) ) ;
INV     gate5172  (.A(II15702), .Z(g13074) ) ;
INV     gate5173  (.A(g12218), .Z(II15705) ) ;
INV     gate5174  (.A(II15705), .Z(g13075) ) ;
INV     gate5175  (.A(g10981), .Z(g13082) ) ;
INV     gate5176  (.A(g6346), .Z(II15717) ) ;
INV     gate5177  (.A(g12012), .Z(g13087) ) ;
INV     gate5178  (.A(g10981), .Z(II15727) ) ;
INV     gate5179  (.A(II15727), .Z(g13096) ) ;
INV     gate5180  (.A(g6692), .Z(II15732) ) ;
INV     gate5181  (.A(g12322), .Z(II15736) ) ;
INV     gate5182  (.A(II15736), .Z(g13101) ) ;
NAND2   gate5183  (.A(g1116), .B(g7304), .Z(g10905) ) ;
INV     gate5184  (.A(g10905), .Z(g13103) ) ;
INV     gate5185  (.A(g10981), .Z(g13106) ) ;
INV     gate5186  (.A(g10476), .Z(g13107) ) ;
NAND2   gate5187  (.A(g1459), .B(g7352), .Z(g10935) ) ;
INV     gate5188  (.A(g10935), .Z(g13116) ) ;
INV     gate5189  (.A(g10981), .Z(g13117) ) ;
AND3    gate5190  (.A(g7475), .B(g7441), .C(g890), .Z(g10632) ) ;
INV     gate5191  (.A(g10632), .Z(g13120) ) ;
INV     gate5192  (.A(g10632), .Z(g13132) ) ;
NAND2   gate5193  (.A(g9483), .B(g1193), .Z(g11330) ) ;
INV     gate5194  (.A(g11330), .Z(g13133) ) ;
AND3    gate5195  (.A(g7704), .B(g5180), .C(g5188), .Z(g10823) ) ;
INV     gate5196  (.A(g10823), .Z(II15765) ) ;
INV     gate5197  (.A(II15765), .Z(g13138) ) ;
INV     gate5198  (.A(g10632), .Z(g13140) ) ;
NAND2   gate5199  (.A(g9536), .B(g1536), .Z(g11374) ) ;
INV     gate5200  (.A(g11374), .Z(g13141) ) ;
INV     gate5201  (.A(g10632), .Z(g13142) ) ;
INV     gate5202  (.A(g10430), .Z(II15773) ) ;
INV     gate5203  (.A(II15773), .Z(g13144) ) ;
INV     gate5204  (.A(g10632), .Z(g13173) ) ;
INV     gate5205  (.A(g10741), .Z(g13174) ) ;
NAND2   gate5206  (.A(g7304), .B(g1116), .Z(g10909) ) ;
INV     gate5207  (.A(g10909), .Z(g13175) ) ;
INV     gate5208  (.A(g10430), .Z(II15782) ) ;
INV     gate5209  (.A(II15782), .Z(g13177) ) ;
INV     gate5210  (.A(g10909), .Z(g13188) ) ;
INV     gate5211  (.A(g10762), .Z(g13189) ) ;
NAND2   gate5212  (.A(g7352), .B(g1459), .Z(g10939) ) ;
INV     gate5213  (.A(g10939), .Z(g13190) ) ;
INV     gate5214  (.A(g10430), .Z(II15788) ) ;
INV     gate5215  (.A(II15788), .Z(g13191) ) ;
INV     gate5216  (.A(g10632), .Z(g13209) ) ;
INV     gate5217  (.A(g10909), .Z(g13215) ) ;
INV     gate5218  (.A(g10939), .Z(g13216) ) ;
AND3    gate5219  (.A(g7246), .B(g7392), .C(II13937), .Z(g10590) ) ;
INV     gate5220  (.A(g10590), .Z(g13222) ) ;
NOR3    gate5221  (.A(g8848), .B(g8993), .C(g376), .Z(g11607) ) ;
INV     gate5222  (.A(g11607), .Z(II15800) ) ;
INV     gate5223  (.A(II15800), .Z(g13223) ) ;
INV     gate5224  (.A(g10632), .Z(g13239) ) ;
INV     gate5225  (.A(g10939), .Z(g13246) ) ;
INV     gate5226  (.A(g10590), .Z(g13249) ) ;
INV     gate5227  (.A(g11128), .Z(II15811) ) ;
INV     gate5228  (.A(II15811), .Z(g13250) ) ;
INV     gate5229  (.A(g11129), .Z(II15814) ) ;
INV     gate5230  (.A(II15814), .Z(g13251) ) ;
INV     gate5231  (.A(g10632), .Z(g13255) ) ;
INV     gate5232  (.A(g11143), .Z(II15821) ) ;
INV     gate5233  (.A(II15821), .Z(g13258) ) ;
INV     gate5234  (.A(g1116), .Z(II15824) ) ;
INV     gate5235  (.A(g10416), .Z(II15831) ) ;
INV     gate5236  (.A(II15831), .Z(g13267) ) ;
INV     gate5237  (.A(g11164), .Z(II15834) ) ;
INV     gate5238  (.A(II15834), .Z(g13271) ) ;
INV     gate5239  (.A(g1459), .Z(II15837) ) ;
NAND2   gate5240  (.A(g6961), .B(g10308), .Z(g10738) ) ;
INV     gate5241  (.A(g10738), .Z(g13278) ) ;
INV     gate5242  (.A(g11181), .Z(II15843) ) ;
INV     gate5243  (.A(II15843), .Z(g13279) ) ;
INV     gate5244  (.A(g11183), .Z(II15846) ) ;
INV     gate5245  (.A(II15846), .Z(g13280) ) ;
NOR2    gate5246  (.A(g7690), .B(g7827), .Z(g10831) ) ;
INV     gate5247  (.A(g10831), .Z(g13297) ) ;
INV     gate5248  (.A(g11215), .Z(II15862) ) ;
INV     gate5249  (.A(II15862), .Z(g13298) ) ;
NOR2    gate5250  (.A(g7701), .B(g7840), .Z(g10862) ) ;
INV     gate5251  (.A(g10862), .Z(g13301) ) ;
INV     gate5252  (.A(g12321), .Z(g13302) ) ;
INV     gate5253  (.A(g11234), .Z(II15869) ) ;
INV     gate5254  (.A(II15869), .Z(g13303) ) ;
INV     gate5255  (.A(g11236), .Z(II15872) ) ;
INV     gate5256  (.A(II15872), .Z(g13304) ) ;
INV     gate5257  (.A(g11048), .Z(g13305) ) ;
INV     gate5258  (.A(g11249), .Z(II15878) ) ;
INV     gate5259  (.A(II15878), .Z(g13311) ) ;
INV     gate5260  (.A(g11048), .Z(g13312) ) ;
NOR3    gate5261  (.A(g1189), .B(g7715), .C(g7749), .Z(g10893) ) ;
INV     gate5262  (.A(g10893), .Z(g13314) ) ;
NOR3    gate5263  (.A(g1532), .B(g7751), .C(g7778), .Z(g10918) ) ;
INV     gate5264  (.A(g10918), .Z(g13322) ) ;
INV     gate5265  (.A(g11048), .Z(g13323) ) ;
INV     gate5266  (.A(g10430), .Z(II15893) ) ;
INV     gate5267  (.A(II15893), .Z(g13329) ) ;
INV     gate5268  (.A(g11048), .Z(g13334) ) ;
INV     gate5269  (.A(g10430), .Z(II15906) ) ;
INV     gate5270  (.A(II15906), .Z(g13350) ) ;
INV     gate5271  (.A(g10430), .Z(II15915) ) ;
INV     gate5272  (.A(II15915), .Z(g13394) ) ;
INV     gate5273  (.A(g12381), .Z(II15918) ) ;
INV     gate5274  (.A(II15918), .Z(g13409) ) ;
INV     gate5275  (.A(g12381), .Z(II15921) ) ;
INV     gate5276  (.A(II15921), .Z(g13410) ) ;
INV     gate5277  (.A(g11963), .Z(g13412) ) ;
OR2     gate5278  (.A(g8359), .B(g8292), .Z(g11737) ) ;
INV     gate5279  (.A(g11737), .Z(g13413) ) ;
INV     gate5280  (.A(g11048), .Z(g13414) ) ;
INV     gate5281  (.A(g10430), .Z(II15929) ) ;
INV     gate5282  (.A(II15929), .Z(g13416) ) ;
INV     gate5283  (.A(g12381), .Z(II15932) ) ;
INV     gate5284  (.A(II15932), .Z(g13431) ) ;
NAND4   gate5285  (.A(g358), .B(g8944), .C(g376), .D(g385), .Z(g11676) ) ;
INV     gate5286  (.A(g11676), .Z(II15937) ) ;
INV     gate5287  (.A(II15937), .Z(g13437) ) ;
INV     gate5288  (.A(g11048), .Z(g13458) ) ;
INV     gate5289  (.A(g12381), .Z(II15942) ) ;
INV     gate5290  (.A(II15942), .Z(g13460) ) ;
INV     gate5291  (.A(g10476), .Z(g13463) ) ;
INV     gate5292  (.A(g11048), .Z(g13474) ) ;
INV     gate5293  (.A(g12381), .Z(II15954) ) ;
INV     gate5294  (.A(II15954), .Z(g13477) ) ;
NOR2    gate5295  (.A(g8431), .B(g8434), .Z(g11270) ) ;
INV     gate5296  (.A(g11270), .Z(g13483) ) ;
INV     gate5297  (.A(g10981), .Z(g13484) ) ;
INV     gate5298  (.A(g10476), .Z(g13485) ) ;
INV     gate5299  (.A(g11912), .Z(g13494) ) ;
NOR2    gate5300  (.A(g8497), .B(g8500), .Z(g11303) ) ;
INV     gate5301  (.A(g11303), .Z(g13504) ) ;
INV     gate5302  (.A(g10981), .Z(g13505) ) ;
NOR2    gate5303  (.A(g8509), .B(g7611), .Z(g10808) ) ;
INV     gate5304  (.A(g10808), .Z(g13506) ) ;
INV     gate5305  (.A(g11290), .Z(II15981) ) ;
INV     gate5306  (.A(II15981), .Z(g13510) ) ;
INV     gate5307  (.A(g12381), .Z(II15987) ) ;
INV     gate5308  (.A(II15987), .Z(g13514) ) ;
NOR2    gate5309  (.A(g8558), .B(g8561), .Z(g11357) ) ;
INV     gate5310  (.A(g11357), .Z(g13521) ) ;
INV     gate5311  (.A(g10981), .Z(g13522) ) ;
AND3    gate5312  (.A(g10295), .B(g3171), .C(g3179), .Z(g12641) ) ;
INV     gate5313  (.A(g12641), .Z(g13530) ) ;
NOR4    gate5314  (.A(g8052), .B(g9197), .C(g9174), .D(g9050), .Z(g11148) ) ;
INV     gate5315  (.A(g11148), .Z(II16010) ) ;
INV     gate5316  (.A(II16010), .Z(g13545) ) ;
AND3    gate5317  (.A(g10323), .B(g3522), .C(g3530), .Z(g12692) ) ;
INV     gate5318  (.A(g12692), .Z(g13555) ) ;
NOR2    gate5319  (.A(g7686), .B(g7836), .Z(g11006) ) ;
INV     gate5320  (.A(g11006), .Z(g13565) ) ;
NAND2   gate5321  (.A(g7845), .B(g7868), .Z(g10951) ) ;
INV     gate5322  (.A(g10951), .Z(g13569) ) ;
NOR4    gate5323  (.A(g8088), .B(g9226), .C(g9200), .D(g9091), .Z(g11171) ) ;
INV     gate5324  (.A(g11171), .Z(II16024) ) ;
INV     gate5325  (.A(II16024), .Z(g13574) ) ;
INV     gate5326  (.A(g12381), .Z(II16028) ) ;
INV     gate5327  (.A(II16028), .Z(g13583) ) ;
AND3    gate5328  (.A(g7121), .B(g3873), .C(g3881), .Z(g12735) ) ;
INV     gate5329  (.A(g12735), .Z(g13584) ) ;
NAND2   gate5330  (.A(g7971), .B(g8133), .Z(g10556) ) ;
INV     gate5331  (.A(g10556), .Z(g13593) ) ;
NOR2    gate5332  (.A(g7693), .B(g7846), .Z(g11012) ) ;
INV     gate5333  (.A(g11012), .Z(g13594) ) ;
INV     gate5334  (.A(g10951), .Z(g13595) ) ;
NAND2   gate5335  (.A(g7867), .B(g7886), .Z(g10971) ) ;
INV     gate5336  (.A(g10971), .Z(g13596) ) ;
INV     gate5337  (.A(g10430), .Z(II16040) ) ;
INV     gate5338  (.A(II16040), .Z(g13605) ) ;
INV     gate5339  (.A(g10556), .Z(g13620) ) ;
NAND2   gate5340  (.A(g7992), .B(g8179), .Z(g10573) ) ;
INV     gate5341  (.A(g10573), .Z(g13621) ) ;
INV     gate5342  (.A(g10951), .Z(g13624) ) ;
INV     gate5343  (.A(g10971), .Z(g13625) ) ;
NOR2    gate5344  (.A(g3061), .B(g8620), .Z(g11273) ) ;
INV     gate5345  (.A(g11273), .Z(g13626) ) ;
INV     gate5346  (.A(g10556), .Z(g13637) ) ;
INV     gate5347  (.A(g10430), .Z(II16057) ) ;
INV     gate5348  (.A(II16057), .Z(g13638) ) ;
INV     gate5349  (.A(g10573), .Z(g13655) ) ;
INV     gate5350  (.A(g10971), .Z(g13663) ) ;
NOR2    gate5351  (.A(g8620), .B(g3057), .Z(g11252) ) ;
INV     gate5352  (.A(g11252), .Z(g13664) ) ;
NOR2    gate5353  (.A(g3412), .B(g8647), .Z(g11306) ) ;
INV     gate5354  (.A(g11306), .Z(g13665) ) ;
INV     gate5355  (.A(g10556), .Z(g13675) ) ;
INV     gate5356  (.A(g10573), .Z(g13679) ) ;
INV     gate5357  (.A(g10430), .Z(II16077) ) ;
INV     gate5358  (.A(II16077), .Z(g13680) ) ;
NOR2    gate5359  (.A(g8647), .B(g3408), .Z(g11280) ) ;
INV     gate5360  (.A(g11280), .Z(g13706) ) ;
NOR2    gate5361  (.A(g3763), .B(g8669), .Z(g11360) ) ;
INV     gate5362  (.A(g11360), .Z(g13707) ) ;
INV     gate5363  (.A(g10573), .Z(g13715) ) ;
INV     gate5364  (.A(g10430), .Z(II16090) ) ;
INV     gate5365  (.A(II16090), .Z(g13716) ) ;
INV     gate5366  (.A(g10951), .Z(g13729) ) ;
NOR2    gate5367  (.A(g8669), .B(g3759), .Z(g11313) ) ;
INV     gate5368  (.A(g11313), .Z(g13736) ) ;
INV     gate5369  (.A(g10430), .Z(II16102) ) ;
INV     gate5370  (.A(II16102), .Z(g13745) ) ;
INV     gate5371  (.A(g10971), .Z(g13763) ) ;
INV     gate5372  (.A(g10430), .Z(II16117) ) ;
INV     gate5373  (.A(II16117), .Z(g13782) ) ;
INV     gate5374  (.A(g11868), .Z(II16120) ) ;
INV     gate5375  (.A(II16120), .Z(g13793) ) ;
INV     gate5376  (.A(g10430), .Z(II16135) ) ;
INV     gate5377  (.A(II16135), .Z(g13809) ) ;
INV     gate5378  (.A(g10430), .Z(II16150) ) ;
INV     gate5379  (.A(II16150), .Z(g13835) ) ;
INV     gate5380  (.A(g11237), .Z(II16160) ) ;
INV     gate5381  (.A(II16160), .Z(g13856) ) ;
INV     gate5382  (.A(g11930), .Z(II16163) ) ;
INV     gate5383  (.A(II16163), .Z(g13857) ) ;
INV     gate5384  (.A(g3321), .Z(II16168) ) ;
NOR2    gate5385  (.A(g8964), .B(g8967), .Z(g11493) ) ;
INV     gate5386  (.A(g11493), .Z(g13868) ) ;
INV     gate5387  (.A(g10831), .Z(g13869) ) ;
NAND2   gate5388  (.A(g10295), .B(g8864), .Z(g11432) ) ;
INV     gate5389  (.A(g11432), .Z(g13876) ) ;
NAND2   gate5390  (.A(II14369), .B(II14370), .Z(g11350) ) ;
INV     gate5391  (.A(g11350), .Z(g13877) ) ;
INV     gate5392  (.A(g3672), .Z(II16181) ) ;
INV     gate5393  (.A(g10862), .Z(g13885) ) ;
INV     gate5394  (.A(g3281), .Z(II16193) ) ;
NAND2   gate5395  (.A(g10323), .B(g8906), .Z(g11480) ) ;
INV     gate5396  (.A(g11480), .Z(g13901) ) ;
NAND2   gate5397  (.A(II14399), .B(II14400), .Z(g11389) ) ;
INV     gate5398  (.A(g11389), .Z(g13902) ) ;
INV     gate5399  (.A(g4023), .Z(II16201) ) ;
INV     gate5400  (.A(g3632), .Z(II16217) ) ;
NAND2   gate5401  (.A(g7121), .B(g8958), .Z(g11534) ) ;
INV     gate5402  (.A(g11534), .Z(g13932) ) ;
NAND2   gate5403  (.A(II14428), .B(II14429), .Z(g11419) ) ;
INV     gate5404  (.A(g11419), .Z(g13933) ) ;
NAND2   gate5405  (.A(g7195), .B(g7115), .Z(g10520) ) ;
INV     gate5406  (.A(g10520), .Z(II16231) ) ;
INV     gate5407  (.A(II16231), .Z(g13943) ) ;
INV     gate5408  (.A(g3983), .Z(II16246) ) ;
INV     gate5409  (.A(g11048), .Z(g13975) ) ;
NAND2   gate5410  (.A(g1221), .B(g7918), .Z(g11130) ) ;
INV     gate5411  (.A(g11130), .Z(g13976) ) ;
NOR3    gate5412  (.A(g7928), .B(g4801), .C(g9030), .Z(g11261) ) ;
INV     gate5413  (.A(g11261), .Z(g13995) ) ;
INV     gate5414  (.A(g11048), .Z(g13999) ) ;
NAND2   gate5415  (.A(g1564), .B(g7948), .Z(g11149) ) ;
INV     gate5416  (.A(g11149), .Z(g14004) ) ;
NOR3    gate5417  (.A(g7953), .B(g4991), .C(g9064), .Z(g11283) ) ;
INV     gate5418  (.A(g11283), .Z(g14029) ) ;
INV     gate5419  (.A(g12107), .Z(II16289) ) ;
INV     gate5420  (.A(II16289), .Z(g14031) ) ;
INV     gate5421  (.A(g11048), .Z(g14032) ) ;
INV     gate5422  (.A(g11048), .Z(g14034) ) ;
INV     gate5423  (.A(g11048), .Z(g14063) ) ;
INV     gate5424  (.A(g11048), .Z(g14065) ) ;
NAND4   gate5425  (.A(g8993), .B(g376), .C(g365), .D(g370), .Z(g11326) ) ;
INV     gate5426  (.A(g11326), .Z(g14095) ) ;
INV     gate5427  (.A(g878), .Z(II16328) ) ;
INV     gate5428  (.A(g881), .Z(II16345) ) ;
INV     gate5429  (.A(g884), .Z(II16357) ) ;
INV     gate5430  (.A(g12381), .Z(g14149) ) ;
INV     gate5431  (.A(g12381), .Z(g14150) ) ;
INV     gate5432  (.A(g11048), .Z(g14166) ) ;
INV     gate5433  (.A(g887), .Z(II16371) ) ;
INV     gate5434  (.A(g12381), .Z(g14169) ) ;
INV     gate5435  (.A(g12076), .Z(g14173) ) ;
INV     gate5436  (.A(g11048), .Z(g14179) ) ;
INV     gate5437  (.A(g12381), .Z(g14183) ) ;
INV     gate5438  (.A(g12381), .Z(g14184) ) ;
NOR2    gate5439  (.A(g7980), .B(g7964), .Z(g11346) ) ;
INV     gate5440  (.A(g11346), .Z(g14186) ) ;
INV     gate5441  (.A(g859), .Z(II16391) ) ;
INV     gate5442  (.A(g12381), .Z(g14191) ) ;
NOR2    gate5443  (.A(g8021), .B(g7985), .Z(g11385) ) ;
INV     gate5444  (.A(g11385), .Z(g14192) ) ;
NOR2    gate5445  (.A(g9721), .B(g9724), .Z(g12160) ) ;
INV     gate5446  (.A(g12160), .Z(g14197) ) ;
INV     gate5447  (.A(g12180), .Z(g14198) ) ;
INV     gate5448  (.A(g869), .Z(II16401) ) ;
INV     gate5449  (.A(g12381), .Z(g14203) ) ;
NAND2   gate5450  (.A(g7753), .B(g7717), .Z(g12155) ) ;
INV     gate5451  (.A(g12155), .Z(g14204) ) ;
INV     gate5452  (.A(g12381), .Z(g14205) ) ;
NOR2    gate5453  (.A(g8059), .B(g8011), .Z(g11563) ) ;
INV     gate5454  (.A(g11563), .Z(g14208) ) ;
NOR2    gate5455  (.A(g8080), .B(g8026), .Z(g11415) ) ;
INV     gate5456  (.A(g11415), .Z(g14209) ) ;
NOR2    gate5457  (.A(g9797), .B(g9800), .Z(g12198) ) ;
INV     gate5458  (.A(g12198), .Z(g14215) ) ;
INV     gate5459  (.A(g875), .Z(II16417) ) ;
INV     gate5460  (.A(g12381), .Z(g14219) ) ;
NOR2    gate5461  (.A(g8114), .B(g8070), .Z(g11618) ) ;
INV     gate5462  (.A(g11618), .Z(g14226) ) ;
NOR2    gate5463  (.A(g9880), .B(g9883), .Z(g12246) ) ;
INV     gate5464  (.A(g12246), .Z(g14231) ) ;
AND2    gate5465  (.A(g8836), .B(g802), .Z(g11083) ) ;
INV     gate5466  (.A(g11083), .Z(g14232) ) ;
NOR2    gate5467  (.A(g8172), .B(g8125), .Z(g11666) ) ;
INV     gate5468  (.A(g11666), .Z(g14237) ) ;
INV     gate5469  (.A(g10823), .Z(g14238) ) ;
NOR2    gate5470  (.A(g9951), .B(g9954), .Z(g12308) ) ;
INV     gate5471  (.A(g12308), .Z(g14251) ) ;
INV     gate5472  (.A(g11165), .Z(II16438) ) ;
INV     gate5473  (.A(II16438), .Z(g14252) ) ;
INV     gate5474  (.A(g12381), .Z(g14255) ) ;
AND3    gate5475  (.A(g7738), .B(g5527), .C(g5535), .Z(g10838) ) ;
INV     gate5476  (.A(g10838), .Z(g14262) ) ;
NOR2    gate5477  (.A(g10019), .B(g10022), .Z(g12358) ) ;
INV     gate5478  (.A(g12358), .Z(g14275) ) ;
INV     gate5479  (.A(g11182), .Z(II16452) ) ;
INV     gate5480  (.A(II16452), .Z(g14276) ) ;
INV     gate5481  (.A(g11845), .Z(II16455) ) ;
INV     gate5482  (.A(II16455), .Z(g14277) ) ;
INV     gate5483  (.A(g10430), .Z(II16460) ) ;
INV     gate5484  (.A(II16460), .Z(g14290) ) ;
AND3    gate5485  (.A(g7766), .B(g5873), .C(g5881), .Z(g10869) ) ;
INV     gate5486  (.A(g10869), .Z(g14297) ) ;
INV     gate5487  (.A(g12760), .Z(II16468) ) ;
INV     gate5488  (.A(II16468), .Z(g14307) ) ;
INV     gate5489  (.A(g12367), .Z(II16471) ) ;
INV     gate5490  (.A(II16471), .Z(g14308) ) ;
INV     gate5491  (.A(g10430), .Z(II16476) ) ;
INV     gate5492  (.A(II16476), .Z(g14314) ) ;
INV     gate5493  (.A(g10430), .Z(II16479) ) ;
INV     gate5494  (.A(II16479), .Z(g14315) ) ;
AND3    gate5495  (.A(g7791), .B(g6219), .C(g6227), .Z(g10874) ) ;
INV     gate5496  (.A(g10874), .Z(g14321) ) ;
INV     gate5497  (.A(g11204), .Z(II16486) ) ;
INV     gate5498  (.A(II16486), .Z(g14330) ) ;
INV     gate5499  (.A(g12793), .Z(II16489) ) ;
INV     gate5500  (.A(II16489), .Z(g14331) ) ;
INV     gate5501  (.A(g12430), .Z(II16492) ) ;
INV     gate5502  (.A(II16492), .Z(g14332) ) ;
INV     gate5503  (.A(g10430), .Z(II16498) ) ;
INV     gate5504  (.A(II16498), .Z(g14336) ) ;
INV     gate5505  (.A(g10430), .Z(II16502) ) ;
INV     gate5506  (.A(II16502), .Z(g14338) ) ;
NOR2    gate5507  (.A(g5073), .B(g9989), .Z(g12163) ) ;
INV     gate5508  (.A(g12163), .Z(g14342) ) ;
AND3    gate5509  (.A(g7812), .B(g6565), .C(g6573), .Z(g10887) ) ;
INV     gate5510  (.A(g10887), .Z(g14348) ) ;
INV     gate5511  (.A(g12181), .Z(g14357) ) ;
INV     gate5512  (.A(g12811), .Z(II16512) ) ;
INV     gate5513  (.A(II16512), .Z(g14358) ) ;
INV     gate5514  (.A(g12477), .Z(II16515) ) ;
INV     gate5515  (.A(II16515), .Z(g14359) ) ;
INV     gate5516  (.A(g10430), .Z(II16521) ) ;
INV     gate5517  (.A(II16521), .Z(g14363) ) ;
INV     gate5518  (.A(g10430), .Z(II16526) ) ;
INV     gate5519  (.A(II16526), .Z(g14366) ) ;
NOR2    gate5520  (.A(g9989), .B(g5069), .Z(g12126) ) ;
INV     gate5521  (.A(g12126), .Z(g14376) ) ;
NOR2    gate5522  (.A(g5417), .B(g10047), .Z(g12201) ) ;
INV     gate5523  (.A(g12201), .Z(g14377) ) ;
INV     gate5524  (.A(g11235), .Z(II16535) ) ;
INV     gate5525  (.A(II16535), .Z(g14383) ) ;
INV     gate5526  (.A(g10417), .Z(II16538) ) ;
INV     gate5527  (.A(II16538), .Z(g14384) ) ;
INV     gate5528  (.A(g11929), .Z(II16541) ) ;
INV     gate5529  (.A(II16541), .Z(g14385) ) ;
INV     gate5530  (.A(g11931), .Z(II16544) ) ;
INV     gate5531  (.A(II16544), .Z(g14386) ) ;
INV     gate5532  (.A(g10430), .Z(II16555) ) ;
INV     gate5533  (.A(II16555), .Z(g14398) ) ;
NOR2    gate5534  (.A(g10047), .B(g5413), .Z(g12170) ) ;
INV     gate5535  (.A(g12170), .Z(g14405) ) ;
NOR2    gate5536  (.A(g5763), .B(g10096), .Z(g12249) ) ;
INV     gate5537  (.A(g12249), .Z(g14406) ) ;
INV     gate5538  (.A(g10429), .Z(II16564) ) ;
INV     gate5539  (.A(II16564), .Z(g14412) ) ;
INV     gate5540  (.A(g3298), .Z(II16575) ) ;
INV     gate5541  (.A(g10981), .Z(II16579) ) ;
INV     gate5542  (.A(II16579), .Z(g14423) ) ;
INV     gate5543  (.A(g11136), .Z(g14424) ) ;
NOR2    gate5544  (.A(g10096), .B(g5759), .Z(g12208) ) ;
INV     gate5545  (.A(g12208), .Z(g14431) ) ;
NOR2    gate5546  (.A(g6109), .B(g10136), .Z(g12311) ) ;
INV     gate5547  (.A(g12311), .Z(g14432) ) ;
INV     gate5548  (.A(g11966), .Z(II16590) ) ;
INV     gate5549  (.A(II16590), .Z(g14441) ) ;
INV     gate5550  (.A(g10498), .Z(II16593) ) ;
INV     gate5551  (.A(II16593), .Z(g14442) ) ;
INV     gate5552  (.A(g12640), .Z(II16596) ) ;
INV     gate5553  (.A(II16596), .Z(g14443) ) ;
INV     gate5554  (.A(g3649), .Z(II16606) ) ;
INV     gate5555  (.A(g10981), .Z(II16610) ) ;
INV     gate5556  (.A(II16610), .Z(g14453) ) ;
INV     gate5557  (.A(g10430), .Z(II16613) ) ;
INV     gate5558  (.A(II16613), .Z(g14454) ) ;
NOR2    gate5559  (.A(g10136), .B(g6105), .Z(g12256) ) ;
INV     gate5560  (.A(g12256), .Z(g14503) ) ;
NOR2    gate5561  (.A(g6455), .B(g10172), .Z(g12361) ) ;
INV     gate5562  (.A(g12361), .Z(g14504) ) ;
INV     gate5563  (.A(g11986), .Z(II16626) ) ;
INV     gate5564  (.A(II16626), .Z(g14509) ) ;
INV     gate5565  (.A(g11987), .Z(II16629) ) ;
INV     gate5566  (.A(II16629), .Z(g14510) ) ;
INV     gate5567  (.A(g4000), .Z(II16639) ) ;
NOR2    gate5568  (.A(g10172), .B(g6451), .Z(g12318) ) ;
INV     gate5569  (.A(g12318), .Z(g14535) ) ;
INV     gate5570  (.A(g10542), .Z(II16651) ) ;
INV     gate5571  (.A(II16651), .Z(g14536) ) ;
NAND4   gate5572  (.A(g2741), .B(g2735), .C(g6856), .D(g2748), .Z(g11405) ) ;
INV     gate5573  (.A(g11405), .Z(g14541) ) ;
INV     gate5574  (.A(g10981), .Z(II16660) ) ;
INV     gate5575  (.A(II16660), .Z(g14543) ) ;
INV     gate5576  (.A(g10981), .Z(II16663) ) ;
INV     gate5577  (.A(II16663), .Z(g14544) ) ;
OR2     gate5578  (.A(g7785), .B(g7202), .Z(g12768) ) ;
INV     gate5579  (.A(g12768), .Z(g14545) ) ;
INV     gate5580  (.A(g12036), .Z(g14562) ) ;
AND2    gate5581  (.A(g7004), .B(g5297), .Z(g10588) ) ;
INV     gate5582  (.A(g10588), .Z(II16676) ) ;
INV     gate5583  (.A(II16676), .Z(g14563) ) ;
INV     gate5584  (.A(g12039), .Z(II16679) ) ;
INV     gate5585  (.A(II16679), .Z(g14564) ) ;
INV     gate5586  (.A(g10981), .Z(II16688) ) ;
INV     gate5587  (.A(II16688), .Z(g14571) ) ;
INV     gate5588  (.A(g12077), .Z(II16698) ) ;
INV     gate5589  (.A(II16698), .Z(g14582) ) ;
INV     gate5590  (.A(g11048), .Z(g14584) ) ;
INV     gate5591  (.A(g10430), .Z(II16709) ) ;
INV     gate5592  (.A(II16709), .Z(g14591) ) ;
INV     gate5593  (.A(g5331), .Z(II16713) ) ;
INV     gate5594  (.A(g12108), .Z(II16724) ) ;
INV     gate5595  (.A(II16724), .Z(g14609) ) ;
NOR2    gate5596  (.A(g9417), .B(g9340), .Z(g12026) ) ;
INV     gate5597  (.A(g12026), .Z(II16733) ) ;
INV     gate5598  (.A(II16733), .Z(g14616) ) ;
NAND2   gate5599  (.A(g7704), .B(g10266), .Z(g12402) ) ;
INV     gate5600  (.A(g12402), .Z(g14630) ) ;
NAND2   gate5601  (.A(II15106), .B(II15107), .Z(g12239) ) ;
INV     gate5602  (.A(g12239), .Z(g14631) ) ;
INV     gate5603  (.A(g5677), .Z(II16741) ) ;
NOR2    gate5604  (.A(g1657), .B(g8139), .Z(g12729) ) ;
INV     gate5605  (.A(g12729), .Z(II16747) ) ;
INV     gate5606  (.A(II16747), .Z(g14639) ) ;
NOR3    gate5607  (.A(g6856), .B(g2748), .C(g9708), .Z(g12377) ) ;
INV     gate5608  (.A(g12377), .Z(II16755) ) ;
INV     gate5609  (.A(II16755), .Z(g14645) ) ;
INV     gate5610  (.A(g5290), .Z(II16762) ) ;
NAND2   gate5611  (.A(g7738), .B(g10281), .Z(g12450) ) ;
INV     gate5612  (.A(g12450), .Z(g14668) ) ;
NAND2   gate5613  (.A(II15148), .B(II15149), .Z(g12301) ) ;
INV     gate5614  (.A(g12301), .Z(g14669) ) ;
INV     gate5615  (.A(g6023), .Z(II16770) ) ;
INV     gate5616  (.A(g12183), .Z(II16775) ) ;
INV     gate5617  (.A(II16775), .Z(g14676) ) ;
INV     gate5618  (.A(g5637), .Z(II16795) ) ;
NAND2   gate5619  (.A(g7766), .B(g10312), .Z(g12512) ) ;
INV     gate5620  (.A(g12512), .Z(g14700) ) ;
NAND2   gate5621  (.A(II15194), .B(II15195), .Z(g12351) ) ;
INV     gate5622  (.A(g12351), .Z(g14701) ) ;
INV     gate5623  (.A(g6369), .Z(II16803) ) ;
INV     gate5624  (.A(g11405), .Z(g14714) ) ;
INV     gate5625  (.A(g5983), .Z(II16821) ) ;
NAND2   gate5626  (.A(g7791), .B(g10341), .Z(g12578) ) ;
INV     gate5627  (.A(g12578), .Z(g14744) ) ;
NAND2   gate5628  (.A(II15242), .B(II15243), .Z(g12423) ) ;
INV     gate5629  (.A(g12423), .Z(g14745) ) ;
INV     gate5630  (.A(g6715), .Z(II16829) ) ;
INV     gate5631  (.A(g11317), .Z(g14753) ) ;
INV     gate5632  (.A(g6329), .Z(II16847) ) ;
NAND2   gate5633  (.A(g7812), .B(g7142), .Z(g12629) ) ;
INV     gate5634  (.A(g12629), .Z(g14785) ) ;
NAND2   gate5635  (.A(II15288), .B(II15289), .Z(g12471) ) ;
INV     gate5636  (.A(g12471), .Z(g14786) ) ;
INV     gate5637  (.A(g10473), .Z(II16855) ) ;
INV     gate5638  (.A(II16855), .Z(g14790) ) ;
INV     gate5639  (.A(g6675), .Z(II16875) ) ;
INV     gate5640  (.A(g11405), .Z(g14833) ) ;
NOR2    gate5641  (.A(g1636), .B(g7308), .Z(g10615) ) ;
INV     gate5642  (.A(g10615), .Z(II16898) ) ;
INV     gate5643  (.A(II16898), .Z(g14873) ) ;
INV     gate5644  (.A(g10582), .Z(II16917) ) ;
INV     gate5645  (.A(II16917), .Z(g14912) ) ;
INV     gate5646  (.A(g13943), .Z(II16969) ) ;
INV     gate5647  (.A(g12857), .Z(II17008) ) ;
INV     gate5648  (.A(II17008), .Z(g15085) ) ;
INV     gate5649  (.A(g14331), .Z(II17094) ) ;
INV     gate5650  (.A(II17094), .Z(g15169) ) ;
INV     gate5651  (.A(g14336), .Z(II17098) ) ;
INV     gate5652  (.A(II17098), .Z(g15171) ) ;
INV     gate5653  (.A(g14338), .Z(II17101) ) ;
INV     gate5654  (.A(II17101), .Z(g15224) ) ;
INV     gate5655  (.A(g12932), .Z(II17104) ) ;
INV     gate5656  (.A(II17104), .Z(g15277) ) ;
NAND2   gate5657  (.A(g7738), .B(g12505), .Z(g14851) ) ;
INV     gate5658  (.A(g14851), .Z(g15344) ) ;
INV     gate5659  (.A(g13782), .Z(II17108) ) ;
INV     gate5660  (.A(II17108), .Z(g15345) ) ;
INV     gate5661  (.A(g13809), .Z(II17111) ) ;
INV     gate5662  (.A(II17111), .Z(g15348) ) ;
INV     gate5663  (.A(g14358), .Z(II17114) ) ;
INV     gate5664  (.A(II17114), .Z(g15371) ) ;
INV     gate5665  (.A(g14363), .Z(II17118) ) ;
INV     gate5666  (.A(II17118), .Z(g15373) ) ;
INV     gate5667  (.A(g14366), .Z(II17121) ) ;
INV     gate5668  (.A(II17121), .Z(g15426) ) ;
NAND2   gate5669  (.A(g7766), .B(g12571), .Z(g14895) ) ;
INV     gate5670  (.A(g14895), .Z(g15479) ) ;
INV     gate5671  (.A(g13809), .Z(II17125) ) ;
INV     gate5672  (.A(II17125), .Z(g15480) ) ;
INV     gate5673  (.A(g13835), .Z(II17128) ) ;
INV     gate5674  (.A(II17128), .Z(g15483) ) ;
INV     gate5675  (.A(g14384), .Z(II17131) ) ;
INV     gate5676  (.A(II17131), .Z(g15506) ) ;
INV     gate5677  (.A(g14398), .Z(II17136) ) ;
INV     gate5678  (.A(II17136), .Z(g15509) ) ;
NAND2   gate5679  (.A(g7791), .B(g12622), .Z(g14943) ) ;
INV     gate5680  (.A(g14943), .Z(g15562) ) ;
INV     gate5681  (.A(g13835), .Z(II17140) ) ;
INV     gate5682  (.A(II17140), .Z(g15563) ) ;
INV     gate5683  (.A(g14412), .Z(II17143) ) ;
INV     gate5684  (.A(II17143), .Z(g15566) ) ;
NAND2   gate5685  (.A(g7812), .B(g12680), .Z(g14984) ) ;
INV     gate5686  (.A(g14984), .Z(g15568) ) ;
INV     gate5687  (.A(g14442), .Z(II17148) ) ;
INV     gate5688  (.A(II17148), .Z(g15569) ) ;
OR2     gate5689  (.A(g11294), .B(g7567), .Z(g13211) ) ;
INV     gate5690  (.A(g13211), .Z(g15571) ) ;
INV     gate5691  (.A(g13605), .Z(II17154) ) ;
INV     gate5692  (.A(II17154), .Z(g15573) ) ;
INV     gate5693  (.A(g13350), .Z(II17159) ) ;
INV     gate5694  (.A(II17159), .Z(g15579) ) ;
OR2     gate5695  (.A(g11336), .B(g7601), .Z(g13242) ) ;
INV     gate5696  (.A(g13242), .Z(g15580) ) ;
INV     gate5697  (.A(g14536), .Z(II17166) ) ;
INV     gate5698  (.A(II17166), .Z(g15588) ) ;
INV     gate5699  (.A(g13716), .Z(II17173) ) ;
INV     gate5700  (.A(II17173), .Z(g15595) ) ;
NOR2    gate5701  (.A(g12822), .B(g12797), .Z(g14914) ) ;
INV     gate5702  (.A(g14914), .Z(g15614) ) ;
INV     gate5703  (.A(g13745), .Z(II17181) ) ;
INV     gate5704  (.A(II17181), .Z(g15615) ) ;
INV     gate5705  (.A(g13782), .Z(II17188) ) ;
INV     gate5706  (.A(II17188), .Z(g15634) ) ;
NOR2    gate5707  (.A(g8347), .B(g10511), .Z(g13202) ) ;
INV     gate5708  (.A(g13202), .Z(g15655) ) ;
INV     gate5709  (.A(g13809), .Z(II17198) ) ;
INV     gate5710  (.A(II17198), .Z(g15656) ) ;
INV     gate5711  (.A(g13835), .Z(II17207) ) ;
INV     gate5712  (.A(II17207), .Z(g15680) ) ;
NAND2   gate5713  (.A(g4082), .B(g10808), .Z(g13217) ) ;
INV     gate5714  (.A(g13217), .Z(g15705) ) ;
INV     gate5715  (.A(g13350), .Z(II17228) ) ;
INV     gate5716  (.A(II17228), .Z(g15714) ) ;
NOR2    gate5717  (.A(g10929), .B(g10905), .Z(g13326) ) ;
INV     gate5718  (.A(g13326), .Z(g15731) ) ;
INV     gate5719  (.A(g13605), .Z(II17249) ) ;
INV     gate5720  (.A(II17249), .Z(g15733) ) ;
NAND2   gate5721  (.A(g10695), .B(g1157), .Z(g13284) ) ;
INV     gate5722  (.A(g13284), .Z(g15739) ) ;
NOR2    gate5723  (.A(g10961), .B(g10935), .Z(g13342) ) ;
INV     gate5724  (.A(g13342), .Z(g15740) ) ;
NAND2   gate5725  (.A(g11117), .B(g8411), .Z(g13121) ) ;
INV     gate5726  (.A(g13121), .Z(g15746) ) ;
NAND2   gate5727  (.A(g1116), .B(g10695), .Z(g13307) ) ;
INV     gate5728  (.A(g13307), .Z(g15747) ) ;
NAND2   gate5729  (.A(g10715), .B(g1500), .Z(g13291) ) ;
INV     gate5730  (.A(g13291), .Z(g15750) ) ;
NAND2   gate5731  (.A(g11134), .B(g8470), .Z(g13134) ) ;
INV     gate5732  (.A(g13134), .Z(g15755) ) ;
NAND2   gate5733  (.A(g1459), .B(g10715), .Z(g13315) ) ;
INV     gate5734  (.A(g13315), .Z(g15756) ) ;
INV     gate5735  (.A(g13605), .Z(II17276) ) ;
INV     gate5736  (.A(II17276), .Z(g15758) ) ;
NOR2    gate5737  (.A(g7841), .B(g10741), .Z(g13110) ) ;
INV     gate5738  (.A(g13110), .Z(g15799) ) ;
OR2     gate5739  (.A(g10776), .B(g8703), .Z(g14044) ) ;
INV     gate5740  (.A(g14044), .Z(II17302) ) ;
INV     gate5741  (.A(II17302), .Z(g15806) ) ;
NOR2    gate5742  (.A(g7863), .B(g10762), .Z(g13125) ) ;
INV     gate5743  (.A(g13125), .Z(g15811) ) ;
OR2     gate5744  (.A(g10776), .B(g8703), .Z(g14078) ) ;
INV     gate5745  (.A(g14078), .Z(II17314) ) ;
INV     gate5746  (.A(II17314), .Z(g15816) ) ;
OR2     gate5747  (.A(g10776), .B(g8703), .Z(g14119) ) ;
INV     gate5748  (.A(g14119), .Z(II17324) ) ;
INV     gate5749  (.A(II17324), .Z(g15824) ) ;
NAND2   gate5750  (.A(g4793), .B(g10831), .Z(g13432) ) ;
INV     gate5751  (.A(g13432), .Z(g15830) ) ;
OR2     gate5752  (.A(g11967), .B(g9479), .Z(g13385) ) ;
INV     gate5753  (.A(g13385), .Z(g15831) ) ;
NAND2   gate5754  (.A(g4983), .B(g10862), .Z(g13469) ) ;
INV     gate5755  (.A(g13469), .Z(g15842) ) ;
INV     gate5756  (.A(g14591), .Z(II17355) ) ;
INV     gate5757  (.A(II17355), .Z(g15862) ) ;
INV     gate5758  (.A(g13638), .Z(II17374) ) ;
INV     gate5759  (.A(II17374), .Z(g15885) ) ;
INV     gate5760  (.A(g13680), .Z(II17392) ) ;
INV     gate5761  (.A(II17392), .Z(g15915) ) ;
INV     gate5762  (.A(g12952), .Z(II17395) ) ;
INV     gate5763  (.A(II17395), .Z(g15932) ) ;
INV     gate5764  (.A(g13394), .Z(II17401) ) ;
INV     gate5765  (.A(II17401), .Z(g15938) ) ;
NOR2    gate5766  (.A(g11245), .B(g4076), .Z(g13806) ) ;
INV     gate5767  (.A(g13806), .Z(II17416) ) ;
INV     gate5768  (.A(II17416), .Z(g15969) ) ;
INV     gate5769  (.A(g13394), .Z(II17420) ) ;
INV     gate5770  (.A(II17420), .Z(g15979) ) ;
INV     gate5771  (.A(g13416), .Z(II17425) ) ;
INV     gate5772  (.A(II17425), .Z(g16000) ) ;
OR2     gate5773  (.A(g9223), .B(g11130), .Z(g13570) ) ;
INV     gate5774  (.A(g13570), .Z(g16030) ) ;
INV     gate5775  (.A(g13416), .Z(II17436) ) ;
INV     gate5776  (.A(II17436), .Z(g16031) ) ;
INV     gate5777  (.A(g13638), .Z(II17442) ) ;
INV     gate5778  (.A(II17442), .Z(g16053) ) ;
OR2     gate5779  (.A(g9247), .B(g11149), .Z(g13597) ) ;
INV     gate5780  (.A(g13597), .Z(g16075) ) ;
INV     gate5781  (.A(g13680), .Z(II17456) ) ;
INV     gate5782  (.A(II17456), .Z(g16077) ) ;
INV     gate5783  (.A(g13530), .Z(g16096) ) ;
INV     gate5784  (.A(g13437), .Z(g16099) ) ;
INV     gate5785  (.A(g13394), .Z(II17471) ) ;
INV     gate5786  (.A(II17471), .Z(g16100) ) ;
INV     gate5787  (.A(g13530), .Z(g16123) ) ;
INV     gate5788  (.A(g13555), .Z(g16124) ) ;
INV     gate5789  (.A(g13437), .Z(g16127) ) ;
INV     gate5790  (.A(g13394), .Z(II17488) ) ;
INV     gate5791  (.A(II17488), .Z(g16129) ) ;
INV     gate5792  (.A(g13416), .Z(II17491) ) ;
INV     gate5793  (.A(II17491), .Z(g16136) ) ;
INV     gate5794  (.A(g13555), .Z(g16158) ) ;
INV     gate5795  (.A(g13584), .Z(g16159) ) ;
INV     gate5796  (.A(g13437), .Z(g16162) ) ;
INV     gate5797  (.A(g13416), .Z(II17507) ) ;
INV     gate5798  (.A(II17507), .Z(g16164) ) ;
INV     gate5799  (.A(g13530), .Z(g16171) ) ;
INV     gate5800  (.A(g13584), .Z(g16172) ) ;
INV     gate5801  (.A(g13437), .Z(g16180) ) ;
NAND2   gate5802  (.A(g1116), .B(g10649), .Z(g13846) ) ;
INV     gate5803  (.A(g13846), .Z(g16182) ) ;
INV     gate5804  (.A(g13555), .Z(g16186) ) ;
INV     gate5805  (.A(g13437), .Z(g16195) ) ;
NAND2   gate5806  (.A(g1459), .B(g10671), .Z(g13861) ) ;
INV     gate5807  (.A(g13861), .Z(g16197) ) ;
INV     gate5808  (.A(g13584), .Z(g16200) ) ;
INV     gate5809  (.A(g13437), .Z(g16206) ) ;
INV     gate5810  (.A(g13437), .Z(g16214) ) ;
INV     gate5811  (.A(g14510), .Z(II17557) ) ;
INV     gate5812  (.A(II17557), .Z(g16216) ) ;
INV     gate5813  (.A(g13437), .Z(g16223) ) ;
INV     gate5814  (.A(g14564), .Z(II17569) ) ;
INV     gate5815  (.A(II17569), .Z(g16228) ) ;
INV     gate5816  (.A(g13437), .Z(g16235) ) ;
INV     gate5817  (.A(g14591), .Z(II17590) ) ;
INV     gate5818  (.A(II17590), .Z(g16249) ) ;
NAND2   gate5819  (.A(g4664), .B(g11006), .Z(g13330) ) ;
INV     gate5820  (.A(g13330), .Z(g16280) ) ;
INV     gate5821  (.A(g13510), .Z(II17609) ) ;
INV     gate5822  (.A(II17609), .Z(g16284) ) ;
INV     gate5823  (.A(g13250), .Z(II17612) ) ;
INV     gate5824  (.A(II17612), .Z(g16285) ) ;
INV     gate5825  (.A(g13251), .Z(II17615) ) ;
INV     gate5826  (.A(II17615), .Z(g16286) ) ;
INV     gate5827  (.A(g13223), .Z(g16289) ) ;
NAND2   gate5828  (.A(g1116), .B(g10666), .Z(g13260) ) ;
INV     gate5829  (.A(g13260), .Z(g16290) ) ;
INV     gate5830  (.A(g14582), .Z(II17626) ) ;
INV     gate5831  (.A(II17626), .Z(g16300) ) ;
NAND2   gate5832  (.A(g4854), .B(g11012), .Z(g13346) ) ;
INV     gate5833  (.A(g13346), .Z(g16305) ) ;
INV     gate5834  (.A(g13258), .Z(II17633) ) ;
INV     gate5835  (.A(II17633), .Z(g16307) ) ;
INV     gate5836  (.A(g14252), .Z(II17636) ) ;
INV     gate5837  (.A(II17636), .Z(g16308) ) ;
INV     gate5838  (.A(g13350), .Z(II17639) ) ;
INV     gate5839  (.A(II17639), .Z(g16309) ) ;
INV     gate5840  (.A(g13223), .Z(g16310) ) ;
NAND2   gate5841  (.A(g1459), .B(g10699), .Z(g13273) ) ;
INV     gate5842  (.A(g13273), .Z(g16311) ) ;
INV     gate5843  (.A(g14454), .Z(g16320) ) ;
INV     gate5844  (.A(g13271), .Z(II17650) ) ;
INV     gate5845  (.A(II17650), .Z(g16322) ) ;
INV     gate5846  (.A(g14276), .Z(II17653) ) ;
INV     gate5847  (.A(II17653), .Z(g16323) ) ;
INV     gate5848  (.A(g13223), .Z(g16325) ) ;
INV     gate5849  (.A(g13394), .Z(II17658) ) ;
INV     gate5850  (.A(II17658), .Z(g16326) ) ;
INV     gate5851  (.A(g13329), .Z(II17661) ) ;
INV     gate5852  (.A(II17661), .Z(g16349) ) ;
NAND2   gate5853  (.A(g11514), .B(g11473), .Z(g14066) ) ;
INV     gate5854  (.A(g14066), .Z(g16423) ) ;
INV     gate5855  (.A(g13279), .Z(II17668) ) ;
INV     gate5856  (.A(II17668), .Z(g16428) ) ;
INV     gate5857  (.A(g13280), .Z(II17671) ) ;
INV     gate5858  (.A(II17671), .Z(g16429) ) ;
INV     gate5859  (.A(g13394), .Z(II17675) ) ;
INV     gate5860  (.A(II17675), .Z(g16431) ) ;
INV     gate5861  (.A(g13416), .Z(II17679) ) ;
INV     gate5862  (.A(II17679), .Z(g16449) ) ;
NAND2   gate5863  (.A(g11566), .B(g8864), .Z(g14098) ) ;
INV     gate5864  (.A(g14098), .Z(g16472) ) ;
NAND2   gate5865  (.A(g11610), .B(g11729), .Z(g13977) ) ;
INV     gate5866  (.A(g13977), .Z(g16473) ) ;
NAND2   gate5867  (.A(g11571), .B(g11527), .Z(g14107) ) ;
INV     gate5868  (.A(g14107), .Z(g16475) ) ;
NAND3   gate5869  (.A(g10831), .B(g4793), .C(g4776), .Z(g13464) ) ;
INV     gate5870  (.A(g13464), .Z(g16482) ) ;
INV     gate5871  (.A(g14330), .Z(II17695) ) ;
INV     gate5872  (.A(II17695), .Z(g16487) ) ;
INV     gate5873  (.A(g13416), .Z(II17699) ) ;
INV     gate5874  (.A(II17699), .Z(g16489) ) ;
INV     gate5875  (.A(g13144), .Z(II17704) ) ;
INV     gate5876  (.A(II17704), .Z(g16508) ) ;
NAND2   gate5877  (.A(g11566), .B(g11729), .Z(g13873) ) ;
INV     gate5878  (.A(g13873), .Z(g16509) ) ;
NAND2   gate5879  (.A(g11610), .B(g11435), .Z(g14008) ) ;
INV     gate5880  (.A(g14008), .Z(g16510) ) ;
NAND2   gate5881  (.A(g11621), .B(g8906), .Z(g14130) ) ;
INV     gate5882  (.A(g14130), .Z(g16511) ) ;
NAND2   gate5883  (.A(g11658), .B(g11747), .Z(g14015) ) ;
INV     gate5884  (.A(g14015), .Z(g16512) ) ;
NAND2   gate5885  (.A(g11626), .B(g11584), .Z(g14139) ) ;
INV     gate5886  (.A(g14139), .Z(g16514) ) ;
NAND3   gate5887  (.A(g10862), .B(g4983), .C(g4966), .Z(g13486) ) ;
INV     gate5888  (.A(g13486), .Z(g16515) ) ;
OR2     gate5889  (.A(g10543), .B(g10565), .Z(g13543) ) ;
INV     gate5890  (.A(g13543), .Z(g16521) ) ;
NAND2   gate5891  (.A(g11566), .B(g11435), .Z(g13889) ) ;
INV     gate5892  (.A(g13889), .Z(g16522) ) ;
NAND2   gate5893  (.A(g11610), .B(g11473), .Z(g14041) ) ;
INV     gate5894  (.A(g14041), .Z(g16523) ) ;
INV     gate5895  (.A(g13177), .Z(II17723) ) ;
INV     gate5896  (.A(II17723), .Z(g16525) ) ;
NAND2   gate5897  (.A(g11621), .B(g11747), .Z(g13898) ) ;
INV     gate5898  (.A(g13898), .Z(g16526) ) ;
NAND2   gate5899  (.A(g11658), .B(g11483), .Z(g14048) ) ;
INV     gate5900  (.A(g14048), .Z(g16527) ) ;
NAND2   gate5901  (.A(g11669), .B(g8958), .Z(g14154) ) ;
INV     gate5902  (.A(g14154), .Z(g16528) ) ;
NAND2   gate5903  (.A(g11697), .B(g11763), .Z(g14055) ) ;
INV     gate5904  (.A(g14055), .Z(g16529) ) ;
INV     gate5905  (.A(g14454), .Z(g16530) ) ;
OR2     gate5906  (.A(g10776), .B(g8703), .Z(g14844) ) ;
INV     gate5907  (.A(g14844), .Z(II17733) ) ;
INV     gate5908  (.A(II17733), .Z(g16533) ) ;
INV     gate5909  (.A(g14912), .Z(II17744) ) ;
INV     gate5910  (.A(II17744), .Z(g16540) ) ;
INV     gate5911  (.A(g13298), .Z(II17747) ) ;
INV     gate5912  (.A(II17747), .Z(g16577) ) ;
INV     gate5913  (.A(g14383), .Z(II17750) ) ;
INV     gate5914  (.A(II17750), .Z(g16578) ) ;
INV     gate5915  (.A(g13267), .Z(g16579) ) ;
INV     gate5916  (.A(g13494), .Z(II17754) ) ;
INV     gate5917  (.A(II17754), .Z(g16580) ) ;
NAND2   gate5918  (.A(g11566), .B(g11473), .Z(g13915) ) ;
INV     gate5919  (.A(g13915), .Z(g16582) ) ;
NAND2   gate5920  (.A(g11653), .B(g8864), .Z(g14069) ) ;
INV     gate5921  (.A(g14069), .Z(g16583) ) ;
NAND2   gate5922  (.A(g11621), .B(g11483), .Z(g13920) ) ;
INV     gate5923  (.A(g13920), .Z(g16584) ) ;
NAND2   gate5924  (.A(g11658), .B(g11527), .Z(g14075) ) ;
INV     gate5925  (.A(g14075), .Z(g16585) ) ;
INV     gate5926  (.A(g13191), .Z(II17763) ) ;
INV     gate5927  (.A(II17763), .Z(g16587) ) ;
NAND2   gate5928  (.A(g11669), .B(g11763), .Z(g13929) ) ;
INV     gate5929  (.A(g13929), .Z(g16588) ) ;
NAND2   gate5930  (.A(g11697), .B(g11537), .Z(g14082) ) ;
INV     gate5931  (.A(g14082), .Z(g16589) ) ;
OR2     gate5932  (.A(g10776), .B(g8703), .Z(g14888) ) ;
INV     gate5933  (.A(g14888), .Z(II17772) ) ;
INV     gate5934  (.A(II17772), .Z(g16594) ) ;
INV     gate5935  (.A(g13303), .Z(II17780) ) ;
INV     gate5936  (.A(II17780), .Z(g16600) ) ;
INV     gate5937  (.A(g13304), .Z(II17783) ) ;
INV     gate5938  (.A(II17783), .Z(g16601) ) ;
NAND2   gate5939  (.A(g11653), .B(g11729), .Z(g14101) ) ;
INV     gate5940  (.A(g14101), .Z(g16602) ) ;
INV     gate5941  (.A(g3267), .Z(II17787) ) ;
NAND2   gate5942  (.A(g11621), .B(g11527), .Z(g13955) ) ;
INV     gate5943  (.A(g13955), .Z(g16605) ) ;
NAND2   gate5944  (.A(g11692), .B(g8906), .Z(g14110) ) ;
INV     gate5945  (.A(g14110), .Z(g16606) ) ;
NAND2   gate5946  (.A(g11669), .B(g11537), .Z(g13960) ) ;
INV     gate5947  (.A(g13960), .Z(g16607) ) ;
NAND2   gate5948  (.A(g11697), .B(g11584), .Z(g14116) ) ;
INV     gate5949  (.A(g14116), .Z(g16608) ) ;
INV     gate5950  (.A(g14454), .Z(g16609) ) ;
OR2     gate5951  (.A(g10776), .B(g8703), .Z(g14936) ) ;
INV     gate5952  (.A(g14936), .Z(II17801) ) ;
INV     gate5953  (.A(II17801), .Z(g16615) ) ;
INV     gate5954  (.A(g13311), .Z(II17808) ) ;
INV     gate5955  (.A(II17808), .Z(g16620) ) ;
NAND2   gate5956  (.A(g11514), .B(g8864), .Z(g14104) ) ;
INV     gate5957  (.A(g14104), .Z(g16622) ) ;
NAND2   gate5958  (.A(g11653), .B(g11435), .Z(g14127) ) ;
INV     gate5959  (.A(g14127), .Z(g16623) ) ;
INV     gate5960  (.A(g3274), .Z(II17814) ) ;
NAND2   gate5961  (.A(g11692), .B(g11747), .Z(g14133) ) ;
INV     gate5962  (.A(g14133), .Z(g16626) ) ;
INV     gate5963  (.A(g3618), .Z(II17819) ) ;
NAND2   gate5964  (.A(g11669), .B(g11584), .Z(g13990) ) ;
INV     gate5965  (.A(g13990), .Z(g16629) ) ;
NAND2   gate5966  (.A(g11715), .B(g8958), .Z(g14142) ) ;
INV     gate5967  (.A(g14142), .Z(g16630) ) ;
INV     gate5968  (.A(g14454), .Z(g16631) ) ;
INV     gate5969  (.A(g14454), .Z(g16632) ) ;
OR2     gate5970  (.A(g10776), .B(g8703), .Z(g14977) ) ;
INV     gate5971  (.A(g14977), .Z(II17834) ) ;
INV     gate5972  (.A(II17834), .Z(g16640) ) ;
INV     gate5973  (.A(g13412), .Z(II17839) ) ;
INV     gate5974  (.A(II17839), .Z(g16643) ) ;
INV     gate5975  (.A(g13051), .Z(II17842) ) ;
INV     gate5976  (.A(II17842), .Z(g16644) ) ;
NAND2   gate5977  (.A(g203), .B(g12812), .Z(g13756) ) ;
INV     gate5978  (.A(g13756), .Z(g16645) ) ;
NAND2   gate5979  (.A(g11514), .B(g11729), .Z(g14005) ) ;
INV     gate5980  (.A(g14005), .Z(g16651) ) ;
NAND2   gate5981  (.A(g11653), .B(g11473), .Z(g13892) ) ;
INV     gate5982  (.A(g13892), .Z(g16652) ) ;
NAND2   gate5983  (.A(g11571), .B(g8906), .Z(g14136) ) ;
INV     gate5984  (.A(g14136), .Z(g16654) ) ;
NAND2   gate5985  (.A(g11692), .B(g11483), .Z(g14151) ) ;
INV     gate5986  (.A(g14151), .Z(g16655) ) ;
INV     gate5987  (.A(g3625), .Z(II17852) ) ;
NAND2   gate5988  (.A(g11715), .B(g11763), .Z(g14157) ) ;
INV     gate5989  (.A(g14157), .Z(g16658) ) ;
INV     gate5990  (.A(g3969), .Z(II17857) ) ;
INV     gate5991  (.A(g14454), .Z(g16661) ) ;
OR2     gate5992  (.A(g10776), .B(g8703), .Z(g15017) ) ;
INV     gate5993  (.A(g15017), .Z(II17873) ) ;
INV     gate5994  (.A(II17873), .Z(g16675) ) ;
INV     gate5995  (.A(g13070), .Z(II17876) ) ;
INV     gate5996  (.A(II17876), .Z(g16676) ) ;
INV     gate5997  (.A(g14386), .Z(II17879) ) ;
INV     gate5998  (.A(II17879), .Z(g16677) ) ;
INV     gate5999  (.A(g13223), .Z(g16680) ) ;
NAND2   gate6000  (.A(g9092), .B(g11858), .Z(g14223) ) ;
INV     gate6001  (.A(g14223), .Z(g16684) ) ;
NAND2   gate6002  (.A(g11514), .B(g11435), .Z(g14038) ) ;
INV     gate6003  (.A(g14038), .Z(g16685) ) ;
INV     gate6004  (.A(g3325), .Z(II17892) ) ;
NAND2   gate6005  (.A(g11571), .B(g11747), .Z(g14045) ) ;
INV     gate6006  (.A(g14045), .Z(g16688) ) ;
NAND2   gate6007  (.A(g11692), .B(g11527), .Z(g13923) ) ;
INV     gate6008  (.A(g13923), .Z(g16689) ) ;
NAND2   gate6009  (.A(g11626), .B(g8958), .Z(g14160) ) ;
INV     gate6010  (.A(g14160), .Z(g16691) ) ;
NAND2   gate6011  (.A(g11715), .B(g11537), .Z(g14170) ) ;
INV     gate6012  (.A(g14170), .Z(g16692) ) ;
INV     gate6013  (.A(g3976), .Z(II17901) ) ;
INV     gate6014  (.A(g14454), .Z(g16695) ) ;
INV     gate6015  (.A(g13087), .Z(II17916) ) ;
INV     gate6016  (.A(II17916), .Z(g16708) ) ;
INV     gate6017  (.A(g14609), .Z(II17919) ) ;
INV     gate6018  (.A(II17919), .Z(g16709) ) ;
INV     gate6019  (.A(g13223), .Z(g16712) ) ;
NAND2   gate6020  (.A(g11610), .B(g8864), .Z(g13948) ) ;
INV     gate6021  (.A(g13948), .Z(g16716) ) ;
NAND2   gate6022  (.A(g10295), .B(g11729), .Z(g13951) ) ;
INV     gate6023  (.A(g13951), .Z(g16717) ) ;
INV     gate6024  (.A(g3310), .Z(II17932) ) ;
NAND2   gate6025  (.A(g9177), .B(g11881), .Z(g14234) ) ;
INV     gate6026  (.A(g14234), .Z(g16720) ) ;
NAND2   gate6027  (.A(g11571), .B(g11483), .Z(g14072) ) ;
INV     gate6028  (.A(g14072), .Z(g16721) ) ;
INV     gate6029  (.A(g3676), .Z(II17938) ) ;
NAND2   gate6030  (.A(g11626), .B(g11763), .Z(g14079) ) ;
INV     gate6031  (.A(g14079), .Z(g16724) ) ;
NAND2   gate6032  (.A(g11715), .B(g11584), .Z(g13963) ) ;
INV     gate6033  (.A(g13963), .Z(g16725) ) ;
INV     gate6034  (.A(g14454), .Z(g16726) ) ;
INV     gate6035  (.A(g14454), .Z(g16727) ) ;
INV     gate6036  (.A(g14562), .Z(II17956) ) ;
INV     gate6037  (.A(II17956), .Z(g16738) ) ;
INV     gate6038  (.A(g13223), .Z(g16739) ) ;
NAND2   gate6039  (.A(g10295), .B(g11435), .Z(g13980) ) ;
INV     gate6040  (.A(g13980), .Z(g16740) ) ;
NAND2   gate6041  (.A(g11658), .B(g8906), .Z(g13983) ) ;
INV     gate6042  (.A(g13983), .Z(g16742) ) ;
NAND2   gate6043  (.A(g10323), .B(g11747), .Z(g13986) ) ;
INV     gate6044  (.A(g13986), .Z(g16743) ) ;
INV     gate6045  (.A(g3661), .Z(II17964) ) ;
NAND2   gate6046  (.A(g9203), .B(g11903), .Z(g14258) ) ;
INV     gate6047  (.A(g14258), .Z(g16746) ) ;
NAND2   gate6048  (.A(g11626), .B(g11537), .Z(g14113) ) ;
INV     gate6049  (.A(g14113), .Z(g16747) ) ;
INV     gate6050  (.A(g4027), .Z(II17970) ) ;
INV     gate6051  (.A(g14454), .Z(g16750) ) ;
INV     gate6052  (.A(g13638), .Z(II17976) ) ;
INV     gate6053  (.A(II17976), .Z(g16752) ) ;
INV     gate6054  (.A(g14173), .Z(II17989) ) ;
INV     gate6055  (.A(II17989), .Z(g16767) ) ;
INV     gate6056  (.A(g13223), .Z(g16768) ) ;
INV     gate6057  (.A(g13530), .Z(g16769) ) ;
NAND2   gate6058  (.A(g10323), .B(g11483), .Z(g14018) ) ;
INV     gate6059  (.A(g14018), .Z(g16771) ) ;
NAND2   gate6060  (.A(g11697), .B(g8958), .Z(g14021) ) ;
INV     gate6061  (.A(g14021), .Z(g16773) ) ;
NAND2   gate6062  (.A(g7121), .B(g11763), .Z(g14024) ) ;
INV     gate6063  (.A(g14024), .Z(g16774) ) ;
INV     gate6064  (.A(g4012), .Z(II17999) ) ;
INV     gate6065  (.A(g13638), .Z(II18003) ) ;
INV     gate6066  (.A(II18003), .Z(g16777) ) ;
INV     gate6067  (.A(g13638), .Z(II18006) ) ;
INV     gate6068  (.A(II18006), .Z(g16782) ) ;
INV     gate6069  (.A(g13680), .Z(II18009) ) ;
INV     gate6070  (.A(II18009), .Z(g16795) ) ;
OR2     gate6071  (.A(g9086), .B(g11048), .Z(g14387) ) ;
INV     gate6072  (.A(g14387), .Z(g16809) ) ;
INV     gate6073  (.A(g13555), .Z(g16812) ) ;
NAND2   gate6074  (.A(g7121), .B(g11537), .Z(g14058) ) ;
INV     gate6075  (.A(g14058), .Z(g16814) ) ;
INV     gate6076  (.A(g13638), .Z(II18028) ) ;
INV     gate6077  (.A(II18028), .Z(g16816) ) ;
INV     gate6078  (.A(g13680), .Z(II18031) ) ;
INV     gate6079  (.A(II18031), .Z(g16821) ) ;
INV     gate6080  (.A(g13680), .Z(II18034) ) ;
INV     gate6081  (.A(II18034), .Z(g16826) ) ;
INV     gate6082  (.A(g13584), .Z(g16853) ) ;
INV     gate6083  (.A(g13638), .Z(II18048) ) ;
INV     gate6084  (.A(II18048), .Z(g16856) ) ;
INV     gate6085  (.A(g13680), .Z(II18051) ) ;
INV     gate6086  (.A(II18051), .Z(g16861) ) ;
INV     gate6087  (.A(g14198), .Z(II18060) ) ;
INV     gate6088  (.A(II18060), .Z(g16872) ) ;
INV     gate6089  (.A(g14357), .Z(II18063) ) ;
INV     gate6090  (.A(II18063), .Z(g16873) ) ;
INV     gate6091  (.A(g3317), .Z(II18066) ) ;
INV     gate6092  (.A(g13680), .Z(II18071) ) ;
INV     gate6093  (.A(II18071), .Z(g16877) ) ;
INV     gate6094  (.A(g13350), .Z(II18078) ) ;
INV     gate6095  (.A(II18078), .Z(g16886) ) ;
INV     gate6096  (.A(g13394), .Z(II18083) ) ;
INV     gate6097  (.A(II18083), .Z(g16897) ) ;
INV     gate6098  (.A(g13856), .Z(II18086) ) ;
INV     gate6099  (.A(II18086), .Z(g16920) ) ;
INV     gate6100  (.A(g13144), .Z(II18089) ) ;
INV     gate6101  (.A(II18089), .Z(g16923) ) ;
INV     gate6102  (.A(g3668), .Z(II18092) ) ;
INV     gate6103  (.A(g13416), .Z(II18101) ) ;
INV     gate6104  (.A(II18101), .Z(g16931) ) ;
INV     gate6105  (.A(g13177), .Z(II18104) ) ;
INV     gate6106  (.A(II18104), .Z(g16954) ) ;
INV     gate6107  (.A(g4019), .Z(II18107) ) ;
INV     gate6108  (.A(g14238), .Z(g16958) ) ;
INV     gate6109  (.A(g14509), .Z(II18114) ) ;
INV     gate6110  (.A(II18114), .Z(g16960) ) ;
INV     gate6111  (.A(g13302), .Z(II18117) ) ;
INV     gate6112  (.A(II18117), .Z(g16963) ) ;
INV     gate6113  (.A(g13350), .Z(II18120) ) ;
INV     gate6114  (.A(II18120), .Z(g16964) ) ;
NOR2    gate6115  (.A(g9839), .B(g12155), .Z(g14291) ) ;
INV     gate6116  (.A(g14291), .Z(g16966) ) ;
INV     gate6117  (.A(g13191), .Z(II18125) ) ;
INV     gate6118  (.A(II18125), .Z(g16967) ) ;
INV     gate6119  (.A(g14238), .Z(g16968) ) ;
INV     gate6120  (.A(g14262), .Z(g16969) ) ;
INV     gate6121  (.A(g13350), .Z(II18131) ) ;
INV     gate6122  (.A(II18131), .Z(g16971) ) ;
INV     gate6123  (.A(g13144), .Z(II18135) ) ;
INV     gate6124  (.A(II18135), .Z(g16987) ) ;
INV     gate6125  (.A(g14277), .Z(II18138) ) ;
INV     gate6126  (.A(II18138), .Z(g17010) ) ;
INV     gate6127  (.A(g14262), .Z(g17013) ) ;
INV     gate6128  (.A(g14297), .Z(g17014) ) ;
INV     gate6129  (.A(g13350), .Z(II18143) ) ;
INV     gate6130  (.A(II18143), .Z(g17015) ) ;
INV     gate6131  (.A(g13437), .Z(g17056) ) ;
OR3     gate6132  (.A(g209), .B(g10685), .C(g301), .Z(g13526) ) ;
INV     gate6133  (.A(g13526), .Z(II18148) ) ;
INV     gate6134  (.A(II18148), .Z(g17058) ) ;
INV     gate6135  (.A(g13144), .Z(II18151) ) ;
INV     gate6136  (.A(II18151), .Z(g17059) ) ;
INV     gate6137  (.A(g13177), .Z(II18154) ) ;
INV     gate6138  (.A(II18154), .Z(g17062) ) ;
INV     gate6139  (.A(g14238), .Z(g17085) ) ;
INV     gate6140  (.A(g14297), .Z(g17086) ) ;
INV     gate6141  (.A(g14321), .Z(g17087) ) ;
INV     gate6142  (.A(g14441), .Z(II18160) ) ;
INV     gate6143  (.A(II18160), .Z(g17088) ) ;
NAND2   gate6144  (.A(g10295), .B(g11473), .Z(g14011) ) ;
INV     gate6145  (.A(g14011), .Z(g17092) ) ;
INV     gate6146  (.A(g13177), .Z(II18165) ) ;
INV     gate6147  (.A(II18165), .Z(g17093) ) ;
INV     gate6148  (.A(g13191), .Z(II18168) ) ;
INV     gate6149  (.A(II18168), .Z(g17096) ) ;
INV     gate6150  (.A(g14262), .Z(g17120) ) ;
INV     gate6151  (.A(g14321), .Z(g17121) ) ;
INV     gate6152  (.A(g14348), .Z(g17122) ) ;
NAND2   gate6153  (.A(g10323), .B(g11527), .Z(g14051) ) ;
INV     gate6154  (.A(g14051), .Z(g17124) ) ;
INV     gate6155  (.A(g13191), .Z(II18177) ) ;
INV     gate6156  (.A(II18177), .Z(g17125) ) ;
INV     gate6157  (.A(g13605), .Z(II18180) ) ;
INV     gate6158  (.A(II18180), .Z(g17128) ) ;
INV     gate6159  (.A(g14297), .Z(g17135) ) ;
INV     gate6160  (.A(g14348), .Z(g17136) ) ;
INV     gate6161  (.A(g14385), .Z(II18191) ) ;
INV     gate6162  (.A(II18191), .Z(g17141) ) ;
NAND2   gate6163  (.A(g7121), .B(g11584), .Z(g14085) ) ;
INV     gate6164  (.A(g14085), .Z(g17144) ) ;
INV     gate6165  (.A(g14321), .Z(g17147) ) ;
INV     gate6166  (.A(g14348), .Z(g17154) ) ;
INV     gate6167  (.A(g14563), .Z(II18205) ) ;
INV     gate6168  (.A(II18205), .Z(g17155) ) ;
INV     gate6169  (.A(g13350), .Z(g17157) ) ;
INV     gate6170  (.A(g12918), .Z(II18214) ) ;
INV     gate6171  (.A(II18214), .Z(g17178) ) ;
INV     gate6172  (.A(g13605), .Z(II18221) ) ;
INV     gate6173  (.A(II18221), .Z(g17183) ) ;
INV     gate6174  (.A(g13793), .Z(II18224) ) ;
INV     gate6175  (.A(II18224), .Z(g17188) ) ;
AND2    gate6176  (.A(g74), .B(g12369), .Z(g14708) ) ;
INV     gate6177  (.A(g14708), .Z(g17189) ) ;
INV     gate6178  (.A(g14639), .Z(II18233) ) ;
INV     gate6179  (.A(II18233), .Z(g17197) ) ;
INV     gate6180  (.A(g13144), .Z(II18238) ) ;
INV     gate6181  (.A(II18238), .Z(g17200) ) ;
INV     gate6182  (.A(g14454), .Z(g17216) ) ;
INV     gate6183  (.A(g14676), .Z(II18245) ) ;
INV     gate6184  (.A(II18245), .Z(g17221) ) ;
INV     gate6185  (.A(g12938), .Z(II18248) ) ;
INV     gate6186  (.A(II18248), .Z(g17224) ) ;
INV     gate6187  (.A(g13177), .Z(II18252) ) ;
INV     gate6188  (.A(II18252), .Z(g17226) ) ;
INV     gate6189  (.A(g14454), .Z(g17242) ) ;
INV     gate6190  (.A(g12946), .Z(II18259) ) ;
INV     gate6191  (.A(II18259), .Z(g17247) ) ;
INV     gate6192  (.A(g13857), .Z(II18262) ) ;
INV     gate6193  (.A(II18262), .Z(g17248) ) ;
INV     gate6194  (.A(g13350), .Z(II18265) ) ;
INV     gate6195  (.A(II18265), .Z(g17249) ) ;
INV     gate6196  (.A(g13191), .Z(II18270) ) ;
INV     gate6197  (.A(II18270), .Z(g17271) ) ;
INV     gate6198  (.A(g1075), .Z(II18276) ) ;
INV     gate6199  (.A(g12951), .Z(II18280) ) ;
INV     gate6200  (.A(II18280), .Z(g17296) ) ;
INV     gate6201  (.A(g14454), .Z(g17301) ) ;
INV     gate6202  (.A(g13638), .Z(II18285) ) ;
INV     gate6203  (.A(II18285), .Z(g17302) ) ;
NAND2   gate6204  (.A(g12492), .B(g12443), .Z(g14876) ) ;
INV     gate6205  (.A(g14876), .Z(g17308) ) ;
INV     gate6206  (.A(g1079), .Z(II18293) ) ;
INV     gate6207  (.A(g1418), .Z(II18297) ) ;
INV     gate6208  (.A(g12976), .Z(II18301) ) ;
INV     gate6209  (.A(II18301), .Z(g17324) ) ;
INV     gate6210  (.A(g14790), .Z(II18304) ) ;
INV     gate6211  (.A(II18304), .Z(g17325) ) ;
INV     gate6212  (.A(g12977), .Z(II18307) ) ;
INV     gate6213  (.A(II18307), .Z(g17326) ) ;
INV     gate6214  (.A(g12978), .Z(II18310) ) ;
INV     gate6215  (.A(II18310), .Z(g17327) ) ;
INV     gate6216  (.A(g13350), .Z(II18313) ) ;
INV     gate6217  (.A(II18313), .Z(g17328) ) ;
INV     gate6218  (.A(g14454), .Z(g17366) ) ;
INV     gate6219  (.A(g13605), .Z(II18320) ) ;
INV     gate6220  (.A(II18320), .Z(g17367) ) ;
INV     gate6221  (.A(g13680), .Z(II18323) ) ;
INV     gate6222  (.A(II18323), .Z(g17384) ) ;
NAND2   gate6223  (.A(g12553), .B(g10266), .Z(g14915) ) ;
INV     gate6224  (.A(g14915), .Z(g17389) ) ;
NAND2   gate6225  (.A(g12593), .B(g12772), .Z(g14755) ) ;
INV     gate6226  (.A(g14755), .Z(g17390) ) ;
NAND2   gate6227  (.A(g12558), .B(g12505), .Z(g14924) ) ;
INV     gate6228  (.A(g14924), .Z(g17392) ) ;
INV     gate6229  (.A(g1083), .Z(II18333) ) ;
INV     gate6230  (.A(g1422), .Z(II18337) ) ;
INV     gate6231  (.A(g14308), .Z(II18341) ) ;
INV     gate6232  (.A(II18341), .Z(g17408) ) ;
INV     gate6233  (.A(g13003), .Z(II18344) ) ;
INV     gate6234  (.A(II18344), .Z(g17409) ) ;
INV     gate6235  (.A(g12955), .Z(g17410) ) ;
INV     gate6236  (.A(g14454), .Z(g17411) ) ;
INV     gate6237  (.A(g13716), .Z(II18350) ) ;
INV     gate6238  (.A(II18350), .Z(g17413) ) ;
NAND2   gate6239  (.A(g12553), .B(g12772), .Z(g14627) ) ;
INV     gate6240  (.A(g14627), .Z(g17414) ) ;
NAND2   gate6241  (.A(g12593), .B(g12405), .Z(g14797) ) ;
INV     gate6242  (.A(g14797), .Z(g17415) ) ;
NAND2   gate6243  (.A(g12604), .B(g10281), .Z(g14956) ) ;
INV     gate6244  (.A(g14956), .Z(g17416) ) ;
NAND2   gate6245  (.A(g12651), .B(g12798), .Z(g14804) ) ;
INV     gate6246  (.A(g14804), .Z(g17417) ) ;
NAND2   gate6247  (.A(g12609), .B(g12571), .Z(g14965) ) ;
INV     gate6248  (.A(g14965), .Z(g17419) ) ;
INV     gate6249  (.A(g1426), .Z(II18360) ) ;
INV     gate6250  (.A(g13009), .Z(II18364) ) ;
INV     gate6251  (.A(II18364), .Z(g17427) ) ;
INV     gate6252  (.A(g13010), .Z(II18367) ) ;
INV     gate6253  (.A(II18367), .Z(g17428) ) ;
INV     gate6254  (.A(g14873), .Z(II18370) ) ;
INV     gate6255  (.A(II18370), .Z(g17429) ) ;
INV     gate6256  (.A(g13011), .Z(II18373) ) ;
INV     gate6257  (.A(II18373), .Z(g17430) ) ;
INV     gate6258  (.A(g14332), .Z(II18376) ) ;
INV     gate6259  (.A(II18376), .Z(g17431) ) ;
INV     gate6260  (.A(g13012), .Z(II18379) ) ;
INV     gate6261  (.A(II18379), .Z(g17432) ) ;
INV     gate6262  (.A(g13350), .Z(II18382) ) ;
INV     gate6263  (.A(II18382), .Z(g17433) ) ;
INV     gate6264  (.A(g12955), .Z(g17465) ) ;
INV     gate6265  (.A(g12983), .Z(g17466) ) ;
NOR2    gate6266  (.A(g12289), .B(g2735), .Z(g14339) ) ;
INV     gate6267  (.A(g14339), .Z(g17467) ) ;
INV     gate6268  (.A(g14454), .Z(g17470) ) ;
INV     gate6269  (.A(g14454), .Z(g17471) ) ;
NAND2   gate6270  (.A(g12553), .B(g12405), .Z(g14656) ) ;
INV     gate6271  (.A(g14656), .Z(g17472) ) ;
NAND2   gate6272  (.A(g12593), .B(g12443), .Z(g14841) ) ;
INV     gate6273  (.A(g14841), .Z(g17473) ) ;
INV     gate6274  (.A(g13745), .Z(II18398) ) ;
INV     gate6275  (.A(II18398), .Z(g17475) ) ;
NAND2   gate6276  (.A(g12604), .B(g12798), .Z(g14665) ) ;
INV     gate6277  (.A(g14665), .Z(g17476) ) ;
NAND2   gate6278  (.A(g12651), .B(g12453), .Z(g14848) ) ;
INV     gate6279  (.A(g14848), .Z(g17477) ) ;
NAND2   gate6280  (.A(g12662), .B(g10312), .Z(g14996) ) ;
INV     gate6281  (.A(g14996), .Z(g17478) ) ;
NAND2   gate6282  (.A(g12700), .B(g12824), .Z(g14855) ) ;
INV     gate6283  (.A(g14855), .Z(g17479) ) ;
NAND2   gate6284  (.A(g12667), .B(g12622), .Z(g15005) ) ;
INV     gate6285  (.A(g15005), .Z(g17481) ) ;
INV     gate6286  (.A(g13017), .Z(II18408) ) ;
INV     gate6287  (.A(II18408), .Z(g17485) ) ;
INV     gate6288  (.A(g13018), .Z(II18411) ) ;
INV     gate6289  (.A(II18411), .Z(g17486) ) ;
INV     gate6290  (.A(g14359), .Z(II18414) ) ;
INV     gate6291  (.A(II18414), .Z(g17487) ) ;
INV     gate6292  (.A(g12955), .Z(g17489) ) ;
INV     gate6293  (.A(g12983), .Z(g17491) ) ;
INV     gate6294  (.A(g14339), .Z(g17494) ) ;
NAND2   gate6295  (.A(g12553), .B(g12443), .Z(g14683) ) ;
INV     gate6296  (.A(g14683), .Z(g17496) ) ;
NAND2   gate6297  (.A(g12646), .B(g10266), .Z(g14879) ) ;
INV     gate6298  (.A(g14879), .Z(g17497) ) ;
NAND2   gate6299  (.A(g12604), .B(g12453), .Z(g14688) ) ;
INV     gate6300  (.A(g14688), .Z(g17498) ) ;
NAND2   gate6301  (.A(g12651), .B(g12505), .Z(g14885) ) ;
INV     gate6302  (.A(g14885), .Z(g17499) ) ;
INV     gate6303  (.A(g13782), .Z(II18434) ) ;
INV     gate6304  (.A(II18434), .Z(g17501) ) ;
NAND2   gate6305  (.A(g12662), .B(g12824), .Z(g14697) ) ;
INV     gate6306  (.A(g14697), .Z(g17502) ) ;
NAND2   gate6307  (.A(g12700), .B(g12515), .Z(g14892) ) ;
INV     gate6308  (.A(g14892), .Z(g17503) ) ;
NAND2   gate6309  (.A(g12711), .B(g10341), .Z(g15021) ) ;
INV     gate6310  (.A(g15021), .Z(g17504) ) ;
NAND2   gate6311  (.A(g12744), .B(g10421), .Z(g14899) ) ;
INV     gate6312  (.A(g14899), .Z(g17505) ) ;
NAND2   gate6313  (.A(g12716), .B(g12680), .Z(g15030) ) ;
INV     gate6314  (.A(g15030), .Z(g17507) ) ;
INV     gate6315  (.A(g13027), .Z(II18443) ) ;
INV     gate6316  (.A(II18443), .Z(g17508) ) ;
INV     gate6317  (.A(g13028), .Z(II18446) ) ;
INV     gate6318  (.A(II18446), .Z(g17509) ) ;
INV     gate6319  (.A(g12983), .Z(g17512) ) ;
NAND2   gate6320  (.A(g12646), .B(g12772), .Z(g14918) ) ;
INV     gate6321  (.A(g14918), .Z(g17518) ) ;
INV     gate6322  (.A(g5276), .Z(II18460) ) ;
NAND2   gate6323  (.A(g12604), .B(g12505), .Z(g14727) ) ;
INV     gate6324  (.A(g14727), .Z(g17521) ) ;
NAND2   gate6325  (.A(g12695), .B(g10281), .Z(g14927) ) ;
INV     gate6326  (.A(g14927), .Z(g17522) ) ;
NAND2   gate6327  (.A(g12662), .B(g12515), .Z(g14732) ) ;
INV     gate6328  (.A(g14732), .Z(g17523) ) ;
NAND2   gate6329  (.A(g12700), .B(g12571), .Z(g14933) ) ;
INV     gate6330  (.A(g14933), .Z(g17524) ) ;
INV     gate6331  (.A(g13809), .Z(II18469) ) ;
INV     gate6332  (.A(II18469), .Z(g17526) ) ;
NAND2   gate6333  (.A(g12711), .B(g10421), .Z(g14741) ) ;
INV     gate6334  (.A(g14741), .Z(g17527) ) ;
NAND2   gate6335  (.A(g12744), .B(g12581), .Z(g14940) ) ;
INV     gate6336  (.A(g14940), .Z(g17528) ) ;
NAND2   gate6337  (.A(g12755), .B(g7142), .Z(g15039) ) ;
INV     gate6338  (.A(g15039), .Z(g17529) ) ;
NAND2   gate6339  (.A(g12785), .B(g10491), .Z(g14947) ) ;
INV     gate6340  (.A(g14947), .Z(g17530) ) ;
INV     gate6341  (.A(g14031), .Z(II18476) ) ;
INV     gate6342  (.A(II18476), .Z(g17531) ) ;
INV     gate6343  (.A(g13041), .Z(II18479) ) ;
INV     gate6344  (.A(II18479), .Z(g17532) ) ;
INV     gate6345  (.A(g13350), .Z(II18482) ) ;
INV     gate6346  (.A(II18482), .Z(g17533) ) ;
OR2     gate6347  (.A(g10278), .B(g12768), .Z(g12911) ) ;
INV     gate6348  (.A(g12911), .Z(g17573) ) ;
NAND2   gate6349  (.A(g12492), .B(g10266), .Z(g14921) ) ;
INV     gate6350  (.A(g14921), .Z(g17575) ) ;
NAND2   gate6351  (.A(g12646), .B(g12405), .Z(g14953) ) ;
INV     gate6352  (.A(g14953), .Z(g17576) ) ;
INV     gate6353  (.A(g5283), .Z(II18504) ) ;
NAND2   gate6354  (.A(g12695), .B(g12798), .Z(g14959) ) ;
INV     gate6355  (.A(g14959), .Z(g17579) ) ;
INV     gate6356  (.A(g5623), .Z(II18509) ) ;
NAND2   gate6357  (.A(g12662), .B(g12571), .Z(g14768) ) ;
INV     gate6358  (.A(g14768), .Z(g17582) ) ;
NAND2   gate6359  (.A(g12739), .B(g10312), .Z(g14968) ) ;
INV     gate6360  (.A(g14968), .Z(g17583) ) ;
NAND2   gate6361  (.A(g12711), .B(g12581), .Z(g14773) ) ;
INV     gate6362  (.A(g14773), .Z(g17584) ) ;
NAND2   gate6363  (.A(g12744), .B(g12622), .Z(g14974) ) ;
INV     gate6364  (.A(g14974), .Z(g17585) ) ;
INV     gate6365  (.A(g13835), .Z(II18518) ) ;
INV     gate6366  (.A(II18518), .Z(g17587) ) ;
NAND2   gate6367  (.A(g12755), .B(g10491), .Z(g14782) ) ;
INV     gate6368  (.A(g14782), .Z(g17588) ) ;
NAND2   gate6369  (.A(g12785), .B(g12632), .Z(g14981) ) ;
INV     gate6370  (.A(g14981), .Z(g17589) ) ;
INV     gate6371  (.A(g14443), .Z(II18523) ) ;
INV     gate6372  (.A(II18523), .Z(g17590) ) ;
INV     gate6373  (.A(g13055), .Z(II18526) ) ;
INV     gate6374  (.A(II18526), .Z(g17591) ) ;
NAND2   gate6375  (.A(g12492), .B(g12772), .Z(g14794) ) ;
INV     gate6376  (.A(g14794), .Z(g17599) ) ;
NAND2   gate6377  (.A(g12646), .B(g12443), .Z(g14659) ) ;
INV     gate6378  (.A(g14659), .Z(g17600) ) ;
NAND2   gate6379  (.A(g12558), .B(g10281), .Z(g14962) ) ;
INV     gate6380  (.A(g14962), .Z(g17602) ) ;
NAND2   gate6381  (.A(g12695), .B(g12453), .Z(g14993) ) ;
INV     gate6382  (.A(g14993), .Z(g17603) ) ;
INV     gate6383  (.A(g5630), .Z(II18555) ) ;
NAND2   gate6384  (.A(g12739), .B(g12824), .Z(g14999) ) ;
INV     gate6385  (.A(g14999), .Z(g17606) ) ;
INV     gate6386  (.A(g5969), .Z(II18560) ) ;
NAND2   gate6387  (.A(g12711), .B(g12622), .Z(g14817) ) ;
INV     gate6388  (.A(g14817), .Z(g17609) ) ;
NAND2   gate6389  (.A(g12780), .B(g10341), .Z(g15008) ) ;
INV     gate6390  (.A(g15008), .Z(g17610) ) ;
NAND2   gate6391  (.A(g12755), .B(g12632), .Z(g14822) ) ;
INV     gate6392  (.A(g14822), .Z(g17611) ) ;
NAND2   gate6393  (.A(g12785), .B(g12680), .Z(g15014) ) ;
INV     gate6394  (.A(g15014), .Z(g17612) ) ;
INV     gate6395  (.A(g13074), .Z(II18571) ) ;
INV     gate6396  (.A(II18571), .Z(g17614) ) ;
INV     gate6397  (.A(g13075), .Z(II18574) ) ;
INV     gate6398  (.A(II18574), .Z(g17615) ) ;
OR2     gate6399  (.A(g10320), .B(g11048), .Z(g14309) ) ;
INV     gate6400  (.A(g14309), .Z(g17616) ) ;
NAND2   gate6401  (.A(g7150), .B(g10515), .Z(g12933) ) ;
INV     gate6402  (.A(g12933), .Z(g17637) ) ;
NAND2   gate6403  (.A(g12492), .B(g12405), .Z(g14838) ) ;
INV     gate6404  (.A(g14838), .Z(g17638) ) ;
INV     gate6405  (.A(g5335), .Z(II18600) ) ;
NAND2   gate6406  (.A(g12558), .B(g12798), .Z(g14845) ) ;
INV     gate6407  (.A(g14845), .Z(g17641) ) ;
NAND2   gate6408  (.A(g12695), .B(g12505), .Z(g14691) ) ;
INV     gate6409  (.A(g14691), .Z(g17642) ) ;
NAND2   gate6410  (.A(g12609), .B(g10312), .Z(g15002) ) ;
INV     gate6411  (.A(g15002), .Z(g17644) ) ;
NAND2   gate6412  (.A(g12739), .B(g12515), .Z(g15018) ) ;
INV     gate6413  (.A(g15018), .Z(g17645) ) ;
INV     gate6414  (.A(g5976), .Z(II18609) ) ;
NAND2   gate6415  (.A(g12780), .B(g10421), .Z(g15024) ) ;
INV     gate6416  (.A(g15024), .Z(g17648) ) ;
INV     gate6417  (.A(g6315), .Z(II18614) ) ;
NAND2   gate6418  (.A(g12755), .B(g12680), .Z(g14868) ) ;
INV     gate6419  (.A(g14868), .Z(g17651) ) ;
NAND2   gate6420  (.A(g12806), .B(g7142), .Z(g15033) ) ;
INV     gate6421  (.A(g15033), .Z(g17652) ) ;
NAND2   gate6422  (.A(g12593), .B(g10266), .Z(g14720) ) ;
INV     gate6423  (.A(g14720), .Z(g17672) ) ;
NAND2   gate6424  (.A(g7704), .B(g12772), .Z(g14723) ) ;
INV     gate6425  (.A(g14723), .Z(g17673) ) ;
INV     gate6426  (.A(g5320), .Z(II18647) ) ;
NAND2   gate6427  (.A(g7167), .B(g10537), .Z(g12941) ) ;
INV     gate6428  (.A(g12941), .Z(g17676) ) ;
NAND2   gate6429  (.A(g12558), .B(g12453), .Z(g14882) ) ;
INV     gate6430  (.A(g14882), .Z(g17677) ) ;
INV     gate6431  (.A(g5681), .Z(II18653) ) ;
NAND2   gate6432  (.A(g12609), .B(g12824), .Z(g14889) ) ;
INV     gate6433  (.A(g14889), .Z(g17680) ) ;
NAND2   gate6434  (.A(g12739), .B(g12571), .Z(g14735) ) ;
INV     gate6435  (.A(g14735), .Z(g17681) ) ;
NAND2   gate6436  (.A(g12667), .B(g10341), .Z(g15027) ) ;
INV     gate6437  (.A(g15027), .Z(g17683) ) ;
NAND2   gate6438  (.A(g12780), .B(g12581), .Z(g15036) ) ;
INV     gate6439  (.A(g15036), .Z(g17684) ) ;
INV     gate6440  (.A(g6322), .Z(II18662) ) ;
NAND2   gate6441  (.A(g12806), .B(g10491), .Z(g15042) ) ;
INV     gate6442  (.A(g15042), .Z(g17687) ) ;
INV     gate6443  (.A(g6661), .Z(II18667) ) ;
INV     gate6444  (.A(g13101), .Z(II18674) ) ;
INV     gate6445  (.A(II18674), .Z(g17691) ) ;
NAND2   gate6446  (.A(g7704), .B(g12405), .Z(g14758) ) ;
INV     gate6447  (.A(g14758), .Z(g17707) ) ;
NAND2   gate6448  (.A(g12651), .B(g10281), .Z(g14761) ) ;
INV     gate6449  (.A(g14761), .Z(g17709) ) ;
NAND2   gate6450  (.A(g7738), .B(g12798), .Z(g14764) ) ;
INV     gate6451  (.A(g14764), .Z(g17710) ) ;
INV     gate6452  (.A(g5666), .Z(II18694) ) ;
NAND2   gate6453  (.A(g7184), .B(g10561), .Z(g12947) ) ;
INV     gate6454  (.A(g12947), .Z(g17713) ) ;
NAND2   gate6455  (.A(g12609), .B(g12515), .Z(g14930) ) ;
INV     gate6456  (.A(g14930), .Z(g17714) ) ;
INV     gate6457  (.A(g6027), .Z(II18700) ) ;
NAND2   gate6458  (.A(g12667), .B(g10421), .Z(g14937) ) ;
INV     gate6459  (.A(g14937), .Z(g17717) ) ;
NAND2   gate6460  (.A(g12780), .B(g12622), .Z(g14776) ) ;
INV     gate6461  (.A(g14776), .Z(g17718) ) ;
NAND2   gate6462  (.A(g12716), .B(g7142), .Z(g15045) ) ;
INV     gate6463  (.A(g15045), .Z(g17720) ) ;
NAND2   gate6464  (.A(g12806), .B(g12632), .Z(g12915) ) ;
INV     gate6465  (.A(g12915), .Z(g17721) ) ;
INV     gate6466  (.A(g6668), .Z(II18709) ) ;
INV     gate6467  (.A(g14238), .Z(g17733) ) ;
NAND2   gate6468  (.A(g7738), .B(g12453), .Z(g14807) ) ;
INV     gate6469  (.A(g14807), .Z(g17735) ) ;
NAND2   gate6470  (.A(g12700), .B(g10312), .Z(g14810) ) ;
INV     gate6471  (.A(g14810), .Z(g17737) ) ;
NAND2   gate6472  (.A(g7766), .B(g12824), .Z(g14813) ) ;
INV     gate6473  (.A(g14813), .Z(g17738) ) ;
INV     gate6474  (.A(g6012), .Z(II18728) ) ;
NAND2   gate6475  (.A(g7209), .B(g10578), .Z(g12972) ) ;
INV     gate6476  (.A(g12972), .Z(g17741) ) ;
NAND2   gate6477  (.A(g12667), .B(g12581), .Z(g14971) ) ;
INV     gate6478  (.A(g14971), .Z(g17742) ) ;
INV     gate6479  (.A(g6373), .Z(II18734) ) ;
NAND2   gate6480  (.A(g12716), .B(g10491), .Z(g14978) ) ;
INV     gate6481  (.A(g14978), .Z(g17745) ) ;
NAND2   gate6482  (.A(g12806), .B(g12680), .Z(g14825) ) ;
INV     gate6483  (.A(g14825), .Z(g17746) ) ;
INV     gate6484  (.A(g14262), .Z(g17754) ) ;
NAND2   gate6485  (.A(g7766), .B(g12515), .Z(g14858) ) ;
INV     gate6486  (.A(g14858), .Z(g17756) ) ;
NAND2   gate6487  (.A(g12744), .B(g10341), .Z(g14861) ) ;
INV     gate6488  (.A(g14861), .Z(g17758) ) ;
NAND2   gate6489  (.A(g7791), .B(g10421), .Z(g14864) ) ;
INV     gate6490  (.A(g14864), .Z(g17759) ) ;
INV     gate6491  (.A(g6358), .Z(II18752) ) ;
NAND2   gate6492  (.A(g7228), .B(g10598), .Z(g13000) ) ;
INV     gate6493  (.A(g13000), .Z(g17762) ) ;
NAND2   gate6494  (.A(g12716), .B(g12632), .Z(g15011) ) ;
INV     gate6495  (.A(g15011), .Z(g17763) ) ;
INV     gate6496  (.A(g6719), .Z(II18758) ) ;
INV     gate6497  (.A(g14297), .Z(g17772) ) ;
NAND2   gate6498  (.A(g7791), .B(g12581), .Z(g14902) ) ;
INV     gate6499  (.A(g14902), .Z(g17774) ) ;
NAND2   gate6500  (.A(g12785), .B(g7142), .Z(g14905) ) ;
INV     gate6501  (.A(g14905), .Z(g17776) ) ;
NAND2   gate6502  (.A(g7812), .B(g10491), .Z(g14908) ) ;
INV     gate6503  (.A(g14908), .Z(g17777) ) ;
INV     gate6504  (.A(g6704), .Z(II18778) ) ;
INV     gate6505  (.A(g13138), .Z(II18788) ) ;
INV     gate6506  (.A(II18788), .Z(g17782) ) ;
INV     gate6507  (.A(g5327), .Z(II18795) ) ;
INV     gate6508  (.A(g14321), .Z(g17789) ) ;
NAND2   gate6509  (.A(g7812), .B(g12632), .Z(g14950) ) ;
INV     gate6510  (.A(g14950), .Z(g17791) ) ;
INV     gate6511  (.A(g13350), .Z(g17794) ) ;
OR2     gate6512  (.A(g8928), .B(g10511), .Z(g12925) ) ;
INV     gate6513  (.A(g12925), .Z(g17811) ) ;
INV     gate6514  (.A(g13716), .Z(II18810) ) ;
INV     gate6515  (.A(II18810), .Z(g17812) ) ;
INV     gate6516  (.A(g5673), .Z(II18813) ) ;
INV     gate6517  (.A(g14348), .Z(g17815) ) ;
INV     gate6518  (.A(g13745), .Z(II18822) ) ;
INV     gate6519  (.A(II18822), .Z(g17818) ) ;
INV     gate6520  (.A(g6019), .Z(II18825) ) ;
INV     gate6521  (.A(g13350), .Z(II18829) ) ;
INV     gate6522  (.A(II18829), .Z(g17821) ) ;
INV     gate6523  (.A(g13782), .Z(II18832) ) ;
INV     gate6524  (.A(II18832), .Z(g17844) ) ;
INV     gate6525  (.A(g6365), .Z(II18835) ) ;
INV     gate6526  (.A(g13716), .Z(II18839) ) ;
INV     gate6527  (.A(II18839), .Z(g17847) ) ;
INV     gate6528  (.A(g13809), .Z(II18842) ) ;
INV     gate6529  (.A(II18842), .Z(g17870) ) ;
INV     gate6530  (.A(g6711), .Z(II18845) ) ;
INV     gate6531  (.A(g14290), .Z(II18849) ) ;
INV     gate6532  (.A(II18849), .Z(g17873) ) ;
INV     gate6533  (.A(g13716), .Z(II18852) ) ;
INV     gate6534  (.A(II18852), .Z(g17926) ) ;
INV     gate6535  (.A(g13745), .Z(II18855) ) ;
INV     gate6536  (.A(II18855), .Z(g17929) ) ;
INV     gate6537  (.A(g13835), .Z(II18858) ) ;
INV     gate6538  (.A(II18858), .Z(g17952) ) ;
INV     gate6539  (.A(g14307), .Z(II18861) ) ;
INV     gate6540  (.A(II18861), .Z(g17953) ) ;
INV     gate6541  (.A(g14314), .Z(II18865) ) ;
INV     gate6542  (.A(II18865), .Z(g17955) ) ;
INV     gate6543  (.A(g14315), .Z(II18868) ) ;
INV     gate6544  (.A(II18868), .Z(g18008) ) ;
NAND2   gate6545  (.A(g7704), .B(g12443), .Z(g14800) ) ;
INV     gate6546  (.A(g14800), .Z(g18061) ) ;
INV     gate6547  (.A(g13745), .Z(II18872) ) ;
INV     gate6548  (.A(II18872), .Z(g18062) ) ;
INV     gate6549  (.A(g13782), .Z(II18875) ) ;
INV     gate6550  (.A(II18875), .Z(g18065) ) ;
INV     gate6551  (.A(g13267), .Z(g18088) ) ;
INV     gate6552  (.A(g13267), .Z(II18879) ) ;
INV     gate6553  (.A(II18879), .Z(g18091) ) ;
INV     gate6554  (.A(g16580), .Z(II18882) ) ;
INV     gate6555  (.A(g16643), .Z(II18885) ) ;
INV     gate6556  (.A(g16644), .Z(II18888) ) ;
INV     gate6557  (.A(g16676), .Z(II18891) ) ;
INV     gate6558  (.A(g16708), .Z(II18894) ) ;
INV     gate6559  (.A(g16738), .Z(II18897) ) ;
INV     gate6560  (.A(g16767), .Z(II18900) ) ;
INV     gate6561  (.A(g16872), .Z(II18903) ) ;
INV     gate6562  (.A(g16963), .Z(II18906) ) ;
INV     gate6563  (.A(g16873), .Z(II18909) ) ;
NOR2    gate6564  (.A(g12834), .B(g13350), .Z(g15050) ) ;
INV     gate6565  (.A(g15050), .Z(II18912) ) ;
INV     gate6566  (.A(II18912), .Z(g18102) ) ;
NOR2    gate6567  (.A(g13350), .B(g6814), .Z(g15060) ) ;
INV     gate6568  (.A(g15060), .Z(II19012) ) ;
INV     gate6569  (.A(II19012), .Z(g18200) ) ;
AND2    gate6570  (.A(g10361), .B(g12955), .Z(g15078) ) ;
INV     gate6571  (.A(g15078), .Z(II19235) ) ;
AND2    gate6572  (.A(g2151), .B(g12955), .Z(g15079) ) ;
INV     gate6573  (.A(g15079), .Z(II19238) ) ;
AND2    gate6574  (.A(g10362), .B(g12983), .Z(g15083) ) ;
INV     gate6575  (.A(g15083), .Z(II19345) ) ;
AND2    gate6576  (.A(g2710), .B(g12983), .Z(g15084) ) ;
INV     gate6577  (.A(g15084), .Z(II19348) ) ;
INV     gate6578  (.A(g15085), .Z(II19384) ) ;
INV     gate6579  (.A(II19384), .Z(g18562) ) ;
NOR2    gate6580  (.A(g6959), .B(g13605), .Z(g15122) ) ;
INV     gate6581  (.A(g15122), .Z(II19484) ) ;
INV     gate6582  (.A(II19484), .Z(g18660) ) ;
OR2     gate6583  (.A(g10363), .B(g13605), .Z(g15125) ) ;
INV     gate6584  (.A(g15125), .Z(II19487) ) ;
INV     gate6585  (.A(II19487), .Z(g18661) ) ;
INV     gate6586  (.A(g16000), .Z(g18827) ) ;
INV     gate6587  (.A(g17955), .Z(g18828) ) ;
INV     gate6588  (.A(g15171), .Z(g18829) ) ;
INV     gate6589  (.A(g18008), .Z(g18830) ) ;
INV     gate6590  (.A(g15224), .Z(g18831) ) ;
INV     gate6591  (.A(g15634), .Z(g18832) ) ;
INV     gate6592  (.A(g17587), .Z(II19661) ) ;
INV     gate6593  (.A(II19661), .Z(g18833) ) ;
INV     gate6594  (.A(g15938), .Z(g18874) ) ;
INV     gate6595  (.A(g15171), .Z(g18875) ) ;
INV     gate6596  (.A(g15373), .Z(g18876) ) ;
INV     gate6597  (.A(g15224), .Z(g18877) ) ;
INV     gate6598  (.A(g15426), .Z(g18878) ) ;
INV     gate6599  (.A(g15656), .Z(g18880) ) ;
INV     gate6600  (.A(g15932), .Z(II19671) ) ;
INV     gate6601  (.A(g15932), .Z(II19674) ) ;
INV     gate6602  (.A(II19674), .Z(g18882) ) ;
INV     gate6603  (.A(g15938), .Z(g18883) ) ;
INV     gate6604  (.A(g15938), .Z(g18884) ) ;
INV     gate6605  (.A(g15979), .Z(g18885) ) ;
INV     gate6606  (.A(g16000), .Z(g18886) ) ;
INV     gate6607  (.A(g15373), .Z(g18887) ) ;
INV     gate6608  (.A(g15426), .Z(g18888) ) ;
INV     gate6609  (.A(g15509), .Z(g18889) ) ;
INV     gate6610  (.A(g16053), .Z(g18891) ) ;
INV     gate6611  (.A(g15680), .Z(g18892) ) ;
INV     gate6612  (.A(g16000), .Z(g18894) ) ;
INV     gate6613  (.A(g16000), .Z(g18895) ) ;
INV     gate6614  (.A(g16031), .Z(g18896) ) ;
INV     gate6615  (.A(g15509), .Z(g18897) ) ;
INV     gate6616  (.A(g15566), .Z(g18898) ) ;
INV     gate6617  (.A(g15758), .Z(g18903) ) ;
INV     gate6618  (.A(g16053), .Z(g18904) ) ;
INV     gate6619  (.A(g16077), .Z(g18905) ) ;
INV     gate6620  (.A(g15979), .Z(g18907) ) ;
INV     gate6621  (.A(g16100), .Z(g18908) ) ;
INV     gate6622  (.A(g15169), .Z(g18911) ) ;
INV     gate6623  (.A(g16053), .Z(g18916) ) ;
INV     gate6624  (.A(g16077), .Z(g18917) ) ;
AND4    gate6625  (.A(g11547), .B(g11592), .C(g6789), .D(II18620), .Z(g17653) ) ;
INV     gate6626  (.A(g17653), .Z(II19704) ) ;
INV     gate6627  (.A(II19704), .Z(g18918) ) ;
INV     gate6628  (.A(g17590), .Z(II19707) ) ;
INV     gate6629  (.A(II19707), .Z(g18926) ) ;
INV     gate6630  (.A(g16100), .Z(g18929) ) ;
OR2     gate6631  (.A(g10819), .B(g13211), .Z(g15789) ) ;
INV     gate6632  (.A(g15789), .Z(g18930) ) ;
INV     gate6633  (.A(g16031), .Z(g18931) ) ;
INV     gate6634  (.A(g16136), .Z(g18932) ) ;
INV     gate6635  (.A(g16053), .Z(g18938) ) ;
INV     gate6636  (.A(g16077), .Z(g18939) ) ;
INV     gate6637  (.A(g17431), .Z(II19719) ) ;
INV     gate6638  (.A(II19719), .Z(g18940) ) ;
INV     gate6639  (.A(g15938), .Z(g18944) ) ;
INV     gate6640  (.A(g16100), .Z(g18945) ) ;
INV     gate6641  (.A(g16100), .Z(g18946) ) ;
INV     gate6642  (.A(g16136), .Z(g18947) ) ;
OR2     gate6643  (.A(g10821), .B(g13242), .Z(g15800) ) ;
INV     gate6644  (.A(g15800), .Z(g18948) ) ;
INV     gate6645  (.A(g16053), .Z(g18952) ) ;
INV     gate6646  (.A(g16077), .Z(g18953) ) ;
INV     gate6647  (.A(g17427), .Z(g18954) ) ;
AND4    gate6648  (.A(g11547), .B(g11592), .C(g6789), .D(II18716), .Z(g17725) ) ;
INV     gate6649  (.A(g17725), .Z(II19734) ) ;
INV     gate6650  (.A(II19734), .Z(g18957) ) ;
INV     gate6651  (.A(g15938), .Z(g18975) ) ;
INV     gate6652  (.A(g16100), .Z(g18976) ) ;
INV     gate6653  (.A(g16100), .Z(g18977) ) ;
INV     gate6654  (.A(g16000), .Z(g18978) ) ;
INV     gate6655  (.A(g16136), .Z(g18979) ) ;
INV     gate6656  (.A(g16136), .Z(g18980) ) ;
INV     gate6657  (.A(g16077), .Z(g18983) ) ;
INV     gate6658  (.A(g17486), .Z(g18984) ) ;
INV     gate6659  (.A(g15979), .Z(g18988) ) ;
INV     gate6660  (.A(g16000), .Z(g18989) ) ;
INV     gate6661  (.A(g16136), .Z(g18990) ) ;
INV     gate6662  (.A(g16136), .Z(g18991) ) ;
INV     gate6663  (.A(g17812), .Z(II19756) ) ;
INV     gate6664  (.A(II19756), .Z(g18997) ) ;
AND4    gate6665  (.A(g6772), .B(g11592), .C(g6789), .D(II18765), .Z(g17767) ) ;
INV     gate6666  (.A(g17767), .Z(II19759) ) ;
INV     gate6667  (.A(II19759), .Z(g19050) ) ;
OR4     gate6668  (.A(g13411), .B(g13384), .C(g13349), .D(g11016), .Z(g15732) ) ;
INV     gate6669  (.A(g15732), .Z(II19762) ) ;
INV     gate6670  (.A(II19762), .Z(g19061) ) ;
INV     gate6671  (.A(g15979), .Z(g19067) ) ;
INV     gate6672  (.A(g16031), .Z(g19068) ) ;
NAND3   gate6673  (.A(g4332), .B(g4322), .C(g13202), .Z(g15591) ) ;
INV     gate6674  (.A(g15591), .Z(g19071) ) ;
INV     gate6675  (.A(g17818), .Z(II19772) ) ;
INV     gate6676  (.A(II19772), .Z(g19074) ) ;
AND4    gate6677  (.A(g6772), .B(g11592), .C(g11640), .D(II18782), .Z(g17780) ) ;
INV     gate6678  (.A(g17780), .Z(II19775) ) ;
INV     gate6679  (.A(II19775), .Z(g19127) ) ;
AND4    gate6680  (.A(g6772), .B(g11592), .C(g6789), .D(II18785), .Z(g17781) ) ;
INV     gate6681  (.A(g17781), .Z(II19778) ) ;
INV     gate6682  (.A(II19778), .Z(g19128) ) ;
INV     gate6683  (.A(g16031), .Z(g19144) ) ;
AND2    gate6684  (.A(g4311), .B(g13202), .Z(g15574) ) ;
INV     gate6685  (.A(g15574), .Z(g19146) ) ;
INV     gate6686  (.A(g17844), .Z(II19786) ) ;
INV     gate6687  (.A(II19786), .Z(g19147) ) ;
AND4    gate6688  (.A(g6772), .B(g11592), .C(g6789), .D(II18803), .Z(g17793) ) ;
INV     gate6689  (.A(g17793), .Z(II19789) ) ;
INV     gate6690  (.A(II19789), .Z(g19200) ) ;
INV     gate6691  (.A(g17367), .Z(g19208) ) ;
INV     gate6692  (.A(g17870), .Z(II19796) ) ;
INV     gate6693  (.A(II19796), .Z(g19210) ) ;
AND4    gate6694  (.A(g11547), .B(g6782), .C(g11640), .D(II18819), .Z(g17817) ) ;
INV     gate6695  (.A(g17817), .Z(II19799) ) ;
INV     gate6696  (.A(II19799), .Z(g19263) ) ;
OR4     gate6697  (.A(g13383), .B(g13345), .C(g13333), .D(g11010), .Z(g15727) ) ;
INV     gate6698  (.A(g15727), .Z(II19802) ) ;
INV     gate6699  (.A(II19802), .Z(g19264) ) ;
INV     gate6700  (.A(g16100), .Z(g19273) ) ;
INV     gate6701  (.A(g17367), .Z(g19276) ) ;
INV     gate6702  (.A(g17952), .Z(II19813) ) ;
INV     gate6703  (.A(II19813), .Z(g19277) ) ;
INV     gate6704  (.A(g17326), .Z(g19330) ) ;
INV     gate6705  (.A(g1056), .Z(II19818) ) ;
INV     gate6706  (.A(g16136), .Z(g19343) ) ;
INV     gate6707  (.A(g17591), .Z(g19345) ) ;
INV     gate6708  (.A(g17367), .Z(g19351) ) ;
INV     gate6709  (.A(g15758), .Z(g19352) ) ;
INV     gate6710  (.A(g16533), .Z(II19831) ) ;
INV     gate6711  (.A(II19831), .Z(g19353) ) ;
NOR2    gate6712  (.A(g10929), .B(g13260), .Z(g16027) ) ;
INV     gate6713  (.A(g16027), .Z(g19355) ) ;
INV     gate6714  (.A(g1399), .Z(II19837) ) ;
INV     gate6715  (.A(g16249), .Z(g19360) ) ;
INV     gate6716  (.A(g16594), .Z(II19843) ) ;
INV     gate6717  (.A(II19843), .Z(g19361) ) ;
NOR2    gate6718  (.A(g10961), .B(g13273), .Z(g16072) ) ;
INV     gate6719  (.A(g16072), .Z(g19362) ) ;
NOR2    gate6720  (.A(g7666), .B(g13217), .Z(g15825) ) ;
INV     gate6721  (.A(g15825), .Z(g19364) ) ;
INV     gate6722  (.A(g16249), .Z(g19365) ) ;
INV     gate6723  (.A(g15885), .Z(g19366) ) ;
INV     gate6724  (.A(g16615), .Z(II19851) ) ;
INV     gate6725  (.A(II19851), .Z(g19367) ) ;
INV     gate6726  (.A(g16326), .Z(g19368) ) ;
AND3    gate6727  (.A(g13314), .B(g1157), .C(g10666), .Z(g15995) ) ;
INV     gate6728  (.A(g15995), .Z(g19369) ) ;
INV     gate6729  (.A(g15915), .Z(g19370) ) ;
INV     gate6730  (.A(g16640), .Z(II19857) ) ;
INV     gate6731  (.A(II19857), .Z(g19371) ) ;
INV     gate6732  (.A(g16449), .Z(g19373) ) ;
AND3    gate6733  (.A(g13322), .B(g1500), .C(g10699), .Z(g16047) ) ;
INV     gate6734  (.A(g16047), .Z(g19374) ) ;
INV     gate6735  (.A(g16675), .Z(II19863) ) ;
INV     gate6736  (.A(II19863), .Z(g19375) ) ;
INV     gate6737  (.A(g17509), .Z(g19376) ) ;
INV     gate6738  (.A(g17327), .Z(g19379) ) ;
INV     gate6739  (.A(g16326), .Z(g19385) ) ;
INV     gate6740  (.A(g16431), .Z(g19386) ) ;
INV     gate6741  (.A(g16431), .Z(g19387) ) ;
INV     gate6742  (.A(g17532), .Z(g19389) ) ;
INV     gate6743  (.A(g16326), .Z(g19394) ) ;
INV     gate6744  (.A(g16431), .Z(g19395) ) ;
INV     gate6745  (.A(g16431), .Z(g19396) ) ;
INV     gate6746  (.A(g16449), .Z(g19397) ) ;
INV     gate6747  (.A(g16489), .Z(g19398) ) ;
INV     gate6748  (.A(g16489), .Z(g19399) ) ;
NOR2    gate6749  (.A(g7913), .B(g13121), .Z(g16268) ) ;
INV     gate6750  (.A(g16268), .Z(g19407) ) ;
NOR2    gate6751  (.A(g10929), .B(g13307), .Z(g16066) ) ;
INV     gate6752  (.A(g16066), .Z(g19408) ) ;
INV     gate6753  (.A(g16431), .Z(g19409) ) ;
INV     gate6754  (.A(g16449), .Z(g19410) ) ;
INV     gate6755  (.A(g16489), .Z(g19411) ) ;
INV     gate6756  (.A(g16489), .Z(g19412) ) ;
INV     gate6757  (.A(g16349), .Z(g19414) ) ;
INV     gate6758  (.A(g15758), .Z(g19415) ) ;
INV     gate6759  (.A(g15885), .Z(g19416) ) ;
INV     gate6760  (.A(g17178), .Z(g19417) ) ;
INV     gate6761  (.A(g16326), .Z(g19421) ) ;
NOR2    gate6762  (.A(g7943), .B(g13134), .Z(g16292) ) ;
INV     gate6763  (.A(g16292), .Z(g19427) ) ;
NOR2    gate6764  (.A(g10961), .B(g13315), .Z(g16090) ) ;
INV     gate6765  (.A(g16090), .Z(g19428) ) ;
INV     gate6766  (.A(g16489), .Z(g19429) ) ;
INV     gate6767  (.A(g16249), .Z(g19431) ) ;
INV     gate6768  (.A(g15885), .Z(g19432) ) ;
INV     gate6769  (.A(g15915), .Z(g19433) ) ;
INV     gate6770  (.A(g16326), .Z(g19434) ) ;
INV     gate6771  (.A(g16449), .Z(g19435) ) ;
INV     gate6772  (.A(g16349), .Z(g19437) ) ;
INV     gate6773  (.A(g16249), .Z(g19438) ) ;
INV     gate6774  (.A(g15885), .Z(g19439) ) ;
INV     gate6775  (.A(g15915), .Z(g19440) ) ;
INV     gate6776  (.A(g16449), .Z(g19443) ) ;
INV     gate6777  (.A(g15915), .Z(g19445) ) ;
INV     gate6778  (.A(g18088), .Z(II19917) ) ;
INV     gate6779  (.A(II19917), .Z(g19446) ) ;
INV     gate6780  (.A(g15938), .Z(g19451) ) ;
INV     gate6781  (.A(g16326), .Z(g19452) ) ;
INV     gate6782  (.A(g16349), .Z(g19454) ) ;
INV     gate6783  (.A(g17408), .Z(II19927) ) ;
INV     gate6784  (.A(II19927), .Z(g19458) ) ;
INV     gate6785  (.A(g15938), .Z(g19468) ) ;
INV     gate6786  (.A(g16326), .Z(g19469) ) ;
INV     gate6787  (.A(g16000), .Z(g19470) ) ;
INV     gate6788  (.A(g16449), .Z(g19471) ) ;
INV     gate6789  (.A(g16349), .Z(g19472) ) ;
INV     gate6790  (.A(g16349), .Z(g19473) ) ;
INV     gate6791  (.A(g16326), .Z(g19476) ) ;
INV     gate6792  (.A(g16431), .Z(g19477) ) ;
INV     gate6793  (.A(g16000), .Z(g19478) ) ;
INV     gate6794  (.A(g16449), .Z(g19479) ) ;
INV     gate6795  (.A(g16349), .Z(g19480) ) ;
INV     gate6796  (.A(g16349), .Z(g19481) ) ;
INV     gate6797  (.A(g16349), .Z(g19482) ) ;
INV     gate6798  (.A(g16449), .Z(g19489) ) ;
INV     gate6799  (.A(g16489), .Z(g19490) ) ;
INV     gate6800  (.A(g16349), .Z(g19491) ) ;
INV     gate6801  (.A(g16349), .Z(g19492) ) ;
INV     gate6802  (.A(g16349), .Z(g19493) ) ;
INV     gate6803  (.A(g16349), .Z(g19494) ) ;
INV     gate6804  (.A(g16752), .Z(g19498) ) ;
INV     gate6805  (.A(g16782), .Z(g19499) ) ;
NAND2   gate6806  (.A(g921), .B(g13110), .Z(g15674) ) ;
INV     gate6807  (.A(g15674), .Z(g19502) ) ;
INV     gate6808  (.A(g16349), .Z(g19503) ) ;
INV     gate6809  (.A(g16349), .Z(g19504) ) ;
INV     gate6810  (.A(g16349), .Z(g19505) ) ;
INV     gate6811  (.A(g16777), .Z(g19517) ) ;
OR2     gate6812  (.A(g7892), .B(g13432), .Z(g16239) ) ;
INV     gate6813  (.A(g16239), .Z(g19518) ) ;
INV     gate6814  (.A(g16795), .Z(g19519) ) ;
INV     gate6815  (.A(g16826), .Z(g19520) ) ;
INV     gate6816  (.A(g16100), .Z(g19523) ) ;
NAND2   gate6817  (.A(g1266), .B(g13125), .Z(g15695) ) ;
INV     gate6818  (.A(g15695), .Z(g19524) ) ;
INV     gate6819  (.A(g16349), .Z(g19526) ) ;
INV     gate6820  (.A(g16349), .Z(g19527) ) ;
INV     gate6821  (.A(g16349), .Z(g19528) ) ;
INV     gate6822  (.A(g16349), .Z(g19529) ) ;
INV     gate6823  (.A(g16816), .Z(g19531) ) ;
INV     gate6824  (.A(g16821), .Z(g19532) ) ;
OR2     gate6825  (.A(g7898), .B(g13469), .Z(g16261) ) ;
INV     gate6826  (.A(g16261), .Z(g19533) ) ;
INV     gate6827  (.A(g15938), .Z(g19537) ) ;
INV     gate6828  (.A(g16100), .Z(g19538) ) ;
INV     gate6829  (.A(g16129), .Z(g19539) ) ;
INV     gate6830  (.A(g16136), .Z(g19541) ) ;
INV     gate6831  (.A(g16349), .Z(g19542) ) ;
INV     gate6832  (.A(g16349), .Z(g19543) ) ;
INV     gate6833  (.A(g16349), .Z(g19544) ) ;
INV     gate6834  (.A(g16856), .Z(g19552) ) ;
INV     gate6835  (.A(g16782), .Z(g19553) ) ;
INV     gate6836  (.A(g16861), .Z(g19554) ) ;
INV     gate6837  (.A(g15938), .Z(g19558) ) ;
INV     gate6838  (.A(g16129), .Z(g19559) ) ;
INV     gate6839  (.A(g16000), .Z(g19565) ) ;
INV     gate6840  (.A(g16136), .Z(g19566) ) ;
INV     gate6841  (.A(g16164), .Z(g19567) ) ;
INV     gate6842  (.A(g16349), .Z(g19569) ) ;
INV     gate6843  (.A(g16349), .Z(g19570) ) ;
INV     gate6844  (.A(g16877), .Z(g19573) ) ;
INV     gate6845  (.A(g16826), .Z(g19574) ) ;
INV     gate6846  (.A(g16129), .Z(g19577) ) ;
INV     gate6847  (.A(g16000), .Z(g19579) ) ;
INV     gate6848  (.A(g16164), .Z(g19580) ) ;
INV     gate6849  (.A(g16349), .Z(g19586) ) ;
AND2    gate6850  (.A(g13296), .B(g13484), .Z(g15706) ) ;
INV     gate6851  (.A(g15706), .Z(II20035) ) ;
INV     gate6852  (.A(II20035), .Z(g19592) ) ;
INV     gate6853  (.A(g16164), .Z(g19600) ) ;
INV     gate6854  (.A(g16349), .Z(g19602) ) ;
INV     gate6855  (.A(g16349), .Z(g19603) ) ;
INV     gate6856  (.A(g17614), .Z(g19606) ) ;
NAND3   gate6857  (.A(g518), .B(g9158), .C(g13223), .Z(g16264) ) ;
INV     gate6858  (.A(g16264), .Z(g19609) ) ;
INV     gate6859  (.A(g16897), .Z(g19612) ) ;
INV     gate6860  (.A(g16349), .Z(g19617) ) ;
INV     gate6861  (.A(g16349), .Z(g19618) ) ;
INV     gate6862  (.A(g17296), .Z(g19620) ) ;
INV     gate6863  (.A(g17409), .Z(g19626) ) ;
INV     gate6864  (.A(g17015), .Z(g19629) ) ;
INV     gate6865  (.A(g16897), .Z(g19630) ) ;
INV     gate6866  (.A(g16931), .Z(g19633) ) ;
INV     gate6867  (.A(g16349), .Z(g19634) ) ;
INV     gate6868  (.A(g16349), .Z(g19635) ) ;
INV     gate6869  (.A(g16987), .Z(g19636) ) ;
INV     gate6870  (.A(g17324), .Z(g19638) ) ;
INV     gate6871  (.A(g17953), .Z(g19644) ) ;
INV     gate6872  (.A(g17015), .Z(g19649) ) ;
INV     gate6873  (.A(g16971), .Z(g19650) ) ;
INV     gate6874  (.A(g16897), .Z(g19652) ) ;
INV     gate6875  (.A(g16897), .Z(g19653) ) ;
INV     gate6876  (.A(g16931), .Z(g19654) ) ;
INV     gate6877  (.A(g16349), .Z(g19657) ) ;
INV     gate6878  (.A(g16987), .Z(g19658) ) ;
INV     gate6879  (.A(g17062), .Z(g19659) ) ;
INV     gate6880  (.A(g17432), .Z(g19662) ) ;
INV     gate6881  (.A(g17188), .Z(g19666) ) ;
INV     gate6882  (.A(g16897), .Z(g19670) ) ;
INV     gate6883  (.A(g16931), .Z(g19672) ) ;
INV     gate6884  (.A(g16931), .Z(g19673) ) ;
INV     gate6885  (.A(g16987), .Z(g19675) ) ;
INV     gate6886  (.A(g17062), .Z(g19676) ) ;
INV     gate6887  (.A(g17096), .Z(g19677) ) ;
INV     gate6888  (.A(g16752), .Z(g19678) ) ;
INV     gate6889  (.A(g16782), .Z(g19679) ) ;
INV     gate6890  (.A(g17015), .Z(g19682) ) ;
INV     gate6891  (.A(g16931), .Z(g19683) ) ;
INV     gate6892  (.A(g16987), .Z(g19685) ) ;
INV     gate6893  (.A(g17062), .Z(g19686) ) ;
INV     gate6894  (.A(g17096), .Z(g19687) ) ;
INV     gate6895  (.A(g16777), .Z(g19688) ) ;
INV     gate6896  (.A(g16795), .Z(g19689) ) ;
INV     gate6897  (.A(g16826), .Z(g19690) ) ;
INV     gate6898  (.A(g16429), .Z(g19694) ) ;
INV     gate6899  (.A(g17015), .Z(g19695) ) ;
INV     gate6900  (.A(g17015), .Z(g19696) ) ;
INV     gate6901  (.A(g16886), .Z(g19697) ) ;
INV     gate6902  (.A(g16971), .Z(g19698) ) ;
NAND4   gate6903  (.A(g13240), .B(g13115), .C(g7903), .D(g13210), .Z(g15737) ) ;
INV     gate6904  (.A(g15737), .Z(II20116) ) ;
INV     gate6905  (.A(II20116), .Z(g19699) ) ;
INV     gate6906  (.A(g16987), .Z(g19709) ) ;
INV     gate6907  (.A(g17059), .Z(g19710) ) ;
INV     gate6908  (.A(g17062), .Z(g19711) ) ;
INV     gate6909  (.A(g17096), .Z(g19712) ) ;
INV     gate6910  (.A(g16816), .Z(g19713) ) ;
INV     gate6911  (.A(g16821), .Z(g19714) ) ;
INV     gate6912  (.A(g17015), .Z(g19718) ) ;
INV     gate6913  (.A(g16897), .Z(g19719) ) ;
NAND4   gate6914  (.A(g13257), .B(g13130), .C(g7922), .D(g13241), .Z(g15748) ) ;
INV     gate6915  (.A(g15748), .Z(II20130) ) ;
INV     gate6916  (.A(II20130), .Z(g19720) ) ;
INV     gate6917  (.A(g17062), .Z(g19730) ) ;
INV     gate6918  (.A(g17093), .Z(g19731) ) ;
INV     gate6919  (.A(g17096), .Z(g19732) ) ;
INV     gate6920  (.A(g16856), .Z(g19733) ) ;
INV     gate6921  (.A(g16861), .Z(g19734) ) ;
INV     gate6922  (.A(g17015), .Z(g19737) ) ;
NOR2    gate6923  (.A(g10929), .B(g13846), .Z(g15992) ) ;
INV     gate6924  (.A(g15992), .Z(g19738) ) ;
INV     gate6925  (.A(g16931), .Z(g19739) ) ;
INV     gate6926  (.A(g16987), .Z(g19741) ) ;
INV     gate6927  (.A(g17096), .Z(g19742) ) ;
INV     gate6928  (.A(g17125), .Z(g19743) ) ;
INV     gate6929  (.A(g15885), .Z(g19744) ) ;
INV     gate6930  (.A(g16877), .Z(g19745) ) ;
INV     gate6931  (.A(g17015), .Z(g19747) ) ;
INV     gate6932  (.A(g17015), .Z(g19748) ) ;
INV     gate6933  (.A(g16326), .Z(g19750) ) ;
NOR2    gate6934  (.A(g10961), .B(g13861), .Z(g16044) ) ;
INV     gate6935  (.A(g16044), .Z(g19751) ) ;
INV     gate6936  (.A(g16987), .Z(g19753) ) ;
INV     gate6937  (.A(g17062), .Z(g19754) ) ;
INV     gate6938  (.A(g15915), .Z(g19755) ) ;
INV     gate6939  (.A(g17224), .Z(g19757) ) ;
INV     gate6940  (.A(g17015), .Z(g19760) ) ;
INV     gate6941  (.A(g17015), .Z(g19761) ) ;
INV     gate6942  (.A(g16326), .Z(g19762) ) ;
INV     gate6943  (.A(g16431), .Z(g19763) ) ;
INV     gate6944  (.A(g16897), .Z(g19765) ) ;
INV     gate6945  (.A(g16449), .Z(g19766) ) ;
INV     gate6946  (.A(g16987), .Z(g19769) ) ;
INV     gate6947  (.A(g17062), .Z(g19770) ) ;
INV     gate6948  (.A(g17096), .Z(g19771) ) ;
INV     gate6949  (.A(g17183), .Z(g19772) ) ;
INV     gate6950  (.A(g17615), .Z(g19773) ) ;
INV     gate6951  (.A(g17015), .Z(g19776) ) ;
INV     gate6952  (.A(g17015), .Z(g19777) ) ;
INV     gate6953  (.A(g16431), .Z(g19779) ) ;
INV     gate6954  (.A(g16449), .Z(g19780) ) ;
INV     gate6955  (.A(g16489), .Z(g19781) ) ;
INV     gate6956  (.A(g16931), .Z(g19783) ) ;
INV     gate6957  (.A(g16987), .Z(g19785) ) ;
INV     gate6958  (.A(g17062), .Z(g19786) ) ;
INV     gate6959  (.A(g17096), .Z(g19787) ) ;
INV     gate6960  (.A(g17015), .Z(g19789) ) ;
INV     gate6961  (.A(g16971), .Z(g19790) ) ;
INV     gate6962  (.A(g16489), .Z(g19794) ) ;
INV     gate6963  (.A(g17200), .Z(g19798) ) ;
INV     gate6964  (.A(g17062), .Z(g19799) ) ;
INV     gate6965  (.A(g17096), .Z(g19800) ) ;
INV     gate6966  (.A(g15862), .Z(II20216) ) ;
INV     gate6967  (.A(II20216), .Z(g19801) ) ;
INV     gate6968  (.A(g17015), .Z(g19852) ) ;
INV     gate6969  (.A(g17226), .Z(g19860) ) ;
INV     gate6970  (.A(g17096), .Z(g19861) ) ;
INV     gate6971  (.A(g17487), .Z(II20233) ) ;
INV     gate6972  (.A(II20233), .Z(g19862) ) ;
INV     gate6973  (.A(g15885), .Z(g19865) ) ;
INV     gate6974  (.A(g16540), .Z(g19866) ) ;
INV     gate6975  (.A(g16540), .Z(g19869) ) ;
INV     gate6976  (.A(g17015), .Z(g19872) ) ;
INV     gate6977  (.A(g17271), .Z(g19878) ) ;
INV     gate6978  (.A(g15915), .Z(g19881) ) ;
INV     gate6979  (.A(g16540), .Z(g19882) ) ;
INV     gate6980  (.A(g17249), .Z(g19885) ) ;
INV     gate6981  (.A(g17200), .Z(g19902) ) ;
INV     gate6982  (.A(g15885), .Z(g19905) ) ;
INV     gate6983  (.A(g16540), .Z(g19908) ) ;
INV     gate6984  (.A(g17328), .Z(g19912) ) ;
INV     gate6985  (.A(g16349), .Z(g19915) ) ;
INV     gate6986  (.A(g17200), .Z(g19930) ) ;
INV     gate6987  (.A(g17200), .Z(g19931) ) ;
INV     gate6988  (.A(g17226), .Z(g19947) ) ;
INV     gate6989  (.A(g15885), .Z(g19950) ) ;
INV     gate6990  (.A(g15915), .Z(g19952) ) ;
INV     gate6991  (.A(g16540), .Z(g19954) ) ;
INV     gate6992  (.A(g16540), .Z(g19957) ) ;
INV     gate6993  (.A(g17433), .Z(g19960) ) ;
INV     gate6994  (.A(g17328), .Z(g19961) ) ;
INV     gate6995  (.A(g16326), .Z(g19963) ) ;
INV     gate6996  (.A(g17200), .Z(g19964) ) ;
INV     gate6997  (.A(g17226), .Z(g19979) ) ;
INV     gate6998  (.A(g17226), .Z(g19980) ) ;
INV     gate6999  (.A(g17271), .Z(g19996) ) ;
INV     gate7000  (.A(g15915), .Z(g19998) ) ;
INV     gate7001  (.A(g17249), .Z(g20004) ) ;
INV     gate7002  (.A(g17433), .Z(g20005) ) ;
INV     gate7003  (.A(g17328), .Z(g20006) ) ;
INV     gate7004  (.A(g16449), .Z(g20008) ) ;
INV     gate7005  (.A(g16349), .Z(g20009) ) ;
INV     gate7006  (.A(g17226), .Z(g20010) ) ;
INV     gate7007  (.A(g17271), .Z(g20025) ) ;
INV     gate7008  (.A(g17271), .Z(g20026) ) ;
INV     gate7009  (.A(g15371), .Z(g20028) ) ;
INV     gate7010  (.A(g16579), .Z(g20033) ) ;
OR2     gate7011  (.A(g182), .B(g13657), .Z(g16430) ) ;
INV     gate7012  (.A(g16430), .Z(g20035) ) ;
INV     gate7013  (.A(g17433), .Z(g20036) ) ;
INV     gate7014  (.A(g17328), .Z(g20037) ) ;
INV     gate7015  (.A(g17328), .Z(g20038) ) ;
INV     gate7016  (.A(g17271), .Z(g20040) ) ;
INV     gate7017  (.A(g15569), .Z(g20041) ) ;
INV     gate7018  (.A(g16540), .Z(g20046) ) ;
INV     gate7019  (.A(g16920), .Z(II20318) ) ;
INV     gate7020  (.A(g16920), .Z(II20321) ) ;
INV     gate7021  (.A(II20321), .Z(g20050) ) ;
INV     gate7022  (.A(g17533), .Z(g20052) ) ;
INV     gate7023  (.A(g17328), .Z(g20053) ) ;
INV     gate7024  (.A(g17328), .Z(g20054) ) ;
INV     gate7025  (.A(g16349), .Z(g20057) ) ;
INV     gate7026  (.A(g16782), .Z(g20058) ) ;
INV     gate7027  (.A(g17302), .Z(g20059) ) ;
INV     gate7028  (.A(g16540), .Z(g20060) ) ;
INV     gate7029  (.A(g17533), .Z(g20064) ) ;
AND3    gate7030  (.A(g14034), .B(g12591), .C(g11185), .Z(g16846) ) ;
INV     gate7031  (.A(g16846), .Z(g20065) ) ;
INV     gate7032  (.A(g17433), .Z(g20066) ) ;
INV     gate7033  (.A(g17328), .Z(g20067) ) ;
OR2     gate7034  (.A(g8796), .B(g13464), .Z(g16173) ) ;
INV     gate7035  (.A(g16173), .Z(g20070) ) ;
INV     gate7036  (.A(g16826), .Z(g20071) ) ;
INV     gate7037  (.A(g17384), .Z(g20072) ) ;
INV     gate7038  (.A(g16540), .Z(g20073) ) ;
INV     gate7039  (.A(g16846), .Z(g20078) ) ;
INV     gate7040  (.A(g17328), .Z(g20079) ) ;
INV     gate7041  (.A(g17328), .Z(g20080) ) ;
OR2     gate7042  (.A(g8822), .B(g13486), .Z(g16187) ) ;
INV     gate7043  (.A(g16187), .Z(g20085) ) ;
AND4    gate7044  (.A(g11547), .B(g11592), .C(g11640), .D(II18568), .Z(g17613) ) ;
INV     gate7045  (.A(g17613), .Z(II20355) ) ;
INV     gate7046  (.A(II20355), .Z(g20086) ) ;
INV     gate7047  (.A(g17249), .Z(g20087) ) ;
INV     gate7048  (.A(g17533), .Z(g20088) ) ;
INV     gate7049  (.A(g17533), .Z(g20089) ) ;
INV     gate7050  (.A(g17433), .Z(g20090) ) ;
INV     gate7051  (.A(g17328), .Z(g20091) ) ;
INV     gate7052  (.A(g16782), .Z(g20096) ) ;
INV     gate7053  (.A(g17691), .Z(g20097) ) ;
AND4    gate7054  (.A(g11547), .B(g11592), .C(g11640), .D(II18671), .Z(g17690) ) ;
INV     gate7055  (.A(g17690), .Z(II20369) ) ;
INV     gate7056  (.A(II20369), .Z(g20100) ) ;
INV     gate7057  (.A(g17533), .Z(g20101) ) ;
INV     gate7058  (.A(g17533), .Z(g20102) ) ;
INV     gate7059  (.A(g17433), .Z(g20103) ) ;
INV     gate7060  (.A(g17433), .Z(g20104) ) ;
INV     gate7061  (.A(g17433), .Z(g20105) ) ;
INV     gate7062  (.A(g17328), .Z(g20106) ) ;
INV     gate7063  (.A(g16897), .Z(g20110) ) ;
INV     gate7064  (.A(g16826), .Z(g20113) ) ;
AND4    gate7065  (.A(g11547), .B(g6782), .C(g11640), .D(II17529), .Z(g16194) ) ;
INV     gate7066  (.A(g16194), .Z(II20385) ) ;
INV     gate7067  (.A(II20385), .Z(g20114) ) ;
AND4    gate7068  (.A(g11547), .B(g11592), .C(g11640), .D(II18713), .Z(g17724) ) ;
INV     gate7069  (.A(g17724), .Z(II20388) ) ;
INV     gate7070  (.A(II20388), .Z(g20127) ) ;
INV     gate7071  (.A(g17533), .Z(g20128) ) ;
INV     gate7072  (.A(g17328), .Z(g20129) ) ;
INV     gate7073  (.A(g17328), .Z(g20130) ) ;
INV     gate7074  (.A(g16931), .Z(g20132) ) ;
AND4    gate7075  (.A(g11547), .B(g6782), .C(g11640), .D(II17542), .Z(g16205) ) ;
INV     gate7076  (.A(g16205), .Z(II20399) ) ;
INV     gate7077  (.A(II20399), .Z(g20136) ) ;
INV     gate7078  (.A(g17533), .Z(g20144) ) ;
INV     gate7079  (.A(g17533), .Z(g20145) ) ;
INV     gate7080  (.A(g17533), .Z(g20146) ) ;
INV     gate7081  (.A(g17328), .Z(g20147) ) ;
INV     gate7082  (.A(g16782), .Z(g20153) ) ;
AND4    gate7083  (.A(g6772), .B(g6782), .C(g11640), .D(II17552), .Z(g16213) ) ;
INV     gate7084  (.A(g16213), .Z(II20412) ) ;
INV     gate7085  (.A(II20412), .Z(g20154) ) ;
INV     gate7086  (.A(g16886), .Z(g20157) ) ;
INV     gate7087  (.A(g16971), .Z(g20158) ) ;
INV     gate7088  (.A(g17533), .Z(g20159) ) ;
INV     gate7089  (.A(g16826), .Z(g20164) ) ;
INV     gate7090  (.A(g16886), .Z(g20166) ) ;
INV     gate7091  (.A(g16971), .Z(g20167) ) ;
INV     gate7092  (.A(g17533), .Z(g20168) ) ;
AND4    gate7093  (.A(g6772), .B(g6782), .C(g11640), .D(II17575), .Z(g16234) ) ;
INV     gate7094  (.A(g16234), .Z(II20433) ) ;
INV     gate7095  (.A(II20433), .Z(g20175) ) ;
INV     gate7096  (.A(g16971), .Z(g20178) ) ;
INV     gate7097  (.A(g17249), .Z(g20179) ) ;
INV     gate7098  (.A(g17533), .Z(g20180) ) ;
INV     gate7099  (.A(g16897), .Z(g20182) ) ;
AND4    gate7100  (.A(g11547), .B(g11592), .C(g6789), .D(II17585), .Z(g16244) ) ;
INV     gate7101  (.A(g16244), .Z(II20447) ) ;
INV     gate7102  (.A(II20447), .Z(g20189) ) ;
INV     gate7103  (.A(g16971), .Z(g20190) ) ;
INV     gate7104  (.A(g17821), .Z(g20191) ) ;
OR2     gate7105  (.A(g9220), .B(g14387), .Z(g17268) ) ;
INV     gate7106  (.A(g17268), .Z(g20192) ) ;
INV     gate7107  (.A(g16897), .Z(g20194) ) ;
INV     gate7108  (.A(g16931), .Z(g20195) ) ;
INV     gate7109  (.A(g16987), .Z(g20197) ) ;
INV     gate7110  (.A(g16578), .Z(g20204) ) ;
INV     gate7111  (.A(g17015), .Z(g20207) ) ;
INV     gate7112  (.A(g17533), .Z(g20208) ) ;
INV     gate7113  (.A(g17821), .Z(g20209) ) ;
INV     gate7114  (.A(g16897), .Z(g20210) ) ;
INV     gate7115  (.A(g16931), .Z(g20211) ) ;
NOR2    gate7116  (.A(g11039), .B(g13480), .Z(g17194) ) ;
INV     gate7117  (.A(g17194), .Z(g20212) ) ;
INV     gate7118  (.A(g17062), .Z(g20213) ) ;
AND4    gate7119  (.A(g11547), .B(g11592), .C(g6789), .D(II17606), .Z(g16283) ) ;
INV     gate7120  (.A(g16283), .Z(II20495) ) ;
INV     gate7121  (.A(II20495), .Z(g20219) ) ;
INV     gate7122  (.A(g17015), .Z(g20229) ) ;
AND2    gate7123  (.A(g14583), .B(g14232), .Z(g16224) ) ;
INV     gate7124  (.A(g16224), .Z(II20499) ) ;
INV     gate7125  (.A(II20499), .Z(g20230) ) ;
INV     gate7126  (.A(g17821), .Z(g20231) ) ;
INV     gate7127  (.A(g16931), .Z(g20232) ) ;
INV     gate7128  (.A(g17873), .Z(g20233) ) ;
INV     gate7129  (.A(g15277), .Z(g20235) ) ;
NOR2    gate7130  (.A(g11107), .B(g13501), .Z(g17213) ) ;
INV     gate7131  (.A(g17213), .Z(g20237) ) ;
INV     gate7132  (.A(g17096), .Z(g20238) ) ;
INV     gate7133  (.A(g17128), .Z(g20239) ) ;
INV     gate7134  (.A(g17847), .Z(g20240) ) ;
INV     gate7135  (.A(g16308), .Z(g20242) ) ;
INV     gate7136  (.A(g17015), .Z(g20247) ) ;
INV     gate7137  (.A(g17821), .Z(g20265) ) ;
INV     gate7138  (.A(g17873), .Z(g20266) ) ;
INV     gate7139  (.A(g17955), .Z(g20267) ) ;
INV     gate7140  (.A(g18008), .Z(g20268) ) ;
NAND3   gate7141  (.A(g14714), .B(g9340), .C(g12378), .Z(g15844) ) ;
INV     gate7142  (.A(g15844), .Z(g20269) ) ;
INV     gate7143  (.A(g15277), .Z(g20270) ) ;
NOR2    gate7144  (.A(g11119), .B(g13518), .Z(g17239) ) ;
INV     gate7145  (.A(g17239), .Z(g20272) ) ;
INV     gate7146  (.A(g17128), .Z(g20273) ) ;
INV     gate7147  (.A(g17847), .Z(g20274) ) ;
INV     gate7148  (.A(g17929), .Z(g20275) ) ;
INV     gate7149  (.A(g16487), .Z(g20277) ) ;
INV     gate7150  (.A(g16309), .Z(II20529) ) ;
INV     gate7151  (.A(II20529), .Z(g20283) ) ;
INV     gate7152  (.A(g17015), .Z(g20320) ) ;
INV     gate7153  (.A(g17821), .Z(g20321) ) ;
INV     gate7154  (.A(g17873), .Z(g20322) ) ;
INV     gate7155  (.A(g17873), .Z(g20323) ) ;
INV     gate7156  (.A(g17955), .Z(g20324) ) ;
INV     gate7157  (.A(g15171), .Z(g20325) ) ;
INV     gate7158  (.A(g18008), .Z(g20326) ) ;
INV     gate7159  (.A(g15224), .Z(g20327) ) ;
NAND3   gate7160  (.A(g14714), .B(g9417), .C(g9340), .Z(g15867) ) ;
INV     gate7161  (.A(g15867), .Z(g20328) ) ;
INV     gate7162  (.A(g15277), .Z(g20329) ) ;
INV     gate7163  (.A(g16508), .Z(II20542) ) ;
INV     gate7164  (.A(II20542), .Z(g20330) ) ;
INV     gate7165  (.A(g17847), .Z(g20372) ) ;
INV     gate7166  (.A(g17929), .Z(g20373) ) ;
INV     gate7167  (.A(g18065), .Z(g20374) ) ;
INV     gate7168  (.A(g17821), .Z(g20379) ) ;
INV     gate7169  (.A(g17955), .Z(g20380) ) ;
INV     gate7170  (.A(g17955), .Z(g20381) ) ;
INV     gate7171  (.A(g15171), .Z(g20382) ) ;
INV     gate7172  (.A(g15373), .Z(g20383) ) ;
INV     gate7173  (.A(g18008), .Z(g20384) ) ;
INV     gate7174  (.A(g18008), .Z(g20385) ) ;
INV     gate7175  (.A(g15224), .Z(g20386) ) ;
INV     gate7176  (.A(g15426), .Z(g20387) ) ;
NAND2   gate7177  (.A(g2729), .B(g14291), .Z(g17297) ) ;
INV     gate7178  (.A(g17297), .Z(g20388) ) ;
INV     gate7179  (.A(g15277), .Z(g20389) ) ;
INV     gate7180  (.A(g16525), .Z(II20562) ) ;
INV     gate7181  (.A(II20562), .Z(g20391) ) ;
INV     gate7182  (.A(g17847), .Z(g20432) ) ;
INV     gate7183  (.A(g17929), .Z(g20433) ) ;
INV     gate7184  (.A(g18065), .Z(g20434) ) ;
INV     gate7185  (.A(g15348), .Z(g20435) ) ;
AND4    gate7186  (.A(g6772), .B(g11592), .C(g6789), .D(II17692), .Z(g16486) ) ;
INV     gate7187  (.A(g16486), .Z(II20569) ) ;
INV     gate7188  (.A(II20569), .Z(g20436) ) ;
INV     gate7189  (.A(g17873), .Z(g20441) ) ;
INV     gate7190  (.A(g15171), .Z(g20442) ) ;
INV     gate7191  (.A(g15171), .Z(g20443) ) ;
INV     gate7192  (.A(g15373), .Z(g20444) ) ;
INV     gate7193  (.A(g15224), .Z(g20445) ) ;
INV     gate7194  (.A(g15224), .Z(g20446) ) ;
INV     gate7195  (.A(g15426), .Z(g20447) ) ;
INV     gate7196  (.A(g15509), .Z(g20448) ) ;
INV     gate7197  (.A(g15277), .Z(g20449) ) ;
INV     gate7198  (.A(g15277), .Z(g20450) ) ;
INV     gate7199  (.A(g15277), .Z(g20451) ) ;
INV     gate7200  (.A(g17200), .Z(g20452) ) ;
INV     gate7201  (.A(g16587), .Z(II20584) ) ;
INV     gate7202  (.A(II20584), .Z(g20453) ) ;
INV     gate7203  (.A(g17847), .Z(g20494) ) ;
INV     gate7204  (.A(g17926), .Z(g20495) ) ;
INV     gate7205  (.A(g17929), .Z(g20496) ) ;
INV     gate7206  (.A(g18065), .Z(g20497) ) ;
INV     gate7207  (.A(g15348), .Z(g20498) ) ;
INV     gate7208  (.A(g15483), .Z(g20499) ) ;
INV     gate7209  (.A(g17873), .Z(g20500) ) ;
INV     gate7210  (.A(g17955), .Z(g20501) ) ;
INV     gate7211  (.A(g15373), .Z(g20502) ) ;
INV     gate7212  (.A(g15373), .Z(g20503) ) ;
INV     gate7213  (.A(g18008), .Z(g20504) ) ;
INV     gate7214  (.A(g15426), .Z(g20505) ) ;
INV     gate7215  (.A(g15426), .Z(g20506) ) ;
INV     gate7216  (.A(g15509), .Z(g20507) ) ;
INV     gate7217  (.A(g15277), .Z(g20508) ) ;
INV     gate7218  (.A(g15277), .Z(g20509) ) ;
INV     gate7219  (.A(g17226), .Z(g20510) ) ;
INV     gate7220  (.A(g17929), .Z(g20511) ) ;
INV     gate7221  (.A(g18062), .Z(g20512) ) ;
INV     gate7222  (.A(g18065), .Z(g20513) ) ;
INV     gate7223  (.A(g15348), .Z(g20514) ) ;
INV     gate7224  (.A(g15483), .Z(g20515) ) ;
AND4    gate7225  (.A(g11547), .B(g6782), .C(g6789), .D(II17741), .Z(g16539) ) ;
INV     gate7226  (.A(g16539), .Z(II20609) ) ;
INV     gate7227  (.A(II20609), .Z(g20516) ) ;
INV     gate7228  (.A(g17821), .Z(g20523) ) ;
INV     gate7229  (.A(g17873), .Z(g20524) ) ;
INV     gate7230  (.A(g17955), .Z(g20525) ) ;
INV     gate7231  (.A(g15171), .Z(g20526) ) ;
INV     gate7232  (.A(g18008), .Z(g20527) ) ;
INV     gate7233  (.A(g15224), .Z(g20528) ) ;
INV     gate7234  (.A(g15509), .Z(g20529) ) ;
INV     gate7235  (.A(g15509), .Z(g20530) ) ;
NAND3   gate7236  (.A(g14833), .B(g9417), .C(g12487), .Z(g15907) ) ;
INV     gate7237  (.A(g15907), .Z(g20531) ) ;
INV     gate7238  (.A(g15277), .Z(g20532) ) ;
INV     gate7239  (.A(g17271), .Z(g20533) ) ;
INV     gate7240  (.A(g17183), .Z(g20534) ) ;
INV     gate7241  (.A(g17847), .Z(g20535) ) ;
INV     gate7242  (.A(g18065), .Z(g20536) ) ;
INV     gate7243  (.A(g15345), .Z(g20537) ) ;
INV     gate7244  (.A(g15348), .Z(g20538) ) ;
INV     gate7245  (.A(g15483), .Z(g20539) ) ;
NOR3    gate7246  (.A(g13437), .B(g11020), .C(g11372), .Z(g16646) ) ;
INV     gate7247  (.A(g16646), .Z(g20540) ) ;
INV     gate7248  (.A(g17821), .Z(g20541) ) ;
INV     gate7249  (.A(g17873), .Z(g20542) ) ;
INV     gate7250  (.A(g17955), .Z(g20543) ) ;
INV     gate7251  (.A(g15171), .Z(g20544) ) ;
INV     gate7252  (.A(g15373), .Z(g20545) ) ;
INV     gate7253  (.A(g18008), .Z(g20546) ) ;
INV     gate7254  (.A(g15224), .Z(g20547) ) ;
INV     gate7255  (.A(g15426), .Z(g20548) ) ;
INV     gate7256  (.A(g15277), .Z(g20549) ) ;
NAND3   gate7257  (.A(g14833), .B(g12543), .C(g12487), .Z(g15864) ) ;
INV     gate7258  (.A(g15864), .Z(g20550) ) ;
INV     gate7259  (.A(g17302), .Z(g20551) ) ;
INV     gate7260  (.A(g17847), .Z(g20552) ) ;
INV     gate7261  (.A(g17929), .Z(g20553) ) ;
INV     gate7262  (.A(g15348), .Z(g20554) ) ;
INV     gate7263  (.A(g15480), .Z(g20555) ) ;
INV     gate7264  (.A(g15483), .Z(g20556) ) ;
INV     gate7265  (.A(g17010), .Z(II20647) ) ;
INV     gate7266  (.A(g17010), .Z(II20650) ) ;
INV     gate7267  (.A(II20650), .Z(g20558) ) ;
INV     gate7268  (.A(g17328), .Z(g20560) ) ;
INV     gate7269  (.A(g17873), .Z(g20561) ) ;
INV     gate7270  (.A(g17955), .Z(g20562) ) ;
INV     gate7271  (.A(g15171), .Z(g20563) ) ;
INV     gate7272  (.A(g15373), .Z(g20564) ) ;
INV     gate7273  (.A(g18008), .Z(g20565) ) ;
INV     gate7274  (.A(g15224), .Z(g20566) ) ;
INV     gate7275  (.A(g15426), .Z(g20567) ) ;
INV     gate7276  (.A(g15509), .Z(g20568) ) ;
INV     gate7277  (.A(g15277), .Z(g20569) ) ;
INV     gate7278  (.A(g15277), .Z(g20570) ) ;
INV     gate7279  (.A(g15277), .Z(g20571) ) ;
NAND3   gate7280  (.A(g14714), .B(g12378), .C(g12337), .Z(g15833) ) ;
INV     gate7281  (.A(g15833), .Z(g20572) ) ;
INV     gate7282  (.A(g17384), .Z(g20573) ) ;
INV     gate7283  (.A(g17847), .Z(g20574) ) ;
INV     gate7284  (.A(g17929), .Z(g20575) ) ;
INV     gate7285  (.A(g18065), .Z(g20576) ) ;
INV     gate7286  (.A(g15483), .Z(g20577) ) ;
INV     gate7287  (.A(g15563), .Z(g20578) ) ;
INV     gate7288  (.A(g17249), .Z(g20579) ) ;
INV     gate7289  (.A(g17328), .Z(g20580) ) ;
INV     gate7290  (.A(g17873), .Z(g20582) ) ;
INV     gate7291  (.A(g17873), .Z(g20583) ) ;
INV     gate7292  (.A(g17873), .Z(g20584) ) ;
INV     gate7293  (.A(g17955), .Z(g20585) ) ;
INV     gate7294  (.A(g15171), .Z(g20586) ) ;
INV     gate7295  (.A(g15373), .Z(g20587) ) ;
INV     gate7296  (.A(g18008), .Z(g20588) ) ;
INV     gate7297  (.A(g15224), .Z(g20589) ) ;
INV     gate7298  (.A(g15426), .Z(g20590) ) ;
INV     gate7299  (.A(g15509), .Z(g20591) ) ;
INV     gate7300  (.A(g15277), .Z(g20592) ) ;
INV     gate7301  (.A(g15277), .Z(g20593) ) ;
INV     gate7302  (.A(g15277), .Z(g20594) ) ;
NAND3   gate7303  (.A(g14833), .B(g9340), .C(g12543), .Z(g15877) ) ;
INV     gate7304  (.A(g15877), .Z(g20595) ) ;
INV     gate7305  (.A(g15733), .Z(II20690) ) ;
INV     gate7306  (.A(II20690), .Z(g20596) ) ;
INV     gate7307  (.A(g17847), .Z(g20597) ) ;
INV     gate7308  (.A(g17929), .Z(g20598) ) ;
INV     gate7309  (.A(g18065), .Z(g20599) ) ;
INV     gate7310  (.A(g15348), .Z(g20600) ) ;
INV     gate7311  (.A(g17433), .Z(g20601) ) ;
INV     gate7312  (.A(g17873), .Z(g20603) ) ;
INV     gate7313  (.A(g17873), .Z(g20604) ) ;
INV     gate7314  (.A(g17955), .Z(g20605) ) ;
INV     gate7315  (.A(g17955), .Z(g20606) ) ;
INV     gate7316  (.A(g17955), .Z(g20607) ) ;
INV     gate7317  (.A(g15171), .Z(g20608) ) ;
INV     gate7318  (.A(g15373), .Z(g20609) ) ;
INV     gate7319  (.A(g18008), .Z(g20610) ) ;
INV     gate7320  (.A(g18008), .Z(g20611) ) ;
INV     gate7321  (.A(g18008), .Z(g20612) ) ;
INV     gate7322  (.A(g15224), .Z(g20613) ) ;
INV     gate7323  (.A(g15426), .Z(g20614) ) ;
INV     gate7324  (.A(g15509), .Z(g20615) ) ;
INV     gate7325  (.A(g15277), .Z(g20616) ) ;
INV     gate7326  (.A(g15277), .Z(g20617) ) ;
INV     gate7327  (.A(g15277), .Z(g20618) ) ;
INV     gate7328  (.A(g15595), .Z(g20622) ) ;
INV     gate7329  (.A(g17929), .Z(g20623) ) ;
INV     gate7330  (.A(g18065), .Z(g20624) ) ;
INV     gate7331  (.A(g15348), .Z(g20625) ) ;
INV     gate7332  (.A(g15483), .Z(g20626) ) ;
INV     gate7333  (.A(g17433), .Z(g20627) ) ;
INV     gate7334  (.A(g17955), .Z(g20629) ) ;
INV     gate7335  (.A(g17955), .Z(g20630) ) ;
INV     gate7336  (.A(g15171), .Z(g20631) ) ;
INV     gate7337  (.A(g15171), .Z(g20632) ) ;
INV     gate7338  (.A(g15171), .Z(g20633) ) ;
INV     gate7339  (.A(g15373), .Z(g20634) ) ;
INV     gate7340  (.A(g18008), .Z(g20635) ) ;
INV     gate7341  (.A(g18008), .Z(g20636) ) ;
INV     gate7342  (.A(g15224), .Z(g20637) ) ;
INV     gate7343  (.A(g15224), .Z(g20638) ) ;
INV     gate7344  (.A(g15224), .Z(g20639) ) ;
INV     gate7345  (.A(g15426), .Z(g20640) ) ;
INV     gate7346  (.A(g15509), .Z(g20641) ) ;
INV     gate7347  (.A(g15277), .Z(g20642) ) ;
NAND3   gate7348  (.A(g14833), .B(g9417), .C(g9340), .Z(g15962) ) ;
INV     gate7349  (.A(g15962), .Z(g20643) ) ;
INV     gate7350  (.A(g15615), .Z(g20648) ) ;
INV     gate7351  (.A(g18065), .Z(g20649) ) ;
INV     gate7352  (.A(g15348), .Z(g20650) ) ;
INV     gate7353  (.A(g15483), .Z(g20651) ) ;
INV     gate7354  (.A(g17141), .Z(II20744) ) ;
INV     gate7355  (.A(g17141), .Z(II20747) ) ;
INV     gate7356  (.A(II20747), .Z(g20653) ) ;
INV     gate7357  (.A(g16677), .Z(II20750) ) ;
INV     gate7358  (.A(g16677), .Z(II20753) ) ;
INV     gate7359  (.A(II20753), .Z(g20655) ) ;
INV     gate7360  (.A(g17249), .Z(g20656) ) ;
INV     gate7361  (.A(g17433), .Z(g20657) ) ;
INV     gate7362  (.A(g17873), .Z(g20659) ) ;
INV     gate7363  (.A(g17873), .Z(g20660) ) ;
INV     gate7364  (.A(g15171), .Z(g20661) ) ;
INV     gate7365  (.A(g15171), .Z(g20662) ) ;
INV     gate7366  (.A(g15373), .Z(g20663) ) ;
INV     gate7367  (.A(g15373), .Z(g20664) ) ;
INV     gate7368  (.A(g15373), .Z(g20665) ) ;
INV     gate7369  (.A(g15224), .Z(g20666) ) ;
INV     gate7370  (.A(g15224), .Z(g20667) ) ;
INV     gate7371  (.A(g15426), .Z(g20668) ) ;
INV     gate7372  (.A(g15426), .Z(g20669) ) ;
INV     gate7373  (.A(g15426), .Z(g20670) ) ;
INV     gate7374  (.A(g15509), .Z(g20671) ) ;
INV     gate7375  (.A(g15277), .Z(g20672) ) ;
INV     gate7376  (.A(g15277), .Z(g20673) ) ;
INV     gate7377  (.A(g15277), .Z(g20674) ) ;
INV     gate7378  (.A(g15634), .Z(g20679) ) ;
INV     gate7379  (.A(g15348), .Z(g20680) ) ;
INV     gate7380  (.A(g15483), .Z(g20681) ) ;
INV     gate7381  (.A(g17155), .Z(II20781) ) ;
INV     gate7382  (.A(II20781), .Z(g20695) ) ;
INV     gate7383  (.A(g17533), .Z(g20696) ) ;
INV     gate7384  (.A(g17433), .Z(g20697) ) ;
INV     gate7385  (.A(g17873), .Z(g20698) ) ;
INV     gate7386  (.A(g17873), .Z(g20699) ) ;
INV     gate7387  (.A(g17873), .Z(g20700) ) ;
INV     gate7388  (.A(g17955), .Z(g20701) ) ;
INV     gate7389  (.A(g17955), .Z(g20702) ) ;
INV     gate7390  (.A(g15373), .Z(g20703) ) ;
INV     gate7391  (.A(g15373), .Z(g20704) ) ;
NOR2    gate7392  (.A(g12435), .B(g12955), .Z(g17694) ) ;
INV     gate7393  (.A(g17694), .Z(II20793) ) ;
INV     gate7394  (.A(II20793), .Z(g20705) ) ;
INV     gate7395  (.A(g18008), .Z(g20706) ) ;
INV     gate7396  (.A(g18008), .Z(g20707) ) ;
INV     gate7397  (.A(g15426), .Z(g20708) ) ;
INV     gate7398  (.A(g15426), .Z(g20709) ) ;
INV     gate7399  (.A(g15509), .Z(g20710) ) ;
INV     gate7400  (.A(g15509), .Z(g20711) ) ;
INV     gate7401  (.A(g15509), .Z(g20712) ) ;
INV     gate7402  (.A(g15277), .Z(g20713) ) ;
INV     gate7403  (.A(g15277), .Z(g20714) ) ;
INV     gate7404  (.A(g15277), .Z(g20715) ) ;
INV     gate7405  (.A(g15277), .Z(g20716) ) ;
INV     gate7406  (.A(g15595), .Z(g20732) ) ;
INV     gate7407  (.A(g15656), .Z(g20737) ) ;
INV     gate7408  (.A(g15483), .Z(g20738) ) ;
INV     gate7409  (.A(g17088), .Z(II20816) ) ;
INV     gate7410  (.A(g17088), .Z(II20819) ) ;
INV     gate7411  (.A(II20819), .Z(g20764) ) ;
NAND3   gate7412  (.A(g562), .B(g14708), .C(g12323), .Z(g17748) ) ;
INV     gate7413  (.A(g17748), .Z(g20765) ) ;
INV     gate7414  (.A(g17433), .Z(g20766) ) ;
INV     gate7415  (.A(g17873), .Z(g20767) ) ;
INV     gate7416  (.A(g17955), .Z(g20768) ) ;
INV     gate7417  (.A(g17955), .Z(g20769) ) ;
INV     gate7418  (.A(g17955), .Z(g20770) ) ;
INV     gate7419  (.A(g15171), .Z(g20771) ) ;
INV     gate7420  (.A(g15171), .Z(g20772) ) ;
NOR2    gate7421  (.A(g14751), .B(g12955), .Z(g17657) ) ;
INV     gate7422  (.A(g17657), .Z(II20830) ) ;
INV     gate7423  (.A(II20830), .Z(g20773) ) ;
INV     gate7424  (.A(g18008), .Z(g20774) ) ;
INV     gate7425  (.A(g18008), .Z(g20775) ) ;
INV     gate7426  (.A(g18008), .Z(g20776) ) ;
INV     gate7427  (.A(g15224), .Z(g20777) ) ;
INV     gate7428  (.A(g15224), .Z(g20778) ) ;
INV     gate7429  (.A(g15509), .Z(g20779) ) ;
INV     gate7430  (.A(g15509), .Z(g20780) ) ;
NOR2    gate7431  (.A(g12486), .B(g12983), .Z(g17727) ) ;
INV     gate7432  (.A(g17727), .Z(II20840) ) ;
INV     gate7433  (.A(II20840), .Z(g20781) ) ;
NAND3   gate7434  (.A(g14714), .B(g9417), .C(g12337), .Z(g15853) ) ;
INV     gate7435  (.A(g15853), .Z(g20782) ) ;
INV     gate7436  (.A(g16923), .Z(II20846) ) ;
INV     gate7437  (.A(II20846), .Z(g20785) ) ;
INV     gate7438  (.A(g15595), .Z(g20852) ) ;
INV     gate7439  (.A(g15595), .Z(g20853) ) ;
INV     gate7440  (.A(g15615), .Z(g20869) ) ;
INV     gate7441  (.A(g15680), .Z(g20874) ) ;
INV     gate7442  (.A(g16960), .Z(II20861) ) ;
INV     gate7443  (.A(g16960), .Z(II20864) ) ;
INV     gate7444  (.A(II20864), .Z(g20900) ) ;
INV     gate7445  (.A(g16216), .Z(II20867) ) ;
INV     gate7446  (.A(g16216), .Z(II20870) ) ;
INV     gate7447  (.A(II20870), .Z(g20902) ) ;
INV     gate7448  (.A(g17249), .Z(g20903) ) ;
INV     gate7449  (.A(g17433), .Z(g20904) ) ;
INV     gate7450  (.A(g17955), .Z(g20909) ) ;
INV     gate7451  (.A(g15171), .Z(g20910) ) ;
INV     gate7452  (.A(g15171), .Z(g20911) ) ;
INV     gate7453  (.A(g15171), .Z(g20912) ) ;
INV     gate7454  (.A(g15373), .Z(g20913) ) ;
INV     gate7455  (.A(g15373), .Z(g20914) ) ;
NOR2    gate7456  (.A(g10179), .B(g12955), .Z(g17619) ) ;
INV     gate7457  (.A(g17619), .Z(II20882) ) ;
INV     gate7458  (.A(II20882), .Z(g20915) ) ;
INV     gate7459  (.A(g18008), .Z(g20916) ) ;
INV     gate7460  (.A(g15224), .Z(g20917) ) ;
INV     gate7461  (.A(g15224), .Z(g20918) ) ;
INV     gate7462  (.A(g15224), .Z(g20919) ) ;
INV     gate7463  (.A(g15426), .Z(g20920) ) ;
INV     gate7464  (.A(g15426), .Z(g20921) ) ;
NOR2    gate7465  (.A(g14792), .B(g12983), .Z(g17700) ) ;
INV     gate7466  (.A(g17700), .Z(II20891) ) ;
INV     gate7467  (.A(II20891), .Z(g20922) ) ;
INV     gate7468  (.A(g15277), .Z(g20923) ) ;
INV     gate7469  (.A(g16954), .Z(II20895) ) ;
INV     gate7470  (.A(II20895), .Z(g20924) ) ;
INV     gate7471  (.A(g15595), .Z(g20978) ) ;
INV     gate7472  (.A(g15615), .Z(g20993) ) ;
INV     gate7473  (.A(g15615), .Z(g20994) ) ;
INV     gate7474  (.A(g15634), .Z(g21010) ) ;
INV     gate7475  (.A(g17197), .Z(II20910) ) ;
INV     gate7476  (.A(II20910), .Z(g21036) ) ;
INV     gate7477  (.A(g16964), .Z(II20913) ) ;
INV     gate7478  (.A(II20913), .Z(g21037) ) ;
INV     gate7479  (.A(g17533), .Z(g21048) ) ;
INV     gate7480  (.A(g17433), .Z(g21049) ) ;
INV     gate7481  (.A(g17873), .Z(g21050) ) ;
INV     gate7482  (.A(g15171), .Z(g21051) ) ;
INV     gate7483  (.A(g15373), .Z(g21052) ) ;
INV     gate7484  (.A(g15373), .Z(g21053) ) ;
INV     gate7485  (.A(g15373), .Z(g21054) ) ;
INV     gate7486  (.A(g15224), .Z(g21055) ) ;
INV     gate7487  (.A(g15426), .Z(g21056) ) ;
INV     gate7488  (.A(g15426), .Z(g21057) ) ;
INV     gate7489  (.A(g15426), .Z(g21058) ) ;
INV     gate7490  (.A(g15509), .Z(g21059) ) ;
INV     gate7491  (.A(g15509), .Z(g21060) ) ;
NOR2    gate7492  (.A(g10205), .B(g12983), .Z(g17663) ) ;
INV     gate7493  (.A(g17663), .Z(II20929) ) ;
INV     gate7494  (.A(II20929), .Z(g21061) ) ;
INV     gate7495  (.A(g15277), .Z(g21068) ) ;
INV     gate7496  (.A(g15277), .Z(g21069) ) ;
INV     gate7497  (.A(g16967), .Z(II20937) ) ;
INV     gate7498  (.A(II20937), .Z(g21070) ) ;
INV     gate7499  (.A(g15615), .Z(g21123) ) ;
INV     gate7500  (.A(g15634), .Z(g21138) ) ;
INV     gate7501  (.A(g15634), .Z(g21139) ) ;
INV     gate7502  (.A(g15656), .Z(g21155) ) ;
INV     gate7503  (.A(g17247), .Z(g21156) ) ;
INV     gate7504  (.A(g17508), .Z(g21160) ) ;
INV     gate7505  (.A(g17782), .Z(II20951) ) ;
INV     gate7506  (.A(II20951), .Z(g21175) ) ;
INV     gate7507  (.A(g16228), .Z(II20954) ) ;
INV     gate7508  (.A(g16228), .Z(II20957) ) ;
INV     gate7509  (.A(II20957), .Z(g21177) ) ;
INV     gate7510  (.A(g17955), .Z(g21178) ) ;
INV     gate7511  (.A(g15373), .Z(g21179) ) ;
INV     gate7512  (.A(g18008), .Z(g21180) ) ;
INV     gate7513  (.A(g15426), .Z(g21181) ) ;
INV     gate7514  (.A(g15509), .Z(g21182) ) ;
INV     gate7515  (.A(g15509), .Z(g21183) ) ;
INV     gate7516  (.A(g15509), .Z(g21184) ) ;
INV     gate7517  (.A(g15277), .Z(g21185) ) ;
INV     gate7518  (.A(g15634), .Z(g21189) ) ;
INV     gate7519  (.A(g15656), .Z(g21204) ) ;
INV     gate7520  (.A(g15656), .Z(g21205) ) ;
INV     gate7521  (.A(g15680), .Z(g21221) ) ;
INV     gate7522  (.A(g17430), .Z(g21222) ) ;
INV     gate7523  (.A(g17428), .Z(g21225) ) ;
INV     gate7524  (.A(g17531), .Z(g21228) ) ;
INV     gate7525  (.A(g16300), .Z(II20982) ) ;
INV     gate7526  (.A(g16300), .Z(II20985) ) ;
INV     gate7527  (.A(II20985), .Z(g21246) ) ;
INV     gate7528  (.A(g15171), .Z(g21247) ) ;
INV     gate7529  (.A(g15224), .Z(g21248) ) ;
INV     gate7530  (.A(g15509), .Z(g21249) ) ;
INV     gate7531  (.A(g15656), .Z(g21252) ) ;
INV     gate7532  (.A(g15680), .Z(g21267) ) ;
INV     gate7533  (.A(g15680), .Z(g21268) ) ;
INV     gate7534  (.A(g15506), .Z(g21269) ) ;
INV     gate7535  (.A(g16709), .Z(II20999) ) ;
INV     gate7536  (.A(g16709), .Z(II21002) ) ;
INV     gate7537  (.A(II21002), .Z(g21271) ) ;
INV     gate7538  (.A(g15579), .Z(II21006) ) ;
INV     gate7539  (.A(II21006), .Z(g21273) ) ;
INV     gate7540  (.A(g15373), .Z(g21274) ) ;
INV     gate7541  (.A(g15426), .Z(g21275) ) ;
INV     gate7542  (.A(g15806), .Z(II21013) ) ;
INV     gate7543  (.A(II21013), .Z(g21278) ) ;
INV     gate7544  (.A(g15680), .Z(g21279) ) ;
INV     gate7545  (.A(g16601), .Z(g21280) ) ;
INV     gate7546  (.A(g16286), .Z(g21281) ) ;
INV     gate7547  (.A(g17325), .Z(II21019) ) ;
INV     gate7548  (.A(II21019), .Z(g21282) ) ;
INV     gate7549  (.A(g15509), .Z(g21286) ) ;
INV     gate7550  (.A(g15816), .Z(II21029) ) ;
INV     gate7551  (.A(II21029), .Z(g21290) ) ;
INV     gate7552  (.A(g16620), .Z(g21291) ) ;
INV     gate7553  (.A(g17221), .Z(II21033) ) ;
INV     gate7554  (.A(g17221), .Z(II21036) ) ;
INV     gate7555  (.A(II21036), .Z(g21293) ) ;
INV     gate7556  (.A(g17533), .Z(g21295) ) ;
INV     gate7557  (.A(g15824), .Z(II21042) ) ;
INV     gate7558  (.A(II21042), .Z(g21297) ) ;
INV     gate7559  (.A(g16600), .Z(g21299) ) ;
INV     gate7560  (.A(g17429), .Z(II21047) ) ;
INV     gate7561  (.A(II21047), .Z(g21300) ) ;
INV     gate7562  (.A(g17367), .Z(g21304) ) ;
INV     gate7563  (.A(g15758), .Z(g21305) ) ;
OR2     gate7564  (.A(g8977), .B(g12925), .Z(g15582) ) ;
INV     gate7565  (.A(g15582), .Z(g21306) ) ;
INV     gate7566  (.A(g17485), .Z(g21308) ) ;
AND4    gate7567  (.A(g6772), .B(g11592), .C(g11640), .D(II18740), .Z(g17747) ) ;
INV     gate7568  (.A(g17747), .Z(II21058) ) ;
INV     gate7569  (.A(II21058), .Z(g21326) ) ;
INV     gate7570  (.A(g16577), .Z(g21329) ) ;
INV     gate7571  (.A(g15573), .Z(II21067) ) ;
INV     gate7572  (.A(II21067), .Z(g21335) ) ;
INV     gate7573  (.A(g17367), .Z(g21336) ) ;
INV     gate7574  (.A(g15758), .Z(g21337) ) ;
AND4    gate7575  (.A(g6772), .B(g11592), .C(g11640), .D(II18762), .Z(g17766) ) ;
INV     gate7576  (.A(g17766), .Z(II21074) ) ;
INV     gate7577  (.A(II21074), .Z(g21340) ) ;
INV     gate7578  (.A(g16428), .Z(g21343) ) ;
INV     gate7579  (.A(g17821), .Z(g21346) ) ;
INV     gate7580  (.A(g15758), .Z(g21349) ) ;
INV     gate7581  (.A(g16322), .Z(g21352) ) ;
INV     gate7582  (.A(g17821), .Z(g21355) ) ;
INV     gate7583  (.A(g16307), .Z(g21358) ) ;
INV     gate7584  (.A(g17873), .Z(g21362) ) ;
INV     gate7585  (.A(g16284), .Z(II21100) ) ;
INV     gate7586  (.A(II21100), .Z(g21366) ) ;
INV     gate7587  (.A(g16285), .Z(g21369) ) ;
INV     gate7588  (.A(g16323), .Z(g21370) ) ;
INV     gate7589  (.A(g17873), .Z(g21379) ) ;
INV     gate7590  (.A(g17955), .Z(g21380) ) ;
INV     gate7591  (.A(g18008), .Z(g21381) ) ;
INV     gate7592  (.A(g17367), .Z(g21383) ) ;
INV     gate7593  (.A(g15714), .Z(II21115) ) ;
INV     gate7594  (.A(II21115), .Z(g21387) ) ;
OR2     gate7595  (.A(g7118), .B(g14309), .Z(g17264) ) ;
INV     gate7596  (.A(g17264), .Z(g21393) ) ;
INV     gate7597  (.A(g17873), .Z(g21395) ) ;
INV     gate7598  (.A(g17955), .Z(g21396) ) ;
INV     gate7599  (.A(g15171), .Z(g21397) ) ;
INV     gate7600  (.A(g18008), .Z(g21398) ) ;
INV     gate7601  (.A(g15224), .Z(g21399) ) ;
INV     gate7602  (.A(g17847), .Z(g21400) ) ;
INV     gate7603  (.A(g17955), .Z(g21406) ) ;
INV     gate7604  (.A(g15171), .Z(g21407) ) ;
INV     gate7605  (.A(g15373), .Z(g21408) ) ;
INV     gate7606  (.A(g18008), .Z(g21409) ) ;
INV     gate7607  (.A(g15224), .Z(g21410) ) ;
INV     gate7608  (.A(g15426), .Z(g21411) ) ;
INV     gate7609  (.A(g15758), .Z(g21412) ) ;
NOR2    gate7610  (.A(g11862), .B(g14194), .Z(g15585) ) ;
INV     gate7611  (.A(g15585), .Z(g21413) ) ;
INV     gate7612  (.A(g17929), .Z(g21414) ) ;
INV     gate7613  (.A(g17821), .Z(g21418) ) ;
INV     gate7614  (.A(g15171), .Z(g21421) ) ;
INV     gate7615  (.A(g15373), .Z(g21422) ) ;
INV     gate7616  (.A(g15224), .Z(g21423) ) ;
INV     gate7617  (.A(g15426), .Z(g21424) ) ;
INV     gate7618  (.A(g15509), .Z(g21425) ) ;
INV     gate7619  (.A(g15277), .Z(g21426) ) ;
INV     gate7620  (.A(g17367), .Z(g21427) ) ;
INV     gate7621  (.A(g15758), .Z(g21428) ) ;
NOR2    gate7622  (.A(g11885), .B(g14212), .Z(g15608) ) ;
INV     gate7623  (.A(g15608), .Z(g21430) ) ;
INV     gate7624  (.A(g18065), .Z(g21431) ) ;
INV     gate7625  (.A(g17248), .Z(g21434) ) ;
AND2    gate7626  (.A(g1075), .B(g13093), .Z(g17292) ) ;
INV     gate7627  (.A(g17292), .Z(II21162) ) ;
INV     gate7628  (.A(II21162), .Z(g21451) ) ;
INV     gate7629  (.A(g15373), .Z(g21454) ) ;
INV     gate7630  (.A(g15426), .Z(g21455) ) ;
INV     gate7631  (.A(g15509), .Z(g21456) ) ;
INV     gate7632  (.A(g17367), .Z(g21457) ) ;
INV     gate7633  (.A(g15758), .Z(g21458) ) ;
NOR2    gate7634  (.A(g11907), .B(g14228), .Z(g15628) ) ;
INV     gate7635  (.A(g15628), .Z(g21460) ) ;
INV     gate7636  (.A(g15348), .Z(g21461) ) ;
INV     gate7637  (.A(g15588), .Z(g21463) ) ;
INV     gate7638  (.A(g15509), .Z(g21466) ) ;
INV     gate7639  (.A(g15758), .Z(g21467) ) ;
INV     gate7640  (.A(g17413), .Z(II21181) ) ;
INV     gate7641  (.A(II21181), .Z(g21468) ) ;
NOR2    gate7642  (.A(g11924), .B(g14248), .Z(g15647) ) ;
INV     gate7643  (.A(g15647), .Z(g21510) ) ;
INV     gate7644  (.A(g15483), .Z(g21511) ) ;
INV     gate7645  (.A(g17475), .Z(II21189) ) ;
INV     gate7646  (.A(II21189), .Z(g21514) ) ;
NOR2    gate7647  (.A(g11945), .B(g14272), .Z(g15669) ) ;
INV     gate7648  (.A(g15669), .Z(g21556) ) ;
INV     gate7649  (.A(g17873), .Z(g21560) ) ;
INV     gate7650  (.A(g15595), .Z(g21561) ) ;
INV     gate7651  (.A(g17501), .Z(II21199) ) ;
INV     gate7652  (.A(II21199), .Z(g21562) ) ;
INV     gate7653  (.A(g15938), .Z(g21604) ) ;
INV     gate7654  (.A(g17873), .Z(g21607) ) ;
INV     gate7655  (.A(g17955), .Z(g21608) ) ;
INV     gate7656  (.A(g18008), .Z(g21609) ) ;
INV     gate7657  (.A(g15615), .Z(g21610) ) ;
INV     gate7658  (.A(g17526), .Z(II21210) ) ;
INV     gate7659  (.A(II21210), .Z(g21611) ) ;
INV     gate7660  (.A(g17663), .Z(g21653) ) ;
INV     gate7661  (.A(g17619), .Z(g21654) ) ;
INV     gate7662  (.A(g17700), .Z(g21656) ) ;
INV     gate7663  (.A(g17657), .Z(g21657) ) ;
INV     gate7664  (.A(g17727), .Z(g21659) ) ;
INV     gate7665  (.A(g17694), .Z(g21660) ) ;
INV     gate7666  (.A(g18091), .Z(II21222) ) ;
INV     gate7667  (.A(II21222), .Z(g21661) ) ;
INV     gate7668  (.A(g16540), .Z(g21662) ) ;
INV     gate7669  (.A(g16540), .Z(II21226) ) ;
INV     gate7670  (.A(II21226), .Z(g21665) ) ;
INV     gate7671  (.A(g16540), .Z(g21666) ) ;
INV     gate7672  (.A(g16540), .Z(II21230) ) ;
INV     gate7673  (.A(II21230), .Z(g21669) ) ;
INV     gate7674  (.A(g16540), .Z(g21670) ) ;
INV     gate7675  (.A(g16540), .Z(II21234) ) ;
INV     gate7676  (.A(II21234), .Z(g21673) ) ;
INV     gate7677  (.A(g16540), .Z(g21674) ) ;
INV     gate7678  (.A(g16540), .Z(II21238) ) ;
INV     gate7679  (.A(II21238), .Z(g21677) ) ;
INV     gate7680  (.A(g16540), .Z(g21678) ) ;
INV     gate7681  (.A(g16540), .Z(II21242) ) ;
INV     gate7682  (.A(II21242), .Z(g21681) ) ;
INV     gate7683  (.A(g16540), .Z(g21682) ) ;
INV     gate7684  (.A(g16540), .Z(II21246) ) ;
INV     gate7685  (.A(II21246), .Z(g21685) ) ;
INV     gate7686  (.A(g16540), .Z(g21686) ) ;
INV     gate7687  (.A(g16540), .Z(II21250) ) ;
INV     gate7688  (.A(II21250), .Z(g21689) ) ;
INV     gate7689  (.A(g16540), .Z(g21690) ) ;
INV     gate7690  (.A(g16540), .Z(II21254) ) ;
INV     gate7691  (.A(II21254), .Z(g21693) ) ;
INV     gate7692  (.A(g16540), .Z(g21694) ) ;
INV     gate7693  (.A(g16540), .Z(II21258) ) ;
INV     gate7694  (.A(II21258), .Z(g21697) ) ;
AND2    gate7695  (.A(g943), .B(g15979), .Z(g18215) ) ;
INV     gate7696  (.A(g18215), .Z(II21285) ) ;
AND2    gate7697  (.A(g967), .B(g15979), .Z(g18216) ) ;
INV     gate7698  (.A(g18216), .Z(II21288) ) ;
AND2    gate7699  (.A(g1287), .B(g16031), .Z(g18273) ) ;
INV     gate7700  (.A(g18273), .Z(II21291) ) ;
AND2    gate7701  (.A(g1311), .B(g16031), .Z(g18274) ) ;
INV     gate7702  (.A(g18274), .Z(II21294) ) ;
AND2    gate7703  (.A(g2975), .B(g16349), .Z(g18597) ) ;
INV     gate7704  (.A(g18597), .Z(II21297) ) ;
AND2    gate7705  (.A(g3003), .B(g16349), .Z(g18598) ) ;
INV     gate7706  (.A(g18598), .Z(II21300) ) ;
AND2    gate7707  (.A(g4737), .B(g16053), .Z(g18695) ) ;
INV     gate7708  (.A(g18695), .Z(II21477) ) ;
AND2    gate7709  (.A(g4741), .B(g16053), .Z(g18696) ) ;
INV     gate7710  (.A(g18696), .Z(II21480) ) ;
AND2    gate7711  (.A(g4927), .B(g16077), .Z(g18726) ) ;
INV     gate7712  (.A(g18726), .Z(II21483) ) ;
AND2    gate7713  (.A(g4931), .B(g16077), .Z(g18727) ) ;
INV     gate7714  (.A(g18727), .Z(II21486) ) ;
INV     gate7715  (.A(g20277), .Z(g22136) ) ;
INV     gate7716  (.A(g21370), .Z(g22137) ) ;
INV     gate7717  (.A(g21370), .Z(g22138) ) ;
INV     gate7718  (.A(g19264), .Z(II21722) ) ;
INV     gate7719  (.A(II21722), .Z(g22139) ) ;
INV     gate7720  (.A(g18997), .Z(g22144) ) ;
INV     gate7721  (.A(g18997), .Z(g22146) ) ;
INV     gate7722  (.A(g18997), .Z(g22147) ) ;
INV     gate7723  (.A(g19074), .Z(g22148) ) ;
INV     gate7724  (.A(g21280), .Z(g22150) ) ;
NOR2    gate7725  (.A(g15979), .B(g962), .Z(g19268) ) ;
INV     gate7726  (.A(g19268), .Z(II21734) ) ;
INV     gate7727  (.A(II21734), .Z(g22151) ) ;
INV     gate7728  (.A(g18997), .Z(g22153) ) ;
INV     gate7729  (.A(g19074), .Z(g22154) ) ;
INV     gate7730  (.A(g19074), .Z(g22155) ) ;
INV     gate7731  (.A(g19147), .Z(g22156) ) ;
NOR2    gate7732  (.A(g16031), .B(g1306), .Z(g19338) ) ;
INV     gate7733  (.A(g19338), .Z(II21744) ) ;
INV     gate7734  (.A(II21744), .Z(g22159) ) ;
INV     gate7735  (.A(g18997), .Z(g22166) ) ;
INV     gate7736  (.A(g19074), .Z(g22167) ) ;
INV     gate7737  (.A(g19147), .Z(g22168) ) ;
INV     gate7738  (.A(g19147), .Z(g22169) ) ;
INV     gate7739  (.A(g19210), .Z(g22170) ) ;
INV     gate7740  (.A(g18882), .Z(g22171) ) ;
INV     gate7741  (.A(g21308), .Z(II21757) ) ;
INV     gate7742  (.A(II21757), .Z(g22173) ) ;
INV     gate7743  (.A(g18997), .Z(g22176) ) ;
INV     gate7744  (.A(g19074), .Z(g22177) ) ;
INV     gate7745  (.A(g19147), .Z(g22178) ) ;
INV     gate7746  (.A(g19210), .Z(g22179) ) ;
INV     gate7747  (.A(g19210), .Z(g22180) ) ;
INV     gate7748  (.A(g19277), .Z(g22181) ) ;
INV     gate7749  (.A(g19620), .Z(II21766) ) ;
INV     gate7750  (.A(II21766), .Z(g22182) ) ;
NOR2    gate7751  (.A(g15979), .B(g13133), .Z(g19402) ) ;
INV     gate7752  (.A(g19402), .Z(II21769) ) ;
INV     gate7753  (.A(II21769), .Z(g22189) ) ;
INV     gate7754  (.A(g19801), .Z(g22192) ) ;
INV     gate7755  (.A(g21308), .Z(II21776) ) ;
INV     gate7756  (.A(II21776), .Z(g22194) ) ;
INV     gate7757  (.A(g19074), .Z(g22197) ) ;
INV     gate7758  (.A(g19147), .Z(g22198) ) ;
INV     gate7759  (.A(g19210), .Z(g22199) ) ;
INV     gate7760  (.A(g19277), .Z(g22200) ) ;
INV     gate7761  (.A(g19277), .Z(g22201) ) ;
INV     gate7762  (.A(g19638), .Z(II21784) ) ;
INV     gate7763  (.A(II21784), .Z(g22202) ) ;
NOR2    gate7764  (.A(g16031), .B(g13141), .Z(g19422) ) ;
INV     gate7765  (.A(g19422), .Z(II21787) ) ;
INV     gate7766  (.A(II21787), .Z(g22207) ) ;
INV     gate7767  (.A(g21308), .Z(II21792) ) ;
INV     gate7768  (.A(II21792), .Z(g22210) ) ;
INV     gate7769  (.A(g19147), .Z(g22213) ) ;
INV     gate7770  (.A(g19210), .Z(g22214) ) ;
INV     gate7771  (.A(g19277), .Z(g22215) ) ;
INV     gate7772  (.A(g21308), .Z(II21802) ) ;
INV     gate7773  (.A(II21802), .Z(g22220) ) ;
INV     gate7774  (.A(g19210), .Z(g22223) ) ;
INV     gate7775  (.A(g19277), .Z(g22224) ) ;
INV     gate7776  (.A(g19801), .Z(g22227) ) ;
INV     gate7777  (.A(g20596), .Z(II21810) ) ;
INV     gate7778  (.A(II21810), .Z(g22228) ) ;
INV     gate7779  (.A(g21308), .Z(II21815) ) ;
INV     gate7780  (.A(II21815), .Z(g22300) ) ;
INV     gate7781  (.A(g19277), .Z(g22303) ) ;
INV     gate7782  (.A(g19801), .Z(g22305) ) ;
AND2    gate7783  (.A(g4322), .B(g15574), .Z(g18935) ) ;
INV     gate7784  (.A(g18935), .Z(g22311) ) ;
INV     gate7785  (.A(g19801), .Z(g22317) ) ;
INV     gate7786  (.A(g19127), .Z(II21831) ) ;
INV     gate7787  (.A(II21831), .Z(g22319) ) ;
INV     gate7788  (.A(g19801), .Z(g22330) ) ;
INV     gate7789  (.A(g19263), .Z(II21838) ) ;
INV     gate7790  (.A(II21838), .Z(g22332) ) ;
INV     gate7791  (.A(g19801), .Z(g22338) ) ;
INV     gate7792  (.A(g19801), .Z(g22339) ) ;
INV     gate7793  (.A(g19801), .Z(g22341) ) ;
INV     gate7794  (.A(g19801), .Z(g22358) ) ;
NAND3   gate7795  (.A(g15969), .B(g10841), .C(g7781), .Z(g19495) ) ;
INV     gate7796  (.A(g19495), .Z(g22359) ) ;
INV     gate7797  (.A(g19620), .Z(II21849) ) ;
INV     gate7798  (.A(II21849), .Z(g22360) ) ;
NAND2   gate7799  (.A(g4087), .B(g15825), .Z(g19506) ) ;
INV     gate7800  (.A(g19506), .Z(g22406) ) ;
NAND3   gate7801  (.A(g15969), .B(g10841), .C(g7781), .Z(g19455) ) ;
INV     gate7802  (.A(g19455), .Z(g22407) ) ;
NAND3   gate7803  (.A(g15969), .B(g10841), .C(g10922), .Z(g19483) ) ;
INV     gate7804  (.A(g19483), .Z(g22408) ) ;
INV     gate7805  (.A(g19638), .Z(II21860) ) ;
INV     gate7806  (.A(II21860), .Z(g22409) ) ;
NAND2   gate7807  (.A(g1199), .B(g15995), .Z(g19597) ) ;
INV     gate7808  (.A(g19597), .Z(g22449) ) ;
INV     gate7809  (.A(g19801), .Z(g22455) ) ;
INV     gate7810  (.A(g19801), .Z(g22456) ) ;
NAND2   gate7811  (.A(g1542), .B(g16047), .Z(g19614) ) ;
INV     gate7812  (.A(g19614), .Z(g22492) ) ;
INV     gate7813  (.A(g19801), .Z(g22493) ) ;
INV     gate7814  (.A(g19801), .Z(g22494) ) ;
INV     gate7815  (.A(g19801), .Z(g22495) ) ;
NAND3   gate7816  (.A(g15969), .B(g10841), .C(g10899), .Z(g19510) ) ;
INV     gate7817  (.A(g19510), .Z(g22496) ) ;
NAND3   gate7818  (.A(g15969), .B(g10841), .C(g10922), .Z(g19513) ) ;
INV     gate7819  (.A(g19513), .Z(g22497) ) ;
INV     gate7820  (.A(g19801), .Z(g22519) ) ;
INV     gate7821  (.A(g19801), .Z(g22520) ) ;
INV     gate7822  (.A(g19801), .Z(g22526) ) ;
NAND3   gate7823  (.A(g15969), .B(g10841), .C(g10884), .Z(g19546) ) ;
INV     gate7824  (.A(g19546), .Z(g22527) ) ;
INV     gate7825  (.A(g19801), .Z(g22528) ) ;
NAND3   gate7826  (.A(g15969), .B(g10841), .C(g10899), .Z(g19549) ) ;
INV     gate7827  (.A(g19549), .Z(g22529) ) ;
INV     gate7828  (.A(g21278), .Z(II21911) ) ;
INV     gate7829  (.A(II21911), .Z(g22541) ) ;
INV     gate7830  (.A(g19801), .Z(g22542) ) ;
INV     gate7831  (.A(g19801), .Z(g22543) ) ;
NAND3   gate7832  (.A(g15969), .B(g10841), .C(g10884), .Z(g19589) ) ;
INV     gate7833  (.A(g19589), .Z(g22544) ) ;
INV     gate7834  (.A(g21290), .Z(II21918) ) ;
INV     gate7835  (.A(II21918), .Z(g22546) ) ;
INV     gate7836  (.A(g21335), .Z(II21922) ) ;
INV     gate7837  (.A(II21922), .Z(g22550) ) ;
INV     gate7838  (.A(g21297), .Z(II21930) ) ;
INV     gate7839  (.A(II21930), .Z(g22592) ) ;
INV     gate7840  (.A(g19801), .Z(g22593) ) ;
INV     gate7841  (.A(g21273), .Z(II21934) ) ;
INV     gate7842  (.A(II21934), .Z(g22594) ) ;
INV     gate7843  (.A(g18918), .Z(II21941) ) ;
INV     gate7844  (.A(II21941), .Z(g22626) ) ;
INV     gate7845  (.A(g19801), .Z(g22635) ) ;
INV     gate7846  (.A(g19389), .Z(g22646) ) ;
INV     gate7847  (.A(g20242), .Z(II21959) ) ;
INV     gate7848  (.A(II21959), .Z(g22647) ) ;
NOR2    gate7849  (.A(g7909), .B(g15674), .Z(g19063) ) ;
INV     gate7850  (.A(g19063), .Z(g22649) ) ;
INV     gate7851  (.A(g21370), .Z(II21969) ) ;
INV     gate7852  (.A(II21969), .Z(g22658) ) ;
NOR2    gate7853  (.A(g7939), .B(g15695), .Z(g19140) ) ;
INV     gate7854  (.A(g19140), .Z(g22660) ) ;
INV     gate7855  (.A(g21156), .Z(g22667) ) ;
INV     gate7856  (.A(g19379), .Z(g22682) ) ;
INV     gate7857  (.A(g20277), .Z(II22000) ) ;
INV     gate7858  (.A(II22000), .Z(g22683) ) ;
INV     gate7859  (.A(g21269), .Z(II22009) ) ;
INV     gate7860  (.A(II22009), .Z(g22698) ) ;
INV     gate7861  (.A(g20436), .Z(g22714) ) ;
NAND2   gate7862  (.A(g13600), .B(g16275), .Z(g19795) ) ;
INV     gate7863  (.A(g19795), .Z(g22716) ) ;
AND2    gate7864  (.A(g16282), .B(g4864), .Z(g20887) ) ;
INV     gate7865  (.A(g20887), .Z(g22718) ) ;
AND2    gate7866  (.A(g15968), .B(g13505), .Z(g19350) ) ;
INV     gate7867  (.A(g19350), .Z(II22024) ) ;
INV     gate7868  (.A(II22024), .Z(g22719) ) ;
INV     gate7869  (.A(g20204), .Z(II22028) ) ;
INV     gate7870  (.A(II22028), .Z(g22721) ) ;
INV     gate7871  (.A(g21387), .Z(II22031) ) ;
INV     gate7872  (.A(II22031), .Z(g22722) ) ;
INV     gate7873  (.A(g20436), .Z(g22756) ) ;
INV     gate7874  (.A(g20330), .Z(g22758) ) ;
NAND2   gate7875  (.A(g13628), .B(g16296), .Z(g19857) ) ;
INV     gate7876  (.A(g19857), .Z(g22759) ) ;
AND2    gate7877  (.A(g16306), .B(g4871), .Z(g21024) ) ;
INV     gate7878  (.A(g21024), .Z(g22761) ) ;
INV     gate7879  (.A(g19330), .Z(II22046) ) ;
INV     gate7880  (.A(II22046), .Z(g22763) ) ;
INV     gate7881  (.A(g20283), .Z(g22830) ) ;
INV     gate7882  (.A(g20330), .Z(g22840) ) ;
INV     gate7883  (.A(g20391), .Z(g22841) ) ;
NAND2   gate7884  (.A(g13667), .B(g16316), .Z(g19875) ) ;
INV     gate7885  (.A(g19875), .Z(g22842) ) ;
AND2    gate7886  (.A(g16321), .B(g4878), .Z(g21163) ) ;
INV     gate7887  (.A(g21163), .Z(g22844) ) ;
AND2    gate7888  (.A(g16238), .B(g4646), .Z(g20682) ) ;
INV     gate7889  (.A(g20682), .Z(g22845) ) ;
INV     gate7890  (.A(g20283), .Z(g22847) ) ;
INV     gate7891  (.A(g20330), .Z(g22854) ) ;
INV     gate7892  (.A(g20391), .Z(g22855) ) ;
INV     gate7893  (.A(g20453), .Z(g22856) ) ;
AND2    gate7894  (.A(g16259), .B(g4674), .Z(g20739) ) ;
INV     gate7895  (.A(g20739), .Z(g22857) ) ;
AND2    gate7896  (.A(g16260), .B(g4836), .Z(g20751) ) ;
INV     gate7897  (.A(g20751), .Z(g22858) ) ;
NOR2    gate7898  (.A(g13661), .B(g16264), .Z(g20000) ) ;
INV     gate7899  (.A(g20000), .Z(g22860) ) ;
INV     gate7900  (.A(g20330), .Z(g22865) ) ;
INV     gate7901  (.A(g20330), .Z(g22866) ) ;
INV     gate7902  (.A(g20391), .Z(g22867) ) ;
INV     gate7903  (.A(g20453), .Z(g22868) ) ;
AND2    gate7904  (.A(g16281), .B(g4681), .Z(g20875) ) ;
INV     gate7905  (.A(g20875), .Z(g22869) ) ;
INV     gate7906  (.A(g20887), .Z(g22870) ) ;
NOR2    gate7907  (.A(g16987), .B(g8058), .Z(g19890) ) ;
INV     gate7908  (.A(g19890), .Z(II22096) ) ;
INV     gate7909  (.A(II22096), .Z(g22881) ) ;
INV     gate7910  (.A(g20391), .Z(g22882) ) ;
INV     gate7911  (.A(g20391), .Z(g22883) ) ;
INV     gate7912  (.A(g20453), .Z(g22884) ) ;
AND2    gate7913  (.A(g16304), .B(g4688), .Z(g21012) ) ;
INV     gate7914  (.A(g21012), .Z(g22896) ) ;
INV     gate7915  (.A(g21024), .Z(g22897) ) ;
INV     gate7916  (.A(g20283), .Z(g22898) ) ;
INV     gate7917  (.A(g20330), .Z(g22903) ) ;
NOR2    gate7918  (.A(g16987), .B(g11205), .Z(g19919) ) ;
INV     gate7919  (.A(g19919), .Z(II22111) ) ;
INV     gate7920  (.A(II22111), .Z(g22904) ) ;
NOR2    gate7921  (.A(g17062), .B(g8113), .Z(g19935) ) ;
INV     gate7922  (.A(g19935), .Z(II22114) ) ;
INV     gate7923  (.A(II22114), .Z(g22905) ) ;
INV     gate7924  (.A(g20453), .Z(g22906) ) ;
INV     gate7925  (.A(g20453), .Z(g22907) ) ;
INV     gate7926  (.A(g21163), .Z(g22919) ) ;
INV     gate7927  (.A(g20330), .Z(g22922) ) ;
INV     gate7928  (.A(g21300), .Z(II22124) ) ;
INV     gate7929  (.A(II22124), .Z(g22923) ) ;
INV     gate7930  (.A(g20391), .Z(g22926) ) ;
NOR2    gate7931  (.A(g17062), .B(g11223), .Z(g19968) ) ;
INV     gate7932  (.A(g19968), .Z(II22128) ) ;
INV     gate7933  (.A(II22128), .Z(g22927) ) ;
NOR2    gate7934  (.A(g17096), .B(g8171), .Z(g19984) ) ;
INV     gate7935  (.A(g19984), .Z(II22131) ) ;
INV     gate7936  (.A(II22131), .Z(g22928) ) ;
INV     gate7937  (.A(g20283), .Z(g22935) ) ;
INV     gate7938  (.A(g20283), .Z(g22936) ) ;
INV     gate7939  (.A(g20189), .Z(II22143) ) ;
INV     gate7940  (.A(II22143), .Z(g22957) ) ;
INV     gate7941  (.A(g20330), .Z(g22973) ) ;
INV     gate7942  (.A(g20330), .Z(g22974) ) ;
INV     gate7943  (.A(g20391), .Z(g22975) ) ;
INV     gate7944  (.A(g21036), .Z(II22149) ) ;
INV     gate7945  (.A(II22149), .Z(g22976) ) ;
INV     gate7946  (.A(g20453), .Z(g22979) ) ;
NOR2    gate7947  (.A(g17096), .B(g11244), .Z(g20014) ) ;
INV     gate7948  (.A(g20014), .Z(II22153) ) ;
INV     gate7949  (.A(II22153), .Z(g22980) ) ;
INV     gate7950  (.A(g20283), .Z(g22981) ) ;
INV     gate7951  (.A(g20330), .Z(g22985) ) ;
INV     gate7952  (.A(g20330), .Z(g22986) ) ;
INV     gate7953  (.A(g20391), .Z(g22987) ) ;
INV     gate7954  (.A(g20391), .Z(g22988) ) ;
INV     gate7955  (.A(g20453), .Z(g22989) ) ;
INV     gate7956  (.A(g20436), .Z(g22994) ) ;
INV     gate7957  (.A(g20330), .Z(g22995) ) ;
INV     gate7958  (.A(g20330), .Z(g22996) ) ;
INV     gate7959  (.A(g20391), .Z(g22997) ) ;
INV     gate7960  (.A(g20391), .Z(g22998) ) ;
INV     gate7961  (.A(g20453), .Z(g22999) ) ;
INV     gate7962  (.A(g20453), .Z(g23000) ) ;
INV     gate7963  (.A(g19801), .Z(g23001) ) ;
INV     gate7964  (.A(g21366), .Z(II22177) ) ;
INV     gate7965  (.A(g21366), .Z(II22180) ) ;
INV     gate7966  (.A(II22180), .Z(g23003) ) ;
INV     gate7967  (.A(g20283), .Z(g23004) ) ;
INV     gate7968  (.A(g20283), .Z(g23005) ) ;
INV     gate7969  (.A(g20330), .Z(g23011) ) ;
INV     gate7970  (.A(g20330), .Z(g23012) ) ;
INV     gate7971  (.A(g20330), .Z(g23013) ) ;
INV     gate7972  (.A(g20391), .Z(g23014) ) ;
INV     gate7973  (.A(g20391), .Z(g23015) ) ;
INV     gate7974  (.A(g20453), .Z(g23016) ) ;
INV     gate7975  (.A(g20453), .Z(g23017) ) ;
INV     gate7976  (.A(g19801), .Z(g23018) ) ;
INV     gate7977  (.A(g19866), .Z(g23019) ) ;
INV     gate7978  (.A(g19869), .Z(g23020) ) ;
INV     gate7979  (.A(g20283), .Z(g23021) ) ;
INV     gate7980  (.A(g20283), .Z(g23022) ) ;
INV     gate7981  (.A(g20391), .Z(g23026) ) ;
INV     gate7982  (.A(g20391), .Z(g23027) ) ;
INV     gate7983  (.A(g20391), .Z(g23028) ) ;
INV     gate7984  (.A(g20453), .Z(g23029) ) ;
INV     gate7985  (.A(g20453), .Z(g23030) ) ;
INV     gate7986  (.A(g19801), .Z(g23031) ) ;
INV     gate7987  (.A(g21463), .Z(II22211) ) ;
INV     gate7988  (.A(II22211), .Z(g23032) ) ;
INV     gate7989  (.A(g19882), .Z(g23041) ) ;
INV     gate7990  (.A(g20283), .Z(g23046) ) ;
INV     gate7991  (.A(g20887), .Z(g23055) ) ;
INV     gate7992  (.A(g20453), .Z(g23057) ) ;
INV     gate7993  (.A(g20453), .Z(g23058) ) ;
INV     gate7994  (.A(g20453), .Z(g23059) ) ;
INV     gate7995  (.A(g19908), .Z(g23060) ) ;
INV     gate7996  (.A(g20283), .Z(g23061) ) ;
INV     gate7997  (.A(g20330), .Z(g23066) ) ;
INV     gate7998  (.A(g21024), .Z(g23082) ) ;
INV     gate7999  (.A(g19954), .Z(g23084) ) ;
INV     gate8000  (.A(g19957), .Z(g23085) ) ;
INV     gate8001  (.A(g20283), .Z(g23086) ) ;
INV     gate8002  (.A(g20086), .Z(II22240) ) ;
INV     gate8003  (.A(II22240), .Z(g23088) ) ;
INV     gate8004  (.A(g20391), .Z(g23111) ) ;
INV     gate8005  (.A(g21163), .Z(g23127) ) ;
INV     gate8006  (.A(g20283), .Z(g23128) ) ;
INV     gate8007  (.A(g20453), .Z(g23138) ) ;
INV     gate8008  (.A(g20283), .Z(g23152) ) ;
INV     gate8009  (.A(g20100), .Z(II22264) ) ;
INV     gate8010  (.A(II22264), .Z(g23154) ) ;
INV     gate8011  (.A(g20046), .Z(g23170) ) ;
INV     gate8012  (.A(g20127), .Z(II22275) ) ;
INV     gate8013  (.A(II22275), .Z(g23172) ) ;
NOR3    gate8014  (.A(g10143), .B(g17748), .C(g12259), .Z(g21389) ) ;
INV     gate8015  (.A(g21389), .Z(g23182) ) ;
INV     gate8016  (.A(g20060), .Z(g23189) ) ;
INV     gate8017  (.A(g19446), .Z(II22286) ) ;
INV     gate8018  (.A(g19446), .Z(II22289) ) ;
INV     gate8019  (.A(II22289), .Z(g23191) ) ;
NAND3   gate8020  (.A(g17056), .B(g14146), .C(g14123), .Z(g20248) ) ;
INV     gate8021  (.A(g20248), .Z(g23192) ) ;
INV     gate8022  (.A(g20785), .Z(g23196) ) ;
INV     gate8023  (.A(g19353), .Z(II22302) ) ;
INV     gate8024  (.A(II22302), .Z(g23202) ) ;
INV     gate8025  (.A(g20073), .Z(g23203) ) ;
INV     gate8026  (.A(g21308), .Z(g23211) ) ;
INV     gate8027  (.A(g20785), .Z(g23214) ) ;
INV     gate8028  (.A(g20785), .Z(g23215) ) ;
INV     gate8029  (.A(g20924), .Z(g23216) ) ;
INV     gate8030  (.A(g19361), .Z(II22316) ) ;
INV     gate8031  (.A(II22316), .Z(g23219) ) ;
INV     gate8032  (.A(g20785), .Z(g23221) ) ;
INV     gate8033  (.A(g20785), .Z(g23222) ) ;
INV     gate8034  (.A(g21308), .Z(g23223) ) ;
INV     gate8035  (.A(g20924), .Z(g23226) ) ;
INV     gate8036  (.A(g20924), .Z(g23227) ) ;
INV     gate8037  (.A(g21070), .Z(g23228) ) ;
INV     gate8038  (.A(g19367), .Z(II22327) ) ;
INV     gate8039  (.A(II22327), .Z(g23230) ) ;
INV     gate8040  (.A(g20050), .Z(g23231) ) ;
INV     gate8041  (.A(g19417), .Z(II22331) ) ;
INV     gate8042  (.A(II22331), .Z(g23232) ) ;
INV     gate8043  (.A(g21037), .Z(g23233) ) ;
AND2    gate8044  (.A(g671), .B(g16846), .Z(g20375) ) ;
INV     gate8045  (.A(g20375), .Z(g23234) ) ;
INV     gate8046  (.A(g20785), .Z(g23235) ) ;
INV     gate8047  (.A(g20785), .Z(g23236) ) ;
INV     gate8048  (.A(g20924), .Z(g23237) ) ;
INV     gate8049  (.A(g20924), .Z(g23238) ) ;
INV     gate8050  (.A(g21308), .Z(g23239) ) ;
INV     gate8051  (.A(g21070), .Z(g23242) ) ;
INV     gate8052  (.A(g21070), .Z(g23243) ) ;
INV     gate8053  (.A(g19371), .Z(II22343) ) ;
INV     gate8054  (.A(II22343), .Z(g23244) ) ;
INV     gate8055  (.A(g20785), .Z(g23245) ) ;
INV     gate8056  (.A(g20785), .Z(g23246) ) ;
INV     gate8057  (.A(g20924), .Z(g23247) ) ;
INV     gate8058  (.A(g20924), .Z(g23248) ) ;
INV     gate8059  (.A(g21070), .Z(g23249) ) ;
INV     gate8060  (.A(g21070), .Z(g23250) ) ;
INV     gate8061  (.A(g19375), .Z(II22353) ) ;
INV     gate8062  (.A(II22353), .Z(g23252) ) ;
INV     gate8063  (.A(g21037), .Z(g23253) ) ;
INV     gate8064  (.A(g20785), .Z(g23256) ) ;
INV     gate8065  (.A(g20924), .Z(g23257) ) ;
INV     gate8066  (.A(g20924), .Z(g23258) ) ;
INV     gate8067  (.A(g21070), .Z(g23259) ) ;
INV     gate8068  (.A(g21070), .Z(g23260) ) ;
INV     gate8069  (.A(g19757), .Z(II22366) ) ;
INV     gate8070  (.A(II22366), .Z(g23263) ) ;
INV     gate8071  (.A(g21037), .Z(g23264) ) ;
INV     gate8072  (.A(g20097), .Z(g23267) ) ;
INV     gate8073  (.A(g20785), .Z(g23270) ) ;
INV     gate8074  (.A(g20785), .Z(g23271) ) ;
INV     gate8075  (.A(g20924), .Z(g23272) ) ;
INV     gate8076  (.A(g21070), .Z(g23273) ) ;
INV     gate8077  (.A(g21070), .Z(g23274) ) ;
INV     gate8078  (.A(g21156), .Z(II22380) ) ;
INV     gate8079  (.A(II22380), .Z(g23277) ) ;
INV     gate8080  (.A(g20283), .Z(g23278) ) ;
INV     gate8081  (.A(g21037), .Z(g23279) ) ;
INV     gate8082  (.A(g20330), .Z(g23282) ) ;
INV     gate8083  (.A(g20785), .Z(g23283) ) ;
INV     gate8084  (.A(g20785), .Z(g23284) ) ;
INV     gate8085  (.A(g20887), .Z(g23285) ) ;
INV     gate8086  (.A(g20924), .Z(g23289) ) ;
INV     gate8087  (.A(g20924), .Z(g23290) ) ;
INV     gate8088  (.A(g21070), .Z(g23291) ) ;
INV     gate8089  (.A(g19620), .Z(II22400) ) ;
INV     gate8090  (.A(II22400), .Z(g23299) ) ;
INV     gate8091  (.A(g20283), .Z(g23300) ) ;
INV     gate8092  (.A(g21037), .Z(g23301) ) ;
INV     gate8093  (.A(g20330), .Z(g23302) ) ;
INV     gate8094  (.A(g20785), .Z(g23303) ) ;
INV     gate8095  (.A(g20785), .Z(g23304) ) ;
INV     gate8096  (.A(g20391), .Z(g23305) ) ;
INV     gate8097  (.A(g20924), .Z(g23306) ) ;
INV     gate8098  (.A(g20924), .Z(g23307) ) ;
INV     gate8099  (.A(g21024), .Z(g23308) ) ;
INV     gate8100  (.A(g21070), .Z(g23312) ) ;
INV     gate8101  (.A(g21070), .Z(g23313) ) ;
INV     gate8102  (.A(g19638), .Z(II22419) ) ;
INV     gate8103  (.A(II22419), .Z(g23320) ) ;
INV     gate8104  (.A(g19330), .Z(II22422) ) ;
INV     gate8105  (.A(II22422), .Z(g23321) ) ;
INV     gate8106  (.A(g19379), .Z(II22425) ) ;
INV     gate8107  (.A(II22425), .Z(g23322) ) ;
INV     gate8108  (.A(g20283), .Z(g23323) ) ;
OR2     gate8109  (.A(g7216), .B(g17264), .Z(g20905) ) ;
INV     gate8110  (.A(g20905), .Z(g23331) ) ;
INV     gate8111  (.A(g20785), .Z(g23332) ) ;
INV     gate8112  (.A(g20785), .Z(g23333) ) ;
INV     gate8113  (.A(g20785), .Z(g23334) ) ;
INV     gate8114  (.A(g20391), .Z(g23335) ) ;
INV     gate8115  (.A(g20924), .Z(g23336) ) ;
INV     gate8116  (.A(g20924), .Z(g23337) ) ;
INV     gate8117  (.A(g20453), .Z(g23338) ) ;
INV     gate8118  (.A(g21070), .Z(g23339) ) ;
INV     gate8119  (.A(g21070), .Z(g23340) ) ;
INV     gate8120  (.A(g21163), .Z(g23341) ) ;
INV     gate8121  (.A(g19626), .Z(II22444) ) ;
INV     gate8122  (.A(II22444), .Z(g23347) ) ;
INV     gate8123  (.A(g20785), .Z(g23350) ) ;
INV     gate8124  (.A(g20924), .Z(g23351) ) ;
INV     gate8125  (.A(g20924), .Z(g23352) ) ;
INV     gate8126  (.A(g20924), .Z(g23353) ) ;
INV     gate8127  (.A(g20453), .Z(g23354) ) ;
INV     gate8128  (.A(g21070), .Z(g23355) ) ;
INV     gate8129  (.A(g21070), .Z(g23356) ) ;
INV     gate8130  (.A(g18954), .Z(II22458) ) ;
INV     gate8131  (.A(II22458), .Z(g23359) ) ;
INV     gate8132  (.A(g21225), .Z(II22461) ) ;
INV     gate8133  (.A(II22461), .Z(g23360) ) ;
INV     gate8134  (.A(g21222), .Z(II22464) ) ;
INV     gate8135  (.A(II22464), .Z(g23361) ) ;
INV     gate8136  (.A(g19662), .Z(II22467) ) ;
INV     gate8137  (.A(II22467), .Z(g23362) ) ;
INV     gate8138  (.A(g21326), .Z(II22470) ) ;
INV     gate8139  (.A(II22470), .Z(g23363) ) ;
INV     gate8140  (.A(g20924), .Z(g23375) ) ;
INV     gate8141  (.A(g21070), .Z(g23376) ) ;
INV     gate8142  (.A(g21070), .Z(g23377) ) ;
INV     gate8143  (.A(g21070), .Z(g23378) ) ;
NAND2   gate8144  (.A(g14317), .B(g17217), .Z(g20619) ) ;
INV     gate8145  (.A(g20619), .Z(g23380) ) ;
INV     gate8146  (.A(g20682), .Z(g23382) ) ;
INV     gate8147  (.A(g21308), .Z(II22485) ) ;
INV     gate8148  (.A(II22485), .Z(g23384) ) ;
INV     gate8149  (.A(g18984), .Z(II22488) ) ;
INV     gate8150  (.A(II22488), .Z(g23385) ) ;
INV     gate8151  (.A(g21070), .Z(g23388) ) ;
INV     gate8152  (.A(g21468), .Z(g23390) ) ;
NAND2   gate8153  (.A(g14344), .B(g17243), .Z(g20645) ) ;
INV     gate8154  (.A(g20645), .Z(g23391) ) ;
INV     gate8155  (.A(g20739), .Z(g23393) ) ;
INV     gate8156  (.A(g21160), .Z(II22499) ) ;
INV     gate8157  (.A(II22499), .Z(g23394) ) ;
INV     gate8158  (.A(g19376), .Z(II22502) ) ;
INV     gate8159  (.A(II22502), .Z(g23395) ) ;
INV     gate8160  (.A(g21468), .Z(g23398) ) ;
INV     gate8161  (.A(g21514), .Z(g23399) ) ;
NAND2   gate8162  (.A(g14379), .B(g17287), .Z(g20676) ) ;
INV     gate8163  (.A(g20676), .Z(g23400) ) ;
INV     gate8164  (.A(g20875), .Z(g23402) ) ;
INV     gate8165  (.A(g19389), .Z(II22512) ) ;
INV     gate8166  (.A(II22512), .Z(g23403) ) ;
INV     gate8167  (.A(g20330), .Z(g23406) ) ;
INV     gate8168  (.A(g21468), .Z(g23408) ) ;
INV     gate8169  (.A(g21514), .Z(g23409) ) ;
INV     gate8170  (.A(g21562), .Z(g23410) ) ;
NAND2   gate8171  (.A(g14408), .B(g17312), .Z(g20734) ) ;
INV     gate8172  (.A(g20734), .Z(g23411) ) ;
INV     gate8173  (.A(g21012), .Z(g23413) ) ;
INV     gate8174  (.A(g19345), .Z(II22525) ) ;
INV     gate8175  (.A(II22525), .Z(g23414) ) ;
INV     gate8176  (.A(g20391), .Z(g23417) ) ;
INV     gate8177  (.A(g21468), .Z(g23418) ) ;
INV     gate8178  (.A(g21468), .Z(g23419) ) ;
INV     gate8179  (.A(g21514), .Z(g23420) ) ;
INV     gate8180  (.A(g21562), .Z(g23421) ) ;
INV     gate8181  (.A(g21611), .Z(g23422) ) ;
NAND2   gate8182  (.A(g14434), .B(g17396), .Z(g20871) ) ;
INV     gate8183  (.A(g20871), .Z(g23423) ) ;
INV     gate8184  (.A(g20751), .Z(g23425) ) ;
INV     gate8185  (.A(g19606), .Z(II22539) ) ;
INV     gate8186  (.A(II22539), .Z(g23426) ) ;
INV     gate8187  (.A(g19773), .Z(II22542) ) ;
INV     gate8188  (.A(II22542), .Z(g23427) ) ;
INV     gate8189  (.A(g20453), .Z(g23429) ) ;
NOR2    gate8190  (.A(g17847), .B(g9299), .Z(g20720) ) ;
INV     gate8191  (.A(g20720), .Z(II22547) ) ;
INV     gate8192  (.A(II22547), .Z(g23430) ) ;
INV     gate8193  (.A(g21514), .Z(g23431) ) ;
INV     gate8194  (.A(g21514), .Z(g23432) ) ;
INV     gate8195  (.A(g21562), .Z(g23433) ) ;
INV     gate8196  (.A(g21611), .Z(g23434) ) ;
INV     gate8197  (.A(g18833), .Z(g23435) ) ;
INV     gate8198  (.A(g20695), .Z(II22557) ) ;
INV     gate8199  (.A(II22557), .Z(g23440) ) ;
INV     gate8200  (.A(g21468), .Z(g23443) ) ;
NOR2    gate8201  (.A(g17847), .B(g12027), .Z(g20841) ) ;
INV     gate8202  (.A(g20841), .Z(II22561) ) ;
INV     gate8203  (.A(II22561), .Z(g23444) ) ;
NOR2    gate8204  (.A(g17929), .B(g9380), .Z(g20857) ) ;
INV     gate8205  (.A(g20857), .Z(II22564) ) ;
INV     gate8206  (.A(II22564), .Z(g23445) ) ;
INV     gate8207  (.A(g21562), .Z(g23446) ) ;
INV     gate8208  (.A(g21562), .Z(g23447) ) ;
INV     gate8209  (.A(g21611), .Z(g23448) ) ;
INV     gate8210  (.A(g18833), .Z(g23449) ) ;
INV     gate8211  (.A(g20097), .Z(II22571) ) ;
INV     gate8212  (.A(II22571), .Z(g23450) ) ;
INV     gate8213  (.A(g21468), .Z(g23452) ) ;
INV     gate8214  (.A(g21282), .Z(II22576) ) ;
INV     gate8215  (.A(II22576), .Z(g23453) ) ;
INV     gate8216  (.A(g21514), .Z(g23456) ) ;
NOR2    gate8217  (.A(g17929), .B(g12065), .Z(g20982) ) ;
INV     gate8218  (.A(g20982), .Z(II22580) ) ;
INV     gate8219  (.A(II22580), .Z(g23457) ) ;
NOR2    gate8220  (.A(g18065), .B(g9450), .Z(g20998) ) ;
INV     gate8221  (.A(g20998), .Z(II22583) ) ;
INV     gate8222  (.A(II22583), .Z(g23458) ) ;
INV     gate8223  (.A(g21611), .Z(g23459) ) ;
INV     gate8224  (.A(g21611), .Z(g23460) ) ;
INV     gate8225  (.A(g18833), .Z(g23461) ) ;
INV     gate8226  (.A(g21340), .Z(II22589) ) ;
INV     gate8227  (.A(II22589), .Z(g23462) ) ;
NOR2    gate8228  (.A(g9547), .B(g17297), .Z(g21062) ) ;
INV     gate8229  (.A(g21062), .Z(g23472) ) ;
INV     gate8230  (.A(g20785), .Z(g23473) ) ;
INV     gate8231  (.A(g21468), .Z(g23476) ) ;
INV     gate8232  (.A(g21468), .Z(g23477) ) ;
INV     gate8233  (.A(g21514), .Z(g23478) ) ;
INV     gate8234  (.A(g21562), .Z(g23479) ) ;
NOR2    gate8235  (.A(g18065), .B(g12099), .Z(g21127) ) ;
INV     gate8236  (.A(g21127), .Z(II22601) ) ;
INV     gate8237  (.A(II22601), .Z(g23480) ) ;
NOR2    gate8238  (.A(g15348), .B(g9517), .Z(g21143) ) ;
INV     gate8239  (.A(g21143), .Z(II22604) ) ;
INV     gate8240  (.A(II22604), .Z(g23481) ) ;
INV     gate8241  (.A(g18833), .Z(g23482) ) ;
INV     gate8242  (.A(g18833), .Z(g23483) ) ;
INV     gate8243  (.A(g20785), .Z(g23485) ) ;
INV     gate8244  (.A(g20785), .Z(g23486) ) ;
INV     gate8245  (.A(g20924), .Z(g23487) ) ;
INV     gate8246  (.A(g21468), .Z(g23488) ) ;
INV     gate8247  (.A(g21468), .Z(g23489) ) ;
INV     gate8248  (.A(g21514), .Z(g23490) ) ;
INV     gate8249  (.A(g21514), .Z(g23491) ) ;
INV     gate8250  (.A(g21562), .Z(g23492) ) ;
INV     gate8251  (.A(g21611), .Z(g23493) ) ;
NOR2    gate8252  (.A(g15348), .B(g12135), .Z(g21193) ) ;
INV     gate8253  (.A(g21193), .Z(II22619) ) ;
INV     gate8254  (.A(II22619), .Z(g23494) ) ;
NOR2    gate8255  (.A(g15483), .B(g9575), .Z(g21209) ) ;
INV     gate8256  (.A(g21209), .Z(II22622) ) ;
INV     gate8257  (.A(II22622), .Z(g23495) ) ;
INV     gate8258  (.A(g20248), .Z(g23496) ) ;
INV     gate8259  (.A(g20785), .Z(g23499) ) ;
INV     gate8260  (.A(g20924), .Z(g23500) ) ;
INV     gate8261  (.A(g20924), .Z(g23501) ) ;
INV     gate8262  (.A(g21070), .Z(g23502) ) ;
INV     gate8263  (.A(g21468), .Z(g23503) ) ;
INV     gate8264  (.A(g21468), .Z(g23504) ) ;
INV     gate8265  (.A(g21514), .Z(g23505) ) ;
INV     gate8266  (.A(g21514), .Z(g23506) ) ;
INV     gate8267  (.A(g21562), .Z(g23507) ) ;
INV     gate8268  (.A(g21562), .Z(g23508) ) ;
INV     gate8269  (.A(g21611), .Z(g23509) ) ;
INV     gate8270  (.A(g18833), .Z(g23510) ) ;
NOR2    gate8271  (.A(g15483), .B(g12179), .Z(g21256) ) ;
INV     gate8272  (.A(g21256), .Z(II22640) ) ;
INV     gate8273  (.A(II22640), .Z(g23511) ) ;
INV     gate8274  (.A(g20248), .Z(g23512) ) ;
INV     gate8275  (.A(g20785), .Z(g23515) ) ;
INV     gate8276  (.A(g20924), .Z(g23516) ) ;
INV     gate8277  (.A(g21070), .Z(g23517) ) ;
INV     gate8278  (.A(g21070), .Z(g23518) ) ;
INV     gate8279  (.A(g21468), .Z(g23519) ) ;
INV     gate8280  (.A(g21468), .Z(g23520) ) ;
INV     gate8281  (.A(g21468), .Z(g23521) ) ;
INV     gate8282  (.A(g21514), .Z(g23522) ) ;
INV     gate8283  (.A(g21514), .Z(g23523) ) ;
INV     gate8284  (.A(g21562), .Z(g23524) ) ;
INV     gate8285  (.A(g21562), .Z(g23525) ) ;
INV     gate8286  (.A(g21611), .Z(g23526) ) ;
INV     gate8287  (.A(g21611), .Z(g23527) ) ;
INV     gate8288  (.A(g18833), .Z(g23528) ) ;
INV     gate8289  (.A(g20558), .Z(g23529) ) ;
INV     gate8290  (.A(g20248), .Z(g23530) ) ;
INV     gate8291  (.A(g21308), .Z(II22665) ) ;
INV     gate8292  (.A(II22665), .Z(g23534) ) ;
INV     gate8293  (.A(g20785), .Z(g23537) ) ;
INV     gate8294  (.A(g20924), .Z(g23538) ) ;
INV     gate8295  (.A(g21070), .Z(g23539) ) ;
INV     gate8296  (.A(g21514), .Z(g23541) ) ;
INV     gate8297  (.A(g21514), .Z(g23542) ) ;
INV     gate8298  (.A(g21514), .Z(g23543) ) ;
INV     gate8299  (.A(g21562), .Z(g23544) ) ;
INV     gate8300  (.A(g21562), .Z(g23545) ) ;
INV     gate8301  (.A(g21611), .Z(g23546) ) ;
INV     gate8302  (.A(g21611), .Z(g23547) ) ;
INV     gate8303  (.A(g18833), .Z(g23548) ) ;
INV     gate8304  (.A(g18833), .Z(g23549) ) ;
INV     gate8305  (.A(g20248), .Z(g23550) ) ;
INV     gate8306  (.A(g21308), .Z(II22692) ) ;
INV     gate8307  (.A(II22692), .Z(g23555) ) ;
INV     gate8308  (.A(g20924), .Z(g23558) ) ;
INV     gate8309  (.A(g21070), .Z(g23559) ) ;
INV     gate8310  (.A(g20682), .Z(g23563) ) ;
INV     gate8311  (.A(g21562), .Z(g23565) ) ;
INV     gate8312  (.A(g21562), .Z(g23566) ) ;
INV     gate8313  (.A(g21562), .Z(g23567) ) ;
INV     gate8314  (.A(g21611), .Z(g23568) ) ;
INV     gate8315  (.A(g21611), .Z(g23569) ) ;
INV     gate8316  (.A(g18833), .Z(g23570) ) ;
INV     gate8317  (.A(g18833), .Z(g23571) ) ;
INV     gate8318  (.A(g20248), .Z(g23573) ) ;
NOR3    gate8319  (.A(g9417), .B(g9340), .C(g17494), .Z(g21250) ) ;
INV     gate8320  (.A(g21250), .Z(II22725) ) ;
INV     gate8321  (.A(II22725), .Z(g23578) ) ;
INV     gate8322  (.A(g21308), .Z(II22729) ) ;
INV     gate8323  (.A(II22729), .Z(g23582) ) ;
INV     gate8324  (.A(g21070), .Z(g23585) ) ;
INV     gate8325  (.A(g21468), .Z(g23589) ) ;
INV     gate8326  (.A(g20739), .Z(g23605) ) ;
INV     gate8327  (.A(g21611), .Z(g23607) ) ;
INV     gate8328  (.A(g21611), .Z(g23608) ) ;
INV     gate8329  (.A(g21611), .Z(g23609) ) ;
INV     gate8330  (.A(g18833), .Z(g23610) ) ;
INV     gate8331  (.A(g18833), .Z(g23611) ) ;
INV     gate8332  (.A(g19458), .Z(II22745) ) ;
INV     gate8333  (.A(g19458), .Z(II22748) ) ;
INV     gate8334  (.A(II22748), .Z(g23613) ) ;
INV     gate8335  (.A(g20248), .Z(g23614) ) ;
NOR3    gate8336  (.A(g9417), .B(g9340), .C(g17467), .Z(g21277) ) ;
INV     gate8337  (.A(g21277), .Z(II22769) ) ;
INV     gate8338  (.A(II22769), .Z(g23620) ) ;
INV     gate8339  (.A(g21514), .Z(g23629) ) ;
INV     gate8340  (.A(g20875), .Z(g23645) ) ;
INV     gate8341  (.A(g18833), .Z(g23647) ) ;
INV     gate8342  (.A(g18833), .Z(g23648) ) ;
INV     gate8343  (.A(g18833), .Z(g23649) ) ;
INV     gate8344  (.A(g20653), .Z(g23650) ) ;
INV     gate8345  (.A(g20655), .Z(g23651) ) ;
INV     gate8346  (.A(g18940), .Z(II22785) ) ;
INV     gate8347  (.A(g18940), .Z(II22788) ) ;
INV     gate8348  (.A(II22788), .Z(g23653) ) ;
INV     gate8349  (.A(g20248), .Z(g23654) ) ;
INV     gate8350  (.A(g21562), .Z(g23665) ) ;
INV     gate8351  (.A(g21012), .Z(g23681) ) ;
INV     gate8352  (.A(g19862), .Z(II22816) ) ;
INV     gate8353  (.A(g19862), .Z(II22819) ) ;
INV     gate8354  (.A(II22819), .Z(g23684) ) ;
INV     gate8355  (.A(g21611), .Z(g23698) ) ;
INV     gate8356  (.A(g20751), .Z(g23714) ) ;
INV     gate8357  (.A(g20764), .Z(g23715) ) ;
INV     gate8358  (.A(g18833), .Z(g23732) ) ;
INV     gate8359  (.A(g20900), .Z(g23745) ) ;
INV     gate8360  (.A(g20902), .Z(g23746) ) ;
INV     gate8361  (.A(g18997), .Z(g23749) ) ;
INV     gate8362  (.A(g18926), .Z(II22886) ) ;
INV     gate8363  (.A(g18926), .Z(II22889) ) ;
INV     gate8364  (.A(II22889), .Z(g23760) ) ;
INV     gate8365  (.A(g21308), .Z(g23764) ) ;
INV     gate8366  (.A(g18997), .Z(g23767) ) ;
INV     gate8367  (.A(g18997), .Z(g23768) ) ;
INV     gate8368  (.A(g19074), .Z(g23769) ) ;
INV     gate8369  (.A(g21177), .Z(g23776) ) ;
INV     gate8370  (.A(g21451), .Z(II22918) ) ;
INV     gate8371  (.A(II22918), .Z(g23777) ) ;
INV     gate8372  (.A(g18997), .Z(g23787) ) ;
INV     gate8373  (.A(g18997), .Z(g23788) ) ;
INV     gate8374  (.A(g21308), .Z(g23789) ) ;
INV     gate8375  (.A(g19074), .Z(g23792) ) ;
INV     gate8376  (.A(g19074), .Z(g23793) ) ;
INV     gate8377  (.A(g19147), .Z(g23794) ) ;
INV     gate8378  (.A(g21246), .Z(g23800) ) ;
INV     gate8379  (.A(g18997), .Z(g23812) ) ;
INV     gate8380  (.A(g18997), .Z(g23813) ) ;
INV     gate8381  (.A(g19074), .Z(g23814) ) ;
INV     gate8382  (.A(g19074), .Z(g23815) ) ;
INV     gate8383  (.A(g21308), .Z(g23816) ) ;
INV     gate8384  (.A(g19147), .Z(g23819) ) ;
INV     gate8385  (.A(g19147), .Z(g23820) ) ;
INV     gate8386  (.A(g19210), .Z(g23821) ) ;
INV     gate8387  (.A(g21175), .Z(II22989) ) ;
INV     gate8388  (.A(II22989), .Z(g23823) ) ;
INV     gate8389  (.A(g21271), .Z(g23824) ) ;
INV     gate8390  (.A(g18997), .Z(g23838) ) ;
INV     gate8391  (.A(g18997), .Z(g23839) ) ;
INV     gate8392  (.A(g19074), .Z(g23840) ) ;
INV     gate8393  (.A(g19074), .Z(g23841) ) ;
INV     gate8394  (.A(g19147), .Z(g23842) ) ;
INV     gate8395  (.A(g19147), .Z(g23843) ) ;
INV     gate8396  (.A(g21308), .Z(g23844) ) ;
INV     gate8397  (.A(g19210), .Z(g23847) ) ;
INV     gate8398  (.A(g19210), .Z(g23848) ) ;
INV     gate8399  (.A(g19277), .Z(g23849) ) ;
INV     gate8400  (.A(g18997), .Z(g23858) ) ;
INV     gate8401  (.A(g19074), .Z(g23859) ) ;
INV     gate8402  (.A(g19074), .Z(g23860) ) ;
INV     gate8403  (.A(g19147), .Z(g23861) ) ;
INV     gate8404  (.A(g19147), .Z(g23862) ) ;
INV     gate8405  (.A(g19210), .Z(g23863) ) ;
INV     gate8406  (.A(g19210), .Z(g23864) ) ;
INV     gate8407  (.A(g21308), .Z(g23865) ) ;
INV     gate8408  (.A(g19277), .Z(g23868) ) ;
INV     gate8409  (.A(g19277), .Z(g23869) ) ;
INV     gate8410  (.A(g21293), .Z(g23870) ) ;
INV     gate8411  (.A(g18997), .Z(g23874) ) ;
INV     gate8412  (.A(g18997), .Z(g23875) ) ;
INV     gate8413  (.A(g19074), .Z(g23876) ) ;
INV     gate8414  (.A(g19147), .Z(g23877) ) ;
INV     gate8415  (.A(g19147), .Z(g23878) ) ;
INV     gate8416  (.A(g19210), .Z(g23879) ) ;
INV     gate8417  (.A(g19210), .Z(g23880) ) ;
INV     gate8418  (.A(g19277), .Z(g23881) ) ;
INV     gate8419  (.A(g19277), .Z(g23882) ) ;
INV     gate8420  (.A(g21468), .Z(g23886) ) ;
INV     gate8421  (.A(g18997), .Z(g23887) ) ;
INV     gate8422  (.A(g18997), .Z(g23888) ) ;
INV     gate8423  (.A(g20682), .Z(g23889) ) ;
INV     gate8424  (.A(g19074), .Z(g23893) ) ;
INV     gate8425  (.A(g19074), .Z(g23894) ) ;
INV     gate8426  (.A(g19147), .Z(g23895) ) ;
INV     gate8427  (.A(g19210), .Z(g23896) ) ;
INV     gate8428  (.A(g19210), .Z(g23897) ) ;
INV     gate8429  (.A(g19277), .Z(g23898) ) ;
INV     gate8430  (.A(g19277), .Z(g23899) ) ;
INV     gate8431  (.A(g21468), .Z(g23902) ) ;
INV     gate8432  (.A(g18997), .Z(g23903) ) ;
INV     gate8433  (.A(g18997), .Z(g23904) ) ;
INV     gate8434  (.A(g21514), .Z(g23905) ) ;
INV     gate8435  (.A(g19074), .Z(g23906) ) ;
INV     gate8436  (.A(g19074), .Z(g23907) ) ;
INV     gate8437  (.A(g20739), .Z(g23908) ) ;
INV     gate8438  (.A(g19147), .Z(g23912) ) ;
INV     gate8439  (.A(g19147), .Z(g23913) ) ;
INV     gate8440  (.A(g19210), .Z(g23914) ) ;
INV     gate8441  (.A(g19277), .Z(g23915) ) ;
INV     gate8442  (.A(g19277), .Z(g23916) ) ;
INV     gate8443  (.A(g18997), .Z(g23922) ) ;
INV     gate8444  (.A(g18997), .Z(g23923) ) ;
INV     gate8445  (.A(g18997), .Z(g23924) ) ;
INV     gate8446  (.A(g21514), .Z(g23925) ) ;
INV     gate8447  (.A(g19074), .Z(g23926) ) ;
INV     gate8448  (.A(g19074), .Z(g23927) ) ;
INV     gate8449  (.A(g21562), .Z(g23928) ) ;
INV     gate8450  (.A(g19147), .Z(g23929) ) ;
INV     gate8451  (.A(g19147), .Z(g23930) ) ;
INV     gate8452  (.A(g20875), .Z(g23931) ) ;
INV     gate8453  (.A(g19210), .Z(g23935) ) ;
INV     gate8454  (.A(g19210), .Z(g23936) ) ;
INV     gate8455  (.A(g19277), .Z(g23937) ) ;
INV     gate8456  (.A(g18997), .Z(g23938) ) ;
INV     gate8457  (.A(g19074), .Z(g23939) ) ;
INV     gate8458  (.A(g19074), .Z(g23940) ) ;
INV     gate8459  (.A(g19074), .Z(g23941) ) ;
INV     gate8460  (.A(g21562), .Z(g23942) ) ;
INV     gate8461  (.A(g19147), .Z(g23943) ) ;
INV     gate8462  (.A(g19147), .Z(g23944) ) ;
INV     gate8463  (.A(g21611), .Z(g23945) ) ;
INV     gate8464  (.A(g19210), .Z(g23946) ) ;
INV     gate8465  (.A(g19210), .Z(g23947) ) ;
INV     gate8466  (.A(g21012), .Z(g23948) ) ;
INV     gate8467  (.A(g19277), .Z(g23952) ) ;
INV     gate8468  (.A(g19277), .Z(g23953) ) ;
INV     gate8469  (.A(g20682), .Z(II23099) ) ;
INV     gate8470  (.A(II23099), .Z(g23954) ) ;
INV     gate8471  (.A(g19074), .Z(g23961) ) ;
INV     gate8472  (.A(g19147), .Z(g23962) ) ;
INV     gate8473  (.A(g19147), .Z(g23963) ) ;
INV     gate8474  (.A(g19147), .Z(g23964) ) ;
INV     gate8475  (.A(g21611), .Z(g23965) ) ;
INV     gate8476  (.A(g19210), .Z(g23966) ) ;
INV     gate8477  (.A(g19210), .Z(g23967) ) ;
INV     gate8478  (.A(g18833), .Z(g23968) ) ;
INV     gate8479  (.A(g19277), .Z(g23969) ) ;
INV     gate8480  (.A(g19277), .Z(g23970) ) ;
INV     gate8481  (.A(g20751), .Z(g23971) ) ;
INV     gate8482  (.A(g19147), .Z(g23982) ) ;
INV     gate8483  (.A(g19210), .Z(g23983) ) ;
INV     gate8484  (.A(g19210), .Z(g23984) ) ;
INV     gate8485  (.A(g19210), .Z(g23985) ) ;
INV     gate8486  (.A(g18833), .Z(g23986) ) ;
INV     gate8487  (.A(g19277), .Z(g23987) ) ;
INV     gate8488  (.A(g19277), .Z(g23988) ) ;
INV     gate8489  (.A(g19210), .Z(g23992) ) ;
INV     gate8490  (.A(g19277), .Z(g23993) ) ;
INV     gate8491  (.A(g19277), .Z(g23994) ) ;
INV     gate8492  (.A(g19277), .Z(g23995) ) ;
INV     gate8493  (.A(g21468), .Z(g23999) ) ;
INV     gate8494  (.A(g19277), .Z(g24000) ) ;
INV     gate8495  (.A(g21514), .Z(g24003) ) ;
INV     gate8496  (.A(g19061), .Z(II23149) ) ;
INV     gate8497  (.A(II23149), .Z(g24005) ) ;
INV     gate8498  (.A(g21562), .Z(g24010) ) ;
INV     gate8499  (.A(g21611), .Z(g24013) ) ;
INV     gate8500  (.A(g18833), .Z(g24017) ) ;
INV     gate8501  (.A(g19968), .Z(g24019) ) ;
INV     gate8502  (.A(g20014), .Z(g24020) ) ;
INV     gate8503  (.A(g20841), .Z(g24021) ) ;
INV     gate8504  (.A(g20982), .Z(g24022) ) ;
INV     gate8505  (.A(g21127), .Z(g24023) ) ;
INV     gate8506  (.A(g21193), .Z(g24024) ) ;
INV     gate8507  (.A(g21256), .Z(g24025) ) ;
INV     gate8508  (.A(g19919), .Z(g24026) ) ;
INV     gate8509  (.A(g20014), .Z(g24027) ) ;
INV     gate8510  (.A(g20841), .Z(g24028) ) ;
INV     gate8511  (.A(g20982), .Z(g24029) ) ;
INV     gate8512  (.A(g21127), .Z(g24030) ) ;
INV     gate8513  (.A(g21193), .Z(g24031) ) ;
INV     gate8514  (.A(g21256), .Z(g24032) ) ;
INV     gate8515  (.A(g19919), .Z(g24033) ) ;
INV     gate8516  (.A(g19968), .Z(g24034) ) ;
INV     gate8517  (.A(g20841), .Z(g24035) ) ;
INV     gate8518  (.A(g20982), .Z(g24036) ) ;
INV     gate8519  (.A(g21127), .Z(g24037) ) ;
INV     gate8520  (.A(g21193), .Z(g24038) ) ;
INV     gate8521  (.A(g21256), .Z(g24039) ) ;
INV     gate8522  (.A(g19919), .Z(g24040) ) ;
INV     gate8523  (.A(g19968), .Z(g24041) ) ;
INV     gate8524  (.A(g20014), .Z(g24042) ) ;
INV     gate8525  (.A(g20982), .Z(g24043) ) ;
INV     gate8526  (.A(g21127), .Z(g24044) ) ;
INV     gate8527  (.A(g21193), .Z(g24045) ) ;
INV     gate8528  (.A(g21256), .Z(g24046) ) ;
INV     gate8529  (.A(g19919), .Z(g24047) ) ;
INV     gate8530  (.A(g19968), .Z(g24048) ) ;
INV     gate8531  (.A(g20014), .Z(g24049) ) ;
INV     gate8532  (.A(g20841), .Z(g24050) ) ;
INV     gate8533  (.A(g21127), .Z(g24051) ) ;
INV     gate8534  (.A(g21193), .Z(g24052) ) ;
INV     gate8535  (.A(g21256), .Z(g24053) ) ;
INV     gate8536  (.A(g19919), .Z(g24054) ) ;
INV     gate8537  (.A(g19968), .Z(g24055) ) ;
INV     gate8538  (.A(g20014), .Z(g24056) ) ;
INV     gate8539  (.A(g20841), .Z(g24057) ) ;
INV     gate8540  (.A(g20982), .Z(g24058) ) ;
INV     gate8541  (.A(g21193), .Z(g24059) ) ;
INV     gate8542  (.A(g21256), .Z(g24060) ) ;
INV     gate8543  (.A(g19919), .Z(g24061) ) ;
INV     gate8544  (.A(g19968), .Z(g24062) ) ;
INV     gate8545  (.A(g20014), .Z(g24063) ) ;
INV     gate8546  (.A(g20841), .Z(g24064) ) ;
INV     gate8547  (.A(g20982), .Z(g24065) ) ;
INV     gate8548  (.A(g21127), .Z(g24066) ) ;
INV     gate8549  (.A(g21256), .Z(g24067) ) ;
INV     gate8550  (.A(g19919), .Z(g24068) ) ;
INV     gate8551  (.A(g19968), .Z(g24069) ) ;
INV     gate8552  (.A(g20014), .Z(g24070) ) ;
INV     gate8553  (.A(g20841), .Z(g24071) ) ;
INV     gate8554  (.A(g20982), .Z(g24072) ) ;
INV     gate8555  (.A(g21127), .Z(g24073) ) ;
INV     gate8556  (.A(g21193), .Z(g24074) ) ;
INV     gate8557  (.A(g19935), .Z(g24075) ) ;
INV     gate8558  (.A(g19984), .Z(g24076) ) ;
INV     gate8559  (.A(g20720), .Z(g24077) ) ;
INV     gate8560  (.A(g20857), .Z(g24078) ) ;
INV     gate8561  (.A(g20998), .Z(g24079) ) ;
INV     gate8562  (.A(g21143), .Z(g24080) ) ;
INV     gate8563  (.A(g21209), .Z(g24081) ) ;
INV     gate8564  (.A(g19890), .Z(g24082) ) ;
INV     gate8565  (.A(g19984), .Z(g24083) ) ;
INV     gate8566  (.A(g20720), .Z(g24084) ) ;
INV     gate8567  (.A(g20857), .Z(g24085) ) ;
INV     gate8568  (.A(g20998), .Z(g24086) ) ;
INV     gate8569  (.A(g21143), .Z(g24087) ) ;
INV     gate8570  (.A(g21209), .Z(g24088) ) ;
INV     gate8571  (.A(g19890), .Z(g24089) ) ;
INV     gate8572  (.A(g19935), .Z(g24090) ) ;
INV     gate8573  (.A(g20720), .Z(g24091) ) ;
INV     gate8574  (.A(g20857), .Z(g24092) ) ;
INV     gate8575  (.A(g20998), .Z(g24093) ) ;
INV     gate8576  (.A(g21143), .Z(g24094) ) ;
INV     gate8577  (.A(g21209), .Z(g24095) ) ;
INV     gate8578  (.A(g19890), .Z(g24096) ) ;
INV     gate8579  (.A(g19935), .Z(g24097) ) ;
INV     gate8580  (.A(g19984), .Z(g24098) ) ;
INV     gate8581  (.A(g20720), .Z(g24099) ) ;
INV     gate8582  (.A(g20857), .Z(g24100) ) ;
INV     gate8583  (.A(g20998), .Z(g24101) ) ;
INV     gate8584  (.A(g21143), .Z(g24102) ) ;
INV     gate8585  (.A(g21209), .Z(g24103) ) ;
INV     gate8586  (.A(g19890), .Z(g24104) ) ;
INV     gate8587  (.A(g19935), .Z(g24105) ) ;
INV     gate8588  (.A(g19984), .Z(g24106) ) ;
INV     gate8589  (.A(g20857), .Z(g24107) ) ;
INV     gate8590  (.A(g20998), .Z(g24108) ) ;
INV     gate8591  (.A(g21143), .Z(g24109) ) ;
INV     gate8592  (.A(g21209), .Z(g24110) ) ;
INV     gate8593  (.A(g19890), .Z(g24111) ) ;
INV     gate8594  (.A(g19935), .Z(g24112) ) ;
INV     gate8595  (.A(g19984), .Z(g24113) ) ;
INV     gate8596  (.A(g20720), .Z(g24114) ) ;
INV     gate8597  (.A(g20998), .Z(g24115) ) ;
INV     gate8598  (.A(g21143), .Z(g24116) ) ;
INV     gate8599  (.A(g21209), .Z(g24117) ) ;
INV     gate8600  (.A(g19890), .Z(g24118) ) ;
INV     gate8601  (.A(g19935), .Z(g24119) ) ;
INV     gate8602  (.A(g19984), .Z(g24120) ) ;
INV     gate8603  (.A(g20720), .Z(g24121) ) ;
INV     gate8604  (.A(g20857), .Z(g24122) ) ;
INV     gate8605  (.A(g21143), .Z(g24123) ) ;
INV     gate8606  (.A(g21209), .Z(g24124) ) ;
INV     gate8607  (.A(g19890), .Z(g24125) ) ;
INV     gate8608  (.A(g19935), .Z(g24126) ) ;
INV     gate8609  (.A(g19984), .Z(g24127) ) ;
INV     gate8610  (.A(g20720), .Z(g24128) ) ;
INV     gate8611  (.A(g20857), .Z(g24129) ) ;
INV     gate8612  (.A(g20998), .Z(g24130) ) ;
INV     gate8613  (.A(g21209), .Z(g24131) ) ;
INV     gate8614  (.A(g19890), .Z(g24132) ) ;
INV     gate8615  (.A(g19935), .Z(g24133) ) ;
INV     gate8616  (.A(g19984), .Z(g24134) ) ;
INV     gate8617  (.A(g20720), .Z(g24135) ) ;
INV     gate8618  (.A(g20857), .Z(g24136) ) ;
INV     gate8619  (.A(g20998), .Z(g24137) ) ;
INV     gate8620  (.A(g21143), .Z(g24138) ) ;
INV     gate8621  (.A(g19422), .Z(g24146) ) ;
INV     gate8622  (.A(g19402), .Z(g24147) ) ;
INV     gate8623  (.A(g19338), .Z(g24149) ) ;
INV     gate8624  (.A(g19268), .Z(g24150) ) ;
INV     gate8625  (.A(g21665), .Z(II23300) ) ;
INV     gate8626  (.A(II23300), .Z(g24152) ) ;
INV     gate8627  (.A(g21669), .Z(II23303) ) ;
INV     gate8628  (.A(II23303), .Z(g24153) ) ;
INV     gate8629  (.A(g21673), .Z(II23306) ) ;
INV     gate8630  (.A(II23306), .Z(g24154) ) ;
INV     gate8631  (.A(g21677), .Z(II23309) ) ;
INV     gate8632  (.A(II23309), .Z(g24155) ) ;
INV     gate8633  (.A(g21681), .Z(II23312) ) ;
INV     gate8634  (.A(II23312), .Z(g24156) ) ;
INV     gate8635  (.A(g21685), .Z(II23315) ) ;
INV     gate8636  (.A(II23315), .Z(g24157) ) ;
INV     gate8637  (.A(g21689), .Z(II23318) ) ;
INV     gate8638  (.A(II23318), .Z(g24158) ) ;
INV     gate8639  (.A(g21693), .Z(II23321) ) ;
INV     gate8640  (.A(II23321), .Z(g24159) ) ;
INV     gate8641  (.A(g21697), .Z(II23324) ) ;
INV     gate8642  (.A(II23324), .Z(g24160) ) ;
INV     gate8643  (.A(g22647), .Z(II23327) ) ;
INV     gate8644  (.A(g22658), .Z(II23330) ) ;
INV     gate8645  (.A(g22683), .Z(II23333) ) ;
INV     gate8646  (.A(g22721), .Z(II23336) ) ;
INV     gate8647  (.A(g23232), .Z(II23339) ) ;
INV     gate8648  (.A(g23299), .Z(II23342) ) ;
INV     gate8649  (.A(g23320), .Z(II23345) ) ;
INV     gate8650  (.A(g23384), .Z(II23348) ) ;
INV     gate8651  (.A(g23263), .Z(II23351) ) ;
INV     gate8652  (.A(g23277), .Z(II23354) ) ;
INV     gate8653  (.A(g23359), .Z(II23357) ) ;
INV     gate8654  (.A(g23360), .Z(II23360) ) ;
INV     gate8655  (.A(g23385), .Z(II23363) ) ;
INV     gate8656  (.A(g23321), .Z(II23366) ) ;
INV     gate8657  (.A(g23347), .Z(II23369) ) ;
INV     gate8658  (.A(g23361), .Z(II23372) ) ;
INV     gate8659  (.A(g23403), .Z(II23375) ) ;
INV     gate8660  (.A(g23426), .Z(II23378) ) ;
INV     gate8661  (.A(g23322), .Z(II23381) ) ;
INV     gate8662  (.A(g23362), .Z(II23384) ) ;
INV     gate8663  (.A(g23394), .Z(II23387) ) ;
INV     gate8664  (.A(g23395), .Z(II23390) ) ;
INV     gate8665  (.A(g23414), .Z(II23393) ) ;
INV     gate8666  (.A(g23427), .Z(II23396) ) ;
INV     gate8667  (.A(g23450), .Z(II23399) ) ;
INV     gate8668  (.A(g22594), .Z(g24356) ) ;
NAND2   gate8669  (.A(g1252), .B(g19140), .Z(g22325) ) ;
INV     gate8670  (.A(g22325), .Z(g24357) ) ;
INV     gate8671  (.A(g22550), .Z(g24358) ) ;
INV     gate8672  (.A(g22550), .Z(g24359) ) ;
INV     gate8673  (.A(g22228), .Z(g24360) ) ;
NAND2   gate8674  (.A(g9104), .B(g20154), .Z(g22885) ) ;
INV     gate8675  (.A(g22885), .Z(g24361) ) ;
INV     gate8676  (.A(g22722), .Z(g24364) ) ;
INV     gate8677  (.A(g22594), .Z(g24365) ) ;
INV     gate8678  (.A(g22594), .Z(g24366) ) ;
INV     gate8679  (.A(g22550), .Z(g24367) ) ;
INV     gate8680  (.A(g22228), .Z(g24368) ) ;
INV     gate8681  (.A(g22885), .Z(g24372) ) ;
NAND2   gate8682  (.A(g9104), .B(g20175), .Z(g22908) ) ;
INV     gate8683  (.A(g22908), .Z(g24373) ) ;
INV     gate8684  (.A(g22722), .Z(g24375) ) ;
INV     gate8685  (.A(g22722), .Z(g24376) ) ;
INV     gate8686  (.A(g22594), .Z(g24377) ) ;
INV     gate8687  (.A(g22550), .Z(g24379) ) ;
INV     gate8688  (.A(g22885), .Z(g24384) ) ;
INV     gate8689  (.A(g22908), .Z(g24385) ) ;
INV     gate8690  (.A(g22594), .Z(g24386) ) ;
INV     gate8691  (.A(g22885), .Z(g24388) ) ;
INV     gate8692  (.A(g22908), .Z(g24389) ) ;
INV     gate8693  (.A(g22228), .Z(g24394) ) ;
INV     gate8694  (.A(g22885), .Z(g24396) ) ;
INV     gate8695  (.A(g22908), .Z(g24397) ) ;
INV     gate8696  (.A(g22908), .Z(g24404) ) ;
INV     gate8697  (.A(g22722), .Z(g24405) ) ;
INV     gate8698  (.A(g22594), .Z(g24407) ) ;
INV     gate8699  (.A(g22171), .Z(g24417) ) ;
INV     gate8700  (.A(g22722), .Z(g24418) ) ;
INV     gate8701  (.A(g22722), .Z(g24419) ) ;
INV     gate8702  (.A(g22722), .Z(g24424) ) ;
INV     gate8703  (.A(g22722), .Z(g24425) ) ;
INV     gate8704  (.A(g22722), .Z(g24426) ) ;
INV     gate8705  (.A(g22722), .Z(g24428) ) ;
INV     gate8706  (.A(g22722), .Z(g24429) ) ;
INV     gate8707  (.A(g22722), .Z(g24431) ) ;
NOR2    gate8708  (.A(g7733), .B(g19506), .Z(g22654) ) ;
INV     gate8709  (.A(g22654), .Z(g24437) ) ;
INV     gate8710  (.A(g22722), .Z(g24438) ) ;
INV     gate8711  (.A(g22722), .Z(g24452) ) ;
INV     gate8712  (.A(g23578), .Z(g24463) ) ;
INV     gate8713  (.A(g23202), .Z(II23671) ) ;
INV     gate8714  (.A(II23671), .Z(g24466) ) ;
INV     gate8715  (.A(g23620), .Z(g24474) ) ;
INV     gate8716  (.A(g23219), .Z(II23680) ) ;
INV     gate8717  (.A(II23680), .Z(g24477) ) ;
INV     gate8718  (.A(g23230), .Z(II23684) ) ;
INV     gate8719  (.A(II23684), .Z(g24481) ) ;
INV     gate8720  (.A(g23244), .Z(II23688) ) ;
INV     gate8721  (.A(II23688), .Z(g24483) ) ;
INV     gate8722  (.A(g23252), .Z(II23694) ) ;
INV     gate8723  (.A(II23694), .Z(g24489) ) ;
INV     gate8724  (.A(g22594), .Z(g24490) ) ;
AND2    gate8725  (.A(g18918), .B(g9104), .Z(g22689) ) ;
INV     gate8726  (.A(g22689), .Z(g24505) ) ;
INV     gate8727  (.A(g23192), .Z(II23711) ) ;
INV     gate8728  (.A(II23711), .Z(g24506) ) ;
INV     gate8729  (.A(g22689), .Z(g24509) ) ;
INV     gate8730  (.A(g22689), .Z(g24515) ) ;
AND2    gate8731  (.A(g20114), .B(g9104), .Z(g22670) ) ;
INV     gate8732  (.A(g22670), .Z(g24516) ) ;
INV     gate8733  (.A(g22689), .Z(g24522) ) ;
AND2    gate8734  (.A(g20136), .B(g9104), .Z(g22876) ) ;
INV     gate8735  (.A(g22876), .Z(g24524) ) ;
INV     gate8736  (.A(g22670), .Z(g24525) ) ;
AND2    gate8737  (.A(g9104), .B(g20219), .Z(g22942) ) ;
INV     gate8738  (.A(g22942), .Z(g24526) ) ;
INV     gate8739  (.A(g22670), .Z(g24527) ) ;
INV     gate8740  (.A(g22876), .Z(g24533) ) ;
INV     gate8741  (.A(g22670), .Z(g24534) ) ;
INV     gate8742  (.A(g22942), .Z(g24535) ) ;
INV     gate8743  (.A(g22942), .Z(g24540) ) ;
INV     gate8744  (.A(g22942), .Z(g24548) ) ;
INV     gate8745  (.A(g22942), .Z(g24560) ) ;
INV     gate8746  (.A(g22942), .Z(g24568) ) ;
INV     gate8747  (.A(g22942), .Z(g24571) ) ;
NAND2   gate8748  (.A(g20887), .B(g10721), .Z(g23067) ) ;
INV     gate8749  (.A(g23067), .Z(g24579) ) ;
NOR2    gate8750  (.A(g16313), .B(g19887), .Z(g23063) ) ;
INV     gate8751  (.A(g23063), .Z(g24585) ) ;
INV     gate8752  (.A(g23067), .Z(g24586) ) ;
NAND2   gate8753  (.A(g21024), .B(g10733), .Z(g23112) ) ;
INV     gate8754  (.A(g23112), .Z(g24587) ) ;
NOR2    gate8755  (.A(g16424), .B(g19932), .Z(g23108) ) ;
INV     gate8756  (.A(g23108), .Z(g24603) ) ;
INV     gate8757  (.A(g23112), .Z(g24604) ) ;
NAND2   gate8758  (.A(g21163), .B(g10756), .Z(g23139) ) ;
INV     gate8759  (.A(g23139), .Z(g24605) ) ;
AND2    gate8760  (.A(g19128), .B(g9104), .Z(g23076) ) ;
INV     gate8761  (.A(g23076), .Z(g24623) ) ;
NOR2    gate8762  (.A(g16476), .B(g19981), .Z(g23135) ) ;
INV     gate8763  (.A(g23135), .Z(g24625) ) ;
INV     gate8764  (.A(g23139), .Z(g24626) ) ;
AND2    gate8765  (.A(g19128), .B(g9104), .Z(g23121) ) ;
INV     gate8766  (.A(g23121), .Z(g24636) ) ;
AND2    gate8767  (.A(g19128), .B(g9104), .Z(g23148) ) ;
INV     gate8768  (.A(g23148), .Z(g24648) ) ;
INV     gate8769  (.A(g23067), .Z(g24655) ) ;
INV     gate8770  (.A(g23067), .Z(g24665) ) ;
INV     gate8771  (.A(g23112), .Z(g24667) ) ;
INV     gate8772  (.A(g23112), .Z(g24683) ) ;
INV     gate8773  (.A(g23139), .Z(g24685) ) ;
NAND2   gate8774  (.A(g482), .B(g20000), .Z(g23047) ) ;
INV     gate8775  (.A(g23047), .Z(g24699) ) ;
INV     gate8776  (.A(g23139), .Z(g24711) ) ;
INV     gate8777  (.A(g22182), .Z(g24718) ) ;
NOR3    gate8778  (.A(g16581), .B(g19462), .C(g10685), .Z(g23042) ) ;
INV     gate8779  (.A(g23042), .Z(g24732) ) ;
INV     gate8780  (.A(g22202), .Z(g24744) ) ;
INV     gate8781  (.A(g22763), .Z(g24756) ) ;
INV     gate8782  (.A(g23003), .Z(g24759) ) ;
INV     gate8783  (.A(g22763), .Z(g24770) ) ;
NAND2   gate8784  (.A(g6875), .B(g20887), .Z(g23286) ) ;
INV     gate8785  (.A(g23286), .Z(g24778) ) ;
NAND2   gate8786  (.A(g6905), .B(g21024), .Z(g23309) ) ;
INV     gate8787  (.A(g23309), .Z(g24789) ) ;
NAND2   gate8788  (.A(g12185), .B(g19462), .Z(g23850) ) ;
INV     gate8789  (.A(g23850), .Z(g24791) ) ;
NAND2   gate8790  (.A(g6928), .B(g21163), .Z(g23342) ) ;
INV     gate8791  (.A(g23342), .Z(g24795) ) ;
INV     gate8792  (.A(g23191), .Z(g24818) ) ;
INV     gate8793  (.A(g22182), .Z(II23998) ) ;
INV     gate8794  (.A(II23998), .Z(g24819) ) ;
NOR3    gate8795  (.A(g10685), .B(g19462), .C(g16488), .Z(g23204) ) ;
INV     gate8796  (.A(g23204), .Z(g24825) ) ;
INV     gate8797  (.A(g22182), .Z(II24008) ) ;
INV     gate8798  (.A(II24008), .Z(g24836) ) ;
AND2    gate8799  (.A(g676), .B(g20375), .Z(g23436) ) ;
INV     gate8800  (.A(g23436), .Z(g24839) ) ;
INV     gate8801  (.A(g22182), .Z(II24022) ) ;
INV     gate8802  (.A(II24022), .Z(g24850) ) ;
INV     gate8803  (.A(g22202), .Z(II24038) ) ;
INV     gate8804  (.A(II24038), .Z(g24866) ) ;
INV     gate8805  (.A(g22182), .Z(II24041) ) ;
INV     gate8806  (.A(II24041), .Z(g24869) ) ;
INV     gate8807  (.A(g23231), .Z(g24891) ) ;
INV     gate8808  (.A(g22202), .Z(II24060) ) ;
INV     gate8809  (.A(II24060), .Z(g24893) ) ;
INV     gate8810  (.A(g22360), .Z(II24078) ) ;
INV     gate8811  (.A(II24078), .Z(g24911) ) ;
INV     gate8812  (.A(g22409), .Z(II24089) ) ;
INV     gate8813  (.A(II24089), .Z(g24920) ) ;
OR2     gate8814  (.A(g9194), .B(g20905), .Z(g23716) ) ;
INV     gate8815  (.A(g23716), .Z(g24960) ) ;
AND3    gate8816  (.A(g9354), .B(g9285), .C(g21287), .Z(g22342) ) ;
INV     gate8817  (.A(g22342), .Z(g24963) ) ;
AND2    gate8818  (.A(g20196), .B(g14219), .Z(g23009) ) ;
INV     gate8819  (.A(g23009), .Z(II24128) ) ;
INV     gate8820  (.A(II24128), .Z(g24964) ) ;
INV     gate8821  (.A(g22763), .Z(g24966) ) ;
NAND2   gate8822  (.A(g20682), .B(g11111), .Z(g23590) ) ;
INV     gate8823  (.A(g23590), .Z(g24971) ) ;
INV     gate8824  (.A(g22342), .Z(g24978) ) ;
AND3    gate8825  (.A(g9354), .B(g7717), .C(g20783), .Z(g22369) ) ;
INV     gate8826  (.A(g22369), .Z(g24979) ) ;
AND3    gate8827  (.A(g9354), .B(g9285), .C(g20784), .Z(g22384) ) ;
INV     gate8828  (.A(g22384), .Z(g24980) ) ;
INV     gate8829  (.A(g22763), .Z(g24981) ) ;
INV     gate8830  (.A(g22763), .Z(g24982) ) ;
NOR2    gate8831  (.A(g17284), .B(g20717), .Z(g23586) ) ;
INV     gate8832  (.A(g23586), .Z(g24985) ) ;
INV     gate8833  (.A(g23590), .Z(g24986) ) ;
NAND2   gate8834  (.A(g20739), .B(g11123), .Z(g23630) ) ;
INV     gate8835  (.A(g23630), .Z(g24987) ) ;
INV     gate8836  (.A(g22369), .Z(g24991) ) ;
AND3    gate8837  (.A(g7753), .B(g9285), .C(g21186), .Z(g22417) ) ;
INV     gate8838  (.A(g22417), .Z(g24992) ) ;
INV     gate8839  (.A(g22384), .Z(g24993) ) ;
AND3    gate8840  (.A(g9354), .B(g7717), .C(g21187), .Z(g22432) ) ;
INV     gate8841  (.A(g22432), .Z(g24994) ) ;
INV     gate8842  (.A(g22763), .Z(g24995) ) ;
INV     gate8843  (.A(g22763), .Z(g24996) ) ;
NOR2    gate8844  (.A(g17309), .B(g20854), .Z(g23626) ) ;
INV     gate8845  (.A(g23626), .Z(g24999) ) ;
INV     gate8846  (.A(g23630), .Z(g25000) ) ;
NAND2   gate8847  (.A(g20875), .B(g11139), .Z(g23666) ) ;
INV     gate8848  (.A(g23666), .Z(g25001) ) ;
INV     gate8849  (.A(g22417), .Z(g25006) ) ;
AND3    gate8850  (.A(g7753), .B(g7717), .C(g21288), .Z(g22457) ) ;
INV     gate8851  (.A(g22457), .Z(g25007) ) ;
INV     gate8852  (.A(g22432), .Z(g25008) ) ;
AND3    gate8853  (.A(g7753), .B(g9285), .C(g21289), .Z(g22472) ) ;
INV     gate8854  (.A(g22472), .Z(g25009) ) ;
INV     gate8855  (.A(g22763), .Z(g25011) ) ;
AND2    gate8856  (.A(g19050), .B(g9104), .Z(g23599) ) ;
INV     gate8857  (.A(g23599), .Z(g25013) ) ;
NOR2    gate8858  (.A(g17393), .B(g20995), .Z(g23662) ) ;
INV     gate8859  (.A(g23662), .Z(g25015) ) ;
INV     gate8860  (.A(g23666), .Z(g25016) ) ;
NAND2   gate8861  (.A(g21012), .B(g11160), .Z(g23699) ) ;
INV     gate8862  (.A(g23699), .Z(g25017) ) ;
INV     gate8863  (.A(g22457), .Z(g25023) ) ;
INV     gate8864  (.A(g22472), .Z(g25024) ) ;
AND3    gate8865  (.A(g7753), .B(g7717), .C(g21334), .Z(g22498) ) ;
INV     gate8866  (.A(g22498), .Z(g25025) ) ;
INV     gate8867  (.A(g22360), .Z(II24191) ) ;
INV     gate8868  (.A(II24191), .Z(g25027) ) ;
AND2    gate8869  (.A(g19050), .B(g9104), .Z(g23639) ) ;
INV     gate8870  (.A(g23639), .Z(g25032) ) ;
NOR2    gate8871  (.A(g17420), .B(g21140), .Z(g23695) ) ;
INV     gate8872  (.A(g23695), .Z(g25034) ) ;
INV     gate8873  (.A(g23699), .Z(g25035) ) ;
NAND2   gate8874  (.A(g20751), .B(g11178), .Z(g23733) ) ;
INV     gate8875  (.A(g23733), .Z(g25036) ) ;
INV     gate8876  (.A(g22498), .Z(g25039) ) ;
AND2    gate8877  (.A(g19050), .B(g9104), .Z(g23675) ) ;
INV     gate8878  (.A(g23675), .Z(g25044) ) ;
NOR2    gate8879  (.A(g17482), .B(g21206), .Z(g23729) ) ;
INV     gate8880  (.A(g23729), .Z(g25046) ) ;
INV     gate8881  (.A(g23733), .Z(g25047) ) ;
INV     gate8882  (.A(g22360), .Z(II24215) ) ;
INV     gate8883  (.A(II24215), .Z(g25051) ) ;
INV     gate8884  (.A(g23590), .Z(g25055) ) ;
AND2    gate8885  (.A(g19050), .B(g9104), .Z(g23708) ) ;
INV     gate8886  (.A(g23708), .Z(g25060) ) ;
INV     gate8887  (.A(g22409), .Z(II24228) ) ;
INV     gate8888  (.A(II24228), .Z(g25064) ) ;
INV     gate8889  (.A(g23590), .Z(g25070) ) ;
INV     gate8890  (.A(g23630), .Z(g25072) ) ;
INV     gate8891  (.A(g23823), .Z(II24237) ) ;
INV     gate8892  (.A(II24237), .Z(g25073) ) ;
AND2    gate8893  (.A(g19128), .B(g9104), .Z(g23742) ) ;
INV     gate8894  (.A(g23742), .Z(g25080) ) ;
INV     gate8895  (.A(g22342), .Z(g25081) ) ;
INV     gate8896  (.A(g22342), .Z(g25082) ) ;
NAND2   gate8897  (.A(g2741), .B(g21062), .Z(g23782) ) ;
INV     gate8898  (.A(g23782), .Z(g25083) ) ;
INV     gate8899  (.A(g23630), .Z(g25090) ) ;
INV     gate8900  (.A(g23666), .Z(g25092) ) ;
INV     gate8901  (.A(g22342), .Z(g25097) ) ;
INV     gate8902  (.A(g22369), .Z(g25098) ) ;
INV     gate8903  (.A(g22369), .Z(g25099) ) ;
INV     gate8904  (.A(g22384), .Z(g25100) ) ;
INV     gate8905  (.A(g22384), .Z(g25101) ) ;
INV     gate8906  (.A(g23666), .Z(g25109) ) ;
INV     gate8907  (.A(g23699), .Z(g25111) ) ;
INV     gate8908  (.A(g23440), .Z(II24278) ) ;
INV     gate8909  (.A(g23440), .Z(II24281) ) ;
INV     gate8910  (.A(II24281), .Z(g25115) ) ;
INV     gate8911  (.A(g22369), .Z(g25116) ) ;
INV     gate8912  (.A(g22417), .Z(g25117) ) ;
INV     gate8913  (.A(g22417), .Z(g25118) ) ;
INV     gate8914  (.A(g22384), .Z(g25119) ) ;
INV     gate8915  (.A(g22432), .Z(g25120) ) ;
INV     gate8916  (.A(g22432), .Z(g25121) ) ;
INV     gate8917  (.A(g23699), .Z(g25131) ) ;
INV     gate8918  (.A(g23733), .Z(g25133) ) ;
INV     gate8919  (.A(g22417), .Z(g25134) ) ;
INV     gate8920  (.A(g22457), .Z(g25135) ) ;
INV     gate8921  (.A(g22457), .Z(g25136) ) ;
INV     gate8922  (.A(g22432), .Z(g25137) ) ;
INV     gate8923  (.A(g22472), .Z(g25138) ) ;
INV     gate8924  (.A(g22472), .Z(g25139) ) ;
INV     gate8925  (.A(g22228), .Z(g25140) ) ;
INV     gate8926  (.A(g23733), .Z(g25153) ) ;
INV     gate8927  (.A(g22457), .Z(g25154) ) ;
INV     gate8928  (.A(g22472), .Z(g25155) ) ;
INV     gate8929  (.A(g22498), .Z(g25156) ) ;
INV     gate8930  (.A(g22498), .Z(g25157) ) ;
INV     gate8931  (.A(g22228), .Z(g25158) ) ;
INV     gate8932  (.A(g22976), .Z(II24331) ) ;
INV     gate8933  (.A(g22976), .Z(II24334) ) ;
INV     gate8934  (.A(II24334), .Z(g25168) ) ;
INV     gate8935  (.A(g22763), .Z(g25169) ) ;
INV     gate8936  (.A(g22498), .Z(g25170) ) ;
INV     gate8937  (.A(g22228), .Z(g25171) ) ;
NAND2   gate8938  (.A(g7004), .B(g20682), .Z(g23890) ) ;
INV     gate8939  (.A(g23890), .Z(g25174) ) ;
INV     gate8940  (.A(g23529), .Z(g25180) ) ;
INV     gate8941  (.A(g22763), .Z(g25182) ) ;
INV     gate8942  (.A(g22763), .Z(g25183) ) ;
INV     gate8943  (.A(g22763), .Z(g25184) ) ;
INV     gate8944  (.A(g22228), .Z(g25185) ) ;
NAND2   gate8945  (.A(g7028), .B(g20739), .Z(g23909) ) ;
INV     gate8946  (.A(g23909), .Z(g25188) ) ;
INV     gate8947  (.A(g22763), .Z(g25193) ) ;
INV     gate8948  (.A(g22763), .Z(g25194) ) ;
INV     gate8949  (.A(g22763), .Z(g25195) ) ;
INV     gate8950  (.A(g22763), .Z(g25196) ) ;
AND2    gate8951  (.A(g9104), .B(g19200), .Z(g23958) ) ;
INV     gate8952  (.A(g23958), .Z(g25197) ) ;
INV     gate8953  (.A(g22228), .Z(g25198) ) ;
NAND2   gate8954  (.A(g7051), .B(g20875), .Z(g23932) ) ;
INV     gate8955  (.A(g23932), .Z(g25202) ) ;
INV     gate8956  (.A(g23613), .Z(g25206) ) ;
INV     gate8957  (.A(g22763), .Z(g25208) ) ;
INV     gate8958  (.A(g22763), .Z(g25209) ) ;
AND2    gate8959  (.A(g9104), .B(g19050), .Z(g23802) ) ;
INV     gate8960  (.A(g23802), .Z(g25210) ) ;
INV     gate8961  (.A(g22763), .Z(g25211) ) ;
INV     gate8962  (.A(g22763), .Z(g25212) ) ;
AND2    gate8963  (.A(g9104), .B(g19200), .Z(g23293) ) ;
INV     gate8964  (.A(g23293), .Z(g25213) ) ;
INV     gate8965  (.A(g22228), .Z(g25214) ) ;
NAND2   gate8966  (.A(g7074), .B(g21012), .Z(g23949) ) ;
INV     gate8967  (.A(g23949), .Z(g25218) ) ;
INV     gate8968  (.A(g23453), .Z(II24393) ) ;
INV     gate8969  (.A(g23453), .Z(II24396) ) ;
INV     gate8970  (.A(II24396), .Z(g25220) ) ;
INV     gate8971  (.A(g23653), .Z(g25221) ) ;
INV     gate8972  (.A(g23954), .Z(II24400) ) ;
INV     gate8973  (.A(II24400), .Z(g25222) ) ;
INV     gate8974  (.A(g22763), .Z(g25224) ) ;
INV     gate8975  (.A(g23802), .Z(g25225) ) ;
INV     gate8976  (.A(g22763), .Z(g25226) ) ;
INV     gate8977  (.A(g22763), .Z(g25227) ) ;
AND2    gate8978  (.A(g9104), .B(g19128), .Z(g23828) ) ;
INV     gate8979  (.A(g23828), .Z(g25228) ) ;
AND2    gate8980  (.A(g9104), .B(g19200), .Z(g23314) ) ;
INV     gate8981  (.A(g23314), .Z(g25230) ) ;
INV     gate8982  (.A(g22228), .Z(g25231) ) ;
INV     gate8983  (.A(g22228), .Z(g25232) ) ;
NAND2   gate8984  (.A(g7097), .B(g20751), .Z(g23972) ) ;
INV     gate8985  (.A(g23972), .Z(g25239) ) ;
INV     gate8986  (.A(g23650), .Z(g25240) ) ;
INV     gate8987  (.A(g23651), .Z(g25241) ) ;
INV     gate8988  (.A(g23684), .Z(g25242) ) ;
INV     gate8989  (.A(g22763), .Z(g25243) ) ;
INV     gate8990  (.A(g23802), .Z(g25244) ) ;
INV     gate8991  (.A(g22763), .Z(g25245) ) ;
INV     gate8992  (.A(g23828), .Z(g25246) ) ;
INV     gate8993  (.A(g22228), .Z(g25248) ) ;
INV     gate8994  (.A(g22228), .Z(g25249) ) ;
INV     gate8995  (.A(g22763), .Z(II24434) ) ;
INV     gate8996  (.A(II24434), .Z(g25250) ) ;
INV     gate8997  (.A(g22923), .Z(II24445) ) ;
INV     gate8998  (.A(g22923), .Z(II24448) ) ;
INV     gate8999  (.A(II24448), .Z(g25260) ) ;
INV     gate9000  (.A(g22763), .Z(g25262) ) ;
INV     gate9001  (.A(g22763), .Z(g25263) ) ;
INV     gate9002  (.A(g23828), .Z(g25264) ) ;
INV     gate9003  (.A(g22541), .Z(II24455) ) ;
INV     gate9004  (.A(II24455), .Z(g25265) ) ;
INV     gate9005  (.A(g22228), .Z(g25266) ) ;
INV     gate9006  (.A(g22228), .Z(g25267) ) ;
INV     gate9007  (.A(g23715), .Z(g25272) ) ;
NAND3   gate9008  (.A(g572), .B(g21389), .C(g12323), .Z(g23978) ) ;
INV     gate9009  (.A(g23978), .Z(g25273) ) ;
INV     gate9010  (.A(g22763), .Z(g25274) ) ;
INV     gate9011  (.A(g22763), .Z(g25282) ) ;
INV     gate9012  (.A(g22763), .Z(g25283) ) ;
INV     gate9013  (.A(g22546), .Z(II24474) ) ;
INV     gate9014  (.A(II24474), .Z(g25284) ) ;
INV     gate9015  (.A(g22228), .Z(g25286) ) ;
INV     gate9016  (.A(g22228), .Z(g25287) ) ;
INV     gate9017  (.A(g22228), .Z(g25288) ) ;
INV     gate9018  (.A(g22228), .Z(g25289) ) ;
INV     gate9019  (.A(g23745), .Z(g25296) ) ;
INV     gate9020  (.A(g23746), .Z(g25297) ) ;
INV     gate9021  (.A(g23760), .Z(g25298) ) ;
INV     gate9022  (.A(g22763), .Z(g25299) ) ;
INV     gate9023  (.A(g22763), .Z(g25307) ) ;
INV     gate9024  (.A(g22763), .Z(g25308) ) ;
INV     gate9025  (.A(g22763), .Z(g25316) ) ;
INV     gate9026  (.A(g22592), .Z(II24497) ) ;
INV     gate9027  (.A(II24497), .Z(g25322) ) ;
INV     gate9028  (.A(g22228), .Z(g25324) ) ;
INV     gate9029  (.A(g22228), .Z(g25325) ) ;
INV     gate9030  (.A(g22228), .Z(g25326) ) ;
AND2    gate9031  (.A(g13202), .B(g19071), .Z(g22161) ) ;
INV     gate9032  (.A(g22161), .Z(g25327) ) ;
INV     gate9033  (.A(g22763), .Z(g25340) ) ;
INV     gate9034  (.A(g22763), .Z(g25348) ) ;
INV     gate9035  (.A(g22763), .Z(g25356) ) ;
INV     gate9036  (.A(g22228), .Z(g25369) ) ;
INV     gate9037  (.A(g22228), .Z(g25370) ) ;
INV     gate9038  (.A(g23776), .Z(g25380) ) ;
INV     gate9039  (.A(g22763), .Z(g25388) ) ;
INV     gate9040  (.A(g22763), .Z(g25399) ) ;
INV     gate9041  (.A(g22228), .Z(g25409) ) ;
INV     gate9042  (.A(g22228), .Z(g25410) ) ;
INV     gate9043  (.A(g23777), .Z(II24558) ) ;
INV     gate9044  (.A(II24558), .Z(g25423) ) ;
INV     gate9045  (.A(g23800), .Z(g25424) ) ;
INV     gate9046  (.A(g22763), .Z(g25438) ) ;
INV     gate9047  (.A(g22228), .Z(g25451) ) ;
INV     gate9048  (.A(g22228), .Z(g25452) ) ;
INV     gate9049  (.A(g23824), .Z(g25465) ) ;
INV     gate9050  (.A(g22228), .Z(g25480) ) ;
INV     gate9051  (.A(g22228), .Z(g25481) ) ;
INV     gate9052  (.A(g22228), .Z(g25505) ) ;
INV     gate9053  (.A(g22228), .Z(g25506) ) ;
INV     gate9054  (.A(g23870), .Z(g25513) ) ;
INV     gate9055  (.A(g22228), .Z(g25517) ) ;
INV     gate9056  (.A(g22550), .Z(g25523) ) ;
INV     gate9057  (.A(g22228), .Z(g25524) ) ;
INV     gate9058  (.A(g22550), .Z(g25525) ) ;
INV     gate9059  (.A(g22594), .Z(g25528) ) ;
INV     gate9060  (.A(g22763), .Z(g25529) ) ;
INV     gate9061  (.A(g22550), .Z(g25533) ) ;
INV     gate9062  (.A(g22763), .Z(g25534) ) ;
INV     gate9063  (.A(g22763), .Z(g25535) ) ;
INV     gate9064  (.A(g22594), .Z(g25538) ) ;
INV     gate9065  (.A(g22763), .Z(g25541) ) ;
INV     gate9066  (.A(g22763), .Z(g25542) ) ;
INV     gate9067  (.A(g22594), .Z(g25544) ) ;
INV     gate9068  (.A(g22550), .Z(g25546) ) ;
INV     gate9069  (.A(g22550), .Z(g25547) ) ;
INV     gate9070  (.A(g22550), .Z(g25548) ) ;
INV     gate9071  (.A(g22763), .Z(g25549) ) ;
INV     gate9072  (.A(g22763), .Z(g25550) ) ;
INV     gate9073  (.A(g22594), .Z(g25552) ) ;
INV     gate9074  (.A(g22550), .Z(g25553) ) ;
INV     gate9075  (.A(g22550), .Z(g25554) ) ;
INV     gate9076  (.A(g22550), .Z(g25555) ) ;
INV     gate9077  (.A(g22763), .Z(g25556) ) ;
INV     gate9078  (.A(g22763), .Z(g25557) ) ;
INV     gate9079  (.A(g22594), .Z(g25558) ) ;
INV     gate9080  (.A(g22550), .Z(g25560) ) ;
INV     gate9081  (.A(g22550), .Z(g25561) ) ;
INV     gate9082  (.A(g22763), .Z(g25562) ) ;
INV     gate9083  (.A(g22594), .Z(g25563) ) ;
NAND2   gate9084  (.A(g907), .B(g19063), .Z(g22312) ) ;
INV     gate9085  (.A(g22312), .Z(g25564) ) ;
INV     gate9086  (.A(g22550), .Z(g25566) ) ;
AND2    gate9087  (.A(g896), .B(g22594), .Z(g24229) ) ;
INV     gate9088  (.A(g24229), .Z(II24759) ) ;
OR2     gate9089  (.A(g22310), .B(g18559), .Z(g24264) ) ;
INV     gate9090  (.A(g24264), .Z(II24781) ) ;
INV     gate9091  (.A(II24781), .Z(g25640) ) ;
OR2     gate9092  (.A(g22316), .B(g18560), .Z(g24265) ) ;
INV     gate9093  (.A(g24265), .Z(II24784) ) ;
INV     gate9094  (.A(II24784), .Z(g25641) ) ;
OR2     gate9095  (.A(g22329), .B(g18561), .Z(g24266) ) ;
INV     gate9096  (.A(g24266), .Z(II24787) ) ;
INV     gate9097  (.A(II24787), .Z(g25642) ) ;
AND2    gate9098  (.A(g4392), .B(g22550), .Z(g24298) ) ;
INV     gate9099  (.A(g24298), .Z(II24839) ) ;
NOR2    gate9100  (.A(g7400), .B(g22312), .Z(g24439) ) ;
INV     gate9101  (.A(g24439), .Z(g25766) ) ;
INV     gate9102  (.A(g25513), .Z(II24920) ) ;
INV     gate9103  (.A(II24920), .Z(g25771) ) ;
NOR2    gate9104  (.A(g7446), .B(g22325), .Z(g24453) ) ;
INV     gate9105  (.A(g24453), .Z(g25773) ) ;
OR2     gate9106  (.A(g22488), .B(g7567), .Z(g24510) ) ;
INV     gate9107  (.A(g24510), .Z(g25781) ) ;
INV     gate9108  (.A(g25250), .Z(g25783) ) ;
OR2     gate9109  (.A(g22517), .B(g7601), .Z(g24518) ) ;
INV     gate9110  (.A(g24518), .Z(g25786) ) ;
INV     gate9111  (.A(g25027), .Z(g25790) ) ;
INV     gate9112  (.A(g25051), .Z(g25820) ) ;
AND2    gate9113  (.A(g10710), .B(g22319), .Z(g24485) ) ;
INV     gate9114  (.A(g24485), .Z(g25830) ) ;
INV     gate9115  (.A(g25064), .Z(g25837) ) ;
INV     gate9116  (.A(g25250), .Z(g25838) ) ;
AND2    gate9117  (.A(g10727), .B(g22332), .Z(g24491) ) ;
INV     gate9118  (.A(g24491), .Z(g25849) ) ;
INV     gate9119  (.A(g25250), .Z(g25869) ) ;
AND2    gate9120  (.A(g22929), .B(g10503), .Z(g25026) ) ;
INV     gate9121  (.A(g25026), .Z(g25882) ) ;
AND2    gate9122  (.A(g22626), .B(g10851), .Z(g24537) ) ;
INV     gate9123  (.A(g24537), .Z(g25886) ) ;
NAND2   gate9124  (.A(g4098), .B(g22654), .Z(g24528) ) ;
INV     gate9125  (.A(g24528), .Z(g25892) ) ;
AND2    gate9126  (.A(g22626), .B(g10851), .Z(g24541) ) ;
INV     gate9127  (.A(g24541), .Z(g25893) ) ;
AND2    gate9128  (.A(g22929), .B(g10419), .Z(g24997) ) ;
INV     gate9129  (.A(g24997), .Z(g25899) ) ;
INV     gate9130  (.A(g24417), .Z(II25005) ) ;
INV     gate9131  (.A(II25005), .Z(g25903) ) ;
AND2    gate9132  (.A(g16288), .B(g23208), .Z(g24484) ) ;
INV     gate9133  (.A(g24484), .Z(II25028) ) ;
INV     gate9134  (.A(II25028), .Z(g25930) ) ;
NOR2    gate9135  (.A(g23498), .B(g23514), .Z(g24575) ) ;
INV     gate9136  (.A(g24575), .Z(g25994) ) ;
INV     gate9137  (.A(g25265), .Z(II25095) ) ;
INV     gate9138  (.A(II25095), .Z(g25997) ) ;
INV     gate9139  (.A(g25284), .Z(II25105) ) ;
INV     gate9140  (.A(II25105), .Z(g26026) ) ;
NAND2   gate9141  (.A(g19916), .B(g23105), .Z(g24804) ) ;
INV     gate9142  (.A(g24804), .Z(g26054) ) ;
INV     gate9143  (.A(g25322), .Z(II25115) ) ;
INV     gate9144  (.A(II25115), .Z(g26055) ) ;
NOR2    gate9145  (.A(g23554), .B(g23581), .Z(g24619) ) ;
INV     gate9146  (.A(g24619), .Z(g26081) ) ;
NAND2   gate9147  (.A(g19965), .B(g23132), .Z(g24809) ) ;
INV     gate9148  (.A(g24809), .Z(g26083) ) ;
NAND2   gate9149  (.A(g20011), .B(g23167), .Z(g24814) ) ;
INV     gate9150  (.A(g24814), .Z(g26093) ) ;
INV     gate9151  (.A(g24911), .Z(II25146) ) ;
INV     gate9152  (.A(II25146), .Z(g26105) ) ;
INV     gate9153  (.A(g24920), .Z(II25161) ) ;
INV     gate9154  (.A(II25161), .Z(g26131) ) ;
INV     gate9155  (.A(g25423), .Z(II25190) ) ;
INV     gate9156  (.A(II25190), .Z(g26187) ) ;
INV     gate9157  (.A(g24759), .Z(g26260) ) ;
NOR3    gate9158  (.A(g8725), .B(g23850), .C(g11083), .Z(g24875) ) ;
INV     gate9159  (.A(g24875), .Z(g26284) ) ;
AND2    gate9160  (.A(g23088), .B(g9104), .Z(g24872) ) ;
INV     gate9161  (.A(g24872), .Z(g26326) ) ;
INV     gate9162  (.A(g24818), .Z(g26337) ) ;
NOR3    gate9163  (.A(g10262), .B(g23978), .C(g12259), .Z(g24953) ) ;
INV     gate9164  (.A(g24953), .Z(g26340) ) ;
OR2     gate9165  (.A(g22151), .B(g22159), .Z(g24641) ) ;
INV     gate9166  (.A(g24641), .Z(II25327) ) ;
INV     gate9167  (.A(II25327), .Z(g26364) ) ;
INV     gate9168  (.A(g24466), .Z(II25351) ) ;
INV     gate9169  (.A(II25351), .Z(g26400) ) ;
OR2     gate9170  (.A(g19345), .B(g24004), .Z(g24374) ) ;
INV     gate9171  (.A(g24374), .Z(II25356) ) ;
INV     gate9172  (.A(II25356), .Z(g26424) ) ;
OR2     gate9173  (.A(g22189), .B(g22207), .Z(g24715) ) ;
INV     gate9174  (.A(g24715), .Z(II25359) ) ;
INV     gate9175  (.A(II25359), .Z(g26483) ) ;
INV     gate9176  (.A(g24477), .Z(II25366) ) ;
INV     gate9177  (.A(II25366), .Z(g26488) ) ;
INV     gate9178  (.A(g24891), .Z(II25369) ) ;
INV     gate9179  (.A(II25369), .Z(g26510) ) ;
NAND2   gate9180  (.A(g20838), .B(g23623), .Z(g25233) ) ;
INV     gate9181  (.A(g25233), .Z(g26518) ) ;
INV     gate9182  (.A(g24481), .Z(II25380) ) ;
INV     gate9183  (.A(II25380), .Z(g26519) ) ;
NAND2   gate9184  (.A(g20979), .B(g23659), .Z(g25255) ) ;
INV     gate9185  (.A(g25255), .Z(g26548) ) ;
INV     gate9186  (.A(g24483), .Z(II25391) ) ;
INV     gate9187  (.A(II25391), .Z(g26549) ) ;
NAND2   gate9188  (.A(g21124), .B(g23692), .Z(g25268) ) ;
INV     gate9189  (.A(g25268), .Z(g26575) ) ;
INV     gate9190  (.A(g24489), .Z(II25399) ) ;
INV     gate9191  (.A(II25399), .Z(g26576) ) ;
NAND2   gate9192  (.A(g21190), .B(g23726), .Z(g25293) ) ;
INV     gate9193  (.A(g25293), .Z(g26605) ) ;
NAND2   gate9194  (.A(g12333), .B(g22342), .Z(g25382) ) ;
INV     gate9195  (.A(g25382), .Z(g26607) ) ;
NAND2   gate9196  (.A(g21253), .B(g23756), .Z(g25334) ) ;
INV     gate9197  (.A(g25334), .Z(g26608) ) ;
NAND2   gate9198  (.A(g12371), .B(g22369), .Z(g25426) ) ;
INV     gate9199  (.A(g25426), .Z(g26614) ) ;
NAND2   gate9200  (.A(g12374), .B(g22384), .Z(g25432) ) ;
INV     gate9201  (.A(g25432), .Z(g26615) ) ;
NAND2   gate9202  (.A(g12432), .B(g22417), .Z(g25467) ) ;
INV     gate9203  (.A(g25467), .Z(g26631) ) ;
NAND2   gate9204  (.A(g12437), .B(g22432), .Z(g25473) ) ;
INV     gate9205  (.A(g25473), .Z(g26632) ) ;
NOR2    gate9206  (.A(g9766), .B(g23782), .Z(g25317) ) ;
INV     gate9207  (.A(g25317), .Z(g26634) ) ;
INV     gate9208  (.A(g25115), .Z(g26648) ) ;
NAND3   gate9209  (.A(g22342), .B(g1648), .C(g8187), .Z(g25337) ) ;
INV     gate9210  (.A(g25337), .Z(g26653) ) ;
NAND2   gate9211  (.A(g22342), .B(g11991), .Z(g25275) ) ;
INV     gate9212  (.A(g25275), .Z(g26654) ) ;
NAND2   gate9213  (.A(g12479), .B(g22457), .Z(g25492) ) ;
INV     gate9214  (.A(g25492), .Z(g26655) ) ;
NAND2   gate9215  (.A(g12483), .B(g22472), .Z(g25495) ) ;
INV     gate9216  (.A(g25495), .Z(g26656) ) ;
INV     gate9217  (.A(g25275), .Z(g26672) ) ;
NAND3   gate9218  (.A(g22369), .B(g1783), .C(g8241), .Z(g25385) ) ;
INV     gate9219  (.A(g25385), .Z(g26679) ) ;
NAND2   gate9220  (.A(g22369), .B(g12018), .Z(g25300) ) ;
INV     gate9221  (.A(g25300), .Z(g26680) ) ;
NAND3   gate9222  (.A(g22384), .B(g2208), .C(g8259), .Z(g25396) ) ;
INV     gate9223  (.A(g25396), .Z(g26681) ) ;
NAND2   gate9224  (.A(g22384), .B(g12021), .Z(g25309) ) ;
INV     gate9225  (.A(g25309), .Z(g26682) ) ;
NAND2   gate9226  (.A(g12540), .B(g22498), .Z(g25514) ) ;
INV     gate9227  (.A(g25514), .Z(g26683) ) ;
INV     gate9228  (.A(g25300), .Z(g26693) ) ;
NAND3   gate9229  (.A(g22417), .B(g1917), .C(g8302), .Z(g25429) ) ;
INV     gate9230  (.A(g25429), .Z(g26700) ) ;
NAND2   gate9231  (.A(g22417), .B(g12047), .Z(g25341) ) ;
INV     gate9232  (.A(g25341), .Z(g26701) ) ;
INV     gate9233  (.A(g25309), .Z(g26702) ) ;
NAND3   gate9234  (.A(g22432), .B(g2342), .C(g8316), .Z(g25435) ) ;
INV     gate9235  (.A(g25435), .Z(g26709) ) ;
NAND2   gate9236  (.A(g22432), .B(g12051), .Z(g25349) ) ;
INV     gate9237  (.A(g25349), .Z(g26710) ) ;
INV     gate9238  (.A(g25168), .Z(g26718) ) ;
INV     gate9239  (.A(g25275), .Z(g26720) ) ;
INV     gate9240  (.A(g25341), .Z(g26724) ) ;
NAND3   gate9241  (.A(g22457), .B(g2051), .C(g8365), .Z(g25470) ) ;
INV     gate9242  (.A(g25470), .Z(g26731) ) ;
NAND2   gate9243  (.A(g22457), .B(g12082), .Z(g25389) ) ;
INV     gate9244  (.A(g25389), .Z(g26732) ) ;
INV     gate9245  (.A(g25349), .Z(g26736) ) ;
NAND3   gate9246  (.A(g22472), .B(g2476), .C(g8373), .Z(g25476) ) ;
INV     gate9247  (.A(g25476), .Z(g26743) ) ;
NAND2   gate9248  (.A(g22472), .B(g12086), .Z(g25400) ) ;
INV     gate9249  (.A(g25400), .Z(g26744) ) ;
INV     gate9250  (.A(g25300), .Z(g26754) ) ;
INV     gate9251  (.A(g25389), .Z(g26758) ) ;
INV     gate9252  (.A(g25309), .Z(g26765) ) ;
INV     gate9253  (.A(g25400), .Z(g26769) ) ;
NAND3   gate9254  (.A(g22498), .B(g2610), .C(g8418), .Z(g25498) ) ;
INV     gate9255  (.A(g25498), .Z(g26776) ) ;
NAND2   gate9256  (.A(g22498), .B(g12122), .Z(g25439) ) ;
INV     gate9257  (.A(g25439), .Z(g26777) ) ;
INV     gate9258  (.A(g25341), .Z(g26784) ) ;
INV     gate9259  (.A(g25349), .Z(g26788) ) ;
INV     gate9260  (.A(g25439), .Z(g26792) ) ;
INV     gate9261  (.A(g25073), .Z(II25511) ) ;
INV     gate9262  (.A(g25073), .Z(II25514) ) ;
INV     gate9263  (.A(II25514), .Z(g26802) ) ;
INV     gate9264  (.A(g25389), .Z(g26803) ) ;
INV     gate9265  (.A(g25400), .Z(g26804) ) ;
INV     gate9266  (.A(g25220), .Z(g26810) ) ;
INV     gate9267  (.A(g25206), .Z(g26811) ) ;
INV     gate9268  (.A(g25439), .Z(g26812) ) ;
INV     gate9269  (.A(g25221), .Z(g26814) ) ;
INV     gate9270  (.A(g25260), .Z(g26816) ) ;
INV     gate9271  (.A(g25242), .Z(g26817) ) ;
INV     gate9272  (.A(g25222), .Z(II25530) ) ;
INV     gate9273  (.A(II25530), .Z(g26818) ) ;
AND2    gate9274  (.A(g11202), .B(g22680), .Z(g25448) ) ;
INV     gate9275  (.A(g25448), .Z(II25534) ) ;
INV     gate9276  (.A(II25534), .Z(g26820) ) ;
INV     gate9277  (.A(g25298), .Z(g26824) ) ;
INV     gate9278  (.A(g25180), .Z(II25541) ) ;
INV     gate9279  (.A(II25541), .Z(g26825) ) ;
INV     gate9280  (.A(g24819), .Z(g26827) ) ;
AND2    gate9281  (.A(g4584), .B(g22161), .Z(g24411) ) ;
INV     gate9282  (.A(g24411), .Z(g26830) ) ;
INV     gate9283  (.A(g24836), .Z(g26831) ) ;
INV     gate9284  (.A(g24850), .Z(g26832) ) ;
INV     gate9285  (.A(g25240), .Z(II25552) ) ;
INV     gate9286  (.A(II25552), .Z(g26834) ) ;
INV     gate9287  (.A(g25241), .Z(II25555) ) ;
INV     gate9288  (.A(II25555), .Z(g26835) ) ;
INV     gate9289  (.A(g24866), .Z(g26836) ) ;
INV     gate9290  (.A(g24869), .Z(g26837) ) ;
INV     gate9291  (.A(g25250), .Z(II25562) ) ;
INV     gate9292  (.A(II25562), .Z(g26840) ) ;
INV     gate9293  (.A(g24893), .Z(g26841) ) ;
INV     gate9294  (.A(g25272), .Z(II25567) ) ;
INV     gate9295  (.A(II25567), .Z(g26843) ) ;
INV     gate9296  (.A(g25296), .Z(II25576) ) ;
INV     gate9297  (.A(II25576), .Z(g26850) ) ;
INV     gate9298  (.A(g25297), .Z(II25579) ) ;
INV     gate9299  (.A(II25579), .Z(g26851) ) ;
NAND2   gate9300  (.A(g22763), .B(g2873), .Z(g25537) ) ;
INV     gate9301  (.A(g25537), .Z(II25586) ) ;
INV     gate9302  (.A(II25586), .Z(g26856) ) ;
INV     gate9303  (.A(g25380), .Z(II25591) ) ;
INV     gate9304  (.A(II25591), .Z(g26859) ) ;
NAND2   gate9305  (.A(g22763), .B(g2868), .Z(g25531) ) ;
INV     gate9306  (.A(g25531), .Z(II25594) ) ;
INV     gate9307  (.A(II25594), .Z(g26860) ) ;
INV     gate9308  (.A(g25424), .Z(II25598) ) ;
INV     gate9309  (.A(II25598), .Z(g26862) ) ;
OR2     gate9310  (.A(g7804), .B(g22669), .Z(g24842) ) ;
INV     gate9311  (.A(g24842), .Z(g26869) ) ;
INV     gate9312  (.A(g25465), .Z(II25606) ) ;
INV     gate9313  (.A(II25606), .Z(g26870) ) ;
INV     gate9314  (.A(g25640), .Z(II25677) ) ;
INV     gate9315  (.A(g25641), .Z(II25680) ) ;
INV     gate9316  (.A(g25642), .Z(II25683) ) ;
OR2     gate9317  (.A(g24812), .B(g21887), .Z(g25688) ) ;
INV     gate9318  (.A(g25688), .Z(II25689) ) ;
INV     gate9319  (.A(II25689), .Z(g26941) ) ;
OR2     gate9320  (.A(g24849), .B(g21888), .Z(g25689) ) ;
INV     gate9321  (.A(g25689), .Z(II25692) ) ;
INV     gate9322  (.A(II25692), .Z(g26942) ) ;
OR2     gate9323  (.A(g24864), .B(g21889), .Z(g25690) ) ;
INV     gate9324  (.A(g25690), .Z(II25695) ) ;
INV     gate9325  (.A(II25695), .Z(g26943) ) ;
INV     gate9326  (.A(g26105), .Z(g26973) ) ;
INV     gate9327  (.A(g26131), .Z(g26987) ) ;
INV     gate9328  (.A(g26105), .Z(g26990) ) ;
INV     gate9329  (.A(g26131), .Z(g27004) ) ;
OR2     gate9330  (.A(g22514), .B(g24510), .Z(g25911) ) ;
INV     gate9331  (.A(g25911), .Z(g27009) ) ;
OR2     gate9332  (.A(g22524), .B(g24518), .Z(g25917) ) ;
INV     gate9333  (.A(g25917), .Z(g27011) ) ;
INV     gate9334  (.A(g25903), .Z(II25743) ) ;
INV     gate9335  (.A(II25743), .Z(g27013) ) ;
NAND2   gate9336  (.A(g914), .B(g24439), .Z(g25888) ) ;
INV     gate9337  (.A(g25888), .Z(g27014) ) ;
INV     gate9338  (.A(g26869), .Z(g27015) ) ;
NAND2   gate9339  (.A(g1259), .B(g24453), .Z(g25895) ) ;
INV     gate9340  (.A(g25895), .Z(g27017) ) ;
AND2    gate9341  (.A(g24401), .B(g13106), .Z(g26823) ) ;
INV     gate9342  (.A(g26823), .Z(II25750) ) ;
INV     gate9343  (.A(II25750), .Z(g27018) ) ;
NOR2    gate9344  (.A(g7680), .B(g24528), .Z(g25932) ) ;
INV     gate9345  (.A(g25932), .Z(g27038) ) ;
INV     gate9346  (.A(g26424), .Z(II25779) ) ;
INV     gate9347  (.A(II25779), .Z(g27051) ) ;
INV     gate9348  (.A(g26424), .Z(II25786) ) ;
INV     gate9349  (.A(II25786), .Z(g27064) ) ;
INV     gate9350  (.A(g26424), .Z(II25790) ) ;
INV     gate9351  (.A(II25790), .Z(g27074) ) ;
OR2     gate9352  (.A(g24433), .B(g10674), .Z(g26673) ) ;
INV     gate9353  (.A(g26673), .Z(g27084) ) ;
OR2     gate9354  (.A(g24444), .B(g10704), .Z(g26694) ) ;
INV     gate9355  (.A(g26694), .Z(g27088) ) ;
OR2     gate9356  (.A(g24447), .B(g10705), .Z(g26703) ) ;
INV     gate9357  (.A(g26703), .Z(g27089) ) ;
OR2     gate9358  (.A(g24457), .B(g10719), .Z(g26725) ) ;
INV     gate9359  (.A(g26725), .Z(g27091) ) ;
OR2     gate9360  (.A(g24460), .B(g10720), .Z(g26737) ) ;
INV     gate9361  (.A(g26737), .Z(g27092) ) ;
OR2     gate9362  (.A(g24468), .B(g7511), .Z(g26759) ) ;
INV     gate9363  (.A(g26759), .Z(g27100) ) ;
OR2     gate9364  (.A(g24471), .B(g10732), .Z(g26770) ) ;
INV     gate9365  (.A(g26770), .Z(g27101) ) ;
OR2     gate9366  (.A(g24478), .B(g7520), .Z(g26793) ) ;
INV     gate9367  (.A(g26793), .Z(g27112) ) ;
INV     gate9368  (.A(g26105), .Z(g27142) ) ;
INV     gate9369  (.A(g26131), .Z(g27155) ) ;
NOR3    gate9370  (.A(g4311), .B(g24380), .C(g24369), .Z(g25851) ) ;
INV     gate9371  (.A(g25851), .Z(II25869) ) ;
INV     gate9372  (.A(II25869), .Z(g27163) ) ;
NOR3    gate9373  (.A(g7166), .B(g24380), .C(g24369), .Z(g25776) ) ;
INV     gate9374  (.A(g25776), .Z(II25882) ) ;
INV     gate9375  (.A(II25882), .Z(g27187) ) ;
NOR2    gate9376  (.A(g23052), .B(g24751), .Z(g26162) ) ;
INV     gate9377  (.A(g26162), .Z(g27237) ) ;
NOR2    gate9378  (.A(g23079), .B(g24766), .Z(g26183) ) ;
INV     gate9379  (.A(g26183), .Z(g27242) ) ;
NOR2    gate9380  (.A(g23124), .B(g24779), .Z(g26209) ) ;
INV     gate9381  (.A(g26209), .Z(g27245) ) ;
NOR2    gate9382  (.A(g8631), .B(g24825), .Z(g26330) ) ;
INV     gate9383  (.A(g26330), .Z(g27279) ) ;
INV     gate9384  (.A(g26818), .Z(II26004) ) ;
INV     gate9385  (.A(II26004), .Z(g27320) ) ;
NAND3   gate9386  (.A(g744), .B(g24875), .C(g11679), .Z(g26352) ) ;
INV     gate9387  (.A(g26352), .Z(g27349) ) ;
OR2     gate9388  (.A(g25504), .B(g25141), .Z(g26365) ) ;
INV     gate9389  (.A(g26365), .Z(II26100) ) ;
INV     gate9390  (.A(II26100), .Z(g27402) ) ;
NAND3   gate9391  (.A(g577), .B(g24953), .C(g12323), .Z(g26382) ) ;
INV     gate9392  (.A(g26382), .Z(g27415) ) ;
INV     gate9393  (.A(g26510), .Z(II26130) ) ;
INV     gate9394  (.A(II26130), .Z(g27438) ) ;
NOR3    gate9395  (.A(g8990), .B(g13756), .C(g24732), .Z(g26598) ) ;
INV     gate9396  (.A(g26598), .Z(g27492) ) ;
INV     gate9397  (.A(g26260), .Z(II26195) ) ;
INV     gate9398  (.A(II26195), .Z(g27527) ) ;
NOR2    gate9399  (.A(g23560), .B(g25144), .Z(g26625) ) ;
INV     gate9400  (.A(g26625), .Z(g27554) ) ;
NOR2    gate9401  (.A(g23602), .B(g25160), .Z(g26645) ) ;
INV     gate9402  (.A(g26645), .Z(g27565) ) ;
NOR2    gate9403  (.A(g23642), .B(g25175), .Z(g26667) ) ;
INV     gate9404  (.A(g26667), .Z(g27573) ) ;
INV     gate9405  (.A(g26081), .Z(g27576) ) ;
NOR2    gate9406  (.A(g23678), .B(g25189), .Z(g26686) ) ;
INV     gate9407  (.A(g26686), .Z(g27583) ) ;
INV     gate9408  (.A(g25994), .Z(g27585) ) ;
NOR2    gate9409  (.A(g23711), .B(g25203), .Z(g26715) ) ;
INV     gate9410  (.A(g26715), .Z(g27592) ) ;
NAND2   gate9411  (.A(g6856), .B(g25317), .Z(g26745) ) ;
INV     gate9412  (.A(g26745), .Z(g27597) ) ;
INV     gate9413  (.A(g26820), .Z(II26296) ) ;
INV     gate9414  (.A(II26296), .Z(g27662) ) ;
INV     gate9415  (.A(g26825), .Z(II26309) ) ;
INV     gate9416  (.A(II26309), .Z(g27675) ) ;
INV     gate9417  (.A(g26648), .Z(g27698) ) ;
INV     gate9418  (.A(g26834), .Z(II26334) ) ;
INV     gate9419  (.A(II26334), .Z(g27708) ) ;
INV     gate9420  (.A(g26835), .Z(II26337) ) ;
INV     gate9421  (.A(II26337), .Z(g27709) ) ;
INV     gate9422  (.A(g26424), .Z(g27730) ) ;
INV     gate9423  (.A(g26843), .Z(II26356) ) ;
INV     gate9424  (.A(II26356), .Z(g27736) ) ;
INV     gate9425  (.A(g26718), .Z(g27737) ) ;
INV     gate9426  (.A(g26850), .Z(II26378) ) ;
INV     gate9427  (.A(II26378), .Z(g27773) ) ;
INV     gate9428  (.A(g26851), .Z(II26381) ) ;
INV     gate9429  (.A(II26381), .Z(g27774) ) ;
INV     gate9430  (.A(g26802), .Z(g27830) ) ;
INV     gate9431  (.A(g26187), .Z(II26406) ) ;
INV     gate9432  (.A(g26187), .Z(II26409) ) ;
INV     gate9433  (.A(II26409), .Z(g27832) ) ;
INV     gate9434  (.A(g26859), .Z(II26427) ) ;
INV     gate9435  (.A(II26427), .Z(g27880) ) ;
INV     gate9436  (.A(g26856), .Z(II26430) ) ;
INV     gate9437  (.A(II26430), .Z(g27881) ) ;
INV     gate9438  (.A(g26810), .Z(g27928) ) ;
INV     gate9439  (.A(g26860), .Z(II26448) ) ;
INV     gate9440  (.A(II26448), .Z(g27929) ) ;
INV     gate9441  (.A(g26862), .Z(II26451) ) ;
INV     gate9442  (.A(II26451), .Z(g27930) ) ;
INV     gate9443  (.A(g26870), .Z(II26466) ) ;
INV     gate9444  (.A(II26466), .Z(g27956) ) ;
INV     gate9445  (.A(g26816), .Z(g27961) ) ;
INV     gate9446  (.A(g25771), .Z(II26479) ) ;
INV     gate9447  (.A(II26479), .Z(g27967) ) ;
INV     gate9448  (.A(g26673), .Z(g27971) ) ;
INV     gate9449  (.A(g26694), .Z(g27975) ) ;
INV     gate9450  (.A(g26703), .Z(g27976) ) ;
INV     gate9451  (.A(g26105), .Z(g27977) ) ;
INV     gate9452  (.A(g26725), .Z(g27983) ) ;
INV     gate9453  (.A(g26737), .Z(g27984) ) ;
INV     gate9454  (.A(g26131), .Z(g27985) ) ;
INV     gate9455  (.A(g26759), .Z(g27989) ) ;
INV     gate9456  (.A(g26770), .Z(g27990) ) ;
AND2    gate9457  (.A(g4593), .B(g24411), .Z(g25852) ) ;
INV     gate9458  (.A(g25852), .Z(g27991) ) ;
INV     gate9459  (.A(g26811), .Z(II26503) ) ;
INV     gate9460  (.A(II26503), .Z(g27993) ) ;
INV     gate9461  (.A(g26793), .Z(g27994) ) ;
INV     gate9462  (.A(g26814), .Z(II26508) ) ;
INV     gate9463  (.A(II26508), .Z(g27996) ) ;
INV     gate9464  (.A(g26817), .Z(II26512) ) ;
INV     gate9465  (.A(II26512), .Z(g27998) ) ;
INV     gate9466  (.A(g26824), .Z(II26516) ) ;
INV     gate9467  (.A(II26516), .Z(g28009) ) ;
INV     gate9468  (.A(g26365), .Z(g28032) ) ;
INV     gate9469  (.A(g26365), .Z(g28033) ) ;
INV     gate9470  (.A(g26365), .Z(g28034) ) ;
INV     gate9471  (.A(g26365), .Z(g28036) ) ;
INV     gate9472  (.A(g26365), .Z(g28037) ) ;
INV     gate9473  (.A(g26365), .Z(g28038) ) ;
INV     gate9474  (.A(g26365), .Z(g28039) ) ;
INV     gate9475  (.A(g26365), .Z(g28040) ) ;
INV     gate9476  (.A(g26941), .Z(II26578) ) ;
INV     gate9477  (.A(g26942), .Z(II26581) ) ;
INV     gate9478  (.A(g26943), .Z(II26584) ) ;
OR3     gate9479  (.A(g26866), .B(g21370), .C(II25736), .Z(g27008) ) ;
INV     gate9480  (.A(g27008), .Z(g28119) ) ;
OR2     gate9481  (.A(g22522), .B(g25911), .Z(g27108) ) ;
INV     gate9482  (.A(g27108), .Z(g28120) ) ;
NOR2    gate9483  (.A(g26712), .B(g26749), .Z(g27093) ) ;
INV     gate9484  (.A(g27093), .Z(g28121) ) ;
OR2     gate9485  (.A(g22537), .B(g25917), .Z(g27122) ) ;
INV     gate9486  (.A(g27122), .Z(g28126) ) ;
NOR2    gate9487  (.A(g26750), .B(g26779), .Z(g27102) ) ;
INV     gate9488  (.A(g27102), .Z(g28127) ) ;
AND2    gate9489  (.A(g25834), .B(g13117), .Z(g27965) ) ;
INV     gate9490  (.A(g27965), .Z(II26638) ) ;
INV     gate9491  (.A(II26638), .Z(g28137) ) ;
INV     gate9492  (.A(g27675), .Z(II26649) ) ;
INV     gate9493  (.A(II26649), .Z(g28142) ) ;
INV     gate9494  (.A(g27576), .Z(II26654) ) ;
INV     gate9495  (.A(II26654), .Z(g28147) ) ;
INV     gate9496  (.A(g27708), .Z(II26664) ) ;
INV     gate9497  (.A(II26664), .Z(g28155) ) ;
INV     gate9498  (.A(g27585), .Z(II26667) ) ;
INV     gate9499  (.A(II26667), .Z(g28156) ) ;
INV     gate9500  (.A(g27709), .Z(II26670) ) ;
INV     gate9501  (.A(II26670), .Z(g28157) ) ;
INV     gate9502  (.A(g27736), .Z(II26676) ) ;
INV     gate9503  (.A(II26676), .Z(g28161) ) ;
INV     gate9504  (.A(g27773), .Z(II26679) ) ;
INV     gate9505  (.A(II26679), .Z(g28162) ) ;
INV     gate9506  (.A(g27774), .Z(II26682) ) ;
INV     gate9507  (.A(II26682), .Z(g28163) ) ;
INV     gate9508  (.A(g27880), .Z(II26687) ) ;
INV     gate9509  (.A(II26687), .Z(g28166) ) ;
INV     gate9510  (.A(g27930), .Z(II26693) ) ;
INV     gate9511  (.A(II26693), .Z(g28173) ) ;
INV     gate9512  (.A(g27956), .Z(II26700) ) ;
INV     gate9513  (.A(II26700), .Z(g28181) ) ;
INV     gate9514  (.A(g27967), .Z(II26705) ) ;
INV     gate9515  (.A(II26705), .Z(g28184) ) ;
NOR3    gate9516  (.A(g22137), .B(g26866), .C(g20277), .Z(g27511) ) ;
INV     gate9517  (.A(g27511), .Z(II26710) ) ;
INV     gate9518  (.A(II26710), .Z(g28187) ) ;
INV     gate9519  (.A(g27064), .Z(g28241) ) ;
INV     gate9520  (.A(g27074), .Z(g28250) ) ;
INV     gate9521  (.A(g27013), .Z(II26785) ) ;
INV     gate9522  (.A(II26785), .Z(g28262) ) ;
AND3    gate9523  (.A(g24688), .B(g26424), .C(g22763), .Z(g27660) ) ;
INV     gate9524  (.A(g27660), .Z(II26799) ) ;
INV     gate9525  (.A(II26799), .Z(g28274) ) ;
NAND2   gate9526  (.A(g24776), .B(g26208), .Z(g27295) ) ;
INV     gate9527  (.A(g27295), .Z(g28294) ) ;
NAND2   gate9528  (.A(g24787), .B(g26235), .Z(g27306) ) ;
INV     gate9529  (.A(g27306), .Z(g28307) ) ;
NAND2   gate9530  (.A(g24793), .B(g26255), .Z(g27317) ) ;
INV     gate9531  (.A(g27317), .Z(g28321) ) ;
NAND3   gate9532  (.A(g287), .B(g26330), .C(g23204), .Z(g27463) ) ;
INV     gate9533  (.A(g27463), .Z(g28325) ) ;
AND2    gate9534  (.A(g255), .B(g26827), .Z(g27414) ) ;
INV     gate9535  (.A(g27414), .Z(g28326) ) ;
INV     gate9536  (.A(g27527), .Z(II26880) ) ;
INV     gate9537  (.A(II26880), .Z(g28367) ) ;
NOR3    gate9538  (.A(g8770), .B(g26352), .C(g11083), .Z(g27528) ) ;
INV     gate9539  (.A(g27528), .Z(g28370) ) ;
INV     gate9540  (.A(g27064), .Z(g28380) ) ;
INV     gate9541  (.A(g27074), .Z(g28399) ) ;
INV     gate9542  (.A(g27015), .Z(II26925) ) ;
INV     gate9543  (.A(II26925), .Z(g28431) ) ;
OR2     gate9544  (.A(g26105), .B(g26131), .Z(g27980) ) ;
INV     gate9545  (.A(g27980), .Z(II26929) ) ;
INV     gate9546  (.A(II26929), .Z(g28436) ) ;
NOR3    gate9547  (.A(g8891), .B(g26382), .C(g12259), .Z(g27629) ) ;
INV     gate9548  (.A(g27629), .Z(g28441) ) ;
AND2    gate9549  (.A(g26337), .B(g20033), .Z(g27599) ) ;
INV     gate9550  (.A(g27599), .Z(II26936) ) ;
INV     gate9551  (.A(II26936), .Z(g28443) ) ;
OR2     gate9552  (.A(g26131), .B(g26105), .Z(g27972) ) ;
INV     gate9553  (.A(g27972), .Z(II26952) ) ;
INV     gate9554  (.A(II26952), .Z(g28463) ) ;
NAND3   gate9555  (.A(g164), .B(g26598), .C(g23042), .Z(g27654) ) ;
INV     gate9556  (.A(g27654), .Z(g28479) ) ;
AND2    gate9557  (.A(g26359), .B(g14191), .Z(g27277) ) ;
INV     gate9558  (.A(g27277), .Z(II26989) ) ;
INV     gate9559  (.A(II26989), .Z(g28508) ) ;
AND4    gate9560  (.A(g22342), .B(g25182), .C(g26424), .D(g26148), .Z(g27700) ) ;
INV     gate9561  (.A(g27700), .Z(g28559) ) ;
AND4    gate9562  (.A(g22369), .B(g25193), .C(g26424), .D(g26166), .Z(g27711) ) ;
INV     gate9563  (.A(g27711), .Z(g28575) ) ;
AND4    gate9564  (.A(g22384), .B(g25195), .C(g26424), .D(g26171), .Z(g27714) ) ;
INV     gate9565  (.A(g27714), .Z(g28579) ) ;
AND4    gate9566  (.A(g22417), .B(g25208), .C(g26424), .D(g26190), .Z(g27724) ) ;
INV     gate9567  (.A(g27724), .Z(g28590) ) ;
AND4    gate9568  (.A(g22432), .B(g25211), .C(g26424), .D(g26195), .Z(g27727) ) ;
INV     gate9569  (.A(g27727), .Z(g28593) ) ;
NOR2    gate9570  (.A(g9492), .B(g26745), .Z(g27717) ) ;
INV     gate9571  (.A(g27717), .Z(g28598) ) ;
AND4    gate9572  (.A(g22457), .B(g25224), .C(g26424), .D(g26213), .Z(g27759) ) ;
INV     gate9573  (.A(g27759), .Z(g28604) ) ;
AND4    gate9574  (.A(g22472), .B(g25226), .C(g26424), .D(g26218), .Z(g27762) ) ;
INV     gate9575  (.A(g27762), .Z(g28606) ) ;
NAND2   gate9576  (.A(g25172), .B(g26666), .Z(g27670) ) ;
INV     gate9577  (.A(g27670), .Z(g28608) ) ;
AND4    gate9578  (.A(g22498), .B(g25245), .C(g26424), .D(g26236), .Z(g27817) ) ;
INV     gate9579  (.A(g27817), .Z(g28615) ) ;
NAND2   gate9580  (.A(g25186), .B(g26685), .Z(g27679) ) ;
INV     gate9581  (.A(g27679), .Z(g28620) ) ;
NAND2   gate9582  (.A(g25200), .B(g26714), .Z(g27687) ) ;
INV     gate9583  (.A(g27687), .Z(g28633) ) ;
NAND2   gate9584  (.A(g25216), .B(g26752), .Z(g27693) ) ;
INV     gate9585  (.A(g27693), .Z(g28648) ) ;
OR2     gate9586  (.A(g17292), .B(g26673), .Z(g27742) ) ;
INV     gate9587  (.A(g27742), .Z(g28656) ) ;
NAND2   gate9588  (.A(g25237), .B(g26782), .Z(g27705) ) ;
INV     gate9589  (.A(g27705), .Z(g28669) ) ;
OR2     gate9590  (.A(g17317), .B(g26694), .Z(g27779) ) ;
INV     gate9591  (.A(g27779), .Z(g28675) ) ;
OR2     gate9592  (.A(g17321), .B(g26703), .Z(g27800) ) ;
INV     gate9593  (.A(g27800), .Z(g28678) ) ;
OR2     gate9594  (.A(g17401), .B(g26725), .Z(g27837) ) ;
INV     gate9595  (.A(g27837), .Z(g28693) ) ;
OR2     gate9596  (.A(g17405), .B(g26737), .Z(g27858) ) ;
INV     gate9597  (.A(g27858), .Z(g28696) ) ;
INV     gate9598  (.A(g27662), .Z(II27192) ) ;
INV     gate9599  (.A(II27192), .Z(g28709) ) ;
OR2     gate9600  (.A(g14438), .B(g26759), .Z(g27886) ) ;
INV     gate9601  (.A(g27886), .Z(g28711) ) ;
OR2     gate9602  (.A(g17424), .B(g26770), .Z(g27907) ) ;
INV     gate9603  (.A(g27907), .Z(g28713) ) ;
OR2     gate9604  (.A(g14506), .B(g26793), .Z(g27937) ) ;
INV     gate9605  (.A(g27937), .Z(g28726) ) ;
INV     gate9606  (.A(g27993), .Z(II27232) ) ;
INV     gate9607  (.A(II27232), .Z(g28752) ) ;
INV     gate9608  (.A(g27320), .Z(II27235) ) ;
INV     gate9609  (.A(g27320), .Z(II27238) ) ;
INV     gate9610  (.A(II27238), .Z(g28754) ) ;
INV     gate9611  (.A(g27996), .Z(II27253) ) ;
INV     gate9612  (.A(II27253), .Z(g28779) ) ;
INV     gate9613  (.A(g27998), .Z(II27271) ) ;
INV     gate9614  (.A(II27271), .Z(g28819) ) ;
INV     gate9615  (.A(g28009), .Z(II27314) ) ;
INV     gate9616  (.A(II27314), .Z(g28917) ) ;
INV     gate9617  (.A(g27832), .Z(g28918) ) ;
INV     gate9618  (.A(g27830), .Z(g28954) ) ;
INV     gate9619  (.A(g27881), .Z(II27368) ) ;
INV     gate9620  (.A(II27368), .Z(g29013) ) ;
INV     gate9621  (.A(g27742), .Z(g29014) ) ;
INV     gate9622  (.A(g27438), .Z(II27385) ) ;
INV     gate9623  (.A(II27385), .Z(g29041) ) ;
INV     gate9624  (.A(g27698), .Z(II27388) ) ;
INV     gate9625  (.A(II27388), .Z(g29042) ) ;
INV     gate9626  (.A(g27929), .Z(II27391) ) ;
INV     gate9627  (.A(II27391), .Z(g29043) ) ;
INV     gate9628  (.A(g27742), .Z(g29044) ) ;
INV     gate9629  (.A(g27779), .Z(g29045) ) ;
INV     gate9630  (.A(g27800), .Z(g29056) ) ;
INV     gate9631  (.A(g27051), .Z(II27401) ) ;
INV     gate9632  (.A(II27401), .Z(g29067) ) ;
INV     gate9633  (.A(g27742), .Z(g29079) ) ;
INV     gate9634  (.A(g27779), .Z(g29080) ) ;
INV     gate9635  (.A(g27837), .Z(g29081) ) ;
INV     gate9636  (.A(g27800), .Z(g29092) ) ;
INV     gate9637  (.A(g27858), .Z(g29093) ) ;
INV     gate9638  (.A(g27779), .Z(g29115) ) ;
INV     gate9639  (.A(g27837), .Z(g29116) ) ;
INV     gate9640  (.A(g27886), .Z(g29117) ) ;
INV     gate9641  (.A(g27800), .Z(g29128) ) ;
INV     gate9642  (.A(g27858), .Z(g29129) ) ;
INV     gate9643  (.A(g27907), .Z(g29130) ) ;
INV     gate9644  (.A(g27737), .Z(II27449) ) ;
INV     gate9645  (.A(II27449), .Z(g29147) ) ;
INV     gate9646  (.A(g27837), .Z(g29149) ) ;
INV     gate9647  (.A(g27886), .Z(g29150) ) ;
INV     gate9648  (.A(g27858), .Z(g29151) ) ;
INV     gate9649  (.A(g27907), .Z(g29152) ) ;
INV     gate9650  (.A(g27937), .Z(g29153) ) ;
INV     gate9651  (.A(g27886), .Z(g29169) ) ;
INV     gate9652  (.A(g27907), .Z(g29170) ) ;
INV     gate9653  (.A(g27937), .Z(g29171) ) ;
AND2    gate9654  (.A(g4601), .B(g25852), .Z(g27020) ) ;
INV     gate9655  (.A(g27020), .Z(g29172) ) ;
INV     gate9656  (.A(g27937), .Z(g29177) ) ;
INV     gate9657  (.A(g27928), .Z(II27481) ) ;
INV     gate9658  (.A(II27481), .Z(g29185) ) ;
NOR2    gate9659  (.A(g7544), .B(g25888), .Z(g27046) ) ;
INV     gate9660  (.A(g27046), .Z(g29190) ) ;
INV     gate9661  (.A(g27511), .Z(II27492) ) ;
INV     gate9662  (.A(II27492), .Z(g29194) ) ;
INV     gate9663  (.A(g27961), .Z(II27495) ) ;
INV     gate9664  (.A(II27495), .Z(g29195) ) ;
NOR2    gate9665  (.A(g7577), .B(g25895), .Z(g27059) ) ;
INV     gate9666  (.A(g27059), .Z(g29196) ) ;
INV     gate9667  (.A(g28187), .Z(II27543) ) ;
INV     gate9668  (.A(g29041), .Z(II27546) ) ;
INV     gate9669  (.A(g28161), .Z(II27549) ) ;
INV     gate9670  (.A(g28162), .Z(II27552) ) ;
INV     gate9671  (.A(g28142), .Z(II27555) ) ;
INV     gate9672  (.A(g28155), .Z(II27558) ) ;
INV     gate9673  (.A(g28163), .Z(II27561) ) ;
INV     gate9674  (.A(g28166), .Z(II27564) ) ;
INV     gate9675  (.A(g28181), .Z(II27567) ) ;
INV     gate9676  (.A(g28262), .Z(II27570) ) ;
INV     gate9677  (.A(g28157), .Z(II27573) ) ;
INV     gate9678  (.A(g28173), .Z(II27576) ) ;
INV     gate9679  (.A(g28184), .Z(II27579) ) ;
AND4    gate9680  (.A(g14438), .B(g25209), .C(g26424), .D(g27469), .Z(g28991) ) ;
INV     gate9681  (.A(g28991), .Z(g29310) ) ;
AND4    gate9682  (.A(g17424), .B(g25212), .C(g26424), .D(g27474), .Z(g28998) ) ;
INV     gate9683  (.A(g28998), .Z(g29311) ) ;
NAND3   gate9684  (.A(g27937), .B(g7490), .C(g7431), .Z(g28877) ) ;
INV     gate9685  (.A(g28877), .Z(g29312) ) ;
INV     gate9686  (.A(g28156), .Z(II27677) ) ;
INV     gate9687  (.A(II27677), .Z(g29317) ) ;
AND4    gate9688  (.A(g14506), .B(g25227), .C(g26424), .D(g27494), .Z(g29029) ) ;
INV     gate9689  (.A(g29029), .Z(g29318) ) ;
NAND2   gate9690  (.A(g925), .B(g27046), .Z(g28167) ) ;
INV     gate9691  (.A(g28167), .Z(g29333) ) ;
INV     gate9692  (.A(g28274), .Z(g29339) ) ;
OR2     gate9693  (.A(g22535), .B(g27108), .Z(g28188) ) ;
INV     gate9694  (.A(g28188), .Z(g29342) ) ;
NAND2   gate9695  (.A(g1270), .B(g27059), .Z(g28174) ) ;
INV     gate9696  (.A(g28174), .Z(g29343) ) ;
OR2     gate9697  (.A(g22540), .B(g27122), .Z(g28194) ) ;
INV     gate9698  (.A(g28194), .Z(g29348) ) ;
AND3    gate9699  (.A(g27163), .B(g22763), .C(g27064), .Z(g28224) ) ;
INV     gate9700  (.A(g28224), .Z(II27713) ) ;
INV     gate9701  (.A(II27713), .Z(g29353) ) ;
AND3    gate9702  (.A(g27187), .B(g22763), .C(g27074), .Z(g28231) ) ;
INV     gate9703  (.A(g28231), .Z(II27718) ) ;
INV     gate9704  (.A(II27718), .Z(g29358) ) ;
INV     gate9705  (.A(g29067), .Z(g29365) ) ;
INV     gate9706  (.A(g28752), .Z(II27730) ) ;
INV     gate9707  (.A(II27730), .Z(g29368) ) ;
INV     gate9708  (.A(g28779), .Z(II27735) ) ;
INV     gate9709  (.A(II27735), .Z(g29371) ) ;
OR2     gate9710  (.A(II26643), .B(II26644), .Z(g28140) ) ;
INV     gate9711  (.A(g28140), .Z(II27738) ) ;
INV     gate9712  (.A(II27738), .Z(g29372) ) ;
INV     gate9713  (.A(g28819), .Z(II27742) ) ;
INV     gate9714  (.A(II27742), .Z(g29374) ) ;
INV     gate9715  (.A(g28917), .Z(II27749) ) ;
INV     gate9716  (.A(II27749), .Z(g29379) ) ;
OR2     gate9717  (.A(g20242), .B(g27511), .Z(g28180) ) ;
INV     gate9718  (.A(g28180), .Z(g29385) ) ;
INV     gate9719  (.A(g28119), .Z(II27758) ) ;
INV     gate9720  (.A(II27758), .Z(g29474) ) ;
INV     gate9721  (.A(g29043), .Z(II27777) ) ;
INV     gate9722  (.A(II27777), .Z(g29491) ) ;
INV     gate9723  (.A(g29013), .Z(II27784) ) ;
INV     gate9724  (.A(II27784), .Z(g29498) ) ;
NAND2   gate9725  (.A(g27051), .B(g4507), .Z(g29186) ) ;
INV     gate9726  (.A(g29186), .Z(g29505) ) ;
NOR3    gate9727  (.A(g9073), .B(g27654), .C(g24732), .Z(g28353) ) ;
INV     gate9728  (.A(g28353), .Z(g29507) ) ;
NOR3    gate9729  (.A(g8575), .B(g27463), .C(g24825), .Z(g28444) ) ;
INV     gate9730  (.A(g28444), .Z(g29597) ) ;
NOR2    gate9731  (.A(g27730), .B(g22763), .Z(g28803) ) ;
INV     gate9732  (.A(g28803), .Z(II27927) ) ;
INV     gate9733  (.A(II27927), .Z(g29653) ) ;
INV     gate9734  (.A(g28803), .Z(II27941) ) ;
INV     gate9735  (.A(II27941), .Z(g29669) ) ;
INV     gate9736  (.A(g28803), .Z(II27954) ) ;
INV     gate9737  (.A(II27954), .Z(g29689) ) ;
NAND4   gate9738  (.A(g27064), .B(g24756), .C(g27163), .D(g19644), .Z(g28336) ) ;
INV     gate9739  (.A(g28336), .Z(g29697) ) ;
NAND3   gate9740  (.A(g758), .B(g27528), .C(g11679), .Z(g28504) ) ;
INV     gate9741  (.A(g28504), .Z(g29707) ) ;
INV     gate9742  (.A(g28803), .Z(II27970) ) ;
INV     gate9743  (.A(II27970), .Z(g29713) ) ;
NAND4   gate9744  (.A(g27074), .B(g24770), .C(g27187), .D(g19644), .Z(g28349) ) ;
INV     gate9745  (.A(g28349), .Z(g29725) ) ;
INV     gate9746  (.A(g28431), .Z(g29744) ) ;
NAND3   gate9747  (.A(g590), .B(g27629), .C(g12323), .Z(g28500) ) ;
INV     gate9748  (.A(g28500), .Z(g29745) ) ;
AND3    gate9749  (.A(g26424), .B(g22763), .C(g27031), .Z(g28153) ) ;
INV     gate9750  (.A(g28153), .Z(II28002) ) ;
INV     gate9751  (.A(II28002), .Z(g29755) ) ;
AND3    gate9752  (.A(g26424), .B(g22763), .C(g27037), .Z(g28158) ) ;
INV     gate9753  (.A(g28158), .Z(II28014) ) ;
INV     gate9754  (.A(II28014), .Z(g29765) ) ;
NAND2   gate9755  (.A(g27064), .B(g13593), .Z(g28363) ) ;
INV     gate9756  (.A(g28363), .Z(g29800) ) ;
NAND2   gate9757  (.A(g27064), .B(g13620), .Z(g28376) ) ;
INV     gate9758  (.A(g28376), .Z(g29811) ) ;
NAND2   gate9759  (.A(g27074), .B(g13621), .Z(g28381) ) ;
INV     gate9760  (.A(g28381), .Z(g29812) ) ;
INV     gate9761  (.A(g29194), .Z(II28062) ) ;
INV     gate9762  (.A(II28062), .Z(g29814) ) ;
NAND2   gate9763  (.A(g27064), .B(g13637), .Z(g28391) ) ;
INV     gate9764  (.A(g28391), .Z(g29846) ) ;
NAND2   gate9765  (.A(g27074), .B(g13655), .Z(g28395) ) ;
INV     gate9766  (.A(g28395), .Z(g29847) ) ;
NAND2   gate9767  (.A(g27064), .B(g13675), .Z(g28406) ) ;
INV     gate9768  (.A(g28406), .Z(g29862) ) ;
NAND2   gate9769  (.A(g27074), .B(g13679), .Z(g28410) ) ;
INV     gate9770  (.A(g28410), .Z(g29863) ) ;
NAND2   gate9771  (.A(g27074), .B(g13715), .Z(g28421) ) ;
INV     gate9772  (.A(g28421), .Z(g29878) ) ;
NAND3   gate9773  (.A(g27742), .B(g7268), .C(g1592), .Z(g28755) ) ;
INV     gate9774  (.A(g28755), .Z(g29893) ) ;
AND2    gate9775  (.A(g27552), .B(g14205), .Z(g28314) ) ;
INV     gate9776  (.A(g28314), .Z(II28128) ) ;
INV     gate9777  (.A(II28128), .Z(g29897) ) ;
NAND3   gate9778  (.A(g27779), .B(g7315), .C(g1728), .Z(g28783) ) ;
INV     gate9779  (.A(g28783), .Z(g29905) ) ;
NAND3   gate9780  (.A(g27800), .B(g7328), .C(g2153), .Z(g28793) ) ;
INV     gate9781  (.A(g28793), .Z(g29906) ) ;
NAND3   gate9782  (.A(g27742), .B(g7308), .C(g1636), .Z(g28780) ) ;
INV     gate9783  (.A(g28780), .Z(g29911) ) ;
NAND3   gate9784  (.A(g27837), .B(g7362), .C(g1862), .Z(g28827) ) ;
INV     gate9785  (.A(g28827), .Z(g29912) ) ;
NAND3   gate9786  (.A(g27858), .B(g7380), .C(g2287), .Z(g28840) ) ;
INV     gate9787  (.A(g28840), .Z(g29913) ) ;
NAND3   gate9788  (.A(g27779), .B(g7356), .C(g1772), .Z(g28824) ) ;
INV     gate9789  (.A(g28824), .Z(g29920) ) ;
NAND3   gate9790  (.A(g27886), .B(g7411), .C(g1996), .Z(g28864) ) ;
INV     gate9791  (.A(g28864), .Z(g29921) ) ;
NAND3   gate9792  (.A(g27800), .B(g7374), .C(g2197), .Z(g28837) ) ;
INV     gate9793  (.A(g28837), .Z(g29922) ) ;
NAND3   gate9794  (.A(g27907), .B(g7424), .C(g2421), .Z(g28874) ) ;
INV     gate9795  (.A(g28874), .Z(g29923) ) ;
NAND3   gate9796  (.A(g27742), .B(g1668), .C(g1592), .Z(g28820) ) ;
INV     gate9797  (.A(g28820), .Z(g29925) ) ;
NAND3   gate9798  (.A(g27837), .B(g7405), .C(g1906), .Z(g28861) ) ;
INV     gate9799  (.A(g28861), .Z(g29927) ) ;
NAND3   gate9800  (.A(g27858), .B(g7418), .C(g2331), .Z(g28871) ) ;
INV     gate9801  (.A(g28871), .Z(g29928) ) ;
NAND3   gate9802  (.A(g27937), .B(g7462), .C(g2555), .Z(g28914) ) ;
INV     gate9803  (.A(g28914), .Z(g29929) ) ;
INV     gate9804  (.A(g28803), .Z(II28162) ) ;
INV     gate9805  (.A(II28162), .Z(g29930) ) ;
NAND3   gate9806  (.A(g27779), .B(g1802), .C(g1728), .Z(g28857) ) ;
INV     gate9807  (.A(g28857), .Z(g29939) ) ;
NAND3   gate9808  (.A(g27886), .B(g7451), .C(g2040), .Z(g28900) ) ;
INV     gate9809  (.A(g28900), .Z(g29941) ) ;
NAND3   gate9810  (.A(g27800), .B(g2227), .C(g2153), .Z(g28867) ) ;
INV     gate9811  (.A(g28867), .Z(g29942) ) ;
NAND3   gate9812  (.A(g27907), .B(g7456), .C(g2465), .Z(g28911) ) ;
INV     gate9813  (.A(g28911), .Z(g29944) ) ;
INV     gate9814  (.A(g28803), .Z(II28174) ) ;
INV     gate9815  (.A(II28174), .Z(g29945) ) ;
NAND3   gate9816  (.A(g27742), .B(g1636), .C(g7252), .Z(g28853) ) ;
INV     gate9817  (.A(g28853), .Z(g29948) ) ;
NAND3   gate9818  (.A(g27837), .B(g1936), .C(g1862), .Z(g28896) ) ;
INV     gate9819  (.A(g28896), .Z(g29950) ) ;
NAND3   gate9820  (.A(g27858), .B(g2361), .C(g2287), .Z(g28907) ) ;
INV     gate9821  (.A(g28907), .Z(g29953) ) ;
NAND3   gate9822  (.A(g27937), .B(g7490), .C(g2599), .Z(g28950) ) ;
INV     gate9823  (.A(g28950), .Z(g29955) ) ;
INV     gate9824  (.A(g28803), .Z(II28185) ) ;
INV     gate9825  (.A(II28185), .Z(g29956) ) ;
NAND3   gate9826  (.A(g27742), .B(g1668), .C(g7268), .Z(g28885) ) ;
INV     gate9827  (.A(g28885), .Z(g29960) ) ;
NAND3   gate9828  (.A(g27779), .B(g1772), .C(g7275), .Z(g28892) ) ;
INV     gate9829  (.A(g28892), .Z(g29961) ) ;
NAND3   gate9830  (.A(g27886), .B(g2070), .C(g1996), .Z(g28931) ) ;
INV     gate9831  (.A(g28931), .Z(g29963) ) ;
NAND3   gate9832  (.A(g27800), .B(g2197), .C(g7280), .Z(g28903) ) ;
INV     gate9833  (.A(g28903), .Z(g29965) ) ;
NAND3   gate9834  (.A(g27907), .B(g2495), .C(g2421), .Z(g28946) ) ;
INV     gate9835  (.A(g28946), .Z(g29967) ) ;
INV     gate9836  (.A(g28803), .Z(II28199) ) ;
INV     gate9837  (.A(II28199), .Z(g29970) ) ;
NAND2   gate9838  (.A(g9586), .B(g27742), .Z(g29018) ) ;
INV     gate9839  (.A(g29018), .Z(g29976) ) ;
NAND3   gate9840  (.A(g27779), .B(g1802), .C(g7315), .Z(g28920) ) ;
INV     gate9841  (.A(g28920), .Z(g29977) ) ;
NAND3   gate9842  (.A(g27837), .B(g1906), .C(g7322), .Z(g28927) ) ;
INV     gate9843  (.A(g28927), .Z(g29978) ) ;
NAND3   gate9844  (.A(g27800), .B(g2227), .C(g7328), .Z(g28935) ) ;
INV     gate9845  (.A(g28935), .Z(g29980) ) ;
NAND3   gate9846  (.A(g27858), .B(g2331), .C(g7335), .Z(g28942) ) ;
INV     gate9847  (.A(g28942), .Z(g29981) ) ;
NAND3   gate9848  (.A(g27937), .B(g2629), .C(g2555), .Z(g28977) ) ;
INV     gate9849  (.A(g28977), .Z(g29983) ) ;
INV     gate9850  (.A(g29018), .Z(g29993) ) ;
NAND2   gate9851  (.A(g9640), .B(g27779), .Z(g29049) ) ;
INV     gate9852  (.A(g29049), .Z(g29994) ) ;
NAND3   gate9853  (.A(g27837), .B(g1936), .C(g7362), .Z(g28955) ) ;
INV     gate9854  (.A(g28955), .Z(g29995) ) ;
NAND3   gate9855  (.A(g27886), .B(g2040), .C(g7369), .Z(g28962) ) ;
INV     gate9856  (.A(g28962), .Z(g29996) ) ;
NAND2   gate9857  (.A(g9649), .B(g27800), .Z(g29060) ) ;
INV     gate9858  (.A(g29060), .Z(g29997) ) ;
NAND3   gate9859  (.A(g27858), .B(g2361), .C(g7380), .Z(g28966) ) ;
INV     gate9860  (.A(g28966), .Z(g29998) ) ;
NAND3   gate9861  (.A(g27907), .B(g2465), .C(g7387), .Z(g28973) ) ;
INV     gate9862  (.A(g28973), .Z(g29999) ) ;
INV     gate9863  (.A(g28709), .Z(II28241) ) ;
INV     gate9864  (.A(II28241), .Z(g30012) ) ;
INV     gate9865  (.A(g29049), .Z(g30016) ) ;
NAND2   gate9866  (.A(g9694), .B(g27837), .Z(g29085) ) ;
INV     gate9867  (.A(g29085), .Z(g30017) ) ;
NAND3   gate9868  (.A(g27886), .B(g2070), .C(g7411), .Z(g28987) ) ;
INV     gate9869  (.A(g28987), .Z(g30018) ) ;
INV     gate9870  (.A(g29060), .Z(g30019) ) ;
NAND2   gate9871  (.A(g9700), .B(g27858), .Z(g29097) ) ;
INV     gate9872  (.A(g29097), .Z(g30020) ) ;
NAND3   gate9873  (.A(g27907), .B(g2495), .C(g7424), .Z(g28994) ) ;
INV     gate9874  (.A(g28994), .Z(g30021) ) ;
NAND3   gate9875  (.A(g27937), .B(g2599), .C(g7431), .Z(g29001) ) ;
INV     gate9876  (.A(g29001), .Z(g30022) ) ;
INV     gate9877  (.A(g29085), .Z(g30036) ) ;
NAND2   gate9878  (.A(g9755), .B(g27886), .Z(g29121) ) ;
INV     gate9879  (.A(g29121), .Z(g30037) ) ;
INV     gate9880  (.A(g29097), .Z(g30038) ) ;
NAND2   gate9881  (.A(g9762), .B(g27907), .Z(g29134) ) ;
INV     gate9882  (.A(g29134), .Z(g30039) ) ;
NAND3   gate9883  (.A(g27937), .B(g2629), .C(g7462), .Z(g29025) ) ;
INV     gate9884  (.A(g29025), .Z(g30040) ) ;
INV     gate9885  (.A(g29018), .Z(g30052) ) ;
INV     gate9886  (.A(g29121), .Z(g30053) ) ;
INV     gate9887  (.A(g29134), .Z(g30054) ) ;
NAND2   gate9888  (.A(g9835), .B(g27937), .Z(g29157) ) ;
INV     gate9889  (.A(g29157), .Z(g30055) ) ;
NAND2   gate9890  (.A(g27742), .B(g9586), .Z(g29015) ) ;
INV     gate9891  (.A(g29015), .Z(g30063) ) ;
INV     gate9892  (.A(g29049), .Z(g30065) ) ;
INV     gate9893  (.A(g29060), .Z(g30067) ) ;
INV     gate9894  (.A(g29157), .Z(g30068) ) ;
INV     gate9895  (.A(g29042), .Z(II28301) ) ;
INV     gate9896  (.A(II28301), .Z(g30072) ) ;
NAND2   gate9897  (.A(g27779), .B(g9640), .Z(g29046) ) ;
INV     gate9898  (.A(g29046), .Z(g30074) ) ;
INV     gate9899  (.A(g29085), .Z(g30076) ) ;
NAND2   gate9900  (.A(g27800), .B(g9649), .Z(g29057) ) ;
INV     gate9901  (.A(g29057), .Z(g30077) ) ;
INV     gate9902  (.A(g29097), .Z(g30079) ) ;
NAND2   gate9903  (.A(g27837), .B(g9694), .Z(g29082) ) ;
INV     gate9904  (.A(g29082), .Z(g30085) ) ;
INV     gate9905  (.A(g29121), .Z(g30087) ) ;
NAND2   gate9906  (.A(g27858), .B(g9700), .Z(g29094) ) ;
INV     gate9907  (.A(g29094), .Z(g30088) ) ;
INV     gate9908  (.A(g29134), .Z(g30090) ) ;
NAND2   gate9909  (.A(g27886), .B(g9755), .Z(g29118) ) ;
INV     gate9910  (.A(g29118), .Z(g30097) ) ;
NAND2   gate9911  (.A(g27907), .B(g9762), .Z(g29131) ) ;
INV     gate9912  (.A(g29131), .Z(g30100) ) ;
INV     gate9913  (.A(g29157), .Z(g30102) ) ;
INV     gate9914  (.A(g29147), .Z(II28336) ) ;
INV     gate9915  (.A(II28336), .Z(g30105) ) ;
NAND2   gate9916  (.A(g27937), .B(g9835), .Z(g29154) ) ;
INV     gate9917  (.A(g29154), .Z(g30113) ) ;
INV     gate9918  (.A(g28367), .Z(II28349) ) ;
INV     gate9919  (.A(II28349), .Z(g30116) ) ;
INV     gate9920  (.A(g28754), .Z(g30142) ) ;
INV     gate9921  (.A(g29185), .Z(II28390) ) ;
INV     gate9922  (.A(II28390), .Z(g30155) ) ;
INV     gate9923  (.A(g29195), .Z(II28419) ) ;
INV     gate9924  (.A(II28419), .Z(g30182) ) ;
AND2    gate9925  (.A(g4608), .B(g27020), .Z(g28144) ) ;
INV     gate9926  (.A(g28144), .Z(g30184) ) ;
AND2    gate9927  (.A(g25869), .B(g27051), .Z(g28114) ) ;
INV     gate9928  (.A(g28114), .Z(II28434) ) ;
INV     gate9929  (.A(II28434), .Z(g30195) ) ;
INV     gate9930  (.A(g28436), .Z(g30206) ) ;
INV     gate9931  (.A(g28443), .Z(II28458) ) ;
INV     gate9932  (.A(II28458), .Z(g30217) ) ;
INV     gate9933  (.A(g28918), .Z(g30218) ) ;
AND2    gate9934  (.A(g27282), .B(g10288), .Z(g28652) ) ;
INV     gate9935  (.A(g28652), .Z(II28480) ) ;
INV     gate9936  (.A(II28480), .Z(g30237) ) ;
INV     gate9937  (.A(g28463), .Z(g30259) ) ;
NAND3   gate9938  (.A(g27742), .B(g7308), .C(g7252), .Z(g28736) ) ;
INV     gate9939  (.A(g28736), .Z(g30292) ) ;
INV     gate9940  (.A(g28954), .Z(II28540) ) ;
INV     gate9941  (.A(II28540), .Z(g30295) ) ;
AND4    gate9942  (.A(g17292), .B(g25169), .C(g26424), .D(g27395), .Z(g28889) ) ;
INV     gate9943  (.A(g28889), .Z(g30296) ) ;
NAND3   gate9944  (.A(g27779), .B(g7356), .C(g7275), .Z(g28758) ) ;
INV     gate9945  (.A(g28758), .Z(g30297) ) ;
NAND3   gate9946  (.A(g27800), .B(g7374), .C(g7280), .Z(g28765) ) ;
INV     gate9947  (.A(g28765), .Z(g30299) ) ;
INV     gate9948  (.A(g28147), .Z(II28548) ) ;
INV     gate9949  (.A(II28548), .Z(g30301) ) ;
AND4    gate9950  (.A(g17317), .B(g25183), .C(g26424), .D(g27416), .Z(g28924) ) ;
INV     gate9951  (.A(g28924), .Z(g30302) ) ;
NAND3   gate9952  (.A(g27837), .B(g7405), .C(g7322), .Z(g28786) ) ;
INV     gate9953  (.A(g28786), .Z(g30303) ) ;
AND4    gate9954  (.A(g17321), .B(g25184), .C(g26424), .D(g27421), .Z(g28939) ) ;
INV     gate9955  (.A(g28939), .Z(g30305) ) ;
NAND3   gate9956  (.A(g27858), .B(g7418), .C(g7335), .Z(g28796) ) ;
INV     gate9957  (.A(g28796), .Z(g30306) ) ;
AND4    gate9958  (.A(g17401), .B(g25194), .C(g26424), .D(g27440), .Z(g28959) ) ;
INV     gate9959  (.A(g28959), .Z(g30309) ) ;
NAND3   gate9960  (.A(g27886), .B(g7451), .C(g7369), .Z(g28830) ) ;
INV     gate9961  (.A(g28830), .Z(g30310) ) ;
AND4    gate9962  (.A(g17405), .B(g25196), .C(g26424), .D(g27445), .Z(g28970) ) ;
INV     gate9963  (.A(g28970), .Z(g30312) ) ;
NAND3   gate9964  (.A(g27907), .B(g7456), .C(g7387), .Z(g28843) ) ;
INV     gate9965  (.A(g28843), .Z(g30313) ) ;
INV     gate9966  (.A(g28274), .Z(g30318) ) ;
INV     gate9967  (.A(g28274), .Z(II28572) ) ;
INV     gate9968  (.A(II28572), .Z(g30321) ) ;
INV     gate9969  (.A(g28431), .Z(g30322) ) ;
INV     gate9970  (.A(g28431), .Z(II28576) ) ;
INV     gate9971  (.A(II28576), .Z(g30325) ) ;
INV     gate9972  (.A(g29474), .Z(II28579) ) ;
INV     gate9973  (.A(g30116), .Z(II28582) ) ;
INV     gate9974  (.A(g30217), .Z(II28585) ) ;
INV     gate9975  (.A(g29368), .Z(II28588) ) ;
INV     gate9976  (.A(g29371), .Z(II28591) ) ;
INV     gate9977  (.A(g29379), .Z(II28594) ) ;
INV     gate9978  (.A(g29374), .Z(II28597) ) ;
INV     gate9979  (.A(g30301), .Z(II28832) ) ;
INV     gate9980  (.A(II28832), .Z(g30565) ) ;
INV     gate9981  (.A(g29930), .Z(g30567) ) ;
INV     gate9982  (.A(g29339), .Z(g30568) ) ;
INV     gate9983  (.A(g29372), .Z(II28838) ) ;
INV     gate9984  (.A(II28838), .Z(g30569) ) ;
INV     gate9985  (.A(g29945), .Z(g30572) ) ;
INV     gate9986  (.A(g29956), .Z(g30578) ) ;
INV     gate9987  (.A(g29317), .Z(II28851) ) ;
INV     gate9988  (.A(II28851), .Z(g30591) ) ;
INV     gate9989  (.A(g29970), .Z(g30593) ) ;
OR2     gate9990  (.A(g28150), .B(g28141), .Z(g29730) ) ;
INV     gate9991  (.A(g29730), .Z(II28866) ) ;
INV     gate9992  (.A(II28866), .Z(g30606) ) ;
INV     gate9993  (.A(g30072), .Z(II28872) ) ;
INV     gate9994  (.A(II28872), .Z(g30610) ) ;
INV     gate9995  (.A(g30105), .Z(II28883) ) ;
INV     gate9996  (.A(II28883), .Z(g30729) ) ;
INV     gate9997  (.A(g30155), .Z(II28897) ) ;
INV     gate9998  (.A(II28897), .Z(g30917) ) ;
INV     gate9999  (.A(g30182), .Z(II28908) ) ;
INV     gate10000  (.A(II28908), .Z(g30928) ) ;
INV     gate10001  (.A(g30322), .Z(II28913) ) ;
INV     gate10002  (.A(II28913), .Z(g30931) ) ;
NAND2   gate10003  (.A(g28363), .B(g13634), .Z(g29657) ) ;
INV     gate10004  (.A(g29657), .Z(g30983) ) ;
NAND2   gate10005  (.A(g28376), .B(g13672), .Z(g29672) ) ;
INV     gate10006  (.A(g29672), .Z(g30989) ) ;
NAND2   gate10007  (.A(g28381), .B(g13676), .Z(g29676) ) ;
INV     gate10008  (.A(g29676), .Z(g30990) ) ;
AND3    gate10009  (.A(g29197), .B(g26424), .C(g22763), .Z(g29987) ) ;
INV     gate10010  (.A(g29987), .Z(II28925) ) ;
INV     gate10011  (.A(II28925), .Z(g30991) ) ;
NAND2   gate10012  (.A(g28391), .B(g13709), .Z(g29694) ) ;
INV     gate10013  (.A(g29694), .Z(g30996) ) ;
NAND2   gate10014  (.A(g28395), .B(g13712), .Z(g29702) ) ;
INV     gate10015  (.A(g29702), .Z(g30997) ) ;
NAND2   gate10016  (.A(g28406), .B(g13739), .Z(g29719) ) ;
INV     gate10017  (.A(g29719), .Z(g30998) ) ;
NAND2   gate10018  (.A(g28410), .B(g13742), .Z(g29722) ) ;
INV     gate10019  (.A(g29722), .Z(g30999) ) ;
NAND2   gate10020  (.A(g28421), .B(g13779), .Z(g29737) ) ;
INV     gate10021  (.A(g29737), .Z(g31000) ) ;
NAND3   gate10022  (.A(g153), .B(g28353), .C(g23042), .Z(g29679) ) ;
INV     gate10023  (.A(g29679), .Z(g31013) ) ;
NAND3   gate10024  (.A(g294), .B(g28444), .C(g23204), .Z(g29778) ) ;
INV     gate10025  (.A(g29778), .Z(g31138) ) ;
NOR3    gate10026  (.A(g28380), .B(g8236), .C(g8354), .Z(g29675) ) ;
INV     gate10027  (.A(g29675), .Z(II29002) ) ;
INV     gate10028  (.A(II29002), .Z(g31189) ) ;
NOR3    gate10029  (.A(g28399), .B(g8284), .C(g8404), .Z(g29705) ) ;
INV     gate10030  (.A(g29705), .Z(II29013) ) ;
INV     gate10031  (.A(II29013), .Z(g31213) ) ;
INV     gate10032  (.A(g29744), .Z(g31227) ) ;
NOR3    gate10033  (.A(g8681), .B(g28504), .C(g11083), .Z(g29916) ) ;
INV     gate10034  (.A(g29916), .Z(g31239) ) ;
NOR3    gate10035  (.A(g8808), .B(g28500), .C(g12259), .Z(g29933) ) ;
INV     gate10036  (.A(g29933), .Z(g31243) ) ;
AND3    gate10037  (.A(g26424), .B(g22763), .C(g28172), .Z(g29382) ) ;
INV     gate10038  (.A(g29382), .Z(II29139) ) ;
INV     gate10039  (.A(II29139), .Z(g31479) ) ;
AND3    gate10040  (.A(g26424), .B(g22763), .C(g28179), .Z(g29384) ) ;
INV     gate10041  (.A(g29384), .Z(II29149) ) ;
INV     gate10042  (.A(II29149), .Z(g31487) ) ;
INV     gate10043  (.A(g30012), .Z(II29182) ) ;
INV     gate10044  (.A(g30012), .Z(II29185) ) ;
INV     gate10045  (.A(II29185), .Z(g31522) ) ;
INV     gate10046  (.A(g30237), .Z(II29199) ) ;
INV     gate10047  (.A(II29199), .Z(g31578) ) ;
INV     gate10048  (.A(g29505), .Z(II29204) ) ;
INV     gate10049  (.A(II29204), .Z(g31596) ) ;
OR2     gate10050  (.A(g28236), .B(g27246), .Z(g30293) ) ;
INV     gate10051  (.A(g30293), .Z(II29207) ) ;
INV     gate10052  (.A(II29207), .Z(g31601) ) ;
INV     gate10053  (.A(g29653), .Z(g31608) ) ;
OR2     gate10054  (.A(g28245), .B(g27251), .Z(g30298) ) ;
INV     gate10055  (.A(g30298), .Z(II29211) ) ;
INV     gate10056  (.A(II29211), .Z(g31609) ) ;
OR2     gate10057  (.A(g28246), .B(g27252), .Z(g30300) ) ;
INV     gate10058  (.A(g30300), .Z(II29214) ) ;
INV     gate10059  (.A(II29214), .Z(g31616) ) ;
INV     gate10060  (.A(g29669), .Z(g31623) ) ;
OR2     gate10061  (.A(g28255), .B(g27259), .Z(g30304) ) ;
INV     gate10062  (.A(g30304), .Z(II29218) ) ;
INV     gate10063  (.A(II29218), .Z(g31624) ) ;
OR2     gate10064  (.A(g28256), .B(g27260), .Z(g30307) ) ;
INV     gate10065  (.A(g30307), .Z(II29221) ) ;
INV     gate10066  (.A(II29221), .Z(g31631) ) ;
INV     gate10067  (.A(g29689), .Z(g31638) ) ;
OR2     gate10068  (.A(g28265), .B(g27265), .Z(g30311) ) ;
INV     gate10069  (.A(g30311), .Z(II29225) ) ;
INV     gate10070  (.A(II29225), .Z(g31639) ) ;
OR2     gate10071  (.A(g28268), .B(g27266), .Z(g30314) ) ;
INV     gate10072  (.A(g30314), .Z(II29228) ) ;
INV     gate10073  (.A(II29228), .Z(g31646) ) ;
INV     gate10074  (.A(g29713), .Z(g31653) ) ;
INV     gate10075  (.A(g30295), .Z(II29233) ) ;
INV     gate10076  (.A(II29233), .Z(g31655) ) ;
INV     gate10077  (.A(g29498), .Z(II29236) ) ;
INV     gate10078  (.A(g29498), .Z(II29239) ) ;
INV     gate10079  (.A(II29239), .Z(g31657) ) ;
OR2     gate10080  (.A(g28284), .B(g27270), .Z(g29313) ) ;
INV     gate10081  (.A(g29313), .Z(II29242) ) ;
INV     gate10082  (.A(II29242), .Z(g31658) ) ;
INV     gate10083  (.A(g29491), .Z(II29245) ) ;
INV     gate10084  (.A(g29491), .Z(II29248) ) ;
INV     gate10085  (.A(II29248), .Z(g31666) ) ;
INV     gate10086  (.A(g30142), .Z(g31667) ) ;
OR2     gate10087  (.A(g28191), .B(g28186), .Z(g30286) ) ;
INV     gate10088  (.A(g30286), .Z(II29337) ) ;
INV     gate10089  (.A(II29337), .Z(g31771) ) ;
INV     gate10090  (.A(g30218), .Z(II29363) ) ;
INV     gate10091  (.A(II29363), .Z(g31791) ) ;
INV     gate10092  (.A(g30321), .Z(II29368) ) ;
INV     gate10093  (.A(II29368), .Z(g31794) ) ;
INV     gate10094  (.A(g30325), .Z(II29371) ) ;
INV     gate10095  (.A(II29371), .Z(g31795) ) ;
INV     gate10096  (.A(g29385), .Z(g31796) ) ;
INV     gate10097  (.A(g29385), .Z(g31797) ) ;
INV     gate10098  (.A(g29385), .Z(g31798) ) ;
INV     gate10099  (.A(g29385), .Z(g31799) ) ;
INV     gate10100  (.A(g29385), .Z(g31800) ) ;
INV     gate10101  (.A(g29385), .Z(g31801) ) ;
INV     gate10102  (.A(g29385), .Z(g31802) ) ;
INV     gate10103  (.A(g29385), .Z(g31803) ) ;
INV     gate10104  (.A(g29385), .Z(g31804) ) ;
INV     gate10105  (.A(g29385), .Z(g31805) ) ;
INV     gate10106  (.A(g29385), .Z(g31806) ) ;
INV     gate10107  (.A(g29385), .Z(g31807) ) ;
INV     gate10108  (.A(g29385), .Z(g31808) ) ;
INV     gate10109  (.A(g29385), .Z(g31809) ) ;
INV     gate10110  (.A(g29385), .Z(g31810) ) ;
INV     gate10111  (.A(g29385), .Z(g31811) ) ;
INV     gate10112  (.A(g29385), .Z(g31812) ) ;
INV     gate10113  (.A(g29385), .Z(g31813) ) ;
INV     gate10114  (.A(g29385), .Z(g31814) ) ;
INV     gate10115  (.A(g29385), .Z(g31815) ) ;
INV     gate10116  (.A(g29385), .Z(g31816) ) ;
INV     gate10117  (.A(g29385), .Z(g31817) ) ;
INV     gate10118  (.A(g29385), .Z(g31818) ) ;
INV     gate10119  (.A(g29385), .Z(g31819) ) ;
INV     gate10120  (.A(g29385), .Z(g31820) ) ;
INV     gate10121  (.A(g29385), .Z(g31821) ) ;
INV     gate10122  (.A(g29385), .Z(g31822) ) ;
INV     gate10123  (.A(g29385), .Z(g31823) ) ;
INV     gate10124  (.A(g29385), .Z(g31824) ) ;
INV     gate10125  (.A(g29385), .Z(g31825) ) ;
INV     gate10126  (.A(g29385), .Z(g31826) ) ;
INV     gate10127  (.A(g29385), .Z(g31827) ) ;
INV     gate10128  (.A(g29385), .Z(g31828) ) ;
INV     gate10129  (.A(g29385), .Z(g31829) ) ;
INV     gate10130  (.A(g29385), .Z(g31830) ) ;
INV     gate10131  (.A(g29385), .Z(g31831) ) ;
INV     gate10132  (.A(g29385), .Z(g31832) ) ;
INV     gate10133  (.A(g29385), .Z(g31833) ) ;
INV     gate10134  (.A(g29385), .Z(g31834) ) ;
INV     gate10135  (.A(g29385), .Z(g31835) ) ;
INV     gate10136  (.A(g29385), .Z(g31836) ) ;
INV     gate10137  (.A(g29385), .Z(g31837) ) ;
INV     gate10138  (.A(g29385), .Z(g31838) ) ;
INV     gate10139  (.A(g29385), .Z(g31839) ) ;
INV     gate10140  (.A(g29385), .Z(g31840) ) ;
INV     gate10141  (.A(g29385), .Z(g31841) ) ;
INV     gate10142  (.A(g29385), .Z(g31842) ) ;
INV     gate10143  (.A(g29385), .Z(g31843) ) ;
INV     gate10144  (.A(g29385), .Z(g31844) ) ;
INV     gate10145  (.A(g29385), .Z(g31845) ) ;
INV     gate10146  (.A(g29385), .Z(g31846) ) ;
INV     gate10147  (.A(g29385), .Z(g31847) ) ;
INV     gate10148  (.A(g29385), .Z(g31848) ) ;
INV     gate10149  (.A(g29385), .Z(g31849) ) ;
INV     gate10150  (.A(g29385), .Z(g31850) ) ;
INV     gate10151  (.A(g29385), .Z(g31851) ) ;
INV     gate10152  (.A(g29385), .Z(g31852) ) ;
INV     gate10153  (.A(g29385), .Z(g31853) ) ;
INV     gate10154  (.A(g29385), .Z(g31854) ) ;
INV     gate10155  (.A(g29385), .Z(g31855) ) ;
INV     gate10156  (.A(g29385), .Z(g31856) ) ;
INV     gate10157  (.A(g29385), .Z(g31857) ) ;
INV     gate10158  (.A(g29385), .Z(g31858) ) ;
INV     gate10159  (.A(g29385), .Z(g31859) ) ;
INV     gate10160  (.A(g30610), .Z(II29438) ) ;
INV     gate10161  (.A(g30917), .Z(II29441) ) ;
INV     gate10162  (.A(g30928), .Z(II29444) ) ;
INV     gate10163  (.A(g30729), .Z(II29447) ) ;
INV     gate10164  (.A(g30991), .Z(g31937) ) ;
INV     gate10165  (.A(g31189), .Z(g31945) ) ;
OR2     gate10166  (.A(II29351), .B(II29352), .Z(g31783) ) ;
INV     gate10167  (.A(g31783), .Z(II29571) ) ;
INV     gate10168  (.A(II29571), .Z(g32015) ) ;
INV     gate10169  (.A(g30565), .Z(II29579) ) ;
INV     gate10170  (.A(II29579), .Z(g32021) ) ;
INV     gate10171  (.A(g30591), .Z(II29582) ) ;
INV     gate10172  (.A(II29582), .Z(g32024) ) ;
INV     gate10173  (.A(g31655), .Z(II29585) ) ;
INV     gate10174  (.A(II29585), .Z(g32027) ) ;
NOR2    gate10175  (.A(g29803), .B(g29835), .Z(g30929) ) ;
INV     gate10176  (.A(g30929), .Z(g32033) ) ;
NOR2    gate10177  (.A(g29836), .B(g29850), .Z(g30934) ) ;
INV     gate10178  (.A(g30934), .Z(g32038) ) ;
NAND3   gate10179  (.A(g27163), .B(g29497), .C(g19644), .Z(g31003) ) ;
INV     gate10180  (.A(g31003), .Z(g32090) ) ;
NAND3   gate10181  (.A(g27187), .B(g29503), .C(g19644), .Z(g31009) ) ;
INV     gate10182  (.A(g31009), .Z(g32099) ) ;
NOR2    gate10183  (.A(g30004), .B(g30026), .Z(g31008) ) ;
INV     gate10184  (.A(g31008), .Z(g32118) ) ;
NOR3    gate10185  (.A(g8033), .B(g29679), .C(g24732), .Z(g31134) ) ;
INV     gate10186  (.A(g31134), .Z(g32137) ) ;
NOR3    gate10187  (.A(g8522), .B(g29778), .C(g24825), .Z(g31233) ) ;
INV     gate10188  (.A(g31233), .Z(g32138) ) ;
INV     gate10189  (.A(g30931), .Z(II29717) ) ;
INV     gate10190  (.A(g30931), .Z(II29720) ) ;
INV     gate10191  (.A(II29720), .Z(g32186) ) ;
NAND3   gate10192  (.A(g767), .B(g29916), .C(g11679), .Z(g31262) ) ;
INV     gate10193  (.A(g31262), .Z(g32192) ) ;
NAND3   gate10194  (.A(g599), .B(g29933), .C(g12323), .Z(g31509) ) ;
INV     gate10195  (.A(g31509), .Z(g32201) ) ;
INV     gate10196  (.A(g31596), .Z(g32318) ) ;
INV     gate10197  (.A(g31522), .Z(g32329) ) ;
INV     gate10198  (.A(g31578), .Z(II29891) ) ;
INV     gate10199  (.A(II29891), .Z(g32363) ) ;
INV     gate10200  (.A(g31771), .Z(II29894) ) ;
INV     gate10201  (.A(II29894), .Z(g32364) ) ;
OR2     gate10202  (.A(g29765), .B(g29755), .Z(g30984) ) ;
INV     gate10203  (.A(g30984), .Z(g32377) ) ;
INV     gate10204  (.A(g31791), .Z(II29909) ) ;
INV     gate10205  (.A(II29909), .Z(g32381) ) ;
INV     gate10206  (.A(g31657), .Z(g32382) ) ;
OR2     gate10207  (.A(g29529), .B(g29520), .Z(g30605) ) ;
INV     gate10208  (.A(g30605), .Z(II29913) ) ;
INV     gate10209  (.A(II29913), .Z(g32383) ) ;
INV     gate10210  (.A(g31666), .Z(g32384) ) ;
NOR2    gate10211  (.A(g16662), .B(g29810), .Z(g30922) ) ;
INV     gate10212  (.A(g30922), .Z(g32393) ) ;
NOR2    gate10213  (.A(g16279), .B(g29718), .Z(g30601) ) ;
INV     gate10214  (.A(g30601), .Z(g32394) ) ;
INV     gate10215  (.A(g30606), .Z(II29936) ) ;
INV     gate10216  (.A(II29936), .Z(g32404) ) ;
INV     gate10217  (.A(g31667), .Z(II29939) ) ;
INV     gate10218  (.A(II29939), .Z(g32407) ) ;
OR2     gate10219  (.A(g29358), .B(g29353), .Z(g31591) ) ;
INV     gate10220  (.A(g31591), .Z(g32415) ) ;
INV     gate10221  (.A(g31213), .Z(g32421) ) ;
INV     gate10222  (.A(g30984), .Z(g32430) ) ;
INV     gate10223  (.A(g30984), .Z(II29961) ) ;
INV     gate10224  (.A(II29961), .Z(g32433) ) ;
INV     gate10225  (.A(g31189), .Z(g32434) ) ;
INV     gate10226  (.A(g31189), .Z(II29965) ) ;
INV     gate10227  (.A(II29965), .Z(g32437) ) ;
INV     gate10228  (.A(g30991), .Z(g32438) ) ;
INV     gate10229  (.A(g30991), .Z(II29969) ) ;
INV     gate10230  (.A(II29969), .Z(g32441) ) ;
INV     gate10231  (.A(g31213), .Z(g32442) ) ;
INV     gate10232  (.A(g31213), .Z(II29973) ) ;
INV     gate10233  (.A(II29973), .Z(g32445) ) ;
INV     gate10234  (.A(g31596), .Z(g32446) ) ;
INV     gate10235  (.A(g31596), .Z(II29977) ) ;
INV     gate10236  (.A(II29977), .Z(g32449) ) ;
INV     gate10237  (.A(g31591), .Z(g32450) ) ;
INV     gate10238  (.A(g31591), .Z(II29981) ) ;
INV     gate10239  (.A(II29981), .Z(g32453) ) ;
AND2    gate10240  (.A(g24952), .B(g29814), .Z(g31376) ) ;
INV     gate10241  (.A(g31376), .Z(g32456) ) ;
AND2    gate10242  (.A(g29814), .B(g22319), .Z(g30735) ) ;
INV     gate10243  (.A(g30735), .Z(g32457) ) ;
AND2    gate10244  (.A(g29814), .B(g22332), .Z(g30825) ) ;
INV     gate10245  (.A(g30825), .Z(g32458) ) ;
AND2    gate10246  (.A(g29814), .B(g25985), .Z(g31070) ) ;
INV     gate10247  (.A(g31070), .Z(g32459) ) ;
AND2    gate10248  (.A(g19128), .B(g29814), .Z(g31194) ) ;
INV     gate10249  (.A(g31194), .Z(g32460) ) ;
AND2    gate10250  (.A(g20154), .B(g29814), .Z(g30614) ) ;
INV     gate10251  (.A(g30614), .Z(g32461) ) ;
AND2    gate10252  (.A(g20175), .B(g29814), .Z(g30673) ) ;
INV     gate10253  (.A(g30673), .Z(g32462) ) ;
AND2    gate10254  (.A(g19050), .B(g29814), .Z(g31566) ) ;
INV     gate10255  (.A(g31566), .Z(g32463) ) ;
INV     gate10256  (.A(g30735), .Z(g32464) ) ;
INV     gate10257  (.A(g30825), .Z(g32465) ) ;
INV     gate10258  (.A(g31070), .Z(g32466) ) ;
INV     gate10259  (.A(g31194), .Z(g32467) ) ;
INV     gate10260  (.A(g30614), .Z(g32468) ) ;
INV     gate10261  (.A(g30673), .Z(g32469) ) ;
INV     gate10262  (.A(g31566), .Z(g32470) ) ;
INV     gate10263  (.A(g31376), .Z(g32471) ) ;
INV     gate10264  (.A(g30825), .Z(g32472) ) ;
INV     gate10265  (.A(g31070), .Z(g32473) ) ;
INV     gate10266  (.A(g31194), .Z(g32474) ) ;
INV     gate10267  (.A(g30614), .Z(g32475) ) ;
INV     gate10268  (.A(g30673), .Z(g32476) ) ;
INV     gate10269  (.A(g31566), .Z(g32477) ) ;
INV     gate10270  (.A(g31376), .Z(g32478) ) ;
INV     gate10271  (.A(g30735), .Z(g32479) ) ;
INV     gate10272  (.A(g31070), .Z(g32480) ) ;
INV     gate10273  (.A(g31194), .Z(g32481) ) ;
INV     gate10274  (.A(g30614), .Z(g32482) ) ;
INV     gate10275  (.A(g30673), .Z(g32483) ) ;
INV     gate10276  (.A(g31566), .Z(g32484) ) ;
INV     gate10277  (.A(g31376), .Z(g32485) ) ;
INV     gate10278  (.A(g30735), .Z(g32486) ) ;
INV     gate10279  (.A(g30825), .Z(g32487) ) ;
INV     gate10280  (.A(g31194), .Z(g32488) ) ;
INV     gate10281  (.A(g30614), .Z(g32489) ) ;
INV     gate10282  (.A(g30673), .Z(g32490) ) ;
INV     gate10283  (.A(g31566), .Z(g32491) ) ;
INV     gate10284  (.A(g31376), .Z(g32492) ) ;
INV     gate10285  (.A(g30735), .Z(g32493) ) ;
INV     gate10286  (.A(g30825), .Z(g32494) ) ;
INV     gate10287  (.A(g31070), .Z(g32495) ) ;
INV     gate10288  (.A(g30614), .Z(g32496) ) ;
INV     gate10289  (.A(g30673), .Z(g32497) ) ;
INV     gate10290  (.A(g31566), .Z(g32498) ) ;
INV     gate10291  (.A(g31376), .Z(g32499) ) ;
INV     gate10292  (.A(g30735), .Z(g32500) ) ;
INV     gate10293  (.A(g30825), .Z(g32501) ) ;
INV     gate10294  (.A(g31070), .Z(g32502) ) ;
INV     gate10295  (.A(g31194), .Z(g32503) ) ;
INV     gate10296  (.A(g30673), .Z(g32504) ) ;
INV     gate10297  (.A(g31566), .Z(g32505) ) ;
INV     gate10298  (.A(g31376), .Z(g32506) ) ;
INV     gate10299  (.A(g30735), .Z(g32507) ) ;
INV     gate10300  (.A(g30825), .Z(g32508) ) ;
INV     gate10301  (.A(g31070), .Z(g32509) ) ;
INV     gate10302  (.A(g31194), .Z(g32510) ) ;
INV     gate10303  (.A(g30614), .Z(g32511) ) ;
INV     gate10304  (.A(g31566), .Z(g32512) ) ;
INV     gate10305  (.A(g31376), .Z(g32513) ) ;
INV     gate10306  (.A(g30735), .Z(g32514) ) ;
INV     gate10307  (.A(g30825), .Z(g32515) ) ;
INV     gate10308  (.A(g31070), .Z(g32516) ) ;
INV     gate10309  (.A(g31194), .Z(g32517) ) ;
INV     gate10310  (.A(g30614), .Z(g32518) ) ;
INV     gate10311  (.A(g30673), .Z(g32519) ) ;
INV     gate10312  (.A(g31376), .Z(g32521) ) ;
INV     gate10313  (.A(g30735), .Z(g32522) ) ;
INV     gate10314  (.A(g30825), .Z(g32523) ) ;
INV     gate10315  (.A(g31070), .Z(g32524) ) ;
AND2    gate10316  (.A(g19128), .B(g29814), .Z(g31170) ) ;
INV     gate10317  (.A(g31170), .Z(g32525) ) ;
INV     gate10318  (.A(g30614), .Z(g32526) ) ;
INV     gate10319  (.A(g30673), .Z(g32527) ) ;
AND2    gate10320  (.A(g19050), .B(g29814), .Z(g31554) ) ;
INV     gate10321  (.A(g31554), .Z(g32528) ) ;
INV     gate10322  (.A(g30735), .Z(g32529) ) ;
INV     gate10323  (.A(g30825), .Z(g32530) ) ;
INV     gate10324  (.A(g31070), .Z(g32531) ) ;
INV     gate10325  (.A(g31170), .Z(g32532) ) ;
INV     gate10326  (.A(g30614), .Z(g32533) ) ;
INV     gate10327  (.A(g30673), .Z(g32534) ) ;
INV     gate10328  (.A(g31554), .Z(g32535) ) ;
INV     gate10329  (.A(g31376), .Z(g32536) ) ;
INV     gate10330  (.A(g30825), .Z(g32537) ) ;
INV     gate10331  (.A(g31070), .Z(g32538) ) ;
INV     gate10332  (.A(g31170), .Z(g32539) ) ;
INV     gate10333  (.A(g30614), .Z(g32540) ) ;
INV     gate10334  (.A(g30673), .Z(g32541) ) ;
INV     gate10335  (.A(g31554), .Z(g32542) ) ;
INV     gate10336  (.A(g31376), .Z(g32543) ) ;
INV     gate10337  (.A(g30735), .Z(g32544) ) ;
INV     gate10338  (.A(g31070), .Z(g32545) ) ;
INV     gate10339  (.A(g31170), .Z(g32546) ) ;
INV     gate10340  (.A(g30614), .Z(g32547) ) ;
INV     gate10341  (.A(g30673), .Z(g32548) ) ;
INV     gate10342  (.A(g31554), .Z(g32549) ) ;
INV     gate10343  (.A(g31376), .Z(g32550) ) ;
INV     gate10344  (.A(g30735), .Z(g32551) ) ;
INV     gate10345  (.A(g30825), .Z(g32552) ) ;
INV     gate10346  (.A(g31170), .Z(g32553) ) ;
INV     gate10347  (.A(g30614), .Z(g32554) ) ;
INV     gate10348  (.A(g30673), .Z(g32555) ) ;
INV     gate10349  (.A(g31554), .Z(g32556) ) ;
INV     gate10350  (.A(g31376), .Z(g32557) ) ;
INV     gate10351  (.A(g30735), .Z(g32558) ) ;
INV     gate10352  (.A(g30825), .Z(g32559) ) ;
INV     gate10353  (.A(g31070), .Z(g32560) ) ;
INV     gate10354  (.A(g30614), .Z(g32561) ) ;
INV     gate10355  (.A(g30673), .Z(g32562) ) ;
INV     gate10356  (.A(g31554), .Z(g32563) ) ;
INV     gate10357  (.A(g31376), .Z(g32564) ) ;
INV     gate10358  (.A(g30735), .Z(g32565) ) ;
INV     gate10359  (.A(g30825), .Z(g32566) ) ;
INV     gate10360  (.A(g31070), .Z(g32567) ) ;
INV     gate10361  (.A(g31170), .Z(g32568) ) ;
INV     gate10362  (.A(g30673), .Z(g32569) ) ;
INV     gate10363  (.A(g31554), .Z(g32570) ) ;
INV     gate10364  (.A(g31376), .Z(g32571) ) ;
INV     gate10365  (.A(g30735), .Z(g32572) ) ;
INV     gate10366  (.A(g30825), .Z(g32573) ) ;
INV     gate10367  (.A(g31070), .Z(g32574) ) ;
INV     gate10368  (.A(g31170), .Z(g32575) ) ;
INV     gate10369  (.A(g30614), .Z(g32576) ) ;
INV     gate10370  (.A(g31554), .Z(g32577) ) ;
INV     gate10371  (.A(g31376), .Z(g32578) ) ;
INV     gate10372  (.A(g30735), .Z(g32579) ) ;
INV     gate10373  (.A(g30825), .Z(g32580) ) ;
INV     gate10374  (.A(g31070), .Z(g32581) ) ;
INV     gate10375  (.A(g31170), .Z(g32582) ) ;
INV     gate10376  (.A(g30614), .Z(g32583) ) ;
INV     gate10377  (.A(g30673), .Z(g32584) ) ;
INV     gate10378  (.A(g31376), .Z(g32586) ) ;
INV     gate10379  (.A(g30735), .Z(g32587) ) ;
INV     gate10380  (.A(g30825), .Z(g32588) ) ;
INV     gate10381  (.A(g31070), .Z(g32589) ) ;
AND2    gate10382  (.A(g19128), .B(g29814), .Z(g31154) ) ;
INV     gate10383  (.A(g31154), .Z(g32590) ) ;
INV     gate10384  (.A(g30614), .Z(g32591) ) ;
INV     gate10385  (.A(g30673), .Z(g32592) ) ;
AND2    gate10386  (.A(g19050), .B(g29814), .Z(g31542) ) ;
INV     gate10387  (.A(g31542), .Z(g32593) ) ;
INV     gate10388  (.A(g30735), .Z(g32594) ) ;
INV     gate10389  (.A(g30825), .Z(g32595) ) ;
INV     gate10390  (.A(g31070), .Z(g32596) ) ;
INV     gate10391  (.A(g31154), .Z(g32597) ) ;
INV     gate10392  (.A(g30614), .Z(g32598) ) ;
INV     gate10393  (.A(g30673), .Z(g32599) ) ;
INV     gate10394  (.A(g31542), .Z(g32600) ) ;
INV     gate10395  (.A(g31376), .Z(g32601) ) ;
INV     gate10396  (.A(g30825), .Z(g32602) ) ;
INV     gate10397  (.A(g31070), .Z(g32603) ) ;
INV     gate10398  (.A(g31154), .Z(g32604) ) ;
INV     gate10399  (.A(g30614), .Z(g32605) ) ;
INV     gate10400  (.A(g30673), .Z(g32606) ) ;
INV     gate10401  (.A(g31542), .Z(g32607) ) ;
INV     gate10402  (.A(g31376), .Z(g32608) ) ;
INV     gate10403  (.A(g30735), .Z(g32609) ) ;
INV     gate10404  (.A(g31070), .Z(g32610) ) ;
INV     gate10405  (.A(g31154), .Z(g32611) ) ;
INV     gate10406  (.A(g30614), .Z(g32612) ) ;
INV     gate10407  (.A(g30673), .Z(g32613) ) ;
INV     gate10408  (.A(g31542), .Z(g32614) ) ;
INV     gate10409  (.A(g31376), .Z(g32615) ) ;
INV     gate10410  (.A(g30735), .Z(g32616) ) ;
INV     gate10411  (.A(g30825), .Z(g32617) ) ;
INV     gate10412  (.A(g31154), .Z(g32618) ) ;
INV     gate10413  (.A(g30614), .Z(g32619) ) ;
INV     gate10414  (.A(g30673), .Z(g32620) ) ;
INV     gate10415  (.A(g31542), .Z(g32621) ) ;
INV     gate10416  (.A(g31376), .Z(g32622) ) ;
INV     gate10417  (.A(g30735), .Z(g32623) ) ;
INV     gate10418  (.A(g30825), .Z(g32624) ) ;
INV     gate10419  (.A(g31070), .Z(g32625) ) ;
INV     gate10420  (.A(g30614), .Z(g32626) ) ;
INV     gate10421  (.A(g30673), .Z(g32627) ) ;
INV     gate10422  (.A(g31542), .Z(g32628) ) ;
INV     gate10423  (.A(g31376), .Z(g32629) ) ;
INV     gate10424  (.A(g30735), .Z(g32630) ) ;
INV     gate10425  (.A(g30825), .Z(g32631) ) ;
INV     gate10426  (.A(g31070), .Z(g32632) ) ;
INV     gate10427  (.A(g31154), .Z(g32633) ) ;
INV     gate10428  (.A(g30673), .Z(g32634) ) ;
INV     gate10429  (.A(g31542), .Z(g32635) ) ;
INV     gate10430  (.A(g31376), .Z(g32636) ) ;
INV     gate10431  (.A(g30735), .Z(g32637) ) ;
INV     gate10432  (.A(g30825), .Z(g32638) ) ;
INV     gate10433  (.A(g31070), .Z(g32639) ) ;
INV     gate10434  (.A(g31154), .Z(g32640) ) ;
INV     gate10435  (.A(g30614), .Z(g32641) ) ;
INV     gate10436  (.A(g31542), .Z(g32642) ) ;
INV     gate10437  (.A(g31376), .Z(g32643) ) ;
INV     gate10438  (.A(g30735), .Z(g32644) ) ;
INV     gate10439  (.A(g30825), .Z(g32645) ) ;
INV     gate10440  (.A(g31070), .Z(g32646) ) ;
INV     gate10441  (.A(g31154), .Z(g32647) ) ;
INV     gate10442  (.A(g30614), .Z(g32648) ) ;
INV     gate10443  (.A(g30673), .Z(g32649) ) ;
INV     gate10444  (.A(g31376), .Z(g32651) ) ;
INV     gate10445  (.A(g30735), .Z(g32652) ) ;
INV     gate10446  (.A(g30825), .Z(g32653) ) ;
INV     gate10447  (.A(g31070), .Z(g32654) ) ;
INV     gate10448  (.A(g30614), .Z(g32655) ) ;
INV     gate10449  (.A(g30673), .Z(g32656) ) ;
AND2    gate10450  (.A(g19050), .B(g29814), .Z(g31528) ) ;
INV     gate10451  (.A(g31528), .Z(g32657) ) ;
AND2    gate10452  (.A(g19128), .B(g29814), .Z(g31579) ) ;
INV     gate10453  (.A(g31579), .Z(g32658) ) ;
INV     gate10454  (.A(g30735), .Z(g32659) ) ;
INV     gate10455  (.A(g30825), .Z(g32660) ) ;
INV     gate10456  (.A(g31070), .Z(g32661) ) ;
INV     gate10457  (.A(g30614), .Z(g32662) ) ;
INV     gate10458  (.A(g30673), .Z(g32663) ) ;
INV     gate10459  (.A(g31528), .Z(g32664) ) ;
INV     gate10460  (.A(g31579), .Z(g32665) ) ;
INV     gate10461  (.A(g31376), .Z(g32666) ) ;
INV     gate10462  (.A(g30825), .Z(g32667) ) ;
INV     gate10463  (.A(g31070), .Z(g32668) ) ;
INV     gate10464  (.A(g30614), .Z(g32669) ) ;
INV     gate10465  (.A(g30673), .Z(g32670) ) ;
INV     gate10466  (.A(g31528), .Z(g32671) ) ;
INV     gate10467  (.A(g31579), .Z(g32672) ) ;
INV     gate10468  (.A(g31376), .Z(g32673) ) ;
INV     gate10469  (.A(g30735), .Z(g32674) ) ;
INV     gate10470  (.A(g31070), .Z(g32675) ) ;
INV     gate10471  (.A(g30614), .Z(g32676) ) ;
INV     gate10472  (.A(g30673), .Z(g32677) ) ;
INV     gate10473  (.A(g31528), .Z(g32678) ) ;
INV     gate10474  (.A(g31579), .Z(g32679) ) ;
INV     gate10475  (.A(g31376), .Z(g32680) ) ;
INV     gate10476  (.A(g30735), .Z(g32681) ) ;
INV     gate10477  (.A(g30825), .Z(g32682) ) ;
INV     gate10478  (.A(g30614), .Z(g32683) ) ;
INV     gate10479  (.A(g30673), .Z(g32684) ) ;
INV     gate10480  (.A(g31528), .Z(g32685) ) ;
INV     gate10481  (.A(g31579), .Z(g32686) ) ;
INV     gate10482  (.A(g31376), .Z(g32687) ) ;
INV     gate10483  (.A(g30735), .Z(g32688) ) ;
INV     gate10484  (.A(g30825), .Z(g32689) ) ;
INV     gate10485  (.A(g31070), .Z(g32690) ) ;
INV     gate10486  (.A(g30673), .Z(g32691) ) ;
INV     gate10487  (.A(g31528), .Z(g32692) ) ;
INV     gate10488  (.A(g31579), .Z(g32693) ) ;
INV     gate10489  (.A(g31376), .Z(g32694) ) ;
INV     gate10490  (.A(g30735), .Z(g32695) ) ;
INV     gate10491  (.A(g30825), .Z(g32696) ) ;
INV     gate10492  (.A(g31070), .Z(g32697) ) ;
INV     gate10493  (.A(g30614), .Z(g32698) ) ;
INV     gate10494  (.A(g31528), .Z(g32699) ) ;
INV     gate10495  (.A(g31579), .Z(g32700) ) ;
INV     gate10496  (.A(g31376), .Z(g32701) ) ;
INV     gate10497  (.A(g30735), .Z(g32702) ) ;
INV     gate10498  (.A(g30825), .Z(g32703) ) ;
INV     gate10499  (.A(g31070), .Z(g32704) ) ;
INV     gate10500  (.A(g30614), .Z(g32705) ) ;
INV     gate10501  (.A(g30673), .Z(g32706) ) ;
INV     gate10502  (.A(g31579), .Z(g32707) ) ;
INV     gate10503  (.A(g31376), .Z(g32708) ) ;
INV     gate10504  (.A(g30735), .Z(g32709) ) ;
INV     gate10505  (.A(g30825), .Z(g32710) ) ;
INV     gate10506  (.A(g31070), .Z(g32711) ) ;
INV     gate10507  (.A(g30614), .Z(g32712) ) ;
INV     gate10508  (.A(g30673), .Z(g32713) ) ;
INV     gate10509  (.A(g31528), .Z(g32714) ) ;
INV     gate10510  (.A(g31376), .Z(g32716) ) ;
INV     gate10511  (.A(g30735), .Z(g32717) ) ;
INV     gate10512  (.A(g30825), .Z(g32718) ) ;
AND2    gate10513  (.A(g29814), .B(g19050), .Z(g31672) ) ;
INV     gate10514  (.A(g31672), .Z(g32719) ) ;
AND2    gate10515  (.A(g29814), .B(g19128), .Z(g31710) ) ;
INV     gate10516  (.A(g31710), .Z(g32720) ) ;
AND2    gate10517  (.A(g26025), .B(g29814), .Z(g31021) ) ;
INV     gate10518  (.A(g31021), .Z(g32721) ) ;
AND2    gate10519  (.A(g22626), .B(g29814), .Z(g30937) ) ;
INV     gate10520  (.A(g30937), .Z(g32722) ) ;
AND2    gate10521  (.A(g19200), .B(g29814), .Z(g31327) ) ;
INV     gate10522  (.A(g31327), .Z(g32723) ) ;
INV     gate10523  (.A(g30735), .Z(g32724) ) ;
INV     gate10524  (.A(g30825), .Z(g32725) ) ;
INV     gate10525  (.A(g31672), .Z(g32726) ) ;
INV     gate10526  (.A(g31710), .Z(g32727) ) ;
INV     gate10527  (.A(g31021), .Z(g32728) ) ;
INV     gate10528  (.A(g30937), .Z(g32729) ) ;
INV     gate10529  (.A(g31327), .Z(g32730) ) ;
INV     gate10530  (.A(g31376), .Z(g32731) ) ;
INV     gate10531  (.A(g30825), .Z(g32732) ) ;
INV     gate10532  (.A(g31672), .Z(g32733) ) ;
INV     gate10533  (.A(g31710), .Z(g32734) ) ;
INV     gate10534  (.A(g31021), .Z(g32735) ) ;
INV     gate10535  (.A(g30937), .Z(g32736) ) ;
INV     gate10536  (.A(g31327), .Z(g32737) ) ;
INV     gate10537  (.A(g31376), .Z(g32738) ) ;
INV     gate10538  (.A(g30735), .Z(g32739) ) ;
INV     gate10539  (.A(g31672), .Z(g32740) ) ;
INV     gate10540  (.A(g31710), .Z(g32741) ) ;
INV     gate10541  (.A(g31021), .Z(g32742) ) ;
INV     gate10542  (.A(g30937), .Z(g32743) ) ;
INV     gate10543  (.A(g31327), .Z(g32744) ) ;
INV     gate10544  (.A(g31376), .Z(g32745) ) ;
INV     gate10545  (.A(g30735), .Z(g32746) ) ;
INV     gate10546  (.A(g30825), .Z(g32747) ) ;
INV     gate10547  (.A(g31710), .Z(g32748) ) ;
INV     gate10548  (.A(g31021), .Z(g32749) ) ;
INV     gate10549  (.A(g30937), .Z(g32750) ) ;
INV     gate10550  (.A(g31327), .Z(g32751) ) ;
INV     gate10551  (.A(g31376), .Z(g32752) ) ;
INV     gate10552  (.A(g30735), .Z(g32753) ) ;
INV     gate10553  (.A(g30825), .Z(g32754) ) ;
INV     gate10554  (.A(g31672), .Z(g32755) ) ;
INV     gate10555  (.A(g31021), .Z(g32756) ) ;
INV     gate10556  (.A(g30937), .Z(g32757) ) ;
INV     gate10557  (.A(g31327), .Z(g32758) ) ;
INV     gate10558  (.A(g31376), .Z(g32759) ) ;
INV     gate10559  (.A(g30735), .Z(g32760) ) ;
INV     gate10560  (.A(g30825), .Z(g32761) ) ;
INV     gate10561  (.A(g31672), .Z(g32762) ) ;
INV     gate10562  (.A(g31710), .Z(g32763) ) ;
INV     gate10563  (.A(g30937), .Z(g32764) ) ;
INV     gate10564  (.A(g31327), .Z(g32765) ) ;
INV     gate10565  (.A(g31376), .Z(g32766) ) ;
INV     gate10566  (.A(g30735), .Z(g32767) ) ;
INV     gate10567  (.A(g30825), .Z(g32768) ) ;
INV     gate10568  (.A(g31672), .Z(g32769) ) ;
INV     gate10569  (.A(g31710), .Z(g32770) ) ;
INV     gate10570  (.A(g31021), .Z(g32771) ) ;
INV     gate10571  (.A(g31327), .Z(g32772) ) ;
INV     gate10572  (.A(g31376), .Z(g32773) ) ;
INV     gate10573  (.A(g30735), .Z(g32774) ) ;
INV     gate10574  (.A(g30825), .Z(g32775) ) ;
INV     gate10575  (.A(g31672), .Z(g32776) ) ;
INV     gate10576  (.A(g31710), .Z(g32777) ) ;
INV     gate10577  (.A(g31021), .Z(g32778) ) ;
INV     gate10578  (.A(g30937), .Z(g32779) ) ;
INV     gate10579  (.A(g31376), .Z(g32781) ) ;
INV     gate10580  (.A(g30735), .Z(g32782) ) ;
INV     gate10581  (.A(g30825), .Z(g32783) ) ;
INV     gate10582  (.A(g31672), .Z(g32784) ) ;
INV     gate10583  (.A(g31710), .Z(g32785) ) ;
INV     gate10584  (.A(g31021), .Z(g32786) ) ;
INV     gate10585  (.A(g30937), .Z(g32787) ) ;
INV     gate10586  (.A(g31327), .Z(g32788) ) ;
INV     gate10587  (.A(g30735), .Z(g32789) ) ;
INV     gate10588  (.A(g30825), .Z(g32790) ) ;
INV     gate10589  (.A(g31672), .Z(g32791) ) ;
INV     gate10590  (.A(g31710), .Z(g32792) ) ;
INV     gate10591  (.A(g31021), .Z(g32793) ) ;
INV     gate10592  (.A(g30937), .Z(g32794) ) ;
INV     gate10593  (.A(g31327), .Z(g32795) ) ;
INV     gate10594  (.A(g31376), .Z(g32796) ) ;
INV     gate10595  (.A(g30825), .Z(g32797) ) ;
INV     gate10596  (.A(g31672), .Z(g32798) ) ;
INV     gate10597  (.A(g31710), .Z(g32799) ) ;
INV     gate10598  (.A(g31021), .Z(g32800) ) ;
INV     gate10599  (.A(g30937), .Z(g32801) ) ;
INV     gate10600  (.A(g31327), .Z(g32802) ) ;
INV     gate10601  (.A(g31376), .Z(g32803) ) ;
INV     gate10602  (.A(g30735), .Z(g32804) ) ;
INV     gate10603  (.A(g31672), .Z(g32805) ) ;
INV     gate10604  (.A(g31710), .Z(g32806) ) ;
INV     gate10605  (.A(g31021), .Z(g32807) ) ;
INV     gate10606  (.A(g30937), .Z(g32808) ) ;
INV     gate10607  (.A(g31327), .Z(g32809) ) ;
INV     gate10608  (.A(g31376), .Z(g32810) ) ;
INV     gate10609  (.A(g30735), .Z(g32811) ) ;
INV     gate10610  (.A(g30825), .Z(g32812) ) ;
INV     gate10611  (.A(g31710), .Z(g32813) ) ;
INV     gate10612  (.A(g31021), .Z(g32814) ) ;
INV     gate10613  (.A(g30937), .Z(g32815) ) ;
INV     gate10614  (.A(g31327), .Z(g32816) ) ;
INV     gate10615  (.A(g31376), .Z(g32817) ) ;
INV     gate10616  (.A(g30735), .Z(g32818) ) ;
INV     gate10617  (.A(g30825), .Z(g32819) ) ;
INV     gate10618  (.A(g31672), .Z(g32820) ) ;
INV     gate10619  (.A(g31021), .Z(g32821) ) ;
INV     gate10620  (.A(g30937), .Z(g32822) ) ;
INV     gate10621  (.A(g31327), .Z(g32823) ) ;
INV     gate10622  (.A(g31376), .Z(g32824) ) ;
INV     gate10623  (.A(g30735), .Z(g32825) ) ;
INV     gate10624  (.A(g30825), .Z(g32826) ) ;
INV     gate10625  (.A(g31672), .Z(g32827) ) ;
INV     gate10626  (.A(g31710), .Z(g32828) ) ;
INV     gate10627  (.A(g30937), .Z(g32829) ) ;
INV     gate10628  (.A(g31327), .Z(g32830) ) ;
INV     gate10629  (.A(g31376), .Z(g32831) ) ;
INV     gate10630  (.A(g30735), .Z(g32832) ) ;
INV     gate10631  (.A(g30825), .Z(g32833) ) ;
INV     gate10632  (.A(g31672), .Z(g32834) ) ;
INV     gate10633  (.A(g31710), .Z(g32835) ) ;
INV     gate10634  (.A(g31021), .Z(g32836) ) ;
INV     gate10635  (.A(g31327), .Z(g32837) ) ;
INV     gate10636  (.A(g31376), .Z(g32838) ) ;
INV     gate10637  (.A(g30735), .Z(g32839) ) ;
INV     gate10638  (.A(g30825), .Z(g32840) ) ;
INV     gate10639  (.A(g31672), .Z(g32841) ) ;
INV     gate10640  (.A(g31710), .Z(g32842) ) ;
INV     gate10641  (.A(g31021), .Z(g32843) ) ;
INV     gate10642  (.A(g30937), .Z(g32844) ) ;
INV     gate10643  (.A(g31376), .Z(g32846) ) ;
INV     gate10644  (.A(g30735), .Z(g32847) ) ;
INV     gate10645  (.A(g30825), .Z(g32848) ) ;
INV     gate10646  (.A(g31021), .Z(g32849) ) ;
INV     gate10647  (.A(g30937), .Z(g32850) ) ;
INV     gate10648  (.A(g31327), .Z(g32851) ) ;
INV     gate10649  (.A(g30614), .Z(g32852) ) ;
INV     gate10650  (.A(g30673), .Z(g32853) ) ;
INV     gate10651  (.A(g30735), .Z(g32854) ) ;
INV     gate10652  (.A(g30825), .Z(g32855) ) ;
INV     gate10653  (.A(g31021), .Z(g32856) ) ;
INV     gate10654  (.A(g30937), .Z(g32857) ) ;
INV     gate10655  (.A(g31327), .Z(g32858) ) ;
INV     gate10656  (.A(g30614), .Z(g32859) ) ;
INV     gate10657  (.A(g30673), .Z(g32860) ) ;
INV     gate10658  (.A(g31376), .Z(g32861) ) ;
INV     gate10659  (.A(g30825), .Z(g32862) ) ;
INV     gate10660  (.A(g31021), .Z(g32863) ) ;
INV     gate10661  (.A(g30937), .Z(g32864) ) ;
INV     gate10662  (.A(g31327), .Z(g32865) ) ;
INV     gate10663  (.A(g30614), .Z(g32866) ) ;
INV     gate10664  (.A(g30673), .Z(g32867) ) ;
INV     gate10665  (.A(g31376), .Z(g32868) ) ;
INV     gate10666  (.A(g30735), .Z(g32869) ) ;
INV     gate10667  (.A(g31021), .Z(g32870) ) ;
INV     gate10668  (.A(g30937), .Z(g32871) ) ;
INV     gate10669  (.A(g31327), .Z(g32872) ) ;
INV     gate10670  (.A(g30614), .Z(g32873) ) ;
INV     gate10671  (.A(g30673), .Z(g32874) ) ;
INV     gate10672  (.A(g31376), .Z(g32875) ) ;
INV     gate10673  (.A(g30735), .Z(g32876) ) ;
INV     gate10674  (.A(g30825), .Z(g32877) ) ;
INV     gate10675  (.A(g30937), .Z(g32878) ) ;
INV     gate10676  (.A(g31327), .Z(g32879) ) ;
INV     gate10677  (.A(g30614), .Z(g32880) ) ;
INV     gate10678  (.A(g30673), .Z(g32881) ) ;
INV     gate10679  (.A(g31376), .Z(g32882) ) ;
INV     gate10680  (.A(g30735), .Z(g32883) ) ;
INV     gate10681  (.A(g30825), .Z(g32884) ) ;
INV     gate10682  (.A(g31021), .Z(g32885) ) ;
INV     gate10683  (.A(g31327), .Z(g32886) ) ;
INV     gate10684  (.A(g30614), .Z(g32887) ) ;
INV     gate10685  (.A(g30673), .Z(g32888) ) ;
INV     gate10686  (.A(g31376), .Z(g32889) ) ;
INV     gate10687  (.A(g30735), .Z(g32890) ) ;
INV     gate10688  (.A(g30825), .Z(g32891) ) ;
INV     gate10689  (.A(g31021), .Z(g32892) ) ;
INV     gate10690  (.A(g30937), .Z(g32893) ) ;
INV     gate10691  (.A(g30614), .Z(g32894) ) ;
INV     gate10692  (.A(g30673), .Z(g32895) ) ;
INV     gate10693  (.A(g31376), .Z(g32896) ) ;
INV     gate10694  (.A(g30735), .Z(g32897) ) ;
INV     gate10695  (.A(g30825), .Z(g32898) ) ;
INV     gate10696  (.A(g31021), .Z(g32899) ) ;
INV     gate10697  (.A(g30937), .Z(g32900) ) ;
INV     gate10698  (.A(g31327), .Z(g32901) ) ;
INV     gate10699  (.A(g30673), .Z(g32902) ) ;
INV     gate10700  (.A(g31376), .Z(g32903) ) ;
INV     gate10701  (.A(g30735), .Z(g32904) ) ;
INV     gate10702  (.A(g30825), .Z(g32905) ) ;
INV     gate10703  (.A(g31021), .Z(g32906) ) ;
INV     gate10704  (.A(g30937), .Z(g32907) ) ;
INV     gate10705  (.A(g31327), .Z(g32908) ) ;
INV     gate10706  (.A(g30614), .Z(g32909) ) ;
INV     gate10707  (.A(g31376), .Z(g32911) ) ;
INV     gate10708  (.A(g30735), .Z(g32912) ) ;
INV     gate10709  (.A(g30825), .Z(g32913) ) ;
INV     gate10710  (.A(g31672), .Z(g32914) ) ;
INV     gate10711  (.A(g31710), .Z(g32915) ) ;
INV     gate10712  (.A(g31021), .Z(g32916) ) ;
INV     gate10713  (.A(g30937), .Z(g32917) ) ;
INV     gate10714  (.A(g31327), .Z(g32918) ) ;
INV     gate10715  (.A(g30735), .Z(g32919) ) ;
INV     gate10716  (.A(g30825), .Z(g32920) ) ;
INV     gate10717  (.A(g31672), .Z(g32921) ) ;
INV     gate10718  (.A(g31710), .Z(g32922) ) ;
INV     gate10719  (.A(g31021), .Z(g32923) ) ;
INV     gate10720  (.A(g30937), .Z(g32924) ) ;
INV     gate10721  (.A(g31327), .Z(g32925) ) ;
INV     gate10722  (.A(g31376), .Z(g32926) ) ;
INV     gate10723  (.A(g30825), .Z(g32927) ) ;
INV     gate10724  (.A(g31672), .Z(g32928) ) ;
INV     gate10725  (.A(g31710), .Z(g32929) ) ;
INV     gate10726  (.A(g31021), .Z(g32930) ) ;
INV     gate10727  (.A(g30937), .Z(g32931) ) ;
INV     gate10728  (.A(g31327), .Z(g32932) ) ;
INV     gate10729  (.A(g31376), .Z(g32933) ) ;
INV     gate10730  (.A(g30735), .Z(g32934) ) ;
INV     gate10731  (.A(g31672), .Z(g32935) ) ;
INV     gate10732  (.A(g31710), .Z(g32936) ) ;
INV     gate10733  (.A(g31021), .Z(g32937) ) ;
INV     gate10734  (.A(g30937), .Z(g32938) ) ;
INV     gate10735  (.A(g31327), .Z(g32939) ) ;
INV     gate10736  (.A(g31376), .Z(g32940) ) ;
INV     gate10737  (.A(g30735), .Z(g32941) ) ;
INV     gate10738  (.A(g30825), .Z(g32942) ) ;
INV     gate10739  (.A(g31710), .Z(g32943) ) ;
INV     gate10740  (.A(g31021), .Z(g32944) ) ;
INV     gate10741  (.A(g30937), .Z(g32945) ) ;
INV     gate10742  (.A(g31327), .Z(g32946) ) ;
INV     gate10743  (.A(g31376), .Z(g32947) ) ;
INV     gate10744  (.A(g30735), .Z(g32948) ) ;
INV     gate10745  (.A(g30825), .Z(g32949) ) ;
INV     gate10746  (.A(g31672), .Z(g32950) ) ;
INV     gate10747  (.A(g31021), .Z(g32951) ) ;
INV     gate10748  (.A(g30937), .Z(g32952) ) ;
INV     gate10749  (.A(g31327), .Z(g32953) ) ;
INV     gate10750  (.A(g31376), .Z(g32954) ) ;
INV     gate10751  (.A(g30735), .Z(g32955) ) ;
INV     gate10752  (.A(g30825), .Z(g32956) ) ;
INV     gate10753  (.A(g31672), .Z(g32957) ) ;
INV     gate10754  (.A(g31710), .Z(g32958) ) ;
INV     gate10755  (.A(g30937), .Z(g32959) ) ;
INV     gate10756  (.A(g31327), .Z(g32960) ) ;
INV     gate10757  (.A(g31376), .Z(g32961) ) ;
INV     gate10758  (.A(g30735), .Z(g32962) ) ;
INV     gate10759  (.A(g30825), .Z(g32963) ) ;
INV     gate10760  (.A(g31672), .Z(g32964) ) ;
INV     gate10761  (.A(g31710), .Z(g32965) ) ;
INV     gate10762  (.A(g31021), .Z(g32966) ) ;
INV     gate10763  (.A(g31327), .Z(g32967) ) ;
INV     gate10764  (.A(g31376), .Z(g32968) ) ;
INV     gate10765  (.A(g30735), .Z(g32969) ) ;
INV     gate10766  (.A(g30825), .Z(g32970) ) ;
INV     gate10767  (.A(g31672), .Z(g32971) ) ;
INV     gate10768  (.A(g31710), .Z(g32972) ) ;
INV     gate10769  (.A(g31021), .Z(g32973) ) ;
INV     gate10770  (.A(g30937), .Z(g32974) ) ;
INV     gate10771  (.A(g32027), .Z(II30537) ) ;
INV     gate10772  (.A(g31945), .Z(g33072) ) ;
INV     gate10773  (.A(g32024), .Z(II30641) ) ;
INV     gate10774  (.A(g32024), .Z(II30644) ) ;
INV     gate10775  (.A(II30644), .Z(g33080) ) ;
INV     gate10776  (.A(g32381), .Z(II30686) ) ;
INV     gate10777  (.A(II30686), .Z(g33120) ) ;
NAND2   gate10778  (.A(g7285), .B(g30573), .Z(g31950) ) ;
INV     gate10779  (.A(g31950), .Z(g33127) ) ;
NAND2   gate10780  (.A(g31003), .B(g13297), .Z(g32057) ) ;
INV     gate10781  (.A(g32057), .Z(g33136) ) ;
NAND2   gate10782  (.A(g31009), .B(g13301), .Z(g32072) ) ;
INV     gate10783  (.A(g32072), .Z(g33142) ) ;
INV     gate10784  (.A(g32363), .Z(II30766) ) ;
INV     gate10785  (.A(II30766), .Z(g33228) ) ;
NOR3    gate10786  (.A(g8859), .B(g31262), .C(g11083), .Z(g32212) ) ;
INV     gate10787  (.A(g32212), .Z(g33246) ) ;
INV     gate10788  (.A(g32186), .Z(g33250) ) ;
NOR3    gate10789  (.A(g9044), .B(g31509), .C(g12259), .Z(g32296) ) ;
INV     gate10790  (.A(g32296), .Z(g33258) ) ;
INV     gate10791  (.A(g32318), .Z(g33326) ) ;
INV     gate10792  (.A(g32383), .Z(II30861) ) ;
INV     gate10793  (.A(II30861), .Z(g33335) ) ;
OR2     gate10794  (.A(g31487), .B(g31479), .Z(g32132) ) ;
INV     gate10795  (.A(g32132), .Z(g33346) ) ;
INV     gate10796  (.A(g32329), .Z(g33354) ) ;
INV     gate10797  (.A(g32377), .Z(g33375) ) ;
INV     gate10798  (.A(g32407), .Z(II30901) ) ;
INV     gate10799  (.A(II30901), .Z(g33377) ) ;
NOR2    gate10800  (.A(g8721), .B(g31294), .Z(g32424) ) ;
INV     gate10801  (.A(g32424), .Z(II30904) ) ;
INV     gate10802  (.A(II30904), .Z(g33378) ) ;
INV     gate10803  (.A(g32033), .Z(g33382) ) ;
INV     gate10804  (.A(g32038), .Z(g33385) ) ;
INV     gate10805  (.A(g32382), .Z(g33388) ) ;
INV     gate10806  (.A(g32384), .Z(g33391) ) ;
NAND2   gate10807  (.A(g30573), .B(g10511), .Z(g31971) ) ;
INV     gate10808  (.A(g31971), .Z(g33413) ) ;
INV     gate10809  (.A(g32415), .Z(g33424) ) ;
NOR2    gate10810  (.A(g31504), .B(g23475), .Z(g32017) ) ;
INV     gate10811  (.A(g32017), .Z(g33426) ) ;
INV     gate10812  (.A(g32421), .Z(g33430) ) ;
INV     gate10813  (.A(g32021), .Z(II30959) ) ;
INV     gate10814  (.A(g32021), .Z(II30962) ) ;
INV     gate10815  (.A(II30962), .Z(g33436) ) ;
INV     gate10816  (.A(g31937), .Z(g33442) ) ;
INV     gate10817  (.A(g32015), .Z(II30971) ) ;
INV     gate10818  (.A(II30971), .Z(g33443) ) ;
INV     gate10819  (.A(g32132), .Z(g33451) ) ;
INV     gate10820  (.A(g32132), .Z(II30980) ) ;
INV     gate10821  (.A(II30980), .Z(g33454) ) ;
INV     gate10822  (.A(g32433), .Z(II30983) ) ;
INV     gate10823  (.A(II30983), .Z(g33455) ) ;
INV     gate10824  (.A(g32437), .Z(II30986) ) ;
INV     gate10825  (.A(II30986), .Z(g33456) ) ;
INV     gate10826  (.A(g32441), .Z(II30989) ) ;
INV     gate10827  (.A(II30989), .Z(g33457) ) ;
INV     gate10828  (.A(g32445), .Z(II30992) ) ;
INV     gate10829  (.A(II30992), .Z(g33458) ) ;
INV     gate10830  (.A(g32449), .Z(II30995) ) ;
INV     gate10831  (.A(II30995), .Z(g33459) ) ;
INV     gate10832  (.A(g32453), .Z(II30998) ) ;
INV     gate10833  (.A(II30998), .Z(g33460) ) ;
INV     gate10834  (.A(g33120), .Z(II31361) ) ;
OR3     gate10835  (.A(g32335), .B(II30760), .C(II30761), .Z(g33219) ) ;
INV     gate10836  (.A(g33219), .Z(II31459) ) ;
INV     gate10837  (.A(II31459), .Z(g33631) ) ;
INV     gate10838  (.A(g33436), .Z(g33635) ) ;
OR2     gate10839  (.A(g31969), .B(g32434), .Z(g33318) ) ;
INV     gate10840  (.A(g33318), .Z(II31463) ) ;
INV     gate10841  (.A(g33318), .Z(II31466) ) ;
INV     gate10842  (.A(II31466), .Z(g33637) ) ;
INV     gate10843  (.A(g33388), .Z(II31469) ) ;
INV     gate10844  (.A(II31469), .Z(g33638) ) ;
OR3     gate10845  (.A(g32328), .B(II30755), .C(II30756), .Z(g33212) ) ;
INV     gate10846  (.A(g33212), .Z(II31474) ) ;
INV     gate10847  (.A(II31474), .Z(g33641) ) ;
INV     gate10848  (.A(g33391), .Z(II31477) ) ;
INV     gate10849  (.A(II31477), .Z(g33645) ) ;
OR3     gate10850  (.A(g32317), .B(II30750), .C(II30751), .Z(g33204) ) ;
INV     gate10851  (.A(g33204), .Z(II31482) ) ;
INV     gate10852  (.A(II31482), .Z(g33648) ) ;
OR3     gate10853  (.A(g32342), .B(II30745), .C(II30746), .Z(g33197) ) ;
INV     gate10854  (.A(g33197), .Z(II31486) ) ;
INV     gate10855  (.A(II31486), .Z(g33653) ) ;
INV     gate10856  (.A(g33080), .Z(g33658) ) ;
OR2     gate10857  (.A(g31995), .B(g30318), .Z(g33283) ) ;
INV     gate10858  (.A(g33283), .Z(II31491) ) ;
INV     gate10859  (.A(g33283), .Z(II31494) ) ;
INV     gate10860  (.A(II31494), .Z(g33660) ) ;
OR3     gate10861  (.A(g32014), .B(II30740), .C(II30741), .Z(g33187) ) ;
INV     gate10862  (.A(g33187), .Z(II31497) ) ;
INV     gate10863  (.A(II31497), .Z(g33661) ) ;
OR3     gate10864  (.A(g32198), .B(II30734), .C(II30735), .Z(g33176) ) ;
INV     gate10865  (.A(g33176), .Z(II31500) ) ;
INV     gate10866  (.A(II31500), .Z(g33665) ) ;
OR3     gate10867  (.A(g32203), .B(II30727), .C(II30728), .Z(g33164) ) ;
INV     gate10868  (.A(g33164), .Z(II31504) ) ;
INV     gate10869  (.A(II31504), .Z(g33670) ) ;
INV     gate10870  (.A(g33187), .Z(II31515) ) ;
INV     gate10871  (.A(II31515), .Z(g33682) ) ;
INV     gate10872  (.A(g33187), .Z(g33686) ) ;
INV     gate10873  (.A(g33187), .Z(II31523) ) ;
INV     gate10874  (.A(II31523), .Z(g33688) ) ;
INV     gate10875  (.A(g33219), .Z(II31528) ) ;
INV     gate10876  (.A(II31528), .Z(g33691) ) ;
INV     gate10877  (.A(g33187), .Z(g33695) ) ;
INV     gate10878  (.A(g33377), .Z(II31535) ) ;
INV     gate10879  (.A(II31535), .Z(g33696) ) ;
INV     gate10880  (.A(g33212), .Z(II31539) ) ;
INV     gate10881  (.A(II31539), .Z(g33698) ) ;
INV     gate10882  (.A(g33219), .Z(II31545) ) ;
INV     gate10883  (.A(II31545), .Z(g33702) ) ;
INV     gate10884  (.A(g33204), .Z(II31550) ) ;
INV     gate10885  (.A(II31550), .Z(g33705) ) ;
INV     gate10886  (.A(g33212), .Z(II31555) ) ;
INV     gate10887  (.A(II31555), .Z(g33708) ) ;
INV     gate10888  (.A(g33197), .Z(II31561) ) ;
INV     gate10889  (.A(II31561), .Z(g33712) ) ;
INV     gate10890  (.A(g33204), .Z(II31564) ) ;
INV     gate10891  (.A(II31564), .Z(g33713) ) ;
INV     gate10892  (.A(g33197), .Z(II31569) ) ;
INV     gate10893  (.A(II31569), .Z(g33716) ) ;
INV     gate10894  (.A(g33164), .Z(II31581) ) ;
INV     gate10895  (.A(II31581), .Z(g33726) ) ;
OR3     gate10896  (.A(g32204), .B(II30717), .C(II30718), .Z(g33149) ) ;
INV     gate10897  (.A(g33149), .Z(II31586) ) ;
INV     gate10898  (.A(II31586), .Z(g33729) ) ;
INV     gate10899  (.A(g33187), .Z(II31597) ) ;
INV     gate10900  (.A(II31597), .Z(g33736) ) ;
INV     gate10901  (.A(g33176), .Z(II31604) ) ;
INV     gate10902  (.A(II31604), .Z(g33744) ) ;
INV     gate10903  (.A(g33164), .Z(II31607) ) ;
INV     gate10904  (.A(II31607), .Z(g33750) ) ;
INV     gate10905  (.A(g33149), .Z(II31610) ) ;
INV     gate10906  (.A(II31610), .Z(g33755) ) ;
INV     gate10907  (.A(g33219), .Z(II31616) ) ;
INV     gate10908  (.A(II31616), .Z(g33761) ) ;
INV     gate10909  (.A(g33212), .Z(II31619) ) ;
INV     gate10910  (.A(II31619), .Z(g33766) ) ;
INV     gate10911  (.A(g33204), .Z(II31622) ) ;
INV     gate10912  (.A(II31622), .Z(g33772) ) ;
INV     gate10913  (.A(g33197), .Z(II31625) ) ;
INV     gate10914  (.A(II31625), .Z(g33778) ) ;
NAND3   gate10915  (.A(g776), .B(g32212), .C(g11679), .Z(g33306) ) ;
INV     gate10916  (.A(g33306), .Z(g33797) ) ;
NAND3   gate10917  (.A(g608), .B(g32296), .C(g12323), .Z(g33299) ) ;
INV     gate10918  (.A(g33299), .Z(g33799) ) ;
INV     gate10919  (.A(g33204), .Z(II31642) ) ;
INV     gate10920  (.A(II31642), .Z(g33800) ) ;
INV     gate10921  (.A(g33250), .Z(g33804) ) ;
INV     gate10922  (.A(g33212), .Z(II31650) ) ;
INV     gate10923  (.A(II31650), .Z(g33806) ) ;
INV     gate10924  (.A(g33219), .Z(II31659) ) ;
INV     gate10925  (.A(II31659), .Z(g33813) ) ;
INV     gate10926  (.A(g33149), .Z(II31672) ) ;
INV     gate10927  (.A(II31672), .Z(g33827) ) ;
INV     gate10928  (.A(g33164), .Z(II31686) ) ;
INV     gate10929  (.A(II31686), .Z(g33839) ) ;
INV     gate10930  (.A(g33176), .Z(II31694) ) ;
INV     gate10931  (.A(II31694), .Z(g33845) ) ;
INV     gate10932  (.A(g33164), .Z(II31701) ) ;
INV     gate10933  (.A(II31701), .Z(g33850) ) ;
OR2     gate10934  (.A(g32336), .B(g32446), .Z(g33076) ) ;
INV     gate10935  (.A(g33076), .Z(II31724) ) ;
INV     gate10936  (.A(g33076), .Z(II31727) ) ;
INV     gate10937  (.A(II31727), .Z(g33875) ) ;
INV     gate10938  (.A(g33346), .Z(g33888) ) ;
INV     gate10939  (.A(g33228), .Z(II31748) ) ;
INV     gate10940  (.A(g33228), .Z(II31751) ) ;
INV     gate10941  (.A(II31751), .Z(g33895) ) ;
INV     gate10942  (.A(g33197), .Z(II31770) ) ;
INV     gate10943  (.A(II31770), .Z(g33912) ) ;
INV     gate10944  (.A(g33204), .Z(II31776) ) ;
INV     gate10945  (.A(II31776), .Z(g33916) ) ;
INV     gate10946  (.A(g33212), .Z(II31779) ) ;
INV     gate10947  (.A(II31779), .Z(g33917) ) ;
INV     gate10948  (.A(g33219), .Z(II31782) ) ;
INV     gate10949  (.A(II31782), .Z(g33918) ) ;
INV     gate10950  (.A(g33197), .Z(II31786) ) ;
INV     gate10951  (.A(II31786), .Z(g33920) ) ;
INV     gate10952  (.A(g33354), .Z(II31791) ) ;
INV     gate10953  (.A(II31791), .Z(g33923) ) ;
INV     gate10954  (.A(g33176), .Z(II31796) ) ;
INV     gate10955  (.A(II31796), .Z(g33926) ) ;
INV     gate10956  (.A(g33164), .Z(II31800) ) ;
INV     gate10957  (.A(II31800), .Z(g33928) ) ;
INV     gate10958  (.A(g33176), .Z(II31803) ) ;
INV     gate10959  (.A(II31803), .Z(g33929) ) ;
INV     gate10960  (.A(g33149), .Z(II31807) ) ;
INV     gate10961  (.A(II31807), .Z(g33931) ) ;
INV     gate10962  (.A(g33164), .Z(II31810) ) ;
INV     gate10963  (.A(II31810), .Z(g33932) ) ;
INV     gate10964  (.A(g33149), .Z(II31814) ) ;
INV     gate10965  (.A(II31814), .Z(g33934) ) ;
OR2     gate10966  (.A(g31936), .B(g32442), .Z(g33323) ) ;
INV     gate10967  (.A(g33323), .Z(II31817) ) ;
INV     gate10968  (.A(g33323), .Z(II31820) ) ;
INV     gate10969  (.A(II31820), .Z(g33936) ) ;
INV     gate10970  (.A(g33149), .Z(II31823) ) ;
INV     gate10971  (.A(II31823), .Z(g33937) ) ;
INV     gate10972  (.A(g33454), .Z(II31829) ) ;
INV     gate10973  (.A(II31829), .Z(g33944) ) ;
INV     gate10974  (.A(g33696), .Z(II31878) ) ;
AND3    gate10975  (.A(g33164), .B(g10710), .C(g22319), .Z(g33674) ) ;
INV     gate10976  (.A(g33674), .Z(g34042) ) ;
AND3    gate10977  (.A(g33164), .B(g10727), .C(g22332), .Z(g33675) ) ;
INV     gate10978  (.A(g33675), .Z(g34044) ) ;
INV     gate10979  (.A(g33637), .Z(g34047) ) ;
AND3    gate10980  (.A(g33149), .B(g10710), .C(g22319), .Z(g33678) ) ;
INV     gate10981  (.A(g33678), .Z(g34049) ) ;
INV     gate10982  (.A(g33635), .Z(g34052) ) ;
AND3    gate10983  (.A(g33149), .B(g10727), .C(g22332), .Z(g33683) ) ;
INV     gate10984  (.A(g33683), .Z(g34053) ) ;
INV     gate10985  (.A(g33660), .Z(g34058) ) ;
INV     gate10986  (.A(g33658), .Z(g34059) ) ;
AND3    gate10987  (.A(g33176), .B(g10710), .C(g22319), .Z(g33704) ) ;
INV     gate10988  (.A(g33704), .Z(g34060) ) ;
AND3    gate10989  (.A(g33176), .B(g10727), .C(g22332), .Z(g33711) ) ;
INV     gate10990  (.A(g33711), .Z(g34062) ) ;
AND3    gate10991  (.A(g22626), .B(g10851), .C(g33187), .Z(g33728) ) ;
INV     gate10992  (.A(g33728), .Z(g34068) ) ;
AND3    gate10993  (.A(g22626), .B(g10851), .C(g33176), .Z(g33725) ) ;
INV     gate10994  (.A(g33725), .Z(g34070) ) ;
INV     gate10995  (.A(g33772), .Z(g34094) ) ;
INV     gate10996  (.A(g33631), .Z(II32051) ) ;
INV     gate10997  (.A(II32051), .Z(g34118) ) ;
INV     gate10998  (.A(g33641), .Z(II32056) ) ;
INV     gate10999  (.A(II32056), .Z(g34121) ) ;
INV     gate11000  (.A(g33648), .Z(II32059) ) ;
INV     gate11001  (.A(II32059), .Z(g34122) ) ;
INV     gate11002  (.A(g33653), .Z(II32062) ) ;
INV     gate11003  (.A(II32062), .Z(g34123) ) ;
AND3    gate11004  (.A(g23088), .B(g33176), .C(g9104), .Z(g33819) ) ;
INV     gate11005  (.A(g33819), .Z(g34124) ) ;
INV     gate11006  (.A(g33661), .Z(II32067) ) ;
INV     gate11007  (.A(II32067), .Z(g34126) ) ;
INV     gate11008  (.A(g33665), .Z(II32071) ) ;
INV     gate11009  (.A(II32071), .Z(g34130) ) ;
INV     gate11010  (.A(g33670), .Z(II32074) ) ;
INV     gate11011  (.A(II32074), .Z(g34131) ) ;
AND3    gate11012  (.A(g23088), .B(g33149), .C(g9104), .Z(g33831) ) ;
INV     gate11013  (.A(g33831), .Z(g34132) ) ;
INV     gate11014  (.A(g33937), .Z(II32079) ) ;
INV     gate11015  (.A(II32079), .Z(g34134) ) ;
INV     gate11016  (.A(g33665), .Z(II32089) ) ;
INV     gate11017  (.A(II32089), .Z(g34142) ) ;
INV     gate11018  (.A(g33670), .Z(II32093) ) ;
INV     gate11019  (.A(II32093), .Z(g34144) ) ;
INV     gate11020  (.A(g33641), .Z(II32096) ) ;
INV     gate11021  (.A(II32096), .Z(g34145) ) ;
NOR3    gate11022  (.A(g8774), .B(g33306), .C(g11083), .Z(g33823) ) ;
INV     gate11023  (.A(g33823), .Z(g34147) ) ;
INV     gate11024  (.A(g33661), .Z(II32103) ) ;
INV     gate11025  (.A(II32103), .Z(g34150) ) ;
INV     gate11026  (.A(g33653), .Z(II32106) ) ;
INV     gate11027  (.A(II32106), .Z(g34151) ) ;
INV     gate11028  (.A(g33631), .Z(II32109) ) ;
INV     gate11029  (.A(II32109), .Z(g34152) ) ;
AND3    gate11030  (.A(g23088), .B(g33219), .C(g9104), .Z(g33907) ) ;
INV     gate11031  (.A(g33907), .Z(g34156) ) ;
INV     gate11032  (.A(g33937), .Z(II32116) ) ;
INV     gate11033  (.A(II32116), .Z(g34159) ) ;
INV     gate11034  (.A(g33648), .Z(II32119) ) ;
INV     gate11035  (.A(II32119), .Z(g34160) ) ;
NOR3    gate11036  (.A(g8854), .B(g33299), .C(g12259), .Z(g33851) ) ;
INV     gate11037  (.A(g33851), .Z(g34161) ) ;
AND3    gate11038  (.A(g23088), .B(g33204), .C(g9104), .Z(g33913) ) ;
INV     gate11039  (.A(g33913), .Z(g34181) ) ;
INV     gate11040  (.A(g33875), .Z(g34188) ) ;
AND3    gate11041  (.A(g33187), .B(g9104), .C(g19200), .Z(g33921) ) ;
INV     gate11042  (.A(g33921), .Z(g34192) ) ;
INV     gate11043  (.A(g33923), .Z(II32150) ) ;
INV     gate11044  (.A(II32150), .Z(g34195) ) ;
AND3    gate11045  (.A(g23088), .B(g33187), .C(g9104), .Z(g33812) ) ;
INV     gate11046  (.A(g33812), .Z(g34197) ) ;
INV     gate11047  (.A(g33895), .Z(g34200) ) ;
OR2     gate11048  (.A(g33379), .B(g32430), .Z(g33791) ) ;
INV     gate11049  (.A(g33791), .Z(II32158) ) ;
INV     gate11050  (.A(g33791), .Z(II32161) ) ;
INV     gate11051  (.A(II32161), .Z(g34202) ) ;
NAND2   gate11052  (.A(g33083), .B(g4369), .Z(g33838) ) ;
INV     gate11053  (.A(g33838), .Z(g34208) ) ;
INV     gate11054  (.A(g33638), .Z(II32170) ) ;
INV     gate11055  (.A(II32170), .Z(g34209) ) ;
INV     gate11056  (.A(g33645), .Z(II32173) ) ;
INV     gate11057  (.A(II32173), .Z(g34210) ) ;
OR2     gate11058  (.A(g33071), .B(g32450), .Z(g33628) ) ;
INV     gate11059  (.A(g33628), .Z(II32192) ) ;
INV     gate11060  (.A(g33628), .Z(II32195) ) ;
INV     gate11061  (.A(II32195), .Z(g34222) ) ;
INV     gate11062  (.A(g33936), .Z(g34229) ) ;
INV     gate11063  (.A(g34118), .Z(II32222) ) ;
INV     gate11064  (.A(II32222), .Z(g34241) ) ;
INV     gate11065  (.A(g34121), .Z(II32225) ) ;
INV     gate11066  (.A(II32225), .Z(g34242) ) ;
INV     gate11067  (.A(g34122), .Z(II32228) ) ;
INV     gate11068  (.A(II32228), .Z(g34243) ) ;
INV     gate11069  (.A(g34123), .Z(II32231) ) ;
INV     gate11070  (.A(II32231), .Z(g34244) ) ;
INV     gate11071  (.A(g34126), .Z(II32234) ) ;
INV     gate11072  (.A(II32234), .Z(g34245) ) ;
INV     gate11073  (.A(g34130), .Z(II32237) ) ;
INV     gate11074  (.A(II32237), .Z(g34246) ) ;
INV     gate11075  (.A(g34131), .Z(II32240) ) ;
INV     gate11076  (.A(II32240), .Z(g34247) ) ;
INV     gate11077  (.A(g34134), .Z(II32243) ) ;
INV     gate11078  (.A(II32243), .Z(g34248) ) ;
INV     gate11079  (.A(g34159), .Z(g34270) ) ;
INV     gate11080  (.A(g34160), .Z(g34271) ) ;
INV     gate11081  (.A(g34229), .Z(g34272) ) ;
INV     gate11082  (.A(g34047), .Z(g34275) ) ;
INV     gate11083  (.A(g34058), .Z(g34276) ) ;
INV     gate11084  (.A(g34195), .Z(II32274) ) ;
INV     gate11085  (.A(II32274), .Z(g34277) ) ;
INV     gate11086  (.A(g34052), .Z(II32284) ) ;
INV     gate11087  (.A(II32284), .Z(g34285) ) ;
INV     gate11088  (.A(g34059), .Z(II32297) ) ;
INV     gate11089  (.A(II32297), .Z(g34296) ) ;
AND3    gate11090  (.A(g22957), .B(g9104), .C(g33750), .Z(g34080) ) ;
INV     gate11091  (.A(g34080), .Z(g34299) ) ;
INV     gate11092  (.A(g34209), .Z(II32305) ) ;
INV     gate11093  (.A(II32305), .Z(g34302) ) ;
INV     gate11094  (.A(g34210), .Z(II32309) ) ;
INV     gate11095  (.A(II32309), .Z(g34304) ) ;
AND3    gate11096  (.A(g33766), .B(g9104), .C(g18957), .Z(g34087) ) ;
INV     gate11097  (.A(g34087), .Z(g34307) ) ;
AND3    gate11098  (.A(g33736), .B(g9104), .C(g18957), .Z(g34088) ) ;
INV     gate11099  (.A(g34088), .Z(g34308) ) ;
AND3    gate11100  (.A(g33772), .B(g9104), .C(g18957), .Z(g34097) ) ;
INV     gate11101  (.A(g34097), .Z(g34311) ) ;
AND3    gate11102  (.A(g33744), .B(g9104), .C(g18957), .Z(g34098) ) ;
INV     gate11103  (.A(g34098), .Z(g34312) ) ;
AND3    gate11104  (.A(g20114), .B(g33766), .C(g9104), .Z(g34086) ) ;
INV     gate11105  (.A(g34086), .Z(g34313) ) ;
AND3    gate11106  (.A(g33761), .B(g9104), .C(g18957), .Z(g34085) ) ;
INV     gate11107  (.A(g34085), .Z(g34315) ) ;
AND3    gate11108  (.A(g20114), .B(g33755), .C(g9104), .Z(g34093) ) ;
INV     gate11109  (.A(g34093), .Z(g34316) ) ;
AND3    gate11110  (.A(g20516), .B(g9104), .C(g33750), .Z(g34115) ) ;
INV     gate11111  (.A(g34115), .Z(g34317) ) ;
AND3    gate11112  (.A(g20516), .B(g9104), .C(g33755), .Z(g34119) ) ;
INV     gate11113  (.A(g34119), .Z(g34320) ) ;
AND3    gate11114  (.A(g33778), .B(g9104), .C(g18957), .Z(g34105) ) ;
INV     gate11115  (.A(g34105), .Z(g34323) ) ;
AND3    gate11116  (.A(g33750), .B(g9104), .C(g18957), .Z(g34092) ) ;
INV     gate11117  (.A(g34092), .Z(g34325) ) ;
AND3    gate11118  (.A(g22957), .B(g9104), .C(g33761), .Z(g34091) ) ;
INV     gate11119  (.A(g34091), .Z(g34326) ) ;
AND3    gate11120  (.A(g22957), .B(g9104), .C(g33766), .Z(g34108) ) ;
INV     gate11121  (.A(g34108), .Z(g34327) ) ;
AND3    gate11122  (.A(g22957), .B(g9104), .C(g33772), .Z(g34096) ) ;
INV     gate11123  (.A(g34096), .Z(g34328) ) ;
AND3    gate11124  (.A(g22957), .B(g9104), .C(g33778), .Z(g34112) ) ;
INV     gate11125  (.A(g34112), .Z(g34336) ) ;
AND3    gate11126  (.A(g22957), .B(g9104), .C(g33736), .Z(g34077) ) ;
INV     gate11127  (.A(g34077), .Z(g34339) ) ;
AND3    gate11128  (.A(g22957), .B(g9104), .C(g33744), .Z(g34089) ) ;
INV     gate11129  (.A(g34089), .Z(g34343) ) ;
AND2    gate11130  (.A(g33804), .B(g31227), .Z(g34169) ) ;
INV     gate11131  (.A(g34169), .Z(II32352) ) ;
INV     gate11132  (.A(II32352), .Z(g34345) ) ;
NAND3   gate11133  (.A(g785), .B(g33823), .C(g11679), .Z(g34162) ) ;
INV     gate11134  (.A(g34162), .Z(g34346) ) ;
NAND3   gate11135  (.A(g617), .B(g33851), .C(g12323), .Z(g34174) ) ;
INV     gate11136  (.A(g34174), .Z(g34351) ) ;
INV     gate11137  (.A(g34208), .Z(II32364) ) ;
INV     gate11138  (.A(II32364), .Z(g34358) ) ;
OR2     gate11139  (.A(g33899), .B(g33451), .Z(g34153) ) ;
INV     gate11140  (.A(g34153), .Z(II32388) ) ;
INV     gate11141  (.A(g34153), .Z(II32391) ) ;
INV     gate11142  (.A(II32391), .Z(g34384) ) ;
INV     gate11143  (.A(g34188), .Z(g34387) ) ;
INV     gate11144  (.A(g34200), .Z(g34391) ) ;
INV     gate11145  (.A(g34202), .Z(g34392) ) ;
INV     gate11146  (.A(g34142), .Z(g34400) ) ;
INV     gate11147  (.A(g34144), .Z(g34408) ) ;
INV     gate11148  (.A(g34145), .Z(g34409) ) ;
INV     gate11149  (.A(g34150), .Z(g34418) ) ;
INV     gate11150  (.A(g34151), .Z(g34419) ) ;
INV     gate11151  (.A(g34152), .Z(g34420) ) ;
INV     gate11152  (.A(g34222), .Z(g34423) ) ;
OR2     gate11153  (.A(g33657), .B(g32438), .Z(g34127) ) ;
INV     gate11154  (.A(g34127), .Z(II32446) ) ;
INV     gate11155  (.A(g34127), .Z(II32449) ) ;
INV     gate11156  (.A(II32449), .Z(g34426) ) ;
INV     gate11157  (.A(g34241), .Z(II32452) ) ;
INV     gate11158  (.A(II32452), .Z(g34427) ) ;
INV     gate11159  (.A(g34242), .Z(II32455) ) ;
INV     gate11160  (.A(II32455), .Z(g34428) ) ;
INV     gate11161  (.A(g34243), .Z(II32458) ) ;
INV     gate11162  (.A(II32458), .Z(g34429) ) ;
INV     gate11163  (.A(g34244), .Z(II32461) ) ;
INV     gate11164  (.A(II32461), .Z(g34430) ) ;
INV     gate11165  (.A(g34245), .Z(II32464) ) ;
INV     gate11166  (.A(II32464), .Z(g34431) ) ;
INV     gate11167  (.A(g34246), .Z(II32467) ) ;
INV     gate11168  (.A(II32467), .Z(g34432) ) ;
INV     gate11169  (.A(g34247), .Z(II32470) ) ;
INV     gate11170  (.A(II32470), .Z(g34433) ) ;
INV     gate11171  (.A(g34248), .Z(II32473) ) ;
INV     gate11172  (.A(II32473), .Z(g34434) ) ;
INV     gate11173  (.A(g34277), .Z(II32476) ) ;
INV     gate11174  (.A(g34302), .Z(II32479) ) ;
INV     gate11175  (.A(g34304), .Z(II32482) ) ;
INV     gate11176  (.A(g34423), .Z(g34471) ) ;
INV     gate11177  (.A(g34285), .Z(II32525) ) ;
INV     gate11178  (.A(II32525), .Z(g34472) ) ;
INV     gate11179  (.A(g34426), .Z(g34473) ) ;
INV     gate11180  (.A(g34296), .Z(II32535) ) ;
INV     gate11181  (.A(II32535), .Z(g34480) ) ;
AND2    gate11182  (.A(g7673), .B(g34068), .Z(g34397) ) ;
INV     gate11183  (.A(g34397), .Z(II32547) ) ;
INV     gate11184  (.A(II32547), .Z(g34490) ) ;
AND2    gate11185  (.A(g7684), .B(g34070), .Z(g34398) ) ;
INV     gate11186  (.A(g34398), .Z(II32550) ) ;
INV     gate11187  (.A(II32550), .Z(g34491) ) ;
INV     gate11188  (.A(g34400), .Z(g34501) ) ;
INV     gate11189  (.A(g34408), .Z(g34504) ) ;
INV     gate11190  (.A(g34409), .Z(g34505) ) ;
INV     gate11191  (.A(g34418), .Z(g34510) ) ;
INV     gate11192  (.A(g34419), .Z(g34511) ) ;
INV     gate11193  (.A(g34420), .Z(g34512) ) ;
INV     gate11194  (.A(g34270), .Z(g34521) ) ;
INV     gate11195  (.A(g34271), .Z(g34522) ) ;
AND2    gate11196  (.A(g11370), .B(g34124), .Z(g34287) ) ;
INV     gate11197  (.A(g34287), .Z(II32591) ) ;
INV     gate11198  (.A(II32591), .Z(g34530) ) ;
AND2    gate11199  (.A(g8679), .B(g34132), .Z(g34298) ) ;
INV     gate11200  (.A(g34298), .Z(II32594) ) ;
INV     gate11201  (.A(II32594), .Z(g34531) ) ;
AND2    gate11202  (.A(g9535), .B(g34156), .Z(g34319) ) ;
INV     gate11203  (.A(g34319), .Z(II32601) ) ;
INV     gate11204  (.A(II32601), .Z(g34536) ) ;
NOR3    gate11205  (.A(g9003), .B(g34162), .C(g11083), .Z(g34354) ) ;
INV     gate11206  (.A(g34354), .Z(g34539) ) ;
INV     gate11207  (.A(g34358), .Z(II32607) ) ;
INV     gate11208  (.A(II32607), .Z(g34540) ) ;
NOR3    gate11209  (.A(g9162), .B(g34174), .C(g12259), .Z(g34359) ) ;
INV     gate11210  (.A(g34359), .Z(g34543) ) ;
AND2    gate11211  (.A(g14511), .B(g34181), .Z(g34329) ) ;
INV     gate11212  (.A(g34329), .Z(II32613) ) ;
INV     gate11213  (.A(II32613), .Z(g34544) ) ;
AND2    gate11214  (.A(g9984), .B(g34192), .Z(g34333) ) ;
INV     gate11215  (.A(g34333), .Z(II32617) ) ;
INV     gate11216  (.A(II32617), .Z(g34549) ) ;
AND2    gate11217  (.A(g8461), .B(g34197), .Z(g34335) ) ;
INV     gate11218  (.A(g34335), .Z(II32621) ) ;
INV     gate11219  (.A(II32621), .Z(g34553) ) ;
INV     gate11220  (.A(g34384), .Z(g34559) ) ;
INV     gate11221  (.A(g34345), .Z(II32639) ) ;
INV     gate11222  (.A(II32639), .Z(g34569) ) ;
INV     gate11223  (.A(g34392), .Z(g34570) ) ;
AND2    gate11224  (.A(g7404), .B(g34042), .Z(g34367) ) ;
INV     gate11225  (.A(g34367), .Z(II32645) ) ;
INV     gate11226  (.A(II32645), .Z(g34573) ) ;
AND2    gate11227  (.A(g7450), .B(g34044), .Z(g34371) ) ;
INV     gate11228  (.A(g34371), .Z(II32648) ) ;
INV     gate11229  (.A(II32648), .Z(g34574) ) ;
AND2    gate11230  (.A(g13077), .B(g34049), .Z(g34375) ) ;
INV     gate11231  (.A(g34375), .Z(II32651) ) ;
INV     gate11232  (.A(II32651), .Z(g34575) ) ;
AND2    gate11233  (.A(g13095), .B(g34053), .Z(g34378) ) ;
INV     gate11234  (.A(g34378), .Z(II32654) ) ;
INV     gate11235  (.A(II32654), .Z(g34576) ) ;
INV     gate11236  (.A(g34391), .Z(II32659) ) ;
INV     gate11237  (.A(II32659), .Z(g34579) ) ;
AND2    gate11238  (.A(g10800), .B(g34060), .Z(g34386) ) ;
INV     gate11239  (.A(g34386), .Z(II32665) ) ;
INV     gate11240  (.A(II32665), .Z(g34583) ) ;
AND2    gate11241  (.A(g10802), .B(g34062), .Z(g34388) ) ;
INV     gate11242  (.A(g34388), .Z(II32671) ) ;
INV     gate11243  (.A(II32671), .Z(g34587) ) ;
INV     gate11244  (.A(g34427), .Z(II32675) ) ;
INV     gate11245  (.A(g34428), .Z(II32678) ) ;
INV     gate11246  (.A(g34429), .Z(II32681) ) ;
INV     gate11247  (.A(g34430), .Z(II32684) ) ;
INV     gate11248  (.A(g34431), .Z(II32687) ) ;
INV     gate11249  (.A(g34432), .Z(II32690) ) ;
INV     gate11250  (.A(g34433), .Z(II32693) ) ;
INV     gate11251  (.A(g34434), .Z(II32696) ) ;
INV     gate11252  (.A(g34569), .Z(II32699) ) ;
INV     gate11253  (.A(g34510), .Z(II32752) ) ;
INV     gate11254  (.A(II32752), .Z(g34648) ) ;
INV     gate11255  (.A(g34511), .Z(II32763) ) ;
INV     gate11256  (.A(II32763), .Z(g34653) ) ;
INV     gate11257  (.A(g34522), .Z(II32766) ) ;
INV     gate11258  (.A(II32766), .Z(g34654) ) ;
INV     gate11259  (.A(g34505), .Z(II32770) ) ;
INV     gate11260  (.A(II32770), .Z(g34656) ) ;
INV     gate11261  (.A(g34512), .Z(II32775) ) ;
INV     gate11262  (.A(II32775), .Z(g34659) ) ;
INV     gate11263  (.A(g34473), .Z(g34660) ) ;
AND2    gate11264  (.A(g27225), .B(g34299), .Z(g34571) ) ;
INV     gate11265  (.A(g34571), .Z(II32782) ) ;
INV     gate11266  (.A(II32782), .Z(g34664) ) ;
AND2    gate11267  (.A(g24577), .B(g34307), .Z(g34577) ) ;
INV     gate11268  (.A(g34577), .Z(II32788) ) ;
INV     gate11269  (.A(II32788), .Z(g34668) ) ;
AND2    gate11270  (.A(g24578), .B(g34308), .Z(g34578) ) ;
INV     gate11271  (.A(g34578), .Z(II32791) ) ;
INV     gate11272  (.A(II32791), .Z(g34669) ) ;
AND2    gate11273  (.A(g29539), .B(g34311), .Z(g34580) ) ;
INV     gate11274  (.A(g34580), .Z(II32794) ) ;
INV     gate11275  (.A(II32794), .Z(g34670) ) ;
AND2    gate11276  (.A(g22864), .B(g34312), .Z(g34581) ) ;
INV     gate11277  (.A(g34581), .Z(II32797) ) ;
INV     gate11278  (.A(II32797), .Z(g34671) ) ;
AND2    gate11279  (.A(g7764), .B(g34313), .Z(g34582) ) ;
INV     gate11280  (.A(g34582), .Z(II32800) ) ;
INV     gate11281  (.A(II32800), .Z(g34672) ) ;
AND2    gate11282  (.A(g24653), .B(g34315), .Z(g34584) ) ;
INV     gate11283  (.A(g34584), .Z(II32803) ) ;
INV     gate11284  (.A(II32803), .Z(g34673) ) ;
AND2    gate11285  (.A(g24705), .B(g34316), .Z(g34585) ) ;
INV     gate11286  (.A(g34585), .Z(II32806) ) ;
INV     gate11287  (.A(II32806), .Z(g34674) ) ;
AND2    gate11288  (.A(g11025), .B(g34317), .Z(g34586) ) ;
INV     gate11289  (.A(g34586), .Z(II32809) ) ;
INV     gate11290  (.A(II32809), .Z(g34675) ) ;
AND2    gate11291  (.A(g26082), .B(g34323), .Z(g34588) ) ;
INV     gate11292  (.A(g34588), .Z(II32812) ) ;
INV     gate11293  (.A(II32812), .Z(g34676) ) ;
AND2    gate11294  (.A(g7834), .B(g34325), .Z(g34470) ) ;
INV     gate11295  (.A(g34470), .Z(II32815) ) ;
INV     gate11296  (.A(II32815), .Z(g34677) ) ;
AND2    gate11297  (.A(g20083), .B(g34326), .Z(g34474) ) ;
INV     gate11298  (.A(g34474), .Z(II32820) ) ;
INV     gate11299  (.A(II32820), .Z(g34680) ) ;
AND2    gate11300  (.A(g27450), .B(g34327), .Z(g34475) ) ;
INV     gate11301  (.A(g34475), .Z(II32824) ) ;
INV     gate11302  (.A(II32824), .Z(g34682) ) ;
AND2    gate11303  (.A(g26344), .B(g34328), .Z(g34477) ) ;
INV     gate11304  (.A(g34477), .Z(II32827) ) ;
INV     gate11305  (.A(II32827), .Z(g34683) ) ;
INV     gate11306  (.A(g34472), .Z(II32834) ) ;
INV     gate11307  (.A(II32834), .Z(g34688) ) ;
AND2    gate11308  (.A(g13888), .B(g34336), .Z(g34498) ) ;
INV     gate11309  (.A(g34498), .Z(II32837) ) ;
INV     gate11310  (.A(II32837), .Z(g34689) ) ;
INV     gate11311  (.A(g34480), .Z(II32840) ) ;
INV     gate11312  (.A(II32840), .Z(g34690) ) ;
AND2    gate11313  (.A(g31288), .B(g34339), .Z(g34499) ) ;
INV     gate11314  (.A(g34499), .Z(II32843) ) ;
INV     gate11315  (.A(II32843), .Z(g34691) ) ;
AND2    gate11316  (.A(g26363), .B(g34343), .Z(g34502) ) ;
INV     gate11317  (.A(g34502), .Z(II32846) ) ;
INV     gate11318  (.A(II32846), .Z(g34692) ) ;
NAND3   gate11319  (.A(g11679), .B(g794), .C(g34354), .Z(g34545) ) ;
INV     gate11320  (.A(g34545), .Z(g34697) ) ;
NAND3   gate11321  (.A(g626), .B(g34359), .C(g12323), .Z(g34550) ) ;
INV     gate11322  (.A(g34550), .Z(g34698) ) ;
INV     gate11323  (.A(g34540), .Z(II32855) ) ;
INV     gate11324  (.A(II32855), .Z(g34699) ) ;
INV     gate11325  (.A(g34559), .Z(g34711) ) ;
INV     gate11326  (.A(g34579), .Z(II32868) ) ;
INV     gate11327  (.A(II32868), .Z(g34712) ) ;
INV     gate11328  (.A(g34521), .Z(II32871) ) ;
INV     gate11329  (.A(II32871), .Z(g34713) ) ;
INV     gate11330  (.A(g34504), .Z(II32874) ) ;
INV     gate11331  (.A(II32874), .Z(g34714) ) ;
INV     gate11332  (.A(g34501), .Z(II32878) ) ;
INV     gate11333  (.A(II32878), .Z(g34716) ) ;
INV     gate11334  (.A(g34688), .Z(II32881) ) ;
INV     gate11335  (.A(g34690), .Z(II32884) ) ;
OR2     gate11336  (.A(g33381), .B(g34572), .Z(g34708) ) ;
INV     gate11337  (.A(g34708), .Z(II32904) ) ;
INV     gate11338  (.A(II32904), .Z(g34736) ) ;
INV     gate11339  (.A(g34712), .Z(II32909) ) ;
INV     gate11340  (.A(II32909), .Z(g34739) ) ;
NAND2   gate11341  (.A(II32757), .B(II32758), .Z(g34650) ) ;
INV     gate11342  (.A(g34650), .Z(II32921) ) ;
INV     gate11343  (.A(II32921), .Z(g34749) ) ;
OR2     gate11344  (.A(g33111), .B(g34492), .Z(g34649) ) ;
INV     gate11345  (.A(g34649), .Z(II32929) ) ;
INV     gate11346  (.A(II32929), .Z(g34755) ) ;
OR2     gate11347  (.A(g33114), .B(g34497), .Z(g34657) ) ;
INV     gate11348  (.A(g34657), .Z(II32935) ) ;
INV     gate11349  (.A(II32935), .Z(g34759) ) ;
OR2     gate11350  (.A(g32028), .B(g34500), .Z(g34663) ) ;
INV     gate11351  (.A(g34663), .Z(II32938) ) ;
INV     gate11352  (.A(II32938), .Z(g34760) ) ;
NOR3    gate11353  (.A(g8899), .B(g34545), .C(g11083), .Z(g34703) ) ;
INV     gate11354  (.A(g34703), .Z(g34766) ) ;
INV     gate11355  (.A(g34659), .Z(II32947) ) ;
INV     gate11356  (.A(II32947), .Z(g34767) ) ;
INV     gate11357  (.A(g34713), .Z(II32950) ) ;
INV     gate11358  (.A(II32950), .Z(g34768) ) ;
INV     gate11359  (.A(g34656), .Z(II32953) ) ;
INV     gate11360  (.A(II32953), .Z(g34769) ) ;
INV     gate11361  (.A(g34654), .Z(II32956) ) ;
INV     gate11362  (.A(II32956), .Z(g34770) ) ;
INV     gate11363  (.A(g34653), .Z(II32960) ) ;
INV     gate11364  (.A(II32960), .Z(g34772) ) ;
INV     gate11365  (.A(g34650), .Z(II32963) ) ;
INV     gate11366  (.A(II32963), .Z(g34773) ) ;
INV     gate11367  (.A(g34648), .Z(II32967) ) ;
INV     gate11368  (.A(II32967), .Z(g34775) ) ;
INV     gate11369  (.A(g34716), .Z(II32970) ) ;
INV     gate11370  (.A(II32970), .Z(g34776) ) ;
INV     gate11371  (.A(g34714), .Z(II32973) ) ;
INV     gate11372  (.A(II32973), .Z(g34777) ) ;
INV     gate11373  (.A(g34699), .Z(II32976) ) ;
INV     gate11374  (.A(II32976), .Z(g34778) ) ;
INV     gate11375  (.A(g34749), .Z(II32982) ) ;
INV     gate11376  (.A(II32982), .Z(g34784) ) ;
INV     gate11377  (.A(g34736), .Z(II32985) ) ;
INV     gate11378  (.A(g34755), .Z(II32988) ) ;
INV     gate11379  (.A(g34759), .Z(II32991) ) ;
INV     gate11380  (.A(g34739), .Z(II32994) ) ;
INV     gate11381  (.A(g34760), .Z(II32997) ) ;
OR2     gate11382  (.A(g33431), .B(g34715), .Z(g34781) ) ;
INV     gate11383  (.A(g34781), .Z(II33020) ) ;
INV     gate11384  (.A(II33020), .Z(g34810) ) ;
OR2     gate11385  (.A(g33110), .B(g34667), .Z(g34783) ) ;
INV     gate11386  (.A(g34783), .Z(II33024) ) ;
INV     gate11387  (.A(II33024), .Z(g34812) ) ;
INV     gate11388  (.A(g34767), .Z(II33027) ) ;
INV     gate11389  (.A(II33027), .Z(g34813) ) ;
INV     gate11390  (.A(g34768), .Z(II33030) ) ;
INV     gate11391  (.A(II33030), .Z(g34816) ) ;
INV     gate11392  (.A(g34769), .Z(II33034) ) ;
INV     gate11393  (.A(II33034), .Z(g34820) ) ;
INV     gate11394  (.A(g34770), .Z(II33037) ) ;
INV     gate11395  (.A(II33037), .Z(g34823) ) ;
INV     gate11396  (.A(g34772), .Z(II33041) ) ;
INV     gate11397  (.A(II33041), .Z(g34827) ) ;
INV     gate11398  (.A(g34775), .Z(II33044) ) ;
INV     gate11399  (.A(II33044), .Z(g34830) ) ;
INV     gate11400  (.A(g34776), .Z(II33047) ) ;
INV     gate11401  (.A(II33047), .Z(g34833) ) ;
INV     gate11402  (.A(g34777), .Z(II33050) ) ;
INV     gate11403  (.A(II33050), .Z(g34836) ) ;
INV     gate11404  (.A(g34778), .Z(II33053) ) ;
INV     gate11405  (.A(g34778), .Z(II33056) ) ;
INV     gate11406  (.A(II33056), .Z(g34840) ) ;
NOR2    gate11407  (.A(g34706), .B(g30003), .Z(g34737) ) ;
INV     gate11408  (.A(g34737), .Z(g34844) ) ;
INV     gate11409  (.A(g34773), .Z(g34845) ) ;
INV     gate11410  (.A(g34784), .Z(II33064) ) ;
INV     gate11411  (.A(II33064), .Z(g34846) ) ;
INV     gate11412  (.A(g34812), .Z(II33067) ) ;
INV     gate11413  (.A(g34810), .Z(II33070) ) ;
OR2     gate11414  (.A(g33924), .B(g34782), .Z(g34843) ) ;
INV     gate11415  (.A(g34843), .Z(II33075) ) ;
INV     gate11416  (.A(II33075), .Z(g34851) ) ;
INV     gate11417  (.A(g34845), .Z(g34852) ) ;
OR2     gate11418  (.A(g33677), .B(g34738), .Z(g34809) ) ;
INV     gate11419  (.A(g34809), .Z(II33079) ) ;
INV     gate11420  (.A(II33079), .Z(g34855) ) ;
INV     gate11421  (.A(g34840), .Z(g34864) ) ;
INV     gate11422  (.A(g34846), .Z(II33103) ) ;
INV     gate11423  (.A(g34855), .Z(II33106) ) ;
INV     gate11424  (.A(g34851), .Z(II33109) ) ;
INV     gate11425  (.A(g34852), .Z(g34883) ) ;
INV     gate11426  (.A(g34852), .Z(II33119) ) ;
INV     gate11427  (.A(II33119), .Z(g34893) ) ;
INV     gate11428  (.A(g34864), .Z(g34910) ) ;
OR2     gate11429  (.A(g34857), .B(g21694), .Z(g34906) ) ;
INV     gate11430  (.A(g34906), .Z(II33131) ) ;
INV     gate11431  (.A(g34906), .Z(II33134) ) ;
INV     gate11432  (.A(II33134), .Z(g34914) ) ;
OR2     gate11433  (.A(g34858), .B(g21666), .Z(g34884) ) ;
INV     gate11434  (.A(g34884), .Z(II33137) ) ;
INV     gate11435  (.A(g34884), .Z(II33140) ) ;
INV     gate11436  (.A(II33140), .Z(g34916) ) ;
OR2     gate11437  (.A(g34859), .B(g21690), .Z(g34903) ) ;
INV     gate11438  (.A(g34903), .Z(II33143) ) ;
INV     gate11439  (.A(g34903), .Z(II33146) ) ;
INV     gate11440  (.A(II33146), .Z(g34918) ) ;
OR2     gate11441  (.A(g34860), .B(g21686), .Z(g34900) ) ;
INV     gate11442  (.A(g34900), .Z(II33149) ) ;
INV     gate11443  (.A(g34900), .Z(II33152) ) ;
INV     gate11444  (.A(II33152), .Z(g34920) ) ;
OR2     gate11445  (.A(g34861), .B(g21682), .Z(g34897) ) ;
INV     gate11446  (.A(g34897), .Z(II33155) ) ;
INV     gate11447  (.A(g34897), .Z(II33158) ) ;
INV     gate11448  (.A(II33158), .Z(g34922) ) ;
OR2     gate11449  (.A(g34862), .B(g21678), .Z(g34894) ) ;
INV     gate11450  (.A(g34894), .Z(II33161) ) ;
INV     gate11451  (.A(g34894), .Z(II33164) ) ;
INV     gate11452  (.A(II33164), .Z(g34924) ) ;
OR2     gate11453  (.A(g34863), .B(g21674), .Z(g34890) ) ;
INV     gate11454  (.A(g34890), .Z(II33167) ) ;
INV     gate11455  (.A(g34890), .Z(II33170) ) ;
INV     gate11456  (.A(II33170), .Z(g34926) ) ;
OR2     gate11457  (.A(g34865), .B(g21670), .Z(g34887) ) ;
INV     gate11458  (.A(g34887), .Z(II33173) ) ;
INV     gate11459  (.A(g34887), .Z(II33176) ) ;
INV     gate11460  (.A(II33176), .Z(g34928) ) ;
INV     gate11461  (.A(g34893), .Z(II33179) ) ;
INV     gate11462  (.A(II33179), .Z(g34929) ) ;
INV     gate11463  (.A(g34910), .Z(II33182) ) ;
INV     gate11464  (.A(II33182), .Z(g34930) ) ;
INV     gate11465  (.A(g34914), .Z(g34932) ) ;
INV     gate11466  (.A(g34916), .Z(g34933) ) ;
INV     gate11467  (.A(g34918), .Z(g34934) ) ;
INV     gate11468  (.A(g34929), .Z(II33189) ) ;
INV     gate11469  (.A(II33189), .Z(g34935) ) ;
INV     gate11470  (.A(g34920), .Z(g34938) ) ;
INV     gate11471  (.A(g34922), .Z(g34939) ) ;
INV     gate11472  (.A(g34924), .Z(g34940) ) ;
INV     gate11473  (.A(g34926), .Z(g34941) ) ;
INV     gate11474  (.A(g34928), .Z(g34942) ) ;
INV     gate11475  (.A(g34930), .Z(II33197) ) ;
INV     gate11476  (.A(II33197), .Z(g34943) ) ;
INV     gate11477  (.A(g34932), .Z(g34944) ) ;
INV     gate11478  (.A(g34933), .Z(g34945) ) ;
INV     gate11479  (.A(g34934), .Z(g34946) ) ;
INV     gate11480  (.A(g34938), .Z(g34947) ) ;
INV     gate11481  (.A(g34939), .Z(g34949) ) ;
INV     gate11482  (.A(g34940), .Z(g34950) ) ;
INV     gate11483  (.A(g34941), .Z(g34951) ) ;
INV     gate11484  (.A(g34942), .Z(g34952) ) ;
INV     gate11485  (.A(g34943), .Z(II33210) ) ;
INV     gate11486  (.A(II33210), .Z(g34954) ) ;
INV     gate11487  (.A(g34954), .Z(II33214) ) ;
AND2    gate11488  (.A(g34931), .B(g34320), .Z(g34955) ) ;
INV     gate11489  (.A(g34955), .Z(II33218) ) ;
INV     gate11490  (.A(II33218), .Z(g34960) ) ;
OR2     gate11491  (.A(g34948), .B(g21662), .Z(g34957) ) ;
INV     gate11492  (.A(g34957), .Z(II33232) ) ;
INV     gate11493  (.A(g34957), .Z(II33235) ) ;
INV     gate11494  (.A(II33235), .Z(g34973) ) ;
INV     gate11495  (.A(g34973), .Z(g34981) ) ;
OR2     gate11496  (.A(g34868), .B(g34961), .Z(g34970) ) ;
INV     gate11497  (.A(g34970), .Z(II33246) ) ;
INV     gate11498  (.A(II33246), .Z(g34982) ) ;
OR2     gate11499  (.A(g34869), .B(g34962), .Z(g34971) ) ;
INV     gate11500  (.A(g34971), .Z(II33249) ) ;
INV     gate11501  (.A(II33249), .Z(g34983) ) ;
OR2     gate11502  (.A(g34870), .B(g34963), .Z(g34974) ) ;
INV     gate11503  (.A(g34974), .Z(II33252) ) ;
INV     gate11504  (.A(II33252), .Z(g34984) ) ;
OR2     gate11505  (.A(g34871), .B(g34964), .Z(g34975) ) ;
INV     gate11506  (.A(g34975), .Z(II33255) ) ;
INV     gate11507  (.A(II33255), .Z(g34985) ) ;
OR2     gate11508  (.A(g34872), .B(g34965), .Z(g34976) ) ;
INV     gate11509  (.A(g34976), .Z(II33258) ) ;
INV     gate11510  (.A(II33258), .Z(g34986) ) ;
OR2     gate11511  (.A(g34873), .B(g34966), .Z(g34977) ) ;
INV     gate11512  (.A(g34977), .Z(II33261) ) ;
INV     gate11513  (.A(II33261), .Z(g34987) ) ;
OR2     gate11514  (.A(g34874), .B(g34967), .Z(g34978) ) ;
INV     gate11515  (.A(g34978), .Z(II33264) ) ;
INV     gate11516  (.A(II33264), .Z(g34988) ) ;
OR2     gate11517  (.A(g34875), .B(g34968), .Z(g34979) ) ;
INV     gate11518  (.A(g34979), .Z(II33267) ) ;
INV     gate11519  (.A(II33267), .Z(g34989) ) ;
INV     gate11520  (.A(g34982), .Z(II33270) ) ;
INV     gate11521  (.A(g34984), .Z(II33273) ) ;
INV     gate11522  (.A(g34985), .Z(II33276) ) ;
INV     gate11523  (.A(g34986), .Z(II33279) ) ;
INV     gate11524  (.A(g34987), .Z(II33282) ) ;
INV     gate11525  (.A(g34988), .Z(II33285) ) ;
INV     gate11526  (.A(g34989), .Z(II33288) ) ;
INV     gate11527  (.A(g34983), .Z(II33291) ) ;
INV     gate11528  (.A(g34981), .Z(g34998) ) ;
OR2     gate11529  (.A(g34953), .B(g34999), .Z(g35000) ) ;
INV     gate11530  (.A(g35000), .Z(II33297) ) ;
INV     gate11531  (.A(II33297), .Z(g35001) ) ;
INV     gate11532  (.A(g35001), .Z(II33300) ) ;
AND2    gate11533  (.A(g452), .B(g392), .Z(g7251) ) ;
AND2    gate11534  (.A(g392), .B(g441), .Z(g7396) ) ;
AND2    gate11535  (.A(g4382), .B(g4438), .Z(g7469) ) ;
AND3    gate11536  (.A(g2145), .B(g2138), .C(g2130), .Z(g7511) ) ;
AND3    gate11537  (.A(g2704), .B(g2697), .C(g2689), .Z(g7520) ) ;
AND2    gate11538  (.A(g4382), .B(g4375), .Z(g7685) ) ;
AND2    gate11539  (.A(g2955), .B(g2950), .Z(g7696) ) ;
AND2    gate11540  (.A(g2965), .B(g2960), .Z(g7763) ) ;
AND3    gate11541  (.A(g723), .B(g822), .C(g817), .Z(g7777) ) ;
AND2    gate11542  (.A(g2975), .B(g2970), .Z(g7804) ) ;
AND2    gate11543  (.A(g4515), .B(g4521), .Z(g8234) ) ;
AND2    gate11544  (.A(g2902), .B(g2907), .Z(g8530) ) ;
AND2    gate11545  (.A(g2917), .B(g2912), .Z(g8583) ) ;
AND2    gate11546  (.A(g2927), .B(g2922), .Z(g8643) ) ;
AND2    gate11547  (.A(g2941), .B(g2936), .Z(g8690) ) ;
AND3    gate11548  (.A(g385), .B(g376), .C(g365), .Z(g8721) ) ;
AND2    gate11549  (.A(g632), .B(g626), .Z(g9217) ) ;
AND2    gate11550  (.A(g305), .B(g324), .Z(g9479) ) ;
AND2    gate11551  (.A(g996), .B(g1157), .Z(g9906) ) ;
AND2    gate11552  (.A(g1178), .B(g1157), .Z(g9967) ) ;
AND2    gate11553  (.A(g1339), .B(g1500), .Z(g9968) ) ;
AND2    gate11554  (.A(g1521), .B(g1500), .Z(g10034) ) ;
AND2    gate11555  (.A(g4358), .B(g4349), .Z(g10290) ) ;
AND3    gate11556  (.A(g7232), .B(g7219), .C(g7258), .Z(II13862) ) ;
AND2    gate11557  (.A(g1233), .B(g9007), .Z(g10501) ) ;
AND2    gate11558  (.A(g1576), .B(g9051), .Z(g10528) ) ;
NAND2   gate11559  (.A(II12469), .B(II12470), .Z(g8238) ) ;
AND2    gate11560  (.A(g8238), .B(g437), .Z(g10543) ) ;
NOR2    gate11561  (.A(g405), .B(g392), .Z(g8182) ) ;
AND2    gate11562  (.A(g8182), .B(g424), .Z(g10565) ) ;
AND3    gate11563  (.A(g7340), .B(g7293), .C(g7261), .Z(II13937) ) ;
AND2    gate11564  (.A(g7998), .B(g174), .Z(g10616) ) ;
AND2    gate11565  (.A(g3080), .B(g7907), .Z(g10619) ) ;
AND2    gate11566  (.A(g8387), .B(g3072), .Z(g10624) ) ;
AND2    gate11567  (.A(g3431), .B(g7926), .Z(g10625) ) ;
AND2    gate11568  (.A(g4057), .B(g7927), .Z(g10626) ) ;
AND2    gate11569  (.A(g3085), .B(g8434), .Z(g10654) ) ;
AND2    gate11570  (.A(g8440), .B(g3423), .Z(g10655) ) ;
AND2    gate11571  (.A(g3782), .B(g7952), .Z(g10656) ) ;
AND2    gate11572  (.A(g8451), .B(g4064), .Z(g10657) ) ;
AND2    gate11573  (.A(g209), .B(g8292), .Z(g10665) ) ;
AND3    gate11574  (.A(g6841), .B(g10200), .C(g2130), .Z(g10674) ) ;
AND2    gate11575  (.A(g3436), .B(g8500), .Z(g10675) ) ;
AND2    gate11576  (.A(g8506), .B(g3774), .Z(g10676) ) ;
AND2    gate11577  (.A(g4141), .B(g7611), .Z(g10677) ) ;
AND2    gate11578  (.A(g7289), .B(g4438), .Z(g10683) ) ;
AND2    gate11579  (.A(g7998), .B(g411), .Z(g10684) ) ;
AND3    gate11580  (.A(g2145), .B(g10200), .C(g2130), .Z(g10704) ) ;
AND3    gate11581  (.A(g6850), .B(g10219), .C(g2689), .Z(g10705) ) ;
AND2    gate11582  (.A(g3338), .B(g8691), .Z(g10706) ) ;
AND2    gate11583  (.A(g3787), .B(g8561), .Z(g10707) ) ;
AND3    gate11584  (.A(g6841), .B(g2138), .C(g2130), .Z(g10719) ) ;
AND3    gate11585  (.A(g2704), .B(g10219), .C(g2689), .Z(g10720) ) ;
AND4    gate11586  (.A(g3288), .B(g6875), .C(g3274), .D(g8481), .Z(g10721) ) ;
AND2    gate11587  (.A(g3689), .B(g8728), .Z(g10724) ) ;
AND3    gate11588  (.A(g6850), .B(g2697), .C(g2689), .Z(g10732) ) ;
AND4    gate11589  (.A(g3639), .B(g6905), .C(g3625), .D(g8542), .Z(g10733) ) ;
AND2    gate11590  (.A(g4040), .B(g8751), .Z(g10736) ) ;
AND4    gate11591  (.A(g3990), .B(g6928), .C(g3976), .D(g8595), .Z(g10756) ) ;
AND2    gate11592  (.A(g4264), .B(g8514), .Z(g10822) ) ;
AND2    gate11593  (.A(g8914), .B(g4258), .Z(g10827) ) ;
AND2    gate11594  (.A(g6888), .B(g7640), .Z(g10828) ) ;
AND2    gate11595  (.A(g7289), .B(g4375), .Z(g10829) ) ;
AND2    gate11596  (.A(g8509), .B(g8567), .Z(g10841) ) ;
AND2    gate11597  (.A(g4269), .B(g8967), .Z(g10856) ) ;
AND2    gate11598  (.A(g3004), .B(g9015), .Z(g10873) ) ;
AND2    gate11599  (.A(g7858), .B(g1135), .Z(g10878) ) ;
AND2    gate11600  (.A(g3355), .B(g9061), .Z(g10883) ) ;
AND2    gate11601  (.A(g7858), .B(g1105), .Z(g10890) ) ;
AND2    gate11602  (.A(g1205), .B(g8654), .Z(g10896) ) ;
AND2    gate11603  (.A(g3706), .B(g9100), .Z(g10898) ) ;
AND2    gate11604  (.A(g7858), .B(g1129), .Z(g10902) ) ;
AND2    gate11605  (.A(g9174), .B(g1087), .Z(g10917) ) ;
AND2    gate11606  (.A(g1548), .B(g8685), .Z(g10921) ) ;
AND2    gate11607  (.A(g7858), .B(g956), .Z(g10925) ) ;
AND2    gate11608  (.A(g9197), .B(g7918), .Z(g10934) ) ;
AND2    gate11609  (.A(g9200), .B(g1430), .Z(g10947) ) ;
AND2    gate11610  (.A(g7880), .B(g1478), .Z(g10948) ) ;
AND2    gate11611  (.A(g9226), .B(g7948), .Z(g10966) ) ;
AND2    gate11612  (.A(g7880), .B(g1448), .Z(g10967) ) ;
AND2    gate11613  (.A(g854), .B(g9582), .Z(g10970) ) ;
AND4    gate11614  (.A(g8567), .B(g8509), .C(g8451), .D(g7650), .Z(g10998) ) ;
AND2    gate11615  (.A(g7880), .B(g1472), .Z(g10999) ) ;
AND2    gate11616  (.A(g7880), .B(g1300), .Z(g11003) ) ;
NOR2    gate11617  (.A(g4709), .B(g4785), .Z(g8933) ) ;
AND2    gate11618  (.A(g4698), .B(g8933), .Z(g11010) ) ;
NOR2    gate11619  (.A(g4899), .B(g4975), .Z(g8984) ) ;
AND2    gate11620  (.A(g4888), .B(g8984), .Z(g11016) ) ;
AND2    gate11621  (.A(g5092), .B(g9036), .Z(g11019) ) ;
AND2    gate11622  (.A(g9669), .B(g5084), .Z(g11023) ) ;
AND2    gate11623  (.A(g5436), .B(g9070), .Z(g11024) ) ;
AND2    gate11624  (.A(g5097), .B(g9724), .Z(g11027) ) ;
AND2    gate11625  (.A(g9730), .B(g5428), .Z(g11028) ) ;
AND2    gate11626  (.A(g5782), .B(g9103), .Z(g11029) ) ;
AND2    gate11627  (.A(g9354), .B(g7717), .Z(g11032) ) ;
AND2    gate11628  (.A(g5441), .B(g9800), .Z(g11035) ) ;
AND2    gate11629  (.A(g9806), .B(g5774), .Z(g11036) ) ;
AND2    gate11630  (.A(g6128), .B(g9184), .Z(g11037) ) ;
AND2    gate11631  (.A(g5343), .B(g10124), .Z(g11044) ) ;
AND2    gate11632  (.A(g5787), .B(g9883), .Z(g11045) ) ;
AND2    gate11633  (.A(g9889), .B(g6120), .Z(g11046) ) ;
AND2    gate11634  (.A(g6474), .B(g9212), .Z(g11047) ) ;
AND4    gate11635  (.A(g5297), .B(g7004), .C(g5283), .D(g9780), .Z(g11111) ) ;
AND2    gate11636  (.A(g5689), .B(g10160), .Z(g11114) ) ;
AND2    gate11637  (.A(g6133), .B(g9954), .Z(g11115) ) ;
AND2    gate11638  (.A(g9960), .B(g6466), .Z(g11116) ) ;
AND4    gate11639  (.A(g5644), .B(g7028), .C(g5630), .D(g9864), .Z(g11123) ) ;
AND2    gate11640  (.A(g6035), .B(g10185), .Z(g11126) ) ;
AND2    gate11641  (.A(g6479), .B(g10022), .Z(g11127) ) ;
AND4    gate11642  (.A(g5990), .B(g7051), .C(g5976), .D(g9935), .Z(g11139) ) ;
AND2    gate11643  (.A(g6381), .B(g10207), .Z(g11142) ) ;
AND4    gate11644  (.A(g225), .B(g8237), .C(g232), .D(g8180), .Z(II14198) ) ;
AND4    gate11645  (.A(g239), .B(g8136), .C(g246), .D(II14198), .Z(g11144) ) ;
AND4    gate11646  (.A(g6336), .B(g7074), .C(g6322), .D(g10003), .Z(g11160) ) ;
AND2    gate11647  (.A(g6727), .B(g10224), .Z(g11163) ) ;
AND4    gate11648  (.A(g8457), .B(g255), .C(g8406), .D(g262), .Z(II14225) ) ;
AND4    gate11649  (.A(g8363), .B(g269), .C(g8296), .D(II14225), .Z(g11166) ) ;
AND4    gate11650  (.A(g6682), .B(g7097), .C(g6668), .D(g10061), .Z(g11178) ) ;
AND2    gate11651  (.A(g8217), .B(g8439), .Z(g11205) ) ;
AND2    gate11652  (.A(g8281), .B(g8505), .Z(g11223) ) ;
AND2    gate11653  (.A(g8346), .B(g8566), .Z(g11244) ) ;
AND2    gate11654  (.A(g5016), .B(g10338), .Z(g11366) ) ;
AND2    gate11655  (.A(g5360), .B(g7139), .Z(g11397) ) ;
AND2    gate11656  (.A(g5706), .B(g7158), .Z(g11427) ) ;
AND2    gate11657  (.A(g6052), .B(g7175), .Z(g11449) ) ;
AND2    gate11658  (.A(g4382), .B(g7495), .Z(g11496) ) ;
AND2    gate11659  (.A(g6398), .B(g7192), .Z(g11497) ) ;
AND2    gate11660  (.A(g7289), .B(g4375), .Z(g11546) ) ;
NAND2   gate11661  (.A(g691), .B(g714), .Z(g8769) ) ;
AND2    gate11662  (.A(g8769), .B(g703), .Z(g11740) ) ;
NOR2    gate11663  (.A(g333), .B(g355), .Z(g7499) ) ;
AND2    gate11664  (.A(g7499), .B(g9155), .Z(g11890) ) ;
AND2    gate11665  (.A(g1668), .B(g7268), .Z(g11893) ) ;
AND2    gate11666  (.A(g1802), .B(g7315), .Z(g11915) ) ;
AND2    gate11667  (.A(g2227), .B(g7328), .Z(g11916) ) ;
AND2    gate11668  (.A(g1936), .B(g7362), .Z(g11937) ) ;
AND2    gate11669  (.A(g2361), .B(g7380), .Z(g11939) ) ;
AND2    gate11670  (.A(g2070), .B(g7411), .Z(g11956) ) ;
AND2    gate11671  (.A(g2495), .B(g7424), .Z(g11960) ) ;
AND2    gate11672  (.A(g311), .B(g7802), .Z(g11967) ) ;
AND2    gate11673  (.A(g2629), .B(g7462), .Z(g11978) ) ;
AND2    gate11674  (.A(g1002), .B(g7567), .Z(g12015) ) ;
AND2    gate11675  (.A(g9499), .B(g9729), .Z(g12027) ) ;
AND2    gate11676  (.A(g1345), .B(g7601), .Z(g12043) ) ;
AND2    gate11677  (.A(g9557), .B(g9805), .Z(g12065) ) ;
AND2    gate11678  (.A(g9619), .B(g9888), .Z(g12099) ) ;
AND2    gate11679  (.A(g9684), .B(g9959), .Z(g12135) ) ;
AND2    gate11680  (.A(g9745), .B(g10027), .Z(g12179) ) ;
AND2    gate11681  (.A(g1178), .B(g7519), .Z(g12186) ) ;
AND2    gate11682  (.A(g1189), .B(g7532), .Z(g12219) ) ;
AND2    gate11683  (.A(g1521), .B(g7535), .Z(g12220) ) ;
AND2    gate11684  (.A(g9480), .B(g640), .Z(g12259) ) ;
AND2    gate11685  (.A(g1532), .B(g7557), .Z(g12284) ) ;
AND2    gate11686  (.A(g8680), .B(g667), .Z(g12527) ) ;
AND2    gate11687  (.A(g9024), .B(g8977), .Z(g12687) ) ;
AND2    gate11688  (.A(g9024), .B(g4349), .Z(g12730) ) ;
AND2    gate11689  (.A(g969), .B(g7567), .Z(g12761) ) ;
AND2    gate11690  (.A(g4358), .B(g8977), .Z(g12762) ) ;
AND2    gate11691  (.A(g1008), .B(g7567), .Z(g12794) ) ;
AND2    gate11692  (.A(g1312), .B(g7601), .Z(g12795) ) ;
AND2    gate11693  (.A(g518), .B(g9158), .Z(g12812) ) ;
AND2    gate11694  (.A(g1351), .B(g7601), .Z(g12817) ) ;
AND2    gate11695  (.A(g1227), .B(g10960), .Z(g12920) ) ;
AND2    gate11696  (.A(g1570), .B(g10980), .Z(g12924) ) ;
AND2    gate11697  (.A(g392), .B(g11048), .Z(g12931) ) ;
AND2    gate11698  (.A(g405), .B(g11048), .Z(g12939) ) ;
AND2    gate11699  (.A(g411), .B(g11048), .Z(g12953) ) ;
AND2    gate11700  (.A(g424), .B(g11048), .Z(g12979) ) ;
AND2    gate11701  (.A(g194), .B(g11737), .Z(g13019) ) ;
AND2    gate11702  (.A(g401), .B(g11048), .Z(g13020) ) ;
AND2    gate11703  (.A(g8431), .B(g11026), .Z(g13025) ) ;
NAND2   gate11704  (.A(II12545), .B(II12546), .Z(g8359) ) ;
AND2    gate11705  (.A(g8359), .B(g11030), .Z(g13029) ) ;
AND2    gate11706  (.A(g429), .B(g11048), .Z(g13030) ) ;
AND2    gate11707  (.A(g8497), .B(g11033), .Z(g13035) ) ;
AND2    gate11708  (.A(g8509), .B(g11034), .Z(g13038) ) ;
AND2    gate11709  (.A(g433), .B(g11048), .Z(g13042) ) ;
AND2    gate11710  (.A(g6870), .B(g11270), .Z(g13046) ) ;
AND2    gate11711  (.A(g8534), .B(g11042), .Z(g13047) ) ;
AND2    gate11712  (.A(g8558), .B(g11043), .Z(g13048) ) ;
AND2    gate11713  (.A(g6900), .B(g11303), .Z(g13059) ) ;
AND2    gate11714  (.A(g8587), .B(g11110), .Z(g13060) ) ;
AND2    gate11715  (.A(g8567), .B(g10808), .Z(g13063) ) ;
AND2    gate11716  (.A(g6923), .B(g11357), .Z(g13080) ) ;
AND2    gate11717  (.A(g8626), .B(g11122), .Z(g13081) ) ;
AND3    gate11718  (.A(g10816), .B(g10812), .C(g10805), .Z(g13156) ) ;
AND2    gate11719  (.A(g6946), .B(g11425), .Z(g13221) ) ;
AND2    gate11720  (.A(g8964), .B(g11316), .Z(g13247) ) ;
NAND2   gate11721  (.A(II14517), .B(II14518), .Z(g11561) ) ;
NAND2   gate11722  (.A(II14481), .B(II14482), .Z(g11511) ) ;
NOR3    gate11723  (.A(g650), .B(g9903), .C(g645), .Z(g11469) ) ;
AND4    gate11724  (.A(g11561), .B(g11511), .C(g11469), .D(g699), .Z(g13252) ) ;
AND2    gate11725  (.A(g9018), .B(g11493), .Z(g13265) ) ;
AND2    gate11726  (.A(g3195), .B(g11432), .Z(g13277) ) ;
AND2    gate11727  (.A(g3546), .B(g11480), .Z(g13282) ) ;
AND2    gate11728  (.A(g1221), .B(g11472), .Z(g13287) ) ;
AND2    gate11729  (.A(g3897), .B(g11534), .Z(g13290) ) ;
AND2    gate11730  (.A(g1564), .B(g11513), .Z(g13294) ) ;
AND2    gate11731  (.A(g437), .B(g11048), .Z(g13299) ) ;
AND2    gate11732  (.A(g441), .B(g11048), .Z(g13306) ) ;
AND2    gate11733  (.A(g475), .B(g11048), .Z(g13313) ) ;
AND4    gate11734  (.A(g4076), .B(g8812), .C(g10658), .D(g8757), .Z(g13319) ) ;
AND2    gate11735  (.A(g417), .B(g11048), .Z(g13320) ) ;
AND2    gate11736  (.A(g847), .B(g11048), .Z(g13321) ) ;
AND2    gate11737  (.A(g854), .B(g11326), .Z(g13324) ) ;
NOR2    gate11738  (.A(g4709), .B(g8796), .Z(g11755) ) ;
AND2    gate11739  (.A(g4743), .B(g11755), .Z(g13333) ) ;
NOR2    gate11740  (.A(g8883), .B(g4785), .Z(g11773) ) ;
AND2    gate11741  (.A(g4754), .B(g11773), .Z(g13345) ) ;
NOR2    gate11742  (.A(g4899), .B(g8822), .Z(g11780) ) ;
AND2    gate11743  (.A(g4933), .B(g11780), .Z(g13349) ) ;
NOR2    gate11744  (.A(g8883), .B(g8796), .Z(g11797) ) ;
AND2    gate11745  (.A(g4765), .B(g11797), .Z(g13383) ) ;
NOR2    gate11746  (.A(g8938), .B(g4975), .Z(g11804) ) ;
AND2    gate11747  (.A(g4944), .B(g11804), .Z(g13384) ) ;
AND2    gate11748  (.A(g703), .B(g11048), .Z(g13393) ) ;
NOR2    gate11749  (.A(g8938), .B(g8822), .Z(g11834) ) ;
AND2    gate11750  (.A(g4955), .B(g11834), .Z(g13411) ) ;
AND2    gate11751  (.A(g837), .B(g11048), .Z(g13415) ) ;
AND2    gate11752  (.A(g9721), .B(g11811), .Z(g13436) ) ;
AND2    gate11753  (.A(g2719), .B(g11819), .Z(g13461) ) ;
AND2    gate11754  (.A(g9797), .B(g11841), .Z(g13473) ) ;
AND2    gate11755  (.A(g6999), .B(g12160), .Z(g13491) ) ;
AND2    gate11756  (.A(g9856), .B(g11865), .Z(g13492) ) ;
AND2    gate11757  (.A(g9880), .B(g11866), .Z(g13493) ) ;
AND2    gate11758  (.A(g2724), .B(g12155), .Z(g13497) ) ;
AND2    gate11759  (.A(g7023), .B(g12198), .Z(g13507) ) ;
AND2    gate11760  (.A(g9927), .B(g11888), .Z(g13508) ) ;
AND2    gate11761  (.A(g9951), .B(g11889), .Z(g13509) ) ;
AND2    gate11762  (.A(g7046), .B(g12246), .Z(g13523) ) ;
AND2    gate11763  (.A(g9995), .B(g11910), .Z(g13524) ) ;
AND2    gate11764  (.A(g10019), .B(g11911), .Z(g13525) ) ;
AND2    gate11765  (.A(g7069), .B(g12308), .Z(g13541) ) ;
AND2    gate11766  (.A(g10053), .B(g11927), .Z(g13542) ) ;
AND2    gate11767  (.A(g4480), .B(g12820), .Z(g13564) ) ;
AND2    gate11768  (.A(g7092), .B(g12358), .Z(g13566) ) ;
AND2    gate11769  (.A(g10102), .B(g11948), .Z(g13567) ) ;
AND2    gate11770  (.A(g4495), .B(g10487), .Z(g13604) ) ;
AND2    gate11771  (.A(g10232), .B(g12228), .Z(g13632) ) ;
AND2    gate11772  (.A(g4567), .B(g10509), .Z(g13633) ) ;
AND2    gate11773  (.A(g278), .B(g11144), .Z(g13656) ) ;
AND2    gate11774  (.A(g4498), .B(g10532), .Z(g13671) ) ;
AND2    gate11775  (.A(g11166), .B(g8608), .Z(g13697) ) ;
AND2    gate11776  (.A(g4501), .B(g10571), .Z(g13737) ) ;
AND2    gate11777  (.A(g8880), .B(g10572), .Z(g13738) ) ;
NAND2   gate11778  (.A(g9842), .B(g3298), .Z(g11409) ) ;
NAND2   gate11779  (.A(g9660), .B(g3274), .Z(g11381) ) ;
AND3    gate11780  (.A(g8691), .B(g11409), .C(g11381), .Z(II16111) ) ;
NAND2   gate11781  (.A(g9599), .B(g3267), .Z(g11441) ) ;
NAND2   gate11782  (.A(g9551), .B(g3310), .Z(g11355) ) ;
NAND2   gate11783  (.A(g9496), .B(g3281), .Z(g11302) ) ;
AND4    gate11784  (.A(g11441), .B(g11355), .C(g11302), .D(II16111), .Z(g13771) ) ;
AND2    gate11785  (.A(g4540), .B(g10597), .Z(g13778) ) ;
NAND2   gate11786  (.A(g9916), .B(g3649), .Z(g11443) ) ;
NAND2   gate11787  (.A(g9713), .B(g3625), .Z(g11411) ) ;
AND3    gate11788  (.A(g8728), .B(g11443), .C(g11411), .Z(II16129) ) ;
NAND2   gate11789  (.A(g9661), .B(g3618), .Z(g11489) ) ;
NAND2   gate11790  (.A(g9600), .B(g3661), .Z(g11394) ) ;
NAND2   gate11791  (.A(g9552), .B(g3632), .Z(g11356) ) ;
AND4    gate11792  (.A(g11489), .B(g11394), .C(g11356), .D(II16129), .Z(g13805) ) ;
AND2    gate11793  (.A(g4504), .B(g10606), .Z(g13807) ) ;
AND2    gate11794  (.A(g4543), .B(g10607), .Z(g13808) ) ;
NAND2   gate11795  (.A(g9982), .B(g4000), .Z(g11491) ) ;
NAND2   gate11796  (.A(g9771), .B(g3976), .Z(g11445) ) ;
AND3    gate11797  (.A(g8751), .B(g11491), .C(g11445), .Z(II16143) ) ;
NAND2   gate11798  (.A(g9714), .B(g3969), .Z(g11543) ) ;
NAND2   gate11799  (.A(g9662), .B(g4012), .Z(g11424) ) ;
NAND2   gate11800  (.A(g9601), .B(g3983), .Z(g11395) ) ;
AND4    gate11801  (.A(g11543), .B(g11424), .C(g11395), .D(II16143), .Z(g13830) ) ;
AND2    gate11802  (.A(g8880), .B(g10612), .Z(g13832) ) ;
AND2    gate11803  (.A(g4546), .B(g10613), .Z(g13833) ) ;
AND2    gate11804  (.A(g4549), .B(g10620), .Z(g13853) ) ;
AND2    gate11805  (.A(g5204), .B(g12402), .Z(g13887) ) ;
AND2    gate11806  (.A(g5551), .B(g12450), .Z(g13912) ) ;
AND2    gate11807  (.A(g5897), .B(g12512), .Z(g13942) ) ;
AND2    gate11808  (.A(g6243), .B(g12578), .Z(g13974) ) ;
AND2    gate11809  (.A(g6589), .B(g12629), .Z(g13998) ) ;
AND2    gate11810  (.A(g8673), .B(g11797), .Z(g14028) ) ;
AND2    gate11811  (.A(g699), .B(g11048), .Z(g14035) ) ;
AND2    gate11812  (.A(g8715), .B(g11834), .Z(g14061) ) ;
AND2    gate11813  (.A(g878), .B(g10632), .Z(g14097) ) ;
AND2    gate11814  (.A(g881), .B(g10632), .Z(g14126) ) ;
AND2    gate11815  (.A(g884), .B(g10632), .Z(g14148) ) ;
AND2    gate11816  (.A(g887), .B(g10632), .Z(g14168) ) ;
AND2    gate11817  (.A(g872), .B(g10632), .Z(g14180) ) ;
AND2    gate11818  (.A(g8686), .B(g11744), .Z(g14185) ) ;
AND2    gate11819  (.A(g859), .B(g10632), .Z(g14190) ) ;
AND2    gate11820  (.A(g7178), .B(g10590), .Z(g14193) ) ;
AND2    gate11821  (.A(g869), .B(g10632), .Z(g14202) ) ;
AND2    gate11822  (.A(g8655), .B(g11790), .Z(g14206) ) ;
AND2    gate11823  (.A(g8639), .B(g11793), .Z(g14207) ) ;
AND2    gate11824  (.A(g4392), .B(g10590), .Z(g14210) ) ;
AND2    gate11825  (.A(g7631), .B(g10608), .Z(g14216) ) ;
AND2    gate11826  (.A(g875), .B(g10632), .Z(g14218) ) ;
AND2    gate11827  (.A(g8612), .B(g11820), .Z(g14220) ) ;
AND2    gate11828  (.A(g8686), .B(g11823), .Z(g14221) ) ;
AND2    gate11829  (.A(g8655), .B(g11826), .Z(g14222) ) ;
AND2    gate11830  (.A(g8639), .B(g11855), .Z(g14233) ) ;
AND2    gate11831  (.A(g2079), .B(g11872), .Z(g14256) ) ;
AND2    gate11832  (.A(g8612), .B(g11878), .Z(g14257) ) ;
AND2    gate11833  (.A(g4507), .B(g10738), .Z(g14261) ) ;
AND2    gate11834  (.A(g1811), .B(g11894), .Z(g14295) ) ;
AND2    gate11835  (.A(g2638), .B(g11897), .Z(g14296) ) ;
AND2    gate11836  (.A(g2370), .B(g11920), .Z(g14316) ) ;
NAND4   gate11837  (.A(g7304), .B(g7661), .C(g979), .D(g1061), .Z(g10726) ) ;
AND2    gate11838  (.A(g1087), .B(g10726), .Z(g14438) ) ;
NAND2   gate11839  (.A(g7512), .B(g5308), .Z(g12341) ) ;
NAND2   gate11840  (.A(g7436), .B(g5283), .Z(g12293) ) ;
AND3    gate11841  (.A(g10124), .B(g12341), .C(g12293), .Z(II16618) ) ;
NAND2   gate11842  (.A(g7393), .B(g5276), .Z(g12411) ) ;
NAND2   gate11843  (.A(g7343), .B(g5320), .Z(g12244) ) ;
NAND2   gate11844  (.A(g7296), .B(g5290), .Z(g12197) ) ;
AND4    gate11845  (.A(g12411), .B(g12244), .C(g12197), .D(II16618), .Z(g14496) ) ;
NAND4   gate11846  (.A(g7352), .B(g7675), .C(g1322), .D(g1404), .Z(g10755) ) ;
AND2    gate11847  (.A(g1430), .B(g10755), .Z(g14506) ) ;
NAND2   gate11848  (.A(g7521), .B(g5654), .Z(g12413) ) ;
NAND2   gate11849  (.A(g7470), .B(g5630), .Z(g12343) ) ;
AND3    gate11850  (.A(g10160), .B(g12413), .C(g12343), .Z(II16646) ) ;
NAND2   gate11851  (.A(g7437), .B(g5623), .Z(g12459) ) ;
NAND2   gate11852  (.A(g7394), .B(g5666), .Z(g12306) ) ;
NAND2   gate11853  (.A(g7344), .B(g5637), .Z(g12245) ) ;
AND4    gate11854  (.A(g12459), .B(g12306), .C(g12245), .D(II16646), .Z(g14528) ) ;
NAND2   gate11855  (.A(g7268), .B(g7308), .Z(g10550) ) ;
NAND2   gate11856  (.A(g1592), .B(g7308), .Z(g10529) ) ;
AND2    gate11857  (.A(g10550), .B(g10529), .Z(g14537) ) ;
NAND2   gate11858  (.A(g7536), .B(g6000), .Z(g12461) ) ;
NAND2   gate11859  (.A(g7496), .B(g5976), .Z(g12415) ) ;
AND3    gate11860  (.A(g10185), .B(g12461), .C(g12415), .Z(II16671) ) ;
NAND2   gate11861  (.A(g7471), .B(g5969), .Z(g12521) ) ;
NAND2   gate11862  (.A(g7438), .B(g6012), .Z(g12356) ) ;
NAND2   gate11863  (.A(g7395), .B(g5983), .Z(g12307) ) ;
AND4    gate11864  (.A(g12521), .B(g12356), .C(g12307), .D(II16671), .Z(g14555) ) ;
NAND2   gate11865  (.A(g8139), .B(g8187), .Z(g11934) ) ;
NAND2   gate11866  (.A(g1624), .B(g8187), .Z(g11952) ) ;
AND2    gate11867  (.A(g11934), .B(g11952), .Z(g14565) ) ;
NAND2   gate11868  (.A(g7315), .B(g7356), .Z(g10566) ) ;
NAND2   gate11869  (.A(g1728), .B(g7356), .Z(g10551) ) ;
AND2    gate11870  (.A(g10566), .B(g10551), .Z(g14566) ) ;
NAND2   gate11871  (.A(g7328), .B(g7374), .Z(g10568) ) ;
NAND2   gate11872  (.A(g2153), .B(g7374), .Z(g10552) ) ;
AND2    gate11873  (.A(g10568), .B(g10552), .Z(g14567) ) ;
NAND2   gate11874  (.A(g7563), .B(g6346), .Z(g12523) ) ;
NAND2   gate11875  (.A(g7513), .B(g6322), .Z(g12463) ) ;
AND3    gate11876  (.A(g10207), .B(g12523), .C(g12463), .Z(II16695) ) ;
NAND2   gate11877  (.A(g7497), .B(g6315), .Z(g12587) ) ;
NAND2   gate11878  (.A(g7472), .B(g6358), .Z(g12428) ) ;
NAND2   gate11879  (.A(g7439), .B(g6329), .Z(g12357) ) ;
AND4    gate11880  (.A(g12587), .B(g12428), .C(g12357), .D(II16695), .Z(g14581) ) ;
AND2    gate11881  (.A(g1141), .B(g10905), .Z(g14585) ) ;
NAND2   gate11882  (.A(g8195), .B(g8241), .Z(g11953) ) ;
NAND2   gate11883  (.A(g1760), .B(g8241), .Z(g11970) ) ;
AND2    gate11884  (.A(g11953), .B(g11970), .Z(g14586) ) ;
NAND2   gate11885  (.A(g7362), .B(g7405), .Z(g10584) ) ;
NAND2   gate11886  (.A(g1862), .B(g7405), .Z(g10567) ) ;
AND2    gate11887  (.A(g10584), .B(g10567), .Z(g14587) ) ;
NAND2   gate11888  (.A(g8205), .B(g8259), .Z(g11957) ) ;
NAND2   gate11889  (.A(g2185), .B(g8259), .Z(g11974) ) ;
AND2    gate11890  (.A(g11957), .B(g11974), .Z(g14588) ) ;
NAND2   gate11891  (.A(g7380), .B(g7418), .Z(g10586) ) ;
NAND2   gate11892  (.A(g2287), .B(g7418), .Z(g10569) ) ;
AND2    gate11893  (.A(g10586), .B(g10569), .Z(g14589) ) ;
NAND2   gate11894  (.A(g7591), .B(g6692), .Z(g12589) ) ;
NAND2   gate11895  (.A(g7522), .B(g6668), .Z(g12525) ) ;
AND3    gate11896  (.A(g10224), .B(g12589), .C(g12525), .Z(II16721) ) ;
NAND2   gate11897  (.A(g7514), .B(g6661), .Z(g12638) ) ;
NAND2   gate11898  (.A(g7498), .B(g6704), .Z(g12476) ) ;
NAND2   gate11899  (.A(g7473), .B(g6675), .Z(g12429) ) ;
AND4    gate11900  (.A(g12638), .B(g12476), .C(g12429), .D(II16721), .Z(g14608) ) ;
AND2    gate11901  (.A(g1484), .B(g10935), .Z(g14610) ) ;
NAND2   gate11902  (.A(g8249), .B(g8302), .Z(g11971) ) ;
NAND2   gate11903  (.A(g1894), .B(g8302), .Z(g11993) ) ;
AND2    gate11904  (.A(g11971), .B(g11993), .Z(g14612) ) ;
NAND2   gate11905  (.A(g7411), .B(g7451), .Z(g10602) ) ;
NAND2   gate11906  (.A(g1996), .B(g7451), .Z(g10585) ) ;
AND2    gate11907  (.A(g10602), .B(g10585), .Z(g14613) ) ;
NAND2   gate11908  (.A(g8267), .B(g8316), .Z(g11975) ) ;
NAND2   gate11909  (.A(g2319), .B(g8316), .Z(g11997) ) ;
AND2    gate11910  (.A(g11975), .B(g11997), .Z(g14614) ) ;
NAND2   gate11911  (.A(g7424), .B(g7456), .Z(g10604) ) ;
NAND2   gate11912  (.A(g2421), .B(g7456), .Z(g10587) ) ;
AND2    gate11913  (.A(g10604), .B(g10587), .Z(g14615) ) ;
NAND2   gate11914  (.A(g8310), .B(g8365), .Z(g11994) ) ;
NAND2   gate11915  (.A(g2028), .B(g8365), .Z(g12020) ) ;
AND2    gate11916  (.A(g11994), .B(g12020), .Z(g14641) ) ;
NAND2   gate11917  (.A(g8324), .B(g8373), .Z(g11998) ) ;
NAND2   gate11918  (.A(g2453), .B(g8373), .Z(g12023) ) ;
AND2    gate11919  (.A(g11998), .B(g12023), .Z(g14643) ) ;
NAND2   gate11920  (.A(g7462), .B(g7490), .Z(g10610) ) ;
NAND2   gate11921  (.A(g2555), .B(g7490), .Z(g10605) ) ;
AND2    gate11922  (.A(g10610), .B(g10605), .Z(g14644) ) ;
AND2    gate11923  (.A(g7178), .B(g10476), .Z(g14654) ) ;
NAND2   gate11924  (.A(g8381), .B(g8418), .Z(g12024) ) ;
NAND2   gate11925  (.A(g2587), .B(g8418), .Z(g12053) ) ;
AND2    gate11926  (.A(g12024), .B(g12053), .Z(g14680) ) ;
AND2    gate11927  (.A(g4392), .B(g10476), .Z(g14681) ) ;
NAND2   gate11928  (.A(g9049), .B(g637), .Z(g12369) ) ;
AND2    gate11929  (.A(g4392), .B(g10830), .Z(g14719) ) ;
AND2    gate11930  (.A(g1146), .B(g10909), .Z(g14791) ) ;
AND2    gate11931  (.A(g1152), .B(g10909), .Z(g14831) ) ;
AND2    gate11932  (.A(g1489), .B(g10939), .Z(g14832) ) ;
AND2    gate11933  (.A(g1099), .B(g10909), .Z(g14874) ) ;
AND2    gate11934  (.A(g1495), .B(g10939), .Z(g14875) ) ;
AND2    gate11935  (.A(g1442), .B(g10939), .Z(g14913) ) ;
NOR2    gate11936  (.A(g10430), .B(g6845), .Z(g12850) ) ;
AND2    gate11937  (.A(g12850), .B(g12955), .Z(g15075) ) ;
AND2    gate11938  (.A(g2130), .B(g12955), .Z(g15076) ) ;
AND2    gate11939  (.A(g2138), .B(g12955), .Z(g15077) ) ;
NOR2    gate11940  (.A(g10430), .B(g6854), .Z(g12855) ) ;
AND2    gate11941  (.A(g12855), .B(g12983), .Z(g15080) ) ;
AND2    gate11942  (.A(g2689), .B(g12983), .Z(g15081) ) ;
AND2    gate11943  (.A(g2697), .B(g12983), .Z(g15082) ) ;
AND2    gate11944  (.A(g4180), .B(g14454), .Z(g15103) ) ;
AND2    gate11945  (.A(g6955), .B(g14454), .Z(g15104) ) ;
AND2    gate11946  (.A(g4235), .B(g14454), .Z(g15105) ) ;
AND2    gate11947  (.A(g4258), .B(g14454), .Z(g15107) ) ;
AND2    gate11948  (.A(g4264), .B(g14454), .Z(g15108) ) ;
AND2    gate11949  (.A(g4269), .B(g14454), .Z(g15109) ) ;
AND2    gate11950  (.A(g4245), .B(g14454), .Z(g15110) ) ;
AND2    gate11951  (.A(g4281), .B(g14454), .Z(g15111) ) ;
AND2    gate11952  (.A(g4284), .B(g14454), .Z(g15112) ) ;
AND2    gate11953  (.A(g4291), .B(g14454), .Z(g15113) ) ;
AND2    gate11954  (.A(g4239), .B(g14454), .Z(g15114) ) ;
AND2    gate11955  (.A(g2946), .B(g14454), .Z(g15115) ) ;
AND2    gate11956  (.A(g4297), .B(g14454), .Z(g15116) ) ;
AND2    gate11957  (.A(g4300), .B(g14454), .Z(g15117) ) ;
AND2    gate11958  (.A(g4253), .B(g14454), .Z(g15118) ) ;
AND2    gate11959  (.A(g4249), .B(g14454), .Z(g15119) ) ;
AND2    gate11960  (.A(g10970), .B(g13305), .Z(g15507) ) ;
AND2    gate11961  (.A(g392), .B(g13312), .Z(g15567) ) ;
AND2    gate11962  (.A(g411), .B(g13334), .Z(g15589) ) ;
AND2    gate11963  (.A(g3139), .B(g13530), .Z(g15590) ) ;
AND2    gate11964  (.A(g471), .B(g13437), .Z(g15611) ) ;
AND2    gate11965  (.A(g3143), .B(g13530), .Z(g15612) ) ;
AND2    gate11966  (.A(g3490), .B(g13555), .Z(g15613) ) ;
AND2    gate11967  (.A(g168), .B(g13437), .Z(g15631) ) ;
AND2    gate11968  (.A(g3494), .B(g13555), .Z(g15632) ) ;
AND2    gate11969  (.A(g3841), .B(g13584), .Z(g15633) ) ;
AND2    gate11970  (.A(g8362), .B(g13413), .Z(g15650) ) ;
AND2    gate11971  (.A(g429), .B(g13414), .Z(g15651) ) ;
AND2    gate11972  (.A(g174), .B(g13437), .Z(g15652) ) ;
AND2    gate11973  (.A(g3119), .B(g13530), .Z(g15653) ) ;
AND2    gate11974  (.A(g3845), .B(g13584), .Z(g15654) ) ;
AND2    gate11975  (.A(g433), .B(g13458), .Z(g15672) ) ;
AND2    gate11976  (.A(g182), .B(g13437), .Z(g15673) ) ;
AND2    gate11977  (.A(g1094), .B(g13846), .Z(g15678) ) ;
AND2    gate11978  (.A(g3470), .B(g13555), .Z(g15679) ) ;
AND2    gate11979  (.A(g269), .B(g13474), .Z(g15693) ) ;
AND2    gate11980  (.A(g457), .B(g13437), .Z(g15694) ) ;
AND2    gate11981  (.A(g1437), .B(g13861), .Z(g15699) ) ;
AND2    gate11982  (.A(g3089), .B(g13483), .Z(g15700) ) ;
AND2    gate11983  (.A(g3821), .B(g13584), .Z(g15701) ) ;
AND2    gate11984  (.A(g452), .B(g13437), .Z(g15703) ) ;
AND2    gate11985  (.A(g3440), .B(g13504), .Z(g15704) ) ;
OR2     gate11986  (.A(g10626), .B(g10657), .Z(g13296) ) ;
AND2    gate11987  (.A(g4082), .B(g13506), .Z(g15707) ) ;
AND2    gate11988  (.A(g460), .B(g13437), .Z(g15711) ) ;
AND2    gate11989  (.A(g3791), .B(g13521), .Z(g15712) ) ;
AND2    gate11990  (.A(g468), .B(g13437), .Z(g15716) ) ;
AND2    gate11991  (.A(g464), .B(g13437), .Z(g15722) ) ;
AND2    gate11992  (.A(g1111), .B(g13260), .Z(g15738) ) ;
AND2    gate11993  (.A(g686), .B(g13223), .Z(g15745) ) ;
AND2    gate11994  (.A(g1454), .B(g13273), .Z(g15749) ) ;
AND2    gate11995  (.A(g3207), .B(g14066), .Z(g15757) ) ;
NAND4   gate11996  (.A(g11396), .B(g8847), .C(g11674), .D(g8803), .Z(g13909) ) ;
AND2    gate11997  (.A(g13909), .B(g11214), .Z(g15779) ) ;
AND2    gate11998  (.A(g3215), .B(g14098), .Z(g15783) ) ;
AND2    gate11999  (.A(g3235), .B(g13977), .Z(g15784) ) ;
AND2    gate12000  (.A(g3558), .B(g14107), .Z(g15785) ) ;
NAND4   gate12001  (.A(g11426), .B(g8889), .C(g11707), .D(g8829), .Z(g13940) ) ;
AND2    gate12002  (.A(g13940), .B(g11233), .Z(g15786) ) ;
AND2    gate12003  (.A(g3219), .B(g13873), .Z(g15793) ) ;
AND2    gate12004  (.A(g3239), .B(g14008), .Z(g15794) ) ;
AND2    gate12005  (.A(g3566), .B(g14130), .Z(g15795) ) ;
AND2    gate12006  (.A(g3586), .B(g14015), .Z(g15796) ) ;
AND2    gate12007  (.A(g3909), .B(g14139), .Z(g15797) ) ;
AND2    gate12008  (.A(g3223), .B(g13889), .Z(g15804) ) ;
AND2    gate12009  (.A(g3243), .B(g14041), .Z(g15805) ) ;
AND2    gate12010  (.A(g3570), .B(g13898), .Z(g15807) ) ;
AND2    gate12011  (.A(g3590), .B(g14048), .Z(g15808) ) ;
AND2    gate12012  (.A(g3917), .B(g14154), .Z(g15809) ) ;
AND2    gate12013  (.A(g3937), .B(g14055), .Z(g15810) ) ;
AND2    gate12014  (.A(g3227), .B(g13915), .Z(g15812) ) ;
AND2    gate12015  (.A(g3247), .B(g14069), .Z(g15813) ) ;
AND2    gate12016  (.A(g3574), .B(g13920), .Z(g15814) ) ;
AND2    gate12017  (.A(g3594), .B(g14075), .Z(g15815) ) ;
AND2    gate12018  (.A(g3921), .B(g13929), .Z(g15817) ) ;
AND2    gate12019  (.A(g3941), .B(g14082), .Z(g15818) ) ;
AND2    gate12020  (.A(g3251), .B(g14101), .Z(g15819) ) ;
AND2    gate12021  (.A(g3578), .B(g13955), .Z(g15820) ) ;
AND2    gate12022  (.A(g3598), .B(g14110), .Z(g15821) ) ;
AND2    gate12023  (.A(g3925), .B(g13960), .Z(g15822) ) ;
AND2    gate12024  (.A(g3945), .B(g14116), .Z(g15823) ) ;
AND2    gate12025  (.A(g3187), .B(g14104), .Z(g15836) ) ;
AND2    gate12026  (.A(g3255), .B(g14127), .Z(g15837) ) ;
AND2    gate12027  (.A(g3602), .B(g14133), .Z(g15838) ) ;
AND2    gate12028  (.A(g3929), .B(g13990), .Z(g15839) ) ;
AND2    gate12029  (.A(g3949), .B(g14142), .Z(g15840) ) ;
AND2    gate12030  (.A(g4273), .B(g13868), .Z(g15841) ) ;
AND2    gate12031  (.A(g3191), .B(g14005), .Z(g15847) ) ;
AND2    gate12032  (.A(g3259), .B(g13892), .Z(g15848) ) ;
AND2    gate12033  (.A(g3538), .B(g14136), .Z(g15849) ) ;
AND2    gate12034  (.A(g3606), .B(g14151), .Z(g15850) ) ;
AND2    gate12035  (.A(g3953), .B(g14157), .Z(g15851) ) ;
OR3     gate12036  (.A(g11184), .B(g9187), .C(g12527), .Z(g13820) ) ;
AND2    gate12037  (.A(g13820), .B(g13223), .Z(g15852) ) ;
AND2    gate12038  (.A(g9056), .B(g14223), .Z(g15856) ) ;
AND2    gate12039  (.A(g3199), .B(g14038), .Z(g15857) ) ;
AND2    gate12040  (.A(g3542), .B(g14045), .Z(g15858) ) ;
AND2    gate12041  (.A(g3610), .B(g13923), .Z(g15859) ) ;
AND2    gate12042  (.A(g3889), .B(g14160), .Z(g15860) ) ;
AND2    gate12043  (.A(g3957), .B(g14170), .Z(g15861) ) ;
OR2     gate12044  (.A(g499), .B(g12527), .Z(g13762) ) ;
AND2    gate12045  (.A(g13762), .B(g13223), .Z(g15863) ) ;
AND2    gate12046  (.A(g3231), .B(g13948), .Z(g15870) ) ;
AND2    gate12047  (.A(g3203), .B(g13951), .Z(g15871) ) ;
AND2    gate12048  (.A(g9095), .B(g14234), .Z(g15872) ) ;
AND2    gate12049  (.A(g3550), .B(g14072), .Z(g15873) ) ;
AND2    gate12050  (.A(g3893), .B(g14079), .Z(g15874) ) ;
AND2    gate12051  (.A(g3961), .B(g13963), .Z(g15875) ) ;
NOR2    gate12052  (.A(g9077), .B(g12527), .Z(g13512) ) ;
AND2    gate12053  (.A(g13512), .B(g13223), .Z(g15876) ) ;
AND2    gate12054  (.A(g3211), .B(g13980), .Z(g15880) ) ;
AND2    gate12055  (.A(g3582), .B(g13983), .Z(g15881) ) ;
AND2    gate12056  (.A(g3554), .B(g13986), .Z(g15882) ) ;
AND2    gate12057  (.A(g9180), .B(g14258), .Z(g15883) ) ;
AND2    gate12058  (.A(g3901), .B(g14113), .Z(g15884) ) ;
AND2    gate12059  (.A(g441), .B(g13975), .Z(g15902) ) ;
NOR2    gate12060  (.A(g9158), .B(g12527), .Z(g13796) ) ;
AND2    gate12061  (.A(g13796), .B(g13223), .Z(g15903) ) ;
AND2    gate12062  (.A(g3111), .B(g13530), .Z(g15911) ) ;
AND2    gate12063  (.A(g3562), .B(g14018), .Z(g15912) ) ;
AND2    gate12064  (.A(g3933), .B(g14021), .Z(g15913) ) ;
AND2    gate12065  (.A(g3905), .B(g14024), .Z(g15914) ) ;
AND2    gate12066  (.A(g475), .B(g13999), .Z(g15936) ) ;
NOR2    gate12067  (.A(g9220), .B(g9166), .Z(g11950) ) ;
AND2    gate12068  (.A(g11950), .B(g14387), .Z(g15937) ) ;
AND2    gate12069  (.A(g3462), .B(g13555), .Z(g15966) ) ;
AND2    gate12070  (.A(g3913), .B(g14058), .Z(g15967) ) ;
AND2    gate12071  (.A(g246), .B(g14032), .Z(g15978) ) ;
NOR2    gate12072  (.A(g8462), .B(g1171), .Z(g10666) ) ;
AND2    gate12073  (.A(g3813), .B(g13584), .Z(g16023) ) ;
AND2    gate12074  (.A(g446), .B(g14063), .Z(g16025) ) ;
AND2    gate12075  (.A(g854), .B(g14065), .Z(g16026) ) ;
NOR2    gate12076  (.A(g8526), .B(g1514), .Z(g10699) ) ;
AND2    gate12077  (.A(g5148), .B(g14238), .Z(g16098) ) ;
AND2    gate12078  (.A(g9491), .B(g14291), .Z(g16122) ) ;
AND2    gate12079  (.A(g5152), .B(g14238), .Z(g16125) ) ;
AND2    gate12080  (.A(g5495), .B(g14262), .Z(g16126) ) ;
NAND4   gate12081  (.A(g12042), .B(g12014), .C(g11990), .D(g11892), .Z(g14333) ) ;
AND2    gate12082  (.A(g14333), .B(g14166), .Z(g16128) ) ;
AND2    gate12083  (.A(g5499), .B(g14262), .Z(g16160) ) ;
AND2    gate12084  (.A(g5841), .B(g14297), .Z(g16161) ) ;
NAND3   gate12085  (.A(g11968), .B(g11933), .C(g11951), .Z(g14254) ) ;
AND2    gate12086  (.A(g14254), .B(g14179), .Z(g16163) ) ;
NAND4   gate12087  (.A(g12196), .B(g9775), .C(g12124), .D(g9663), .Z(g14596) ) ;
AND2    gate12088  (.A(g14596), .B(g11779), .Z(g16176) ) ;
AND2    gate12089  (.A(g5128), .B(g14238), .Z(g16177) ) ;
AND2    gate12090  (.A(g5845), .B(g14297), .Z(g16178) ) ;
AND2    gate12091  (.A(g6187), .B(g14321), .Z(g16179) ) ;
AND2    gate12092  (.A(g9285), .B(g14183), .Z(g16184) ) ;
AND2    gate12093  (.A(g3263), .B(g14011), .Z(g16185) ) ;
NAND4   gate12094  (.A(g12232), .B(g9852), .C(g12159), .D(g9715), .Z(g14626) ) ;
AND2    gate12095  (.A(g14626), .B(g11810), .Z(g16190) ) ;
AND2    gate12096  (.A(g5475), .B(g14262), .Z(g16191) ) ;
AND2    gate12097  (.A(g6191), .B(g14321), .Z(g16192) ) ;
AND2    gate12098  (.A(g6533), .B(g14348), .Z(g16193) ) ;
AND3    gate12099  (.A(g13156), .B(g11450), .C(g6756), .Z(II17529) ) ;
AND2    gate12100  (.A(g3614), .B(g14051), .Z(g16199) ) ;
AND2    gate12101  (.A(g86), .B(g14197), .Z(g16202) ) ;
AND2    gate12102  (.A(g5821), .B(g14297), .Z(g16203) ) ;
AND2    gate12103  (.A(g6537), .B(g14348), .Z(g16204) ) ;
AND3    gate12104  (.A(g13156), .B(g6767), .C(g6756), .Z(II17542) ) ;
AND2    gate12105  (.A(g9839), .B(g14204), .Z(g16207) ) ;
AND2    gate12106  (.A(g3965), .B(g14085), .Z(g16208) ) ;
AND2    gate12107  (.A(g5445), .B(g14215), .Z(g16211) ) ;
AND2    gate12108  (.A(g6167), .B(g14321), .Z(g16212) ) ;
AND3    gate12109  (.A(g13156), .B(g11450), .C(g11498), .Z(II17552) ) ;
AND2    gate12110  (.A(g5791), .B(g14231), .Z(g16221) ) ;
AND2    gate12111  (.A(g6513), .B(g14348), .Z(g16222) ) ;
OR2     gate12112  (.A(g10685), .B(g542), .Z(g14583) ) ;
AND2    gate12113  (.A(g6137), .B(g14251), .Z(g16233) ) ;
AND3    gate12114  (.A(g13156), .B(g11450), .C(g6756), .Z(II17575) ) ;
AND2    gate12115  (.A(g6483), .B(g14275), .Z(g16243) ) ;
NOR3    gate12116  (.A(g10816), .B(g10812), .C(g10805), .Z(g14988) ) ;
AND3    gate12117  (.A(g14988), .B(g11450), .C(g11498), .Z(II17585) ) ;
NOR3    gate12118  (.A(g562), .B(g12259), .C(g9217), .Z(g14278) ) ;
AND2    gate12119  (.A(g14278), .B(g14708), .Z(g16245) ) ;
AND2    gate12120  (.A(g4512), .B(g14424), .Z(g16279) ) ;
AND3    gate12121  (.A(g14988), .B(g11450), .C(g6756), .Z(II17606) ) ;
AND2    gate12122  (.A(g4527), .B(g12921), .Z(g16303) ) ;
OR2     gate12123  (.A(g7251), .B(g10616), .Z(g13657) ) ;
AND2    gate12124  (.A(g13657), .B(g182), .Z(g16324) ) ;
NAND2   gate12125  (.A(g11172), .B(g8388), .Z(g13627) ) ;
AND2    gate12126  (.A(g8216), .B(g13627), .Z(g16422) ) ;
AND2    gate12127  (.A(g5216), .B(g14876), .Z(g16427) ) ;
NAND2   gate12128  (.A(g11190), .B(g8441), .Z(g13666) ) ;
AND2    gate12129  (.A(g8280), .B(g13666), .Z(g16474) ) ;
AND2    gate12130  (.A(g5224), .B(g14915), .Z(g16483) ) ;
AND2    gate12131  (.A(g5244), .B(g14755), .Z(g16484) ) ;
AND2    gate12132  (.A(g5563), .B(g14924), .Z(g16485) ) ;
AND3    gate12133  (.A(g14988), .B(g11450), .C(g6756), .Z(II17692) ) ;
NAND2   gate12134  (.A(g11200), .B(g8507), .Z(g13708) ) ;
AND2    gate12135  (.A(g8345), .B(g13708), .Z(g16513) ) ;
AND2    gate12136  (.A(g5228), .B(g14627), .Z(g16516) ) ;
AND2    gate12137  (.A(g5248), .B(g14797), .Z(g16517) ) ;
AND2    gate12138  (.A(g5571), .B(g14956), .Z(g16518) ) ;
AND2    gate12139  (.A(g5591), .B(g14804), .Z(g16519) ) ;
AND2    gate12140  (.A(g5909), .B(g14965), .Z(g16520) ) ;
AND2    gate12141  (.A(g5232), .B(g14656), .Z(g16531) ) ;
AND2    gate12142  (.A(g5252), .B(g14841), .Z(g16532) ) ;
AND2    gate12143  (.A(g5575), .B(g14665), .Z(g16534) ) ;
AND2    gate12144  (.A(g5595), .B(g14848), .Z(g16535) ) ;
AND2    gate12145  (.A(g5917), .B(g14996), .Z(g16536) ) ;
AND2    gate12146  (.A(g5937), .B(g14855), .Z(g16537) ) ;
AND2    gate12147  (.A(g6255), .B(g15005), .Z(g16538) ) ;
AND3    gate12148  (.A(g14988), .B(g11450), .C(g11498), .Z(II17741) ) ;
AND2    gate12149  (.A(g5236), .B(g14683), .Z(g16590) ) ;
AND2    gate12150  (.A(g5256), .B(g14879), .Z(g16591) ) ;
AND2    gate12151  (.A(g5579), .B(g14688), .Z(g16592) ) ;
AND2    gate12152  (.A(g5599), .B(g14885), .Z(g16593) ) ;
AND2    gate12153  (.A(g5921), .B(g14697), .Z(g16595) ) ;
AND2    gate12154  (.A(g5941), .B(g14892), .Z(g16596) ) ;
AND2    gate12155  (.A(g6263), .B(g15021), .Z(g16597) ) ;
AND2    gate12156  (.A(g6283), .B(g14899), .Z(g16598) ) ;
AND2    gate12157  (.A(g6601), .B(g15030), .Z(g16599) ) ;
AND2    gate12158  (.A(g5260), .B(g14918), .Z(g16610) ) ;
AND2    gate12159  (.A(g5583), .B(g14727), .Z(g16611) ) ;
AND2    gate12160  (.A(g5603), .B(g14927), .Z(g16612) ) ;
AND2    gate12161  (.A(g5925), .B(g14732), .Z(g16613) ) ;
AND2    gate12162  (.A(g5945), .B(g14933), .Z(g16614) ) ;
AND2    gate12163  (.A(g6267), .B(g14741), .Z(g16616) ) ;
AND2    gate12164  (.A(g6287), .B(g14940), .Z(g16617) ) ;
AND2    gate12165  (.A(g6609), .B(g15039), .Z(g16618) ) ;
AND2    gate12166  (.A(g6629), .B(g14947), .Z(g16619) ) ;
NAND2   gate12167  (.A(g11251), .B(g8340), .Z(g13821) ) ;
AND2    gate12168  (.A(g8278), .B(g13821), .Z(g16621) ) ;
AND2    gate12169  (.A(g5196), .B(g14921), .Z(g16633) ) ;
AND2    gate12170  (.A(g5264), .B(g14953), .Z(g16634) ) ;
AND2    gate12171  (.A(g5607), .B(g14959), .Z(g16635) ) ;
AND2    gate12172  (.A(g5929), .B(g14768), .Z(g16636) ) ;
AND2    gate12173  (.A(g5949), .B(g14968), .Z(g16637) ) ;
AND2    gate12174  (.A(g6271), .B(g14773), .Z(g16638) ) ;
AND2    gate12175  (.A(g6291), .B(g14974), .Z(g16639) ) ;
AND2    gate12176  (.A(g6613), .B(g14782), .Z(g16641) ) ;
AND2    gate12177  (.A(g6633), .B(g14981), .Z(g16642) ) ;
NAND2   gate12178  (.A(g11279), .B(g8396), .Z(g13850) ) ;
AND2    gate12179  (.A(g8343), .B(g13850), .Z(g16653) ) ;
AND2    gate12180  (.A(g4552), .B(g14753), .Z(g16662) ) ;
AND2    gate12181  (.A(g5200), .B(g14794), .Z(g16666) ) ;
AND2    gate12182  (.A(g5268), .B(g14659), .Z(g16667) ) ;
AND2    gate12183  (.A(g5543), .B(g14962), .Z(g16668) ) ;
AND2    gate12184  (.A(g5611), .B(g14993), .Z(g16669) ) ;
AND2    gate12185  (.A(g5953), .B(g14999), .Z(g16670) ) ;
AND2    gate12186  (.A(g6275), .B(g14817), .Z(g16671) ) ;
AND2    gate12187  (.A(g6295), .B(g15008), .Z(g16672) ) ;
AND2    gate12188  (.A(g6617), .B(g14822), .Z(g16673) ) ;
AND2    gate12189  (.A(g6637), .B(g15014), .Z(g16674) ) ;
NAND2   gate12190  (.A(g11312), .B(g8449), .Z(g13867) ) ;
AND2    gate12191  (.A(g8399), .B(g13867), .Z(g16690) ) ;
AND2    gate12192  (.A(g7134), .B(g12933), .Z(g16699) ) ;
AND2    gate12193  (.A(g5208), .B(g14838), .Z(g16700) ) ;
AND2    gate12194  (.A(g5547), .B(g14845), .Z(g16701) ) ;
AND2    gate12195  (.A(g5615), .B(g14691), .Z(g16702) ) ;
AND2    gate12196  (.A(g5889), .B(g15002), .Z(g16703) ) ;
AND2    gate12197  (.A(g5957), .B(g15018), .Z(g16704) ) ;
AND2    gate12198  (.A(g6299), .B(g15024), .Z(g16705) ) ;
AND2    gate12199  (.A(g6621), .B(g14868), .Z(g16706) ) ;
AND2    gate12200  (.A(g6641), .B(g15033), .Z(g16707) ) ;
AND2    gate12201  (.A(g5240), .B(g14720), .Z(g16729) ) ;
AND2    gate12202  (.A(g5212), .B(g14723), .Z(g16730) ) ;
AND2    gate12203  (.A(g7153), .B(g12941), .Z(g16731) ) ;
AND2    gate12204  (.A(g5555), .B(g14882), .Z(g16732) ) ;
AND2    gate12205  (.A(g5893), .B(g14889), .Z(g16733) ) ;
AND2    gate12206  (.A(g5961), .B(g14735), .Z(g16734) ) ;
AND2    gate12207  (.A(g6235), .B(g15027), .Z(g16735) ) ;
AND2    gate12208  (.A(g6303), .B(g15036), .Z(g16736) ) ;
AND2    gate12209  (.A(g6645), .B(g15042), .Z(g16737) ) ;
OR2     gate12210  (.A(g11496), .B(g11546), .Z(g13155) ) ;
AND2    gate12211  (.A(g13155), .B(g13065), .Z(g16751) ) ;
AND2    gate12212  (.A(g5220), .B(g14758), .Z(g16758) ) ;
AND2    gate12213  (.A(g5587), .B(g14761), .Z(g16759) ) ;
AND2    gate12214  (.A(g5559), .B(g14764), .Z(g16760) ) ;
AND2    gate12215  (.A(g7170), .B(g12947), .Z(g16761) ) ;
AND2    gate12216  (.A(g5901), .B(g14930), .Z(g16762) ) ;
AND2    gate12217  (.A(g6239), .B(g14937), .Z(g16763) ) ;
AND2    gate12218  (.A(g6307), .B(g14776), .Z(g16764) ) ;
AND2    gate12219  (.A(g6581), .B(g15045), .Z(g16765) ) ;
AND2    gate12220  (.A(g6649), .B(g12915), .Z(g16766) ) ;
AND2    gate12221  (.A(g5120), .B(g14238), .Z(g16801) ) ;
AND2    gate12222  (.A(g5567), .B(g14807), .Z(g16802) ) ;
AND2    gate12223  (.A(g5933), .B(g14810), .Z(g16803) ) ;
AND2    gate12224  (.A(g5905), .B(g14813), .Z(g16804) ) ;
AND2    gate12225  (.A(g7187), .B(g12972), .Z(g16805) ) ;
AND2    gate12226  (.A(g6247), .B(g14971), .Z(g16806) ) ;
AND2    gate12227  (.A(g6585), .B(g14978), .Z(g16807) ) ;
AND2    gate12228  (.A(g6653), .B(g14825), .Z(g16808) ) ;
AND2    gate12229  (.A(g5467), .B(g14262), .Z(g16840) ) ;
AND2    gate12230  (.A(g5913), .B(g14858), .Z(g16841) ) ;
AND2    gate12231  (.A(g6279), .B(g14861), .Z(g16842) ) ;
AND2    gate12232  (.A(g6251), .B(g14864), .Z(g16843) ) ;
AND2    gate12233  (.A(g7212), .B(g13000), .Z(g16844) ) ;
AND2    gate12234  (.A(g6593), .B(g15011), .Z(g16845) ) ;
NOR2    gate12235  (.A(g504), .B(g9040), .Z(g12591) ) ;
NOR3    gate12236  (.A(g8038), .B(g8183), .C(g6804), .Z(g11185) ) ;
AND2    gate12237  (.A(g4392), .B(g13107), .Z(g16855) ) ;
AND2    gate12238  (.A(g5813), .B(g14297), .Z(g16868) ) ;
AND2    gate12239  (.A(g6259), .B(g14902), .Z(g16869) ) ;
AND2    gate12240  (.A(g6625), .B(g14905), .Z(g16870) ) ;
AND2    gate12241  (.A(g6597), .B(g14908), .Z(g16871) ) ;
AND2    gate12242  (.A(g6159), .B(g14321), .Z(g16884) ) ;
AND2    gate12243  (.A(g6605), .B(g14950), .Z(g16885) ) ;
AND2    gate12244  (.A(g262), .B(g13120), .Z(g16896) ) ;
AND2    gate12245  (.A(g6505), .B(g14348), .Z(g16929) ) ;
AND2    gate12246  (.A(g239), .B(g13132), .Z(g16930) ) ;
AND2    gate12247  (.A(g13064), .B(g10418), .Z(g16957) ) ;
AND2    gate12248  (.A(g269), .B(g13140), .Z(g16965) ) ;
AND2    gate12249  (.A(g246), .B(g13142), .Z(g16986) ) ;
AND2    gate12250  (.A(g446), .B(g13173), .Z(g17057) ) ;
AND2    gate12251  (.A(g8659), .B(g12940), .Z(g17091) ) ;
AND2    gate12252  (.A(g5272), .B(g14800), .Z(g17119) ) ;
AND2    gate12253  (.A(g225), .B(g13209), .Z(g17123) ) ;
AND2    gate12254  (.A(g10683), .B(g13222), .Z(g17133) ) ;
AND2    gate12255  (.A(g5619), .B(g14851), .Z(g17134) ) ;
AND2    gate12256  (.A(g255), .B(g13239), .Z(g17138) ) ;
AND2    gate12257  (.A(g8635), .B(g12967), .Z(g17139) ) ;
AND2    gate12258  (.A(g8616), .B(g12968), .Z(g17140) ) ;
AND2    gate12259  (.A(g7469), .B(g13249), .Z(g17145) ) ;
AND2    gate12260  (.A(g5965), .B(g14895), .Z(g17146) ) ;
AND2    gate12261  (.A(g232), .B(g13255), .Z(g17149) ) ;
AND2    gate12262  (.A(g8579), .B(g12995), .Z(g17150) ) ;
AND2    gate12263  (.A(g8659), .B(g12996), .Z(g17151) ) ;
AND2    gate12264  (.A(g8635), .B(g12997), .Z(g17152) ) ;
AND2    gate12265  (.A(g6311), .B(g14943), .Z(g17153) ) ;
AND2    gate12266  (.A(g305), .B(g13385), .Z(g17156) ) ;
AND2    gate12267  (.A(g8616), .B(g13008), .Z(g17176) ) ;
AND2    gate12268  (.A(g6657), .B(g14984), .Z(g17177) ) ;
AND2    gate12269  (.A(g1041), .B(g13211), .Z(g17179) ) ;
AND2    gate12270  (.A(g1945), .B(g13014), .Z(g17181) ) ;
AND2    gate12271  (.A(g8579), .B(g13016), .Z(g17182) ) ;
AND2    gate12272  (.A(g1384), .B(g13242), .Z(g17191) ) ;
AND2    gate12273  (.A(g1677), .B(g13022), .Z(g17192) ) ;
AND2    gate12274  (.A(g2504), .B(g13023), .Z(g17193) ) ;
AND2    gate12275  (.A(g2236), .B(g13034), .Z(g17199) ) ;
NAND4   gate12276  (.A(g10649), .B(g7661), .C(g979), .D(g1061), .Z(g13093) ) ;
NAND2   gate12277  (.A(g11961), .B(g9670), .Z(g14343) ) ;
AND2    gate12278  (.A(g9498), .B(g14343), .Z(g17307) ) ;
NAND4   gate12279  (.A(g10666), .B(g7661), .C(g979), .D(g1061), .Z(g13124) ) ;
AND2    gate12280  (.A(g1079), .B(g13124), .Z(g17317) ) ;
NAND4   gate12281  (.A(g10671), .B(g7675), .C(g1322), .D(g1404), .Z(g13105) ) ;
AND2    gate12282  (.A(g1418), .B(g13105), .Z(g17321) ) ;
AND2    gate12283  (.A(g7650), .B(g13036), .Z(g17365) ) ;
NAND2   gate12284  (.A(g11979), .B(g9731), .Z(g14378) ) ;
AND2    gate12285  (.A(g9556), .B(g14378), .Z(g17391) ) ;
NAND4   gate12286  (.A(g10695), .B(g7661), .C(g979), .D(g1061), .Z(g13143) ) ;
AND2    gate12287  (.A(g1083), .B(g13143), .Z(g17401) ) ;
NAND4   gate12288  (.A(g10699), .B(g7675), .C(g1322), .D(g1404), .Z(g13137) ) ;
AND2    gate12289  (.A(g1422), .B(g13137), .Z(g17405) ) ;
NAND2   gate12290  (.A(g12008), .B(g9807), .Z(g14407) ) ;
AND2    gate12291  (.A(g9618), .B(g14407), .Z(g17418) ) ;
NAND4   gate12292  (.A(g10715), .B(g7675), .C(g1322), .D(g1404), .Z(g13176) ) ;
AND2    gate12293  (.A(g1426), .B(g13176), .Z(g17424) ) ;
AND2    gate12294  (.A(g4076), .B(g13217), .Z(g17469) ) ;
NAND2   gate12295  (.A(g12035), .B(g9890), .Z(g14433) ) ;
AND2    gate12296  (.A(g9683), .B(g14433), .Z(g17480) ) ;
NAND2   gate12297  (.A(g12073), .B(g9961), .Z(g14505) ) ;
AND2    gate12298  (.A(g9744), .B(g14505), .Z(g17506) ) ;
NAND2   gate12299  (.A(g12125), .B(g9613), .Z(g14546) ) ;
AND2    gate12300  (.A(g9554), .B(g14546), .Z(g17574) ) ;
NAND2   gate12301  (.A(g12169), .B(g9678), .Z(g14572) ) ;
AND2    gate12302  (.A(g9616), .B(g14572), .Z(g17601) ) ;
AND3    gate12303  (.A(g13156), .B(g11450), .C(g11498), .Z(II18568) ) ;
NAND2   gate12304  (.A(II12270), .B(II12271), .Z(g7885) ) ;
AND2    gate12305  (.A(g7885), .B(g13326), .Z(g17617) ) ;
AND2    gate12306  (.A(g10829), .B(g13463), .Z(g17636) ) ;
NAND2   gate12307  (.A(g12207), .B(g9739), .Z(g14599) ) ;
AND2    gate12308  (.A(g9681), .B(g14599), .Z(g17643) ) ;
AND3    gate12309  (.A(g13156), .B(g11450), .C(g11498), .Z(II18620) ) ;
AND2    gate12310  (.A(g962), .B(g13284), .Z(g17654) ) ;
NAND2   gate12311  (.A(II12288), .B(II12289), .Z(g7897) ) ;
AND2    gate12312  (.A(g7897), .B(g13342), .Z(g17655) ) ;
AND2    gate12313  (.A(g7685), .B(g13485), .Z(g17671) ) ;
NAND2   gate12314  (.A(g12255), .B(g9815), .Z(g14637) ) ;
AND2    gate12315  (.A(g9742), .B(g14637), .Z(g17682) ) ;
AND3    gate12316  (.A(g13156), .B(g11450), .C(g6756), .Z(II18671) ) ;
AND2    gate12317  (.A(g1124), .B(g13307), .Z(g17692) ) ;
AND2    gate12318  (.A(g1306), .B(g13291), .Z(g17693) ) ;
NAND2   gate12319  (.A(g12317), .B(g9898), .Z(g14675) ) ;
AND2    gate12320  (.A(g9818), .B(g14675), .Z(g17719) ) ;
AND3    gate12321  (.A(g13156), .B(g6767), .C(g6756), .Z(II18713) ) ;
AND3    gate12322  (.A(g13156), .B(g11450), .C(g6756), .Z(II18716) ) ;
AND2    gate12323  (.A(g1467), .B(g13315), .Z(g17726) ) ;
AND3    gate12324  (.A(g13156), .B(g11450), .C(g11498), .Z(II18740) ) ;
AND2    gate12325  (.A(g7841), .B(g13174), .Z(g17752) ) ;
NAND2   gate12326  (.A(g10916), .B(g1099), .Z(g13281) ) ;
AND2    gate12327  (.A(g13281), .B(g13175), .Z(g17753) ) ;
AND3    gate12328  (.A(g13156), .B(g6767), .C(g11498), .Z(II18762) ) ;
AND3    gate12329  (.A(g13156), .B(g11450), .C(g11498), .Z(II18765) ) ;
NOR2    gate12330  (.A(g7841), .B(g10741), .Z(g13325) ) ;
AND2    gate12331  (.A(g13325), .B(g10741), .Z(g17768) ) ;
AND2    gate12332  (.A(g1146), .B(g13188), .Z(g17769) ) ;
AND2    gate12333  (.A(g7863), .B(g13189), .Z(g17770) ) ;
NAND2   gate12334  (.A(g10946), .B(g1442), .Z(g13288) ) ;
AND2    gate12335  (.A(g13288), .B(g13190), .Z(g17771) ) ;
AND3    gate12336  (.A(g13156), .B(g11450), .C(g6756), .Z(II18782) ) ;
AND3    gate12337  (.A(g13156), .B(g6767), .C(g11498), .Z(II18785) ) ;
AND2    gate12338  (.A(g7851), .B(g13110), .Z(g17783) ) ;
AND2    gate12339  (.A(g1152), .B(g13215), .Z(g17784) ) ;
NOR2    gate12340  (.A(g7863), .B(g10762), .Z(g13341) ) ;
AND2    gate12341  (.A(g13341), .B(g10762), .Z(g17785) ) ;
AND2    gate12342  (.A(g1489), .B(g13216), .Z(g17786) ) ;
AND3    gate12343  (.A(g13156), .B(g11450), .C(g6756), .Z(II18803) ) ;
AND2    gate12344  (.A(g7873), .B(g13125), .Z(g17809) ) ;
AND2    gate12345  (.A(g1495), .B(g13246), .Z(g17810) ) ;
AND3    gate12346  (.A(g13156), .B(g11450), .C(g11498), .Z(II18819) ) ;
AND2    gate12347  (.A(g401), .B(g17015), .Z(g18103) ) ;
AND2    gate12348  (.A(g392), .B(g17015), .Z(g18104) ) ;
AND2    gate12349  (.A(g417), .B(g17015), .Z(g18105) ) ;
AND2    gate12350  (.A(g411), .B(g17015), .Z(g18106) ) ;
AND2    gate12351  (.A(g429), .B(g17015), .Z(g18107) ) ;
AND2    gate12352  (.A(g433), .B(g17015), .Z(g18108) ) ;
AND2    gate12353  (.A(g437), .B(g17015), .Z(g18109) ) ;
AND2    gate12354  (.A(g441), .B(g17015), .Z(g18110) ) ;
AND2    gate12355  (.A(g174), .B(g17015), .Z(g18111) ) ;
AND2    gate12356  (.A(g182), .B(g17015), .Z(g18112) ) ;
AND2    gate12357  (.A(g405), .B(g17015), .Z(g18113) ) ;
AND2    gate12358  (.A(g452), .B(g17015), .Z(g18114) ) ;
AND2    gate12359  (.A(g460), .B(g17015), .Z(g18115) ) ;
AND2    gate12360  (.A(g168), .B(g17015), .Z(g18116) ) ;
AND2    gate12361  (.A(g464), .B(g17015), .Z(g18117) ) ;
AND2    gate12362  (.A(g471), .B(g17015), .Z(g18118) ) ;
AND2    gate12363  (.A(g475), .B(g17015), .Z(g18119) ) ;
AND2    gate12364  (.A(g457), .B(g17015), .Z(g18120) ) ;
AND2    gate12365  (.A(g424), .B(g17015), .Z(g18121) ) ;
NOR2    gate12366  (.A(g12835), .B(g13350), .Z(g15052) ) ;
AND2    gate12367  (.A(g15052), .B(g17015), .Z(g18122) ) ;
AND2    gate12368  (.A(g479), .B(g16886), .Z(g18123) ) ;
AND2    gate12369  (.A(g102), .B(g16886), .Z(g18124) ) ;
NOR2    gate12370  (.A(g12836), .B(g13350), .Z(g15053) ) ;
AND2    gate12371  (.A(g15053), .B(g16886), .Z(g18125) ) ;
NOR2    gate12372  (.A(g12837), .B(g13350), .Z(g15054) ) ;
AND2    gate12373  (.A(g15054), .B(g16971), .Z(g18126) ) ;
AND2    gate12374  (.A(g499), .B(g16971), .Z(g18127) ) ;
AND2    gate12375  (.A(g504), .B(g16971), .Z(g18128) ) ;
AND2    gate12376  (.A(g518), .B(g16971), .Z(g18129) ) ;
AND2    gate12377  (.A(g528), .B(g16971), .Z(g18130) ) ;
AND2    gate12378  (.A(g482), .B(g16971), .Z(g18131) ) ;
AND2    gate12379  (.A(g513), .B(g16971), .Z(g18132) ) ;
NOR2    gate12380  (.A(g6808), .B(g13350), .Z(g15055) ) ;
AND2    gate12381  (.A(g15055), .B(g17249), .Z(g18133) ) ;
AND2    gate12382  (.A(g534), .B(g17249), .Z(g18134) ) ;
AND2    gate12383  (.A(g136), .B(g17249), .Z(g18135) ) ;
AND2    gate12384  (.A(g550), .B(g17249), .Z(g18136) ) ;
AND2    gate12385  (.A(g538), .B(g17249), .Z(g18137) ) ;
AND2    gate12386  (.A(g546), .B(g17249), .Z(g18138) ) ;
AND2    gate12387  (.A(g542), .B(g17249), .Z(g18139) ) ;
AND2    gate12388  (.A(g559), .B(g17533), .Z(g18140) ) ;
AND2    gate12389  (.A(g568), .B(g17533), .Z(g18141) ) ;
AND2    gate12390  (.A(g577), .B(g17533), .Z(g18142) ) ;
AND2    gate12391  (.A(g586), .B(g17533), .Z(g18143) ) ;
AND2    gate12392  (.A(g590), .B(g17533), .Z(g18144) ) ;
AND2    gate12393  (.A(g582), .B(g17533), .Z(g18145) ) ;
AND2    gate12394  (.A(g595), .B(g17533), .Z(g18146) ) ;
AND2    gate12395  (.A(g599), .B(g17533), .Z(g18147) ) ;
AND2    gate12396  (.A(g562), .B(g17533), .Z(g18148) ) ;
AND2    gate12397  (.A(g608), .B(g17533), .Z(g18149) ) ;
AND2    gate12398  (.A(g604), .B(g17533), .Z(g18150) ) ;
AND2    gate12399  (.A(g617), .B(g17533), .Z(g18151) ) ;
AND2    gate12400  (.A(g613), .B(g17533), .Z(g18152) ) ;
AND2    gate12401  (.A(g626), .B(g17533), .Z(g18153) ) ;
AND2    gate12402  (.A(g622), .B(g17533), .Z(g18154) ) ;
NOR2    gate12403  (.A(g6809), .B(g13350), .Z(g15056) ) ;
AND2    gate12404  (.A(g15056), .B(g17533), .Z(g18155) ) ;
AND2    gate12405  (.A(g572), .B(g17533), .Z(g18156) ) ;
NOR2    gate12406  (.A(g6810), .B(g13350), .Z(g15057) ) ;
AND2    gate12407  (.A(g15057), .B(g17433), .Z(g18157) ) ;
AND2    gate12408  (.A(g667), .B(g17433), .Z(g18158) ) ;
AND2    gate12409  (.A(g671), .B(g17433), .Z(g18159) ) ;
AND2    gate12410  (.A(g645), .B(g17433), .Z(g18160) ) ;
AND2    gate12411  (.A(g691), .B(g17433), .Z(g18161) ) ;
AND2    gate12412  (.A(g686), .B(g17433), .Z(g18162) ) ;
AND2    gate12413  (.A(g79), .B(g17433), .Z(g18163) ) ;
AND2    gate12414  (.A(g699), .B(g17433), .Z(g18164) ) ;
AND2    gate12415  (.A(g650), .B(g17433), .Z(g18165) ) ;
AND2    gate12416  (.A(g655), .B(g17433), .Z(g18166) ) ;
AND2    gate12417  (.A(g718), .B(g17433), .Z(g18167) ) ;
AND2    gate12418  (.A(g681), .B(g17433), .Z(g18168) ) ;
AND2    gate12419  (.A(g676), .B(g17433), .Z(g18169) ) ;
AND2    gate12420  (.A(g661), .B(g17433), .Z(g18170) ) ;
AND2    gate12421  (.A(g728), .B(g17433), .Z(g18171) ) ;
NOR2    gate12422  (.A(g12838), .B(g13350), .Z(g15058) ) ;
AND2    gate12423  (.A(g15058), .B(g17328), .Z(g18172) ) ;
AND2    gate12424  (.A(g736), .B(g17328), .Z(g18173) ) ;
AND2    gate12425  (.A(g739), .B(g17328), .Z(g18174) ) ;
AND2    gate12426  (.A(g744), .B(g17328), .Z(g18175) ) ;
AND2    gate12427  (.A(g732), .B(g17328), .Z(g18176) ) ;
AND2    gate12428  (.A(g749), .B(g17328), .Z(g18177) ) ;
AND2    gate12429  (.A(g758), .B(g17328), .Z(g18178) ) ;
AND2    gate12430  (.A(g763), .B(g17328), .Z(g18179) ) ;
AND2    gate12431  (.A(g767), .B(g17328), .Z(g18180) ) ;
AND2    gate12432  (.A(g772), .B(g17328), .Z(g18181) ) ;
AND2    gate12433  (.A(g776), .B(g17328), .Z(g18182) ) ;
AND2    gate12434  (.A(g781), .B(g17328), .Z(g18183) ) ;
AND2    gate12435  (.A(g785), .B(g17328), .Z(g18184) ) ;
AND2    gate12436  (.A(g790), .B(g17328), .Z(g18185) ) ;
AND2    gate12437  (.A(g753), .B(g17328), .Z(g18186) ) ;
AND2    gate12438  (.A(g794), .B(g17328), .Z(g18187) ) ;
AND2    gate12439  (.A(g807), .B(g17328), .Z(g18188) ) ;
AND2    gate12440  (.A(g812), .B(g17821), .Z(g18189) ) ;
AND2    gate12441  (.A(g822), .B(g17821), .Z(g18190) ) ;
AND2    gate12442  (.A(g827), .B(g17821), .Z(g18191) ) ;
AND2    gate12443  (.A(g817), .B(g17821), .Z(g18192) ) ;
AND2    gate12444  (.A(g837), .B(g17821), .Z(g18193) ) ;
AND2    gate12445  (.A(g843), .B(g17821), .Z(g18194) ) ;
AND2    gate12446  (.A(g847), .B(g17821), .Z(g18195) ) ;
AND2    gate12447  (.A(g703), .B(g17821), .Z(g18196) ) ;
AND2    gate12448  (.A(g854), .B(g17821), .Z(g18197) ) ;
NOR2    gate12449  (.A(g12839), .B(g13350), .Z(g15059) ) ;
AND2    gate12450  (.A(g15059), .B(g17821), .Z(g18198) ) ;
AND2    gate12451  (.A(g832), .B(g17821), .Z(g18199) ) ;
NOR2    gate12452  (.A(g6815), .B(g13394), .Z(g15061) ) ;
AND2    gate12453  (.A(g15061), .B(g15938), .Z(g18201) ) ;
AND2    gate12454  (.A(g907), .B(g15938), .Z(g18202) ) ;
AND2    gate12455  (.A(g911), .B(g15938), .Z(g18203) ) ;
AND2    gate12456  (.A(g914), .B(g15938), .Z(g18204) ) ;
AND2    gate12457  (.A(g904), .B(g15938), .Z(g18205) ) ;
AND2    gate12458  (.A(g918), .B(g15938), .Z(g18206) ) ;
AND2    gate12459  (.A(g925), .B(g15938), .Z(g18207) ) ;
AND2    gate12460  (.A(g930), .B(g15938), .Z(g18208) ) ;
AND2    gate12461  (.A(g921), .B(g15938), .Z(g18209) ) ;
AND2    gate12462  (.A(g936), .B(g15938), .Z(g18210) ) ;
NOR2    gate12463  (.A(g6817), .B(g13394), .Z(g15062) ) ;
AND2    gate12464  (.A(g15062), .B(g15979), .Z(g18211) ) ;
AND2    gate12465  (.A(g947), .B(g15979), .Z(g18212) ) ;
AND2    gate12466  (.A(g952), .B(g15979), .Z(g18213) ) ;
AND2    gate12467  (.A(g939), .B(g15979), .Z(g18214) ) ;
NOR2    gate12468  (.A(g6818), .B(g13394), .Z(g15063) ) ;
AND2    gate12469  (.A(g15063), .B(g16100), .Z(g18217) ) ;
AND2    gate12470  (.A(g1008), .B(g16100), .Z(g18218) ) ;
AND2    gate12471  (.A(g969), .B(g16100), .Z(g18219) ) ;
AND2    gate12472  (.A(g1002), .B(g16100), .Z(g18220) ) ;
AND2    gate12473  (.A(g1018), .B(g16100), .Z(g18221) ) ;
AND2    gate12474  (.A(g1024), .B(g16100), .Z(g18222) ) ;
AND2    gate12475  (.A(g1030), .B(g16100), .Z(g18223) ) ;
AND2    gate12476  (.A(g1036), .B(g16100), .Z(g18224) ) ;
AND2    gate12477  (.A(g1041), .B(g16100), .Z(g18225) ) ;
NOR2    gate12478  (.A(g6820), .B(g13394), .Z(g15064) ) ;
AND2    gate12479  (.A(g15064), .B(g16129), .Z(g18226) ) ;
AND2    gate12480  (.A(g1052), .B(g16129), .Z(g18227) ) ;
AND2    gate12481  (.A(g1061), .B(g16129), .Z(g18228) ) ;
AND2    gate12482  (.A(g1099), .B(g16326), .Z(g18229) ) ;
AND2    gate12483  (.A(g1111), .B(g16326), .Z(g18230) ) ;
AND2    gate12484  (.A(g1105), .B(g16326), .Z(g18231) ) ;
AND2    gate12485  (.A(g1124), .B(g16326), .Z(g18232) ) ;
AND2    gate12486  (.A(g1094), .B(g16326), .Z(g18233) ) ;
AND2    gate12487  (.A(g1129), .B(g16326), .Z(g18234) ) ;
AND2    gate12488  (.A(g1141), .B(g16326), .Z(g18235) ) ;
NOR2    gate12489  (.A(g13394), .B(g12840), .Z(g15065) ) ;
AND2    gate12490  (.A(g15065), .B(g16326), .Z(g18236) ) ;
AND2    gate12491  (.A(g1146), .B(g16326), .Z(g18237) ) ;
AND2    gate12492  (.A(g1152), .B(g16326), .Z(g18238) ) ;
AND2    gate12493  (.A(g1135), .B(g16326), .Z(g18239) ) ;
NOR2    gate12494  (.A(g12841), .B(g13394), .Z(g15066) ) ;
AND2    gate12495  (.A(g15066), .B(g16431), .Z(g18240) ) ;
AND2    gate12496  (.A(g1183), .B(g16431), .Z(g18241) ) ;
AND2    gate12497  (.A(g962), .B(g16431), .Z(g18242) ) ;
AND2    gate12498  (.A(g1189), .B(g16431), .Z(g18243) ) ;
AND2    gate12499  (.A(g1171), .B(g16431), .Z(g18244) ) ;
AND2    gate12500  (.A(g1193), .B(g16431), .Z(g18245) ) ;
AND2    gate12501  (.A(g1199), .B(g16431), .Z(g18246) ) ;
AND2    gate12502  (.A(g1178), .B(g16431), .Z(g18247) ) ;
NOR2    gate12503  (.A(g12842), .B(g13394), .Z(g15067) ) ;
AND2    gate12504  (.A(g15067), .B(g16897), .Z(g18248) ) ;
AND2    gate12505  (.A(g1216), .B(g16897), .Z(g18249) ) ;
AND2    gate12506  (.A(g6821), .B(g16897), .Z(g18250) ) ;
AND2    gate12507  (.A(g996), .B(g16897), .Z(g18251) ) ;
AND2    gate12508  (.A(g990), .B(g16897), .Z(g18252) ) ;
AND2    gate12509  (.A(g1211), .B(g16897), .Z(g18253) ) ;
AND2    gate12510  (.A(g1236), .B(g16897), .Z(g18254) ) ;
AND2    gate12511  (.A(g1087), .B(g16897), .Z(g18255) ) ;
AND2    gate12512  (.A(g1242), .B(g16897), .Z(g18256) ) ;
AND2    gate12513  (.A(g1205), .B(g16897), .Z(g18257) ) ;
AND2    gate12514  (.A(g1221), .B(g16897), .Z(g18258) ) ;
NOR2    gate12515  (.A(g6826), .B(g13416), .Z(g15068) ) ;
AND2    gate12516  (.A(g15068), .B(g16000), .Z(g18259) ) ;
AND2    gate12517  (.A(g1252), .B(g16000), .Z(g18260) ) ;
AND2    gate12518  (.A(g1256), .B(g16000), .Z(g18261) ) ;
AND2    gate12519  (.A(g1259), .B(g16000), .Z(g18262) ) ;
AND2    gate12520  (.A(g1249), .B(g16000), .Z(g18263) ) ;
AND2    gate12521  (.A(g1263), .B(g16000), .Z(g18264) ) ;
AND2    gate12522  (.A(g1270), .B(g16000), .Z(g18265) ) ;
AND2    gate12523  (.A(g1274), .B(g16000), .Z(g18266) ) ;
AND2    gate12524  (.A(g1266), .B(g16000), .Z(g18267) ) ;
AND2    gate12525  (.A(g1280), .B(g16000), .Z(g18268) ) ;
NOR2    gate12526  (.A(g6828), .B(g13416), .Z(g15069) ) ;
AND2    gate12527  (.A(g15069), .B(g16031), .Z(g18269) ) ;
AND2    gate12528  (.A(g1291), .B(g16031), .Z(g18270) ) ;
AND2    gate12529  (.A(g1296), .B(g16031), .Z(g18271) ) ;
AND2    gate12530  (.A(g1283), .B(g16031), .Z(g18272) ) ;
NOR2    gate12531  (.A(g6829), .B(g13416), .Z(g15070) ) ;
AND2    gate12532  (.A(g15070), .B(g16136), .Z(g18275) ) ;
AND2    gate12533  (.A(g1351), .B(g16136), .Z(g18276) ) ;
AND2    gate12534  (.A(g1312), .B(g16136), .Z(g18277) ) ;
AND2    gate12535  (.A(g1345), .B(g16136), .Z(g18278) ) ;
AND2    gate12536  (.A(g1361), .B(g16136), .Z(g18279) ) ;
AND2    gate12537  (.A(g1367), .B(g16136), .Z(g18280) ) ;
AND2    gate12538  (.A(g1373), .B(g16136), .Z(g18281) ) ;
AND2    gate12539  (.A(g1379), .B(g16136), .Z(g18282) ) ;
AND2    gate12540  (.A(g1384), .B(g16136), .Z(g18283) ) ;
NOR2    gate12541  (.A(g6831), .B(g13416), .Z(g15071) ) ;
AND2    gate12542  (.A(g15071), .B(g16164), .Z(g18284) ) ;
AND2    gate12543  (.A(g1395), .B(g16164), .Z(g18285) ) ;
AND2    gate12544  (.A(g1404), .B(g16164), .Z(g18286) ) ;
AND2    gate12545  (.A(g1442), .B(g16449), .Z(g18287) ) ;
AND2    gate12546  (.A(g1454), .B(g16449), .Z(g18288) ) ;
AND2    gate12547  (.A(g1448), .B(g16449), .Z(g18289) ) ;
AND2    gate12548  (.A(g1467), .B(g16449), .Z(g18290) ) ;
AND2    gate12549  (.A(g1437), .B(g16449), .Z(g18291) ) ;
AND2    gate12550  (.A(g1472), .B(g16449), .Z(g18292) ) ;
AND2    gate12551  (.A(g1484), .B(g16449), .Z(g18293) ) ;
NOR2    gate12552  (.A(g13416), .B(g12843), .Z(g15072) ) ;
AND2    gate12553  (.A(g15072), .B(g16449), .Z(g18294) ) ;
AND2    gate12554  (.A(g1489), .B(g16449), .Z(g18295) ) ;
AND2    gate12555  (.A(g1495), .B(g16449), .Z(g18296) ) ;
AND2    gate12556  (.A(g1478), .B(g16449), .Z(g18297) ) ;
NOR2    gate12557  (.A(g12844), .B(g13416), .Z(g15073) ) ;
AND2    gate12558  (.A(g15073), .B(g16489), .Z(g18298) ) ;
AND2    gate12559  (.A(g1526), .B(g16489), .Z(g18299) ) ;
AND2    gate12560  (.A(g1306), .B(g16489), .Z(g18300) ) ;
AND2    gate12561  (.A(g1532), .B(g16489), .Z(g18301) ) ;
AND2    gate12562  (.A(g1514), .B(g16489), .Z(g18302) ) ;
AND2    gate12563  (.A(g1536), .B(g16489), .Z(g18303) ) ;
AND2    gate12564  (.A(g1542), .B(g16489), .Z(g18304) ) ;
AND2    gate12565  (.A(g1521), .B(g16489), .Z(g18305) ) ;
NOR2    gate12566  (.A(g12845), .B(g13416), .Z(g15074) ) ;
AND2    gate12567  (.A(g15074), .B(g16931), .Z(g18306) ) ;
AND2    gate12568  (.A(g1559), .B(g16931), .Z(g18307) ) ;
AND2    gate12569  (.A(g6832), .B(g16931), .Z(g18308) ) ;
AND2    gate12570  (.A(g1339), .B(g16931), .Z(g18309) ) ;
AND2    gate12571  (.A(g1333), .B(g16931), .Z(g18310) ) ;
AND2    gate12572  (.A(g1554), .B(g16931), .Z(g18311) ) ;
AND2    gate12573  (.A(g1579), .B(g16931), .Z(g18312) ) ;
AND2    gate12574  (.A(g1430), .B(g16931), .Z(g18313) ) ;
AND2    gate12575  (.A(g1585), .B(g16931), .Z(g18314) ) ;
AND2    gate12576  (.A(g1548), .B(g16931), .Z(g18315) ) ;
AND2    gate12577  (.A(g1564), .B(g16931), .Z(g18316) ) ;
NOR2    gate12578  (.A(g6837), .B(g10430), .Z(g12846) ) ;
AND2    gate12579  (.A(g12846), .B(g17873), .Z(g18317) ) ;
AND2    gate12580  (.A(g1604), .B(g17873), .Z(g18318) ) ;
AND2    gate12581  (.A(g1600), .B(g17873), .Z(g18319) ) ;
AND2    gate12582  (.A(g1616), .B(g17873), .Z(g18320) ) ;
AND2    gate12583  (.A(g1620), .B(g17873), .Z(g18321) ) ;
AND2    gate12584  (.A(g1608), .B(g17873), .Z(g18322) ) ;
AND2    gate12585  (.A(g1632), .B(g17873), .Z(g18323) ) ;
AND2    gate12586  (.A(g1644), .B(g17873), .Z(g18324) ) ;
AND2    gate12587  (.A(g1624), .B(g17873), .Z(g18325) ) ;
AND2    gate12588  (.A(g1664), .B(g17873), .Z(g18326) ) ;
AND2    gate12589  (.A(g1636), .B(g17873), .Z(g18327) ) ;
AND2    gate12590  (.A(g1657), .B(g17873), .Z(g18328) ) ;
AND2    gate12591  (.A(g1612), .B(g17873), .Z(g18329) ) ;
AND2    gate12592  (.A(g1668), .B(g17873), .Z(g18330) ) ;
AND2    gate12593  (.A(g1682), .B(g17873), .Z(g18331) ) ;
AND2    gate12594  (.A(g1677), .B(g17873), .Z(g18332) ) ;
AND2    gate12595  (.A(g1691), .B(g17873), .Z(g18333) ) ;
AND2    gate12596  (.A(g1696), .B(g17873), .Z(g18334) ) ;
AND2    gate12597  (.A(g1687), .B(g17873), .Z(g18335) ) ;
AND2    gate12598  (.A(g1700), .B(g17873), .Z(g18336) ) ;
AND2    gate12599  (.A(g1706), .B(g17873), .Z(g18337) ) ;
AND2    gate12600  (.A(g1710), .B(g17873), .Z(g18338) ) ;
AND2    gate12601  (.A(g1714), .B(g17873), .Z(g18339) ) ;
AND2    gate12602  (.A(g1720), .B(g17873), .Z(g18340) ) ;
AND2    gate12603  (.A(g1648), .B(g17873), .Z(g18341) ) ;
AND2    gate12604  (.A(g1592), .B(g17873), .Z(g18342) ) ;
NOR2    gate12605  (.A(g6838), .B(g10430), .Z(g12847) ) ;
AND2    gate12606  (.A(g12847), .B(g17955), .Z(g18343) ) ;
AND2    gate12607  (.A(g1740), .B(g17955), .Z(g18344) ) ;
AND2    gate12608  (.A(g1736), .B(g17955), .Z(g18345) ) ;
AND2    gate12609  (.A(g1752), .B(g17955), .Z(g18346) ) ;
AND2    gate12610  (.A(g1756), .B(g17955), .Z(g18347) ) ;
AND2    gate12611  (.A(g1744), .B(g17955), .Z(g18348) ) ;
AND2    gate12612  (.A(g1768), .B(g17955), .Z(g18349) ) ;
AND2    gate12613  (.A(g1779), .B(g17955), .Z(g18350) ) ;
AND2    gate12614  (.A(g1760), .B(g17955), .Z(g18351) ) ;
AND2    gate12615  (.A(g1798), .B(g17955), .Z(g18352) ) ;
AND2    gate12616  (.A(g1772), .B(g17955), .Z(g18353) ) ;
AND2    gate12617  (.A(g1792), .B(g17955), .Z(g18354) ) ;
AND2    gate12618  (.A(g1748), .B(g17955), .Z(g18355) ) ;
AND2    gate12619  (.A(g1802), .B(g17955), .Z(g18356) ) ;
AND2    gate12620  (.A(g1816), .B(g17955), .Z(g18357) ) ;
AND2    gate12621  (.A(g1811), .B(g17955), .Z(g18358) ) ;
AND2    gate12622  (.A(g1825), .B(g17955), .Z(g18359) ) ;
AND2    gate12623  (.A(g1830), .B(g17955), .Z(g18360) ) ;
AND2    gate12624  (.A(g1821), .B(g17955), .Z(g18361) ) ;
AND2    gate12625  (.A(g1834), .B(g17955), .Z(g18362) ) ;
AND2    gate12626  (.A(g1840), .B(g17955), .Z(g18363) ) ;
AND2    gate12627  (.A(g1844), .B(g17955), .Z(g18364) ) ;
AND2    gate12628  (.A(g1848), .B(g17955), .Z(g18365) ) ;
AND2    gate12629  (.A(g1854), .B(g17955), .Z(g18366) ) ;
AND2    gate12630  (.A(g1783), .B(g17955), .Z(g18367) ) ;
AND2    gate12631  (.A(g1728), .B(g17955), .Z(g18368) ) ;
NOR2    gate12632  (.A(g6839), .B(g10430), .Z(g12848) ) ;
AND2    gate12633  (.A(g12848), .B(g15171), .Z(g18369) ) ;
AND2    gate12634  (.A(g1874), .B(g15171), .Z(g18370) ) ;
AND2    gate12635  (.A(g1870), .B(g15171), .Z(g18371) ) ;
AND2    gate12636  (.A(g1886), .B(g15171), .Z(g18372) ) ;
AND2    gate12637  (.A(g1890), .B(g15171), .Z(g18373) ) ;
AND2    gate12638  (.A(g1878), .B(g15171), .Z(g18374) ) ;
AND2    gate12639  (.A(g1902), .B(g15171), .Z(g18375) ) ;
AND2    gate12640  (.A(g1913), .B(g15171), .Z(g18376) ) ;
AND2    gate12641  (.A(g1894), .B(g15171), .Z(g18377) ) ;
AND2    gate12642  (.A(g1932), .B(g15171), .Z(g18378) ) ;
AND2    gate12643  (.A(g1906), .B(g15171), .Z(g18379) ) ;
AND2    gate12644  (.A(g1926), .B(g15171), .Z(g18380) ) ;
AND2    gate12645  (.A(g1882), .B(g15171), .Z(g18381) ) ;
AND2    gate12646  (.A(g1936), .B(g15171), .Z(g18382) ) ;
AND2    gate12647  (.A(g1950), .B(g15171), .Z(g18383) ) ;
AND2    gate12648  (.A(g1945), .B(g15171), .Z(g18384) ) ;
AND2    gate12649  (.A(g1959), .B(g15171), .Z(g18385) ) ;
AND2    gate12650  (.A(g1964), .B(g15171), .Z(g18386) ) ;
AND2    gate12651  (.A(g1955), .B(g15171), .Z(g18387) ) ;
AND2    gate12652  (.A(g1968), .B(g15171), .Z(g18388) ) ;
AND2    gate12653  (.A(g1974), .B(g15171), .Z(g18389) ) ;
AND2    gate12654  (.A(g1978), .B(g15171), .Z(g18390) ) ;
AND2    gate12655  (.A(g1982), .B(g15171), .Z(g18391) ) ;
AND2    gate12656  (.A(g1988), .B(g15171), .Z(g18392) ) ;
AND2    gate12657  (.A(g1917), .B(g15171), .Z(g18393) ) ;
AND2    gate12658  (.A(g1862), .B(g15171), .Z(g18394) ) ;
NOR2    gate12659  (.A(g6840), .B(g10430), .Z(g12849) ) ;
AND2    gate12660  (.A(g12849), .B(g15373), .Z(g18395) ) ;
AND2    gate12661  (.A(g2008), .B(g15373), .Z(g18396) ) ;
AND2    gate12662  (.A(g2004), .B(g15373), .Z(g18397) ) ;
AND2    gate12663  (.A(g2020), .B(g15373), .Z(g18398) ) ;
AND2    gate12664  (.A(g2024), .B(g15373), .Z(g18399) ) ;
AND2    gate12665  (.A(g2012), .B(g15373), .Z(g18400) ) ;
AND2    gate12666  (.A(g2036), .B(g15373), .Z(g18401) ) ;
AND2    gate12667  (.A(g2047), .B(g15373), .Z(g18402) ) ;
AND2    gate12668  (.A(g2028), .B(g15373), .Z(g18403) ) ;
AND2    gate12669  (.A(g2066), .B(g15373), .Z(g18404) ) ;
AND2    gate12670  (.A(g2040), .B(g15373), .Z(g18405) ) ;
AND2    gate12671  (.A(g2060), .B(g15373), .Z(g18406) ) ;
AND2    gate12672  (.A(g2016), .B(g15373), .Z(g18407) ) ;
AND2    gate12673  (.A(g2070), .B(g15373), .Z(g18408) ) ;
AND2    gate12674  (.A(g2084), .B(g15373), .Z(g18409) ) ;
AND2    gate12675  (.A(g2079), .B(g15373), .Z(g18410) ) ;
AND2    gate12676  (.A(g2093), .B(g15373), .Z(g18411) ) ;
AND2    gate12677  (.A(g2098), .B(g15373), .Z(g18412) ) ;
AND2    gate12678  (.A(g2089), .B(g15373), .Z(g18413) ) ;
AND2    gate12679  (.A(g2102), .B(g15373), .Z(g18414) ) ;
AND2    gate12680  (.A(g2108), .B(g15373), .Z(g18415) ) ;
AND2    gate12681  (.A(g2112), .B(g15373), .Z(g18416) ) ;
AND2    gate12682  (.A(g2116), .B(g15373), .Z(g18417) ) ;
AND2    gate12683  (.A(g2122), .B(g15373), .Z(g18418) ) ;
AND2    gate12684  (.A(g2051), .B(g15373), .Z(g18419) ) ;
AND2    gate12685  (.A(g1996), .B(g15373), .Z(g18420) ) ;
NOR2    gate12686  (.A(g6846), .B(g10430), .Z(g12851) ) ;
AND2    gate12687  (.A(g12851), .B(g18008), .Z(g18423) ) ;
AND2    gate12688  (.A(g2165), .B(g18008), .Z(g18424) ) ;
AND2    gate12689  (.A(g2161), .B(g18008), .Z(g18425) ) ;
AND2    gate12690  (.A(g2177), .B(g18008), .Z(g18426) ) ;
AND2    gate12691  (.A(g2181), .B(g18008), .Z(g18427) ) ;
AND2    gate12692  (.A(g2169), .B(g18008), .Z(g18428) ) ;
AND2    gate12693  (.A(g2193), .B(g18008), .Z(g18429) ) ;
AND2    gate12694  (.A(g2204), .B(g18008), .Z(g18430) ) ;
AND2    gate12695  (.A(g2185), .B(g18008), .Z(g18431) ) ;
AND2    gate12696  (.A(g2223), .B(g18008), .Z(g18432) ) ;
AND2    gate12697  (.A(g2197), .B(g18008), .Z(g18433) ) ;
AND2    gate12698  (.A(g2217), .B(g18008), .Z(g18434) ) ;
AND2    gate12699  (.A(g2173), .B(g18008), .Z(g18435) ) ;
AND2    gate12700  (.A(g2227), .B(g18008), .Z(g18436) ) ;
AND2    gate12701  (.A(g2241), .B(g18008), .Z(g18437) ) ;
AND2    gate12702  (.A(g2236), .B(g18008), .Z(g18438) ) ;
AND2    gate12703  (.A(g2250), .B(g18008), .Z(g18439) ) ;
AND2    gate12704  (.A(g2255), .B(g18008), .Z(g18440) ) ;
AND2    gate12705  (.A(g2246), .B(g18008), .Z(g18441) ) ;
AND2    gate12706  (.A(g2259), .B(g18008), .Z(g18442) ) ;
AND2    gate12707  (.A(g2265), .B(g18008), .Z(g18443) ) ;
AND2    gate12708  (.A(g2269), .B(g18008), .Z(g18444) ) ;
AND2    gate12709  (.A(g2273), .B(g18008), .Z(g18445) ) ;
AND2    gate12710  (.A(g2279), .B(g18008), .Z(g18446) ) ;
AND2    gate12711  (.A(g2208), .B(g18008), .Z(g18447) ) ;
AND2    gate12712  (.A(g2153), .B(g18008), .Z(g18448) ) ;
NOR2    gate12713  (.A(g6847), .B(g10430), .Z(g12852) ) ;
AND2    gate12714  (.A(g12852), .B(g15224), .Z(g18449) ) ;
AND2    gate12715  (.A(g2299), .B(g15224), .Z(g18450) ) ;
AND2    gate12716  (.A(g2295), .B(g15224), .Z(g18451) ) ;
AND2    gate12717  (.A(g2311), .B(g15224), .Z(g18452) ) ;
AND2    gate12718  (.A(g2315), .B(g15224), .Z(g18453) ) ;
AND2    gate12719  (.A(g2303), .B(g15224), .Z(g18454) ) ;
AND2    gate12720  (.A(g2327), .B(g15224), .Z(g18455) ) ;
AND2    gate12721  (.A(g2338), .B(g15224), .Z(g18456) ) ;
AND2    gate12722  (.A(g2319), .B(g15224), .Z(g18457) ) ;
AND2    gate12723  (.A(g2357), .B(g15224), .Z(g18458) ) ;
AND2    gate12724  (.A(g2331), .B(g15224), .Z(g18459) ) ;
AND2    gate12725  (.A(g2351), .B(g15224), .Z(g18460) ) ;
AND2    gate12726  (.A(g2307), .B(g15224), .Z(g18461) ) ;
AND2    gate12727  (.A(g2361), .B(g15224), .Z(g18462) ) ;
AND2    gate12728  (.A(g2375), .B(g15224), .Z(g18463) ) ;
AND2    gate12729  (.A(g2370), .B(g15224), .Z(g18464) ) ;
AND2    gate12730  (.A(g2384), .B(g15224), .Z(g18465) ) ;
AND2    gate12731  (.A(g2389), .B(g15224), .Z(g18466) ) ;
AND2    gate12732  (.A(g2380), .B(g15224), .Z(g18467) ) ;
AND2    gate12733  (.A(g2393), .B(g15224), .Z(g18468) ) ;
AND2    gate12734  (.A(g2399), .B(g15224), .Z(g18469) ) ;
AND2    gate12735  (.A(g2403), .B(g15224), .Z(g18470) ) ;
AND2    gate12736  (.A(g2407), .B(g15224), .Z(g18471) ) ;
AND2    gate12737  (.A(g2413), .B(g15224), .Z(g18472) ) ;
AND2    gate12738  (.A(g2342), .B(g15224), .Z(g18473) ) ;
AND2    gate12739  (.A(g2287), .B(g15224), .Z(g18474) ) ;
NOR2    gate12740  (.A(g6848), .B(g10430), .Z(g12853) ) ;
AND2    gate12741  (.A(g12853), .B(g15426), .Z(g18475) ) ;
AND2    gate12742  (.A(g2433), .B(g15426), .Z(g18476) ) ;
AND2    gate12743  (.A(g2429), .B(g15426), .Z(g18477) ) ;
AND2    gate12744  (.A(g2445), .B(g15426), .Z(g18478) ) ;
AND2    gate12745  (.A(g2449), .B(g15426), .Z(g18479) ) ;
AND2    gate12746  (.A(g2437), .B(g15426), .Z(g18480) ) ;
AND2    gate12747  (.A(g2461), .B(g15426), .Z(g18481) ) ;
AND2    gate12748  (.A(g2472), .B(g15426), .Z(g18482) ) ;
AND2    gate12749  (.A(g2453), .B(g15426), .Z(g18483) ) ;
AND2    gate12750  (.A(g2491), .B(g15426), .Z(g18484) ) ;
AND2    gate12751  (.A(g2465), .B(g15426), .Z(g18485) ) ;
AND2    gate12752  (.A(g2485), .B(g15426), .Z(g18486) ) ;
AND2    gate12753  (.A(g2441), .B(g15426), .Z(g18487) ) ;
AND2    gate12754  (.A(g2495), .B(g15426), .Z(g18488) ) ;
AND2    gate12755  (.A(g2509), .B(g15426), .Z(g18489) ) ;
AND2    gate12756  (.A(g2504), .B(g15426), .Z(g18490) ) ;
AND2    gate12757  (.A(g2518), .B(g15426), .Z(g18491) ) ;
AND2    gate12758  (.A(g2523), .B(g15426), .Z(g18492) ) ;
AND2    gate12759  (.A(g2514), .B(g15426), .Z(g18493) ) ;
AND2    gate12760  (.A(g2527), .B(g15426), .Z(g18494) ) ;
AND2    gate12761  (.A(g2533), .B(g15426), .Z(g18495) ) ;
AND2    gate12762  (.A(g2537), .B(g15426), .Z(g18496) ) ;
AND2    gate12763  (.A(g2541), .B(g15426), .Z(g18497) ) ;
AND2    gate12764  (.A(g2547), .B(g15426), .Z(g18498) ) ;
AND2    gate12765  (.A(g2476), .B(g15426), .Z(g18499) ) ;
AND2    gate12766  (.A(g2421), .B(g15426), .Z(g18500) ) ;
NOR2    gate12767  (.A(g6849), .B(g10430), .Z(g12854) ) ;
AND2    gate12768  (.A(g12854), .B(g15509), .Z(g18501) ) ;
AND2    gate12769  (.A(g2567), .B(g15509), .Z(g18502) ) ;
AND2    gate12770  (.A(g2563), .B(g15509), .Z(g18503) ) ;
AND2    gate12771  (.A(g2579), .B(g15509), .Z(g18504) ) ;
AND2    gate12772  (.A(g2583), .B(g15509), .Z(g18505) ) ;
AND2    gate12773  (.A(g2571), .B(g15509), .Z(g18506) ) ;
AND2    gate12774  (.A(g2595), .B(g15509), .Z(g18507) ) ;
AND2    gate12775  (.A(g2606), .B(g15509), .Z(g18508) ) ;
AND2    gate12776  (.A(g2587), .B(g15509), .Z(g18509) ) ;
AND2    gate12777  (.A(g2625), .B(g15509), .Z(g18510) ) ;
AND2    gate12778  (.A(g2599), .B(g15509), .Z(g18511) ) ;
AND2    gate12779  (.A(g2619), .B(g15509), .Z(g18512) ) ;
AND2    gate12780  (.A(g2575), .B(g15509), .Z(g18513) ) ;
AND2    gate12781  (.A(g2629), .B(g15509), .Z(g18514) ) ;
AND2    gate12782  (.A(g2643), .B(g15509), .Z(g18515) ) ;
AND2    gate12783  (.A(g2638), .B(g15509), .Z(g18516) ) ;
AND2    gate12784  (.A(g2652), .B(g15509), .Z(g18517) ) ;
AND2    gate12785  (.A(g2657), .B(g15509), .Z(g18518) ) ;
AND2    gate12786  (.A(g2648), .B(g15509), .Z(g18519) ) ;
AND2    gate12787  (.A(g2661), .B(g15509), .Z(g18520) ) ;
AND2    gate12788  (.A(g2667), .B(g15509), .Z(g18521) ) ;
AND2    gate12789  (.A(g2671), .B(g15509), .Z(g18522) ) ;
AND2    gate12790  (.A(g2675), .B(g15509), .Z(g18523) ) ;
AND2    gate12791  (.A(g2681), .B(g15509), .Z(g18524) ) ;
AND2    gate12792  (.A(g2610), .B(g15509), .Z(g18525) ) ;
AND2    gate12793  (.A(g2555), .B(g15509), .Z(g18526) ) ;
AND2    gate12794  (.A(g2712), .B(g15277), .Z(g18529) ) ;
AND2    gate12795  (.A(g2715), .B(g15277), .Z(g18530) ) ;
AND2    gate12796  (.A(g2719), .B(g15277), .Z(g18531) ) ;
AND2    gate12797  (.A(g2724), .B(g15277), .Z(g18532) ) ;
AND2    gate12798  (.A(g2729), .B(g15277), .Z(g18533) ) ;
AND2    gate12799  (.A(g2735), .B(g15277), .Z(g18534) ) ;
AND2    gate12800  (.A(g2741), .B(g15277), .Z(g18535) ) ;
AND2    gate12801  (.A(g2748), .B(g15277), .Z(g18536) ) ;
AND2    gate12802  (.A(g6856), .B(g15277), .Z(g18537) ) ;
AND2    gate12803  (.A(g2759), .B(g15277), .Z(g18538) ) ;
AND2    gate12804  (.A(g2763), .B(g15277), .Z(g18539) ) ;
AND2    gate12805  (.A(g2775), .B(g15277), .Z(g18540) ) ;
AND2    gate12806  (.A(g2767), .B(g15277), .Z(g18541) ) ;
AND2    gate12807  (.A(g2787), .B(g15277), .Z(g18542) ) ;
AND2    gate12808  (.A(g2779), .B(g15277), .Z(g18543) ) ;
AND2    gate12809  (.A(g2791), .B(g15277), .Z(g18544) ) ;
AND2    gate12810  (.A(g2783), .B(g15277), .Z(g18545) ) ;
AND2    gate12811  (.A(g2795), .B(g15277), .Z(g18546) ) ;
AND2    gate12812  (.A(g121), .B(g15277), .Z(g18547) ) ;
AND2    gate12813  (.A(g2807), .B(g15277), .Z(g18548) ) ;
AND2    gate12814  (.A(g2799), .B(g15277), .Z(g18549) ) ;
AND2    gate12815  (.A(g2819), .B(g15277), .Z(g18550) ) ;
AND2    gate12816  (.A(g2811), .B(g15277), .Z(g18551) ) ;
AND2    gate12817  (.A(g2815), .B(g15277), .Z(g18552) ) ;
AND2    gate12818  (.A(g2827), .B(g15277), .Z(g18553) ) ;
AND2    gate12819  (.A(g2831), .B(g15277), .Z(g18554) ) ;
AND2    gate12820  (.A(g2834), .B(g15277), .Z(g18555) ) ;
AND2    gate12821  (.A(g2823), .B(g15277), .Z(g18556) ) ;
AND2    gate12822  (.A(g2771), .B(g15277), .Z(g18557) ) ;
AND2    gate12823  (.A(g2803), .B(g15277), .Z(g18558) ) ;
NOR2    gate12824  (.A(g10430), .B(g6855), .Z(g12856) ) ;
AND2    gate12825  (.A(g12856), .B(g15277), .Z(g18559) ) ;
AND2    gate12826  (.A(g2837), .B(g15277), .Z(g18560) ) ;
AND2    gate12827  (.A(g2841), .B(g15277), .Z(g18561) ) ;
AND2    gate12828  (.A(g2890), .B(g16349), .Z(g18563) ) ;
AND2    gate12829  (.A(g2844), .B(g16349), .Z(g18564) ) ;
AND2    gate12830  (.A(g2852), .B(g16349), .Z(g18565) ) ;
AND2    gate12831  (.A(g2860), .B(g16349), .Z(g18566) ) ;
AND2    gate12832  (.A(g2894), .B(g16349), .Z(g18567) ) ;
AND2    gate12833  (.A(g37), .B(g16349), .Z(g18568) ) ;
AND2    gate12834  (.A(g94), .B(g16349), .Z(g18569) ) ;
AND2    gate12835  (.A(g2848), .B(g16349), .Z(g18570) ) ;
AND2    gate12836  (.A(g2856), .B(g16349), .Z(g18571) ) ;
AND2    gate12837  (.A(g2864), .B(g16349), .Z(g18572) ) ;
AND2    gate12838  (.A(g2898), .B(g16349), .Z(g18573) ) ;
AND2    gate12839  (.A(g2882), .B(g16349), .Z(g18574) ) ;
AND2    gate12840  (.A(g2878), .B(g16349), .Z(g18575) ) ;
AND2    gate12841  (.A(g2868), .B(g16349), .Z(g18576) ) ;
AND2    gate12842  (.A(g2988), .B(g16349), .Z(g18577) ) ;
AND2    gate12843  (.A(g2873), .B(g16349), .Z(g18578) ) ;
AND2    gate12844  (.A(g2984), .B(g16349), .Z(g18579) ) ;
AND2    gate12845  (.A(g2907), .B(g16349), .Z(g18580) ) ;
AND2    gate12846  (.A(g2912), .B(g16349), .Z(g18581) ) ;
AND2    gate12847  (.A(g2922), .B(g16349), .Z(g18582) ) ;
AND2    gate12848  (.A(g2936), .B(g16349), .Z(g18583) ) ;
AND2    gate12849  (.A(g2950), .B(g16349), .Z(g18584) ) ;
AND2    gate12850  (.A(g2960), .B(g16349), .Z(g18585) ) ;
AND2    gate12851  (.A(g2886), .B(g16349), .Z(g18586) ) ;
AND2    gate12852  (.A(g2980), .B(g16349), .Z(g18587) ) ;
AND2    gate12853  (.A(g2970), .B(g16349), .Z(g18588) ) ;
AND2    gate12854  (.A(g2902), .B(g16349), .Z(g18589) ) ;
AND2    gate12855  (.A(g2917), .B(g16349), .Z(g18590) ) ;
AND2    gate12856  (.A(g2965), .B(g16349), .Z(g18591) ) ;
AND2    gate12857  (.A(g2994), .B(g16349), .Z(g18592) ) ;
AND2    gate12858  (.A(g2999), .B(g16349), .Z(g18593) ) ;
NOR2    gate12859  (.A(g10365), .B(g10430), .Z(g12858) ) ;
AND2    gate12860  (.A(g12858), .B(g16349), .Z(g18594) ) ;
AND2    gate12861  (.A(g2927), .B(g16349), .Z(g18595) ) ;
AND2    gate12862  (.A(g2941), .B(g16349), .Z(g18596) ) ;
AND2    gate12863  (.A(g2955), .B(g16349), .Z(g18599) ) ;
AND2    gate12864  (.A(g3111), .B(g16987), .Z(g18600) ) ;
AND2    gate12865  (.A(g3106), .B(g16987), .Z(g18601) ) ;
AND2    gate12866  (.A(g3115), .B(g16987), .Z(g18602) ) ;
AND2    gate12867  (.A(g3119), .B(g16987), .Z(g18603) ) ;
AND2    gate12868  (.A(g3125), .B(g16987), .Z(g18604) ) ;
AND2    gate12869  (.A(g3129), .B(g16987), .Z(g18605) ) ;
AND2    gate12870  (.A(g3133), .B(g16987), .Z(g18606) ) ;
AND2    gate12871  (.A(g3139), .B(g16987), .Z(g18607) ) ;
NOR2    gate12872  (.A(g12860), .B(g13144), .Z(g15087) ) ;
AND2    gate12873  (.A(g15087), .B(g16987), .Z(g18608) ) ;
AND2    gate12874  (.A(g3147), .B(g16987), .Z(g18609) ) ;
NOR2    gate12875  (.A(g13144), .B(g6874), .Z(g15088) ) ;
AND2    gate12876  (.A(g15088), .B(g17059), .Z(g18610) ) ;
NOR2    gate12877  (.A(g13144), .B(g12862), .Z(g15090) ) ;
AND2    gate12878  (.A(g15090), .B(g17200), .Z(g18611) ) ;
AND2    gate12879  (.A(g3329), .B(g17200), .Z(g18612) ) ;
AND2    gate12880  (.A(g3338), .B(g17200), .Z(g18613) ) ;
AND2    gate12881  (.A(g3343), .B(g17200), .Z(g18614) ) ;
AND2    gate12882  (.A(g3347), .B(g17200), .Z(g18615) ) ;
AND2    gate12883  (.A(g6875), .B(g17200), .Z(g18616) ) ;
AND2    gate12884  (.A(g3462), .B(g17062), .Z(g18617) ) ;
AND2    gate12885  (.A(g3457), .B(g17062), .Z(g18618) ) ;
AND2    gate12886  (.A(g3466), .B(g17062), .Z(g18619) ) ;
AND2    gate12887  (.A(g3470), .B(g17062), .Z(g18620) ) ;
AND2    gate12888  (.A(g3476), .B(g17062), .Z(g18621) ) ;
AND2    gate12889  (.A(g3480), .B(g17062), .Z(g18622) ) ;
AND2    gate12890  (.A(g3484), .B(g17062), .Z(g18623) ) ;
AND2    gate12891  (.A(g3490), .B(g17062), .Z(g18624) ) ;
NOR2    gate12892  (.A(g12864), .B(g13177), .Z(g15092) ) ;
AND2    gate12893  (.A(g15092), .B(g17062), .Z(g18625) ) ;
AND2    gate12894  (.A(g3498), .B(g17062), .Z(g18626) ) ;
NOR2    gate12895  (.A(g13177), .B(g6904), .Z(g15093) ) ;
AND2    gate12896  (.A(g15093), .B(g17093), .Z(g18627) ) ;
NOR2    gate12897  (.A(g13177), .B(g12866), .Z(g15095) ) ;
AND2    gate12898  (.A(g15095), .B(g17226), .Z(g18628) ) ;
AND2    gate12899  (.A(g3680), .B(g17226), .Z(g18629) ) ;
AND2    gate12900  (.A(g3689), .B(g17226), .Z(g18630) ) ;
AND2    gate12901  (.A(g3694), .B(g17226), .Z(g18631) ) ;
AND2    gate12902  (.A(g3698), .B(g17226), .Z(g18632) ) ;
AND2    gate12903  (.A(g6905), .B(g17226), .Z(g18633) ) ;
AND2    gate12904  (.A(g3813), .B(g17096), .Z(g18634) ) ;
AND2    gate12905  (.A(g3808), .B(g17096), .Z(g18635) ) ;
AND2    gate12906  (.A(g3817), .B(g17096), .Z(g18636) ) ;
AND2    gate12907  (.A(g3821), .B(g17096), .Z(g18637) ) ;
AND2    gate12908  (.A(g3827), .B(g17096), .Z(g18638) ) ;
AND2    gate12909  (.A(g3831), .B(g17096), .Z(g18639) ) ;
AND2    gate12910  (.A(g3835), .B(g17096), .Z(g18640) ) ;
AND2    gate12911  (.A(g3841), .B(g17096), .Z(g18641) ) ;
NOR2    gate12912  (.A(g12868), .B(g13191), .Z(g15097) ) ;
AND2    gate12913  (.A(g15097), .B(g17096), .Z(g18642) ) ;
AND2    gate12914  (.A(g3849), .B(g17096), .Z(g18643) ) ;
NOR2    gate12915  (.A(g13191), .B(g6927), .Z(g15098) ) ;
AND2    gate12916  (.A(g15098), .B(g17125), .Z(g18644) ) ;
NOR2    gate12917  (.A(g13191), .B(g12870), .Z(g15100) ) ;
AND2    gate12918  (.A(g15100), .B(g17271), .Z(g18645) ) ;
AND2    gate12919  (.A(g4031), .B(g17271), .Z(g18646) ) ;
AND2    gate12920  (.A(g4040), .B(g17271), .Z(g18647) ) ;
AND2    gate12921  (.A(g4045), .B(g17271), .Z(g18648) ) ;
AND2    gate12922  (.A(g4049), .B(g17271), .Z(g18649) ) ;
AND2    gate12923  (.A(g6928), .B(g17271), .Z(g18650) ) ;
NOR2    gate12924  (.A(g14591), .B(g6954), .Z(g15102) ) ;
AND2    gate12925  (.A(g15102), .B(g16249), .Z(g18651) ) ;
AND2    gate12926  (.A(g4172), .B(g16249), .Z(g18652) ) ;
AND2    gate12927  (.A(g4176), .B(g16249), .Z(g18653) ) ;
AND2    gate12928  (.A(g4146), .B(g16249), .Z(g18654) ) ;
NOR2    gate12929  (.A(g12872), .B(g10430), .Z(g15106) ) ;
AND2    gate12930  (.A(g15106), .B(g14454), .Z(g18655) ) ;
NOR2    gate12931  (.A(g12873), .B(g13605), .Z(g15120) ) ;
AND2    gate12932  (.A(g15120), .B(g17128), .Z(g18656) ) ;
AND2    gate12933  (.A(g4308), .B(g17128), .Z(g18657) ) ;
NOR2    gate12934  (.A(g12874), .B(g13605), .Z(g15121) ) ;
AND2    gate12935  (.A(g15121), .B(g17183), .Z(g18658) ) ;
AND2    gate12936  (.A(g4366), .B(g17183), .Z(g18659) ) ;
NOR2    gate12937  (.A(g12878), .B(g13605), .Z(g15126) ) ;
AND2    gate12938  (.A(g15126), .B(g17367), .Z(g18662) ) ;
AND2    gate12939  (.A(g4311), .B(g17367), .Z(g18663) ) ;
AND2    gate12940  (.A(g4332), .B(g17367), .Z(g18664) ) ;
AND2    gate12941  (.A(g4584), .B(g17367), .Z(g18665) ) ;
AND2    gate12942  (.A(g4593), .B(g17367), .Z(g18666) ) ;
AND2    gate12943  (.A(g4601), .B(g17367), .Z(g18667) ) ;
AND2    gate12944  (.A(g4322), .B(g17367), .Z(g18668) ) ;
AND2    gate12945  (.A(g4608), .B(g17367), .Z(g18669) ) ;
AND2    gate12946  (.A(g4621), .B(g15758), .Z(g18670) ) ;
AND2    gate12947  (.A(g4628), .B(g15758), .Z(g18671) ) ;
NOR2    gate12948  (.A(g12879), .B(g13605), .Z(g15127) ) ;
AND2    gate12949  (.A(g15127), .B(g15758), .Z(g18672) ) ;
AND2    gate12950  (.A(g4643), .B(g15758), .Z(g18673) ) ;
AND2    gate12951  (.A(g4340), .B(g15758), .Z(g18674) ) ;
AND2    gate12952  (.A(g4349), .B(g15758), .Z(g18675) ) ;
AND2    gate12953  (.A(g4358), .B(g15758), .Z(g18676) ) ;
AND2    gate12954  (.A(g4639), .B(g15758), .Z(g18677) ) ;
AND2    gate12955  (.A(g66), .B(g15758), .Z(g18678) ) ;
AND2    gate12956  (.A(g4633), .B(g15758), .Z(g18679) ) ;
NOR2    gate12957  (.A(g13638), .B(g12880), .Z(g15128) ) ;
AND2    gate12958  (.A(g15128), .B(g15885), .Z(g18680) ) ;
AND2    gate12959  (.A(g4653), .B(g15885), .Z(g18681) ) ;
AND2    gate12960  (.A(g4646), .B(g15885), .Z(g18682) ) ;
AND2    gate12961  (.A(g4674), .B(g15885), .Z(g18683) ) ;
AND2    gate12962  (.A(g4681), .B(g15885), .Z(g18684) ) ;
AND2    gate12963  (.A(g4688), .B(g15885), .Z(g18685) ) ;
AND2    gate12964  (.A(g4659), .B(g15885), .Z(g18686) ) ;
AND2    gate12965  (.A(g4664), .B(g15885), .Z(g18687) ) ;
AND2    gate12966  (.A(g4704), .B(g16752), .Z(g18688) ) ;
NOR2    gate12967  (.A(g6984), .B(g13638), .Z(g15129) ) ;
AND2    gate12968  (.A(g15129), .B(g16752), .Z(g18689) ) ;
NOR2    gate12969  (.A(g13638), .B(g6985), .Z(g15130) ) ;
AND2    gate12970  (.A(g15130), .B(g16053), .Z(g18690) ) ;
AND2    gate12971  (.A(g4727), .B(g16053), .Z(g18691) ) ;
AND2    gate12972  (.A(g4732), .B(g16053), .Z(g18692) ) ;
AND2    gate12973  (.A(g4717), .B(g16053), .Z(g18693) ) ;
AND2    gate12974  (.A(g4722), .B(g16053), .Z(g18694) ) ;
AND2    gate12975  (.A(g4749), .B(g16777), .Z(g18697) ) ;
NOR2    gate12976  (.A(g12881), .B(g13638), .Z(g15131) ) ;
AND2    gate12977  (.A(g15131), .B(g16777), .Z(g18698) ) ;
AND2    gate12978  (.A(g4760), .B(g16816), .Z(g18699) ) ;
NOR2    gate12979  (.A(g12882), .B(g13638), .Z(g15132) ) ;
AND2    gate12980  (.A(g15132), .B(g16816), .Z(g18700) ) ;
AND2    gate12981  (.A(g4771), .B(g16856), .Z(g18701) ) ;
NOR2    gate12982  (.A(g12883), .B(g13638), .Z(g15133) ) ;
AND2    gate12983  (.A(g15133), .B(g16856), .Z(g18702) ) ;
AND2    gate12984  (.A(g4776), .B(g16782), .Z(g18703) ) ;
AND2    gate12985  (.A(g4793), .B(g16782), .Z(g18704) ) ;
AND2    gate12986  (.A(g4801), .B(g16782), .Z(g18705) ) ;
AND2    gate12987  (.A(g4785), .B(g16782), .Z(g18706) ) ;
NOR2    gate12988  (.A(g13638), .B(g12884), .Z(g15134) ) ;
AND2    gate12989  (.A(g15134), .B(g16782), .Z(g18707) ) ;
AND2    gate12990  (.A(g4818), .B(g16782), .Z(g18708) ) ;
AND2    gate12991  (.A(g59), .B(g17302), .Z(g18709) ) ;
NOR2    gate12992  (.A(g6990), .B(g13638), .Z(g15135) ) ;
AND2    gate12993  (.A(g15135), .B(g17302), .Z(g18710) ) ;
NOR2    gate12994  (.A(g13680), .B(g12885), .Z(g15136) ) ;
AND2    gate12995  (.A(g15136), .B(g15915), .Z(g18711) ) ;
AND2    gate12996  (.A(g4843), .B(g15915), .Z(g18712) ) ;
AND2    gate12997  (.A(g4836), .B(g15915), .Z(g18713) ) ;
AND2    gate12998  (.A(g4864), .B(g15915), .Z(g18714) ) ;
AND2    gate12999  (.A(g4871), .B(g15915), .Z(g18715) ) ;
AND2    gate13000  (.A(g4878), .B(g15915), .Z(g18716) ) ;
AND2    gate13001  (.A(g4849), .B(g15915), .Z(g18717) ) ;
AND2    gate13002  (.A(g4854), .B(g15915), .Z(g18718) ) ;
AND2    gate13003  (.A(g4894), .B(g16795), .Z(g18719) ) ;
NOR2    gate13004  (.A(g6992), .B(g13680), .Z(g15137) ) ;
AND2    gate13005  (.A(g15137), .B(g16795), .Z(g18720) ) ;
NOR2    gate13006  (.A(g13680), .B(g6993), .Z(g15138) ) ;
AND2    gate13007  (.A(g15138), .B(g16077), .Z(g18721) ) ;
AND2    gate13008  (.A(g4917), .B(g16077), .Z(g18722) ) ;
AND2    gate13009  (.A(g4922), .B(g16077), .Z(g18723) ) ;
AND2    gate13010  (.A(g4907), .B(g16077), .Z(g18724) ) ;
AND2    gate13011  (.A(g4912), .B(g16077), .Z(g18725) ) ;
AND2    gate13012  (.A(g4939), .B(g16821), .Z(g18728) ) ;
NOR2    gate13013  (.A(g12886), .B(g13680), .Z(g15139) ) ;
AND2    gate13014  (.A(g15139), .B(g16821), .Z(g18729) ) ;
AND2    gate13015  (.A(g4950), .B(g16861), .Z(g18730) ) ;
NOR2    gate13016  (.A(g12887), .B(g13680), .Z(g15140) ) ;
AND2    gate13017  (.A(g15140), .B(g16861), .Z(g18731) ) ;
AND2    gate13018  (.A(g4961), .B(g16877), .Z(g18732) ) ;
NOR2    gate13019  (.A(g12888), .B(g13680), .Z(g15141) ) ;
AND2    gate13020  (.A(g15141), .B(g16877), .Z(g18733) ) ;
AND2    gate13021  (.A(g4966), .B(g16826), .Z(g18734) ) ;
AND2    gate13022  (.A(g4983), .B(g16826), .Z(g18735) ) ;
AND2    gate13023  (.A(g4991), .B(g16826), .Z(g18736) ) ;
AND2    gate13024  (.A(g4975), .B(g16826), .Z(g18737) ) ;
NOR2    gate13025  (.A(g13680), .B(g12889), .Z(g15142) ) ;
AND2    gate13026  (.A(g15142), .B(g16826), .Z(g18738) ) ;
AND2    gate13027  (.A(g5008), .B(g16826), .Z(g18739) ) ;
AND2    gate13028  (.A(g4572), .B(g17384), .Z(g18740) ) ;
NOR2    gate13029  (.A(g6998), .B(g13680), .Z(g15143) ) ;
AND2    gate13030  (.A(g15143), .B(g17384), .Z(g18741) ) ;
AND2    gate13031  (.A(g5120), .B(g17847), .Z(g18742) ) ;
AND2    gate13032  (.A(g5115), .B(g17847), .Z(g18743) ) ;
AND2    gate13033  (.A(g5124), .B(g17847), .Z(g18744) ) ;
AND2    gate13034  (.A(g5128), .B(g17847), .Z(g18745) ) ;
AND2    gate13035  (.A(g5134), .B(g17847), .Z(g18746) ) ;
AND2    gate13036  (.A(g5138), .B(g17847), .Z(g18747) ) ;
AND2    gate13037  (.A(g5142), .B(g17847), .Z(g18748) ) ;
AND2    gate13038  (.A(g5148), .B(g17847), .Z(g18749) ) ;
NOR2    gate13039  (.A(g12891), .B(g13716), .Z(g15145) ) ;
AND2    gate13040  (.A(g15145), .B(g17847), .Z(g18750) ) ;
AND2    gate13041  (.A(g5156), .B(g17847), .Z(g18751) ) ;
NOR2    gate13042  (.A(g13716), .B(g7003), .Z(g15146) ) ;
AND2    gate13043  (.A(g15146), .B(g17926), .Z(g18752) ) ;
NOR2    gate13044  (.A(g13716), .B(g12893), .Z(g15148) ) ;
AND2    gate13045  (.A(g15148), .B(g15595), .Z(g18753) ) ;
AND2    gate13046  (.A(g5339), .B(g15595), .Z(g18754) ) ;
AND2    gate13047  (.A(g5343), .B(g15595), .Z(g18755) ) ;
AND2    gate13048  (.A(g5348), .B(g15595), .Z(g18756) ) ;
AND2    gate13049  (.A(g5352), .B(g15595), .Z(g18757) ) ;
AND2    gate13050  (.A(g7004), .B(g15595), .Z(g18758) ) ;
AND2    gate13051  (.A(g5467), .B(g17929), .Z(g18759) ) ;
AND2    gate13052  (.A(g5462), .B(g17929), .Z(g18760) ) ;
AND2    gate13053  (.A(g5471), .B(g17929), .Z(g18761) ) ;
AND2    gate13054  (.A(g5475), .B(g17929), .Z(g18762) ) ;
AND2    gate13055  (.A(g5481), .B(g17929), .Z(g18763) ) ;
AND2    gate13056  (.A(g5485), .B(g17929), .Z(g18764) ) ;
AND2    gate13057  (.A(g5489), .B(g17929), .Z(g18765) ) ;
AND2    gate13058  (.A(g5495), .B(g17929), .Z(g18766) ) ;
NOR2    gate13059  (.A(g12895), .B(g13745), .Z(g15150) ) ;
AND2    gate13060  (.A(g15150), .B(g17929), .Z(g18767) ) ;
AND2    gate13061  (.A(g5503), .B(g17929), .Z(g18768) ) ;
NOR2    gate13062  (.A(g13745), .B(g7027), .Z(g15151) ) ;
AND2    gate13063  (.A(g15151), .B(g18062), .Z(g18769) ) ;
NOR2    gate13064  (.A(g13745), .B(g12897), .Z(g15153) ) ;
AND2    gate13065  (.A(g15153), .B(g15615), .Z(g18770) ) ;
AND2    gate13066  (.A(g5685), .B(g15615), .Z(g18771) ) ;
AND2    gate13067  (.A(g5689), .B(g15615), .Z(g18772) ) ;
AND2    gate13068  (.A(g5694), .B(g15615), .Z(g18773) ) ;
AND2    gate13069  (.A(g5698), .B(g15615), .Z(g18774) ) ;
AND2    gate13070  (.A(g7028), .B(g15615), .Z(g18775) ) ;
AND2    gate13071  (.A(g5813), .B(g18065), .Z(g18776) ) ;
AND2    gate13072  (.A(g5808), .B(g18065), .Z(g18777) ) ;
AND2    gate13073  (.A(g5817), .B(g18065), .Z(g18778) ) ;
AND2    gate13074  (.A(g5821), .B(g18065), .Z(g18779) ) ;
AND2    gate13075  (.A(g5827), .B(g18065), .Z(g18780) ) ;
AND2    gate13076  (.A(g5831), .B(g18065), .Z(g18781) ) ;
AND2    gate13077  (.A(g5835), .B(g18065), .Z(g18782) ) ;
AND2    gate13078  (.A(g5841), .B(g18065), .Z(g18783) ) ;
NOR2    gate13079  (.A(g12899), .B(g13782), .Z(g15155) ) ;
AND2    gate13080  (.A(g15155), .B(g18065), .Z(g18784) ) ;
AND2    gate13081  (.A(g5849), .B(g18065), .Z(g18785) ) ;
NOR2    gate13082  (.A(g13782), .B(g7050), .Z(g15156) ) ;
AND2    gate13083  (.A(g15156), .B(g15345), .Z(g18786) ) ;
NOR2    gate13084  (.A(g13782), .B(g12901), .Z(g15158) ) ;
AND2    gate13085  (.A(g15158), .B(g15634), .Z(g18787) ) ;
AND2    gate13086  (.A(g6031), .B(g15634), .Z(g18788) ) ;
AND2    gate13087  (.A(g6035), .B(g15634), .Z(g18789) ) ;
AND2    gate13088  (.A(g6040), .B(g15634), .Z(g18790) ) ;
AND2    gate13089  (.A(g6044), .B(g15634), .Z(g18791) ) ;
AND2    gate13090  (.A(g7051), .B(g15634), .Z(g18792) ) ;
AND2    gate13091  (.A(g6159), .B(g15348), .Z(g18793) ) ;
AND2    gate13092  (.A(g6154), .B(g15348), .Z(g18794) ) ;
AND2    gate13093  (.A(g6163), .B(g15348), .Z(g18795) ) ;
AND2    gate13094  (.A(g6167), .B(g15348), .Z(g18796) ) ;
AND2    gate13095  (.A(g6173), .B(g15348), .Z(g18797) ) ;
AND2    gate13096  (.A(g6177), .B(g15348), .Z(g18798) ) ;
AND2    gate13097  (.A(g6181), .B(g15348), .Z(g18799) ) ;
AND2    gate13098  (.A(g6187), .B(g15348), .Z(g18800) ) ;
NOR2    gate13099  (.A(g12903), .B(g13809), .Z(g15160) ) ;
AND2    gate13100  (.A(g15160), .B(g15348), .Z(g18801) ) ;
AND2    gate13101  (.A(g6195), .B(g15348), .Z(g18802) ) ;
NOR2    gate13102  (.A(g13809), .B(g7073), .Z(g15161) ) ;
AND2    gate13103  (.A(g15161), .B(g15480), .Z(g18803) ) ;
NOR2    gate13104  (.A(g13809), .B(g12905), .Z(g15163) ) ;
AND2    gate13105  (.A(g15163), .B(g15656), .Z(g18804) ) ;
AND2    gate13106  (.A(g6377), .B(g15656), .Z(g18805) ) ;
AND2    gate13107  (.A(g6381), .B(g15656), .Z(g18806) ) ;
AND2    gate13108  (.A(g6386), .B(g15656), .Z(g18807) ) ;
AND2    gate13109  (.A(g6390), .B(g15656), .Z(g18808) ) ;
AND2    gate13110  (.A(g7074), .B(g15656), .Z(g18809) ) ;
AND2    gate13111  (.A(g6505), .B(g15483), .Z(g18810) ) ;
AND2    gate13112  (.A(g6500), .B(g15483), .Z(g18811) ) ;
AND2    gate13113  (.A(g6509), .B(g15483), .Z(g18812) ) ;
AND2    gate13114  (.A(g6513), .B(g15483), .Z(g18813) ) ;
AND2    gate13115  (.A(g6519), .B(g15483), .Z(g18814) ) ;
AND2    gate13116  (.A(g6523), .B(g15483), .Z(g18815) ) ;
AND2    gate13117  (.A(g6527), .B(g15483), .Z(g18816) ) ;
AND2    gate13118  (.A(g6533), .B(g15483), .Z(g18817) ) ;
NOR2    gate13119  (.A(g12907), .B(g13835), .Z(g15165) ) ;
AND2    gate13120  (.A(g15165), .B(g15483), .Z(g18818) ) ;
AND2    gate13121  (.A(g6541), .B(g15483), .Z(g18819) ) ;
NOR2    gate13122  (.A(g13835), .B(g7096), .Z(g15166) ) ;
AND2    gate13123  (.A(g15166), .B(g15563), .Z(g18820) ) ;
NOR2    gate13124  (.A(g13835), .B(g12909), .Z(g15168) ) ;
AND2    gate13125  (.A(g15168), .B(g15680), .Z(g18821) ) ;
AND2    gate13126  (.A(g6723), .B(g15680), .Z(g18822) ) ;
AND2    gate13127  (.A(g6727), .B(g15680), .Z(g18823) ) ;
AND2    gate13128  (.A(g6732), .B(g15680), .Z(g18824) ) ;
AND2    gate13129  (.A(g6736), .B(g15680), .Z(g18825) ) ;
AND2    gate13130  (.A(g7097), .B(g15680), .Z(g18826) ) ;
NOR2    gate13131  (.A(g14541), .B(g12123), .Z(g17625) ) ;
AND2    gate13132  (.A(g10158), .B(g17625), .Z(g18890) ) ;
NOR2    gate13133  (.A(g1211), .B(g13545), .Z(g16215) ) ;
AND2    gate13134  (.A(g16215), .B(g16030), .Z(g18893) ) ;
NOR2    gate13135  (.A(g8046), .B(g12527), .Z(g13568) ) ;
AND2    gate13136  (.A(g13568), .B(g16264), .Z(g18906) ) ;
NOR2    gate13137  (.A(g8052), .B(g13545), .Z(g16226) ) ;
AND2    gate13138  (.A(g16226), .B(g13570), .Z(g18909) ) ;
NOR2    gate13139  (.A(g1554), .B(g13574), .Z(g16227) ) ;
AND2    gate13140  (.A(g16227), .B(g16075), .Z(g18910) ) ;
NOR2    gate13141  (.A(g8088), .B(g13574), .Z(g16237) ) ;
AND2    gate13142  (.A(g16237), .B(g13597), .Z(g18933) ) ;
AND2    gate13143  (.A(g3133), .B(g16096), .Z(g18934) ) ;
AND2    gate13144  (.A(g269), .B(g16099), .Z(g18943) ) ;
AND2    gate13145  (.A(g10183), .B(g17625), .Z(g18949) ) ;
NAND2   gate13146  (.A(II14258), .B(II14259), .Z(g11193) ) ;
AND2    gate13147  (.A(g11193), .B(g16123), .Z(g18950) ) ;
AND2    gate13148  (.A(g3484), .B(g16124), .Z(g18951) ) ;
AND2    gate13149  (.A(g174), .B(g16127), .Z(g18974) ) ;
NAND2   gate13150  (.A(II14276), .B(II14277), .Z(g11206) ) ;
AND2    gate13151  (.A(g11206), .B(g16158), .Z(g18981) ) ;
AND2    gate13152  (.A(g3835), .B(g16159), .Z(g18982) ) ;
AND2    gate13153  (.A(g182), .B(g16162), .Z(g18987) ) ;
AND2    gate13154  (.A(g8341), .B(g16171), .Z(g18992) ) ;
NAND2   gate13155  (.A(II14290), .B(II14291), .Z(g11224) ) ;
AND2    gate13156  (.A(g11224), .B(g16172), .Z(g18993) ) ;
AND2    gate13157  (.A(g446), .B(g16180), .Z(g19062) ) ;
AND2    gate13158  (.A(g8397), .B(g16186), .Z(g19069) ) ;
AND2    gate13159  (.A(g452), .B(g16195), .Z(g19139) ) ;
AND2    gate13160  (.A(g8450), .B(g16200), .Z(g19145) ) ;
AND2    gate13161  (.A(g460), .B(g16206), .Z(g19206) ) ;
NAND2   gate13162  (.A(II12204), .B(II12205), .Z(g7803) ) ;
AND2    gate13163  (.A(g7803), .B(g15992), .Z(g19207) ) ;
AND2    gate13164  (.A(g246), .B(g16214), .Z(g19266) ) ;
NAND2   gate13165  (.A(II12218), .B(II12219), .Z(g7823) ) ;
AND2    gate13166  (.A(g7823), .B(g16044), .Z(g19275) ) ;
AND2    gate13167  (.A(g464), .B(g16223), .Z(g19333) ) ;
OR2     gate13168  (.A(g13038), .B(g10677), .Z(g15968) ) ;
AND2    gate13169  (.A(g471), .B(g16235), .Z(g19354) ) ;
AND2    gate13170  (.A(g686), .B(g16289), .Z(g19372) ) ;
NAND3   gate13171  (.A(g10685), .B(g13252), .C(g703), .Z(g16893) ) ;
AND2    gate13172  (.A(g16893), .B(g13223), .Z(g19383) ) ;
AND2    gate13173  (.A(g667), .B(g16310), .Z(g19384) ) ;
AND2    gate13174  (.A(g691), .B(g16325), .Z(g19393) ) ;
NAND2   gate13175  (.A(g10147), .B(g10110), .Z(g11708) ) ;
AND2    gate13176  (.A(g11708), .B(g16846), .Z(g19461) ) ;
NAND2   gate13177  (.A(g554), .B(g807), .Z(g7850) ) ;
OR3     gate13178  (.A(g11741), .B(g11721), .C(g753), .Z(g14182) ) ;
NAND3   gate13179  (.A(g11741), .B(g11721), .C(g753), .Z(g14177) ) ;
AND4    gate13180  (.A(g7850), .B(g14182), .C(g14177), .D(g16646), .Z(g19462) ) ;
AND2    gate13181  (.A(g499), .B(g16680), .Z(g19487) ) ;
AND2    gate13182  (.A(g504), .B(g16712), .Z(g19500) ) ;
NAND2   gate13183  (.A(g13319), .B(g10998), .Z(g16097) ) ;
AND2    gate13184  (.A(g7824), .B(g16097), .Z(g19516) ) ;
AND2    gate13185  (.A(g513), .B(g16739), .Z(g19521) ) ;
AND2    gate13186  (.A(g518), .B(g16768), .Z(g19536) ) ;
NAND2   gate13187  (.A(II17380), .B(II17381), .Z(g15904) ) ;
AND2    gate13188  (.A(g1124), .B(g15904), .Z(g19540) ) ;
AND2    gate13189  (.A(g3147), .B(g16769), .Z(g19545) ) ;
NOR2    gate13190  (.A(g843), .B(g9166), .Z(g11932) ) ;
AND2    gate13191  (.A(g11932), .B(g16809), .Z(g19556) ) ;
NAND3   gate13192  (.A(g7903), .B(g7479), .C(g13256), .Z(g15832) ) ;
AND3    gate13193  (.A(g15832), .B(g1157), .C(g10893), .Z(g19560) ) ;
NOR2    gate13194  (.A(g1216), .B(g13545), .Z(g17175) ) ;
AND2    gate13195  (.A(g17175), .B(g13976), .Z(g19564) ) ;
NAND2   gate13196  (.A(II17405), .B(II17406), .Z(g15959) ) ;
AND2    gate13197  (.A(g1467), .B(g15959), .Z(g19568) ) ;
AND2    gate13198  (.A(g3498), .B(g16812), .Z(g19571) ) ;
NOR2    gate13199  (.A(g9223), .B(g13545), .Z(g16183) ) ;
AND2    gate13200  (.A(g16183), .B(g11130), .Z(g19578) ) ;
NAND3   gate13201  (.A(g7922), .B(g7503), .C(g13264), .Z(g15843) ) ;
AND3    gate13202  (.A(g15843), .B(g1500), .C(g10918), .Z(g19581) ) ;
NOR2    gate13203  (.A(g1559), .B(g13574), .Z(g17180) ) ;
AND2    gate13204  (.A(g17180), .B(g14004), .Z(g19585) ) ;
AND2    gate13205  (.A(g3849), .B(g16853), .Z(g19588) ) ;
NOR2    gate13206  (.A(g7197), .B(g9166), .Z(g11913) ) ;
AND2    gate13207  (.A(g11913), .B(g17268), .Z(g19594) ) ;
NAND2   gate13208  (.A(II17884), .B(II17885), .Z(g16681) ) ;
AND2    gate13209  (.A(g1094), .B(g16681), .Z(g19596) ) ;
NOR2    gate13210  (.A(g9247), .B(g13574), .Z(g16198) ) ;
AND2    gate13211  (.A(g16198), .B(g11149), .Z(g19601) ) ;
NAND2   gate13212  (.A(II17447), .B(II17448), .Z(g16069) ) ;
AND2    gate13213  (.A(g1141), .B(g16069), .Z(g19610) ) ;
NAND2   gate13214  (.A(II17924), .B(II17925), .Z(g16713) ) ;
AND2    gate13215  (.A(g1437), .B(g16713), .Z(g19613) ) ;
NAND2   gate13216  (.A(II17461), .B(II17462), .Z(g16093) ) ;
AND2    gate13217  (.A(g1484), .B(g16093), .Z(g19631) ) ;
AND2    gate13218  (.A(g5142), .B(g16958), .Z(g19637) ) ;
NAND2   gate13219  (.A(II17475), .B(II17476), .Z(g16119) ) ;
AND2    gate13220  (.A(g1111), .B(g16119), .Z(g19651) ) ;
AND2    gate13221  (.A(g2729), .B(g16966), .Z(g19655) ) ;
AND2    gate13222  (.A(g2807), .B(g15844), .Z(g19656) ) ;
NAND2   gate13223  (.A(II14854), .B(II14855), .Z(g12001) ) ;
AND2    gate13224  (.A(g12001), .B(g16968), .Z(g19660) ) ;
AND2    gate13225  (.A(g5489), .B(g16969), .Z(g19661) ) ;
NAND2   gate13226  (.A(II17495), .B(II17496), .Z(g16155) ) ;
AND2    gate13227  (.A(g1454), .B(g16155), .Z(g19671) ) ;
AND2    gate13228  (.A(g2819), .B(g15867), .Z(g19674) ) ;
NAND2   gate13229  (.A(II14884), .B(II14885), .Z(g12028) ) ;
AND2    gate13230  (.A(g12028), .B(g17013), .Z(g19680) ) ;
AND2    gate13231  (.A(g5835), .B(g17014), .Z(g19681) ) ;
AND2    gate13232  (.A(g2735), .B(g17297), .Z(g19684) ) ;
AND2    gate13233  (.A(g9614), .B(g17085), .Z(g19691) ) ;
NAND2   gate13234  (.A(II14924), .B(II14925), .Z(g12066) ) ;
AND2    gate13235  (.A(g12066), .B(g17086), .Z(g19692) ) ;
AND2    gate13236  (.A(g6181), .B(g17087), .Z(g19693) ) ;
AND2    gate13237  (.A(g9679), .B(g17120), .Z(g19715) ) ;
NAND2   gate13238  (.A(II14956), .B(II14957), .Z(g12100) ) ;
AND2    gate13239  (.A(g12100), .B(g17121), .Z(g19716) ) ;
AND2    gate13240  (.A(g6527), .B(g17122), .Z(g19717) ) ;
AND2    gate13241  (.A(g9740), .B(g17135), .Z(g19735) ) ;
NAND2   gate13242  (.A(II14992), .B(II14993), .Z(g12136) ) ;
AND2    gate13243  (.A(g12136), .B(g17136), .Z(g19736) ) ;
AND2    gate13244  (.A(g2783), .B(g15907), .Z(g19740) ) ;
AND2    gate13245  (.A(g9816), .B(g17147), .Z(g19746) ) ;
AND2    gate13246  (.A(g732), .B(g16646), .Z(g19749) ) ;
AND2    gate13247  (.A(g2771), .B(g15864), .Z(g19752) ) ;
AND2    gate13248  (.A(g9899), .B(g17154), .Z(g19756) ) ;
OR2     gate13249  (.A(g13461), .B(g11032), .Z(g16810) ) ;
AND2    gate13250  (.A(g16810), .B(g14203), .Z(g19767) ) ;
AND2    gate13251  (.A(g2803), .B(g15833), .Z(g19768) ) ;
AND2    gate13252  (.A(g2775), .B(g15877), .Z(g19784) ) ;
AND2    gate13253  (.A(g9983), .B(g17216), .Z(g19788) ) ;
NOR3    gate13254  (.A(g10032), .B(g12259), .C(g9217), .Z(g14253) ) ;
AND2    gate13255  (.A(g14253), .B(g17189), .Z(g19791) ) ;
AND2    gate13256  (.A(g2787), .B(g15962), .Z(g19855) ) ;
NOR2    gate13257  (.A(g10143), .B(g12259), .Z(g14707) ) ;
AND2    gate13258  (.A(g14707), .B(g17748), .Z(g19911) ) ;
AND2    gate13259  (.A(g2815), .B(g15853), .Z(g19914) ) ;
NOR2    gate13260  (.A(g13221), .B(g10828), .Z(g17515) ) ;
AND2    gate13261  (.A(g17515), .B(g16320), .Z(g19948) ) ;
NAND2   gate13262  (.A(g13551), .B(g13545), .Z(g16291) ) ;
AND4    gate13263  (.A(g16291), .B(g9007), .C(g8954), .D(g8903), .Z(g20056) ) ;
NAND2   gate13264  (.A(g13580), .B(g13574), .Z(g16312) ) ;
AND4    gate13265  (.A(g16312), .B(g9051), .C(g9011), .D(g8955), .Z(g20069) ) ;
NAND2   gate13266  (.A(II14531), .B(II14532), .Z(g11591) ) ;
AND2    gate13267  (.A(g11591), .B(g16609), .Z(g20084) ) ;
NOR2    gate13268  (.A(g817), .B(g14279), .Z(g15372) ) ;
AND2    gate13269  (.A(g15372), .B(g14584), .Z(g20093) ) ;
AND2    gate13270  (.A(g8872), .B(g16631), .Z(g20094) ) ;
NAND2   gate13271  (.A(II12849), .B(II12850), .Z(g8873) ) ;
AND2    gate13272  (.A(g8873), .B(g16632), .Z(g20095) ) ;
NOR2    gate13273  (.A(g10320), .B(g14279), .Z(g15508) ) ;
AND2    gate13274  (.A(g15508), .B(g11048), .Z(g20108) ) ;
NOR2    gate13275  (.A(g832), .B(g14279), .Z(g17954) ) ;
AND2    gate13276  (.A(g17954), .B(g17616), .Z(g20109) ) ;
OR2     gate13277  (.A(g10822), .B(g10827), .Z(g13540) ) ;
AND2    gate13278  (.A(g13540), .B(g16661), .Z(g20112) ) ;
NOR2    gate13279  (.A(g7118), .B(g14279), .Z(g15170) ) ;
AND2    gate13280  (.A(g15170), .B(g14309), .Z(g20131) ) ;
OR2     gate13281  (.A(g13247), .B(g10856), .Z(g16258) ) ;
AND2    gate13282  (.A(g16258), .B(g16695), .Z(g20135) ) ;
NAND2   gate13283  (.A(II14498), .B(II14499), .Z(g11545) ) ;
AND2    gate13284  (.A(g11545), .B(g16727), .Z(g20152) ) ;
NAND2   gate13285  (.A(II12729), .B(II12730), .Z(g8737) ) ;
AND2    gate13286  (.A(g8737), .B(g16750), .Z(g20162) ) ;
AND2    gate13287  (.A(g5156), .B(g17733), .Z(g20165) ) ;
NOR2    gate13288  (.A(g14719), .B(g12490), .Z(g16479) ) ;
AND2    gate13289  (.A(g16479), .B(g10476), .Z(g20171) ) ;
AND2    gate13290  (.A(g5503), .B(g17754), .Z(g20174) ) ;
AND2    gate13291  (.A(g5849), .B(g17772), .Z(g20188) ) ;
NOR2    gate13292  (.A(g7216), .B(g14279), .Z(g15578) ) ;
AND2    gate13293  (.A(g15578), .B(g17264), .Z(g20193) ) ;
AND2    gate13294  (.A(g6195), .B(g17789), .Z(g20203) ) ;
AND2    gate13295  (.A(g16479), .B(g10476), .Z(g20215) ) ;
AND2    gate13296  (.A(g6541), .B(g17815), .Z(g20218) ) ;
AND2    gate13297  (.A(g336), .B(g15831), .Z(g20559) ) ;
NOR2    gate13298  (.A(g1041), .B(g7479), .Z(g10801) ) ;
AND2    gate13299  (.A(g10801), .B(g15571), .Z(g20581) ) ;
NOR2    gate13300  (.A(g1384), .B(g7503), .Z(g10803) ) ;
AND2    gate13301  (.A(g10803), .B(g15580), .Z(g20602) ) ;
AND2    gate13302  (.A(g1046), .B(g15789), .Z(g20628) ) ;
AND2    gate13303  (.A(g1389), .B(g15800), .Z(g20658) ) ;
NAND3   gate13304  (.A(g4698), .B(g13883), .C(g12054), .Z(g16238) ) ;
NAND3   gate13305  (.A(g4743), .B(g13908), .C(g12054), .Z(g16259) ) ;
NAND3   gate13306  (.A(g4888), .B(g13910), .C(g12088), .Z(g16260) ) ;
NAND3   gate13307  (.A(g4754), .B(g13937), .C(g12054), .Z(g16281) ) ;
NAND3   gate13308  (.A(g4933), .B(g13939), .C(g12088), .Z(g16282) ) ;
NOR2    gate13309  (.A(g4294), .B(g4297), .Z(g10123) ) ;
AND2    gate13310  (.A(g10123), .B(g17301), .Z(g20977) ) ;
NAND3   gate13311  (.A(g4765), .B(g13970), .C(g12054), .Z(g16304) ) ;
NAND3   gate13312  (.A(g4944), .B(g13971), .C(g12088), .Z(g16306) ) ;
AND2    gate13313  (.A(g10043), .B(g17625), .Z(g21066) ) ;
AND2    gate13314  (.A(g10085), .B(g17625), .Z(g21067) ) ;
NAND3   gate13315  (.A(g4955), .B(g13996), .C(g12088), .Z(g16321) ) ;
AND2    gate13316  (.A(g7666), .B(g15705), .Z(g21188) ) ;
OR2     gate13317  (.A(g11448), .B(g8913), .Z(g13969) ) ;
AND2    gate13318  (.A(g13969), .B(g17470), .Z(g21251) ) ;
AND2    gate13319  (.A(g10157), .B(g17625), .Z(g21276) ) ;
NAND2   gate13320  (.A(II12241), .B(II12242), .Z(g7857) ) ;
AND2    gate13321  (.A(g7857), .B(g16027), .Z(g21285) ) ;
NAND2   gate13322  (.A(II12262), .B(II12263), .Z(g7879) ) ;
AND2    gate13323  (.A(g7879), .B(g16072), .Z(g21296) ) ;
AND2    gate13324  (.A(g7697), .B(g15825), .Z(g21298) ) ;
AND2    gate13325  (.A(g956), .B(g15731), .Z(g21302) ) ;
AND2    gate13326  (.A(g10120), .B(g17625), .Z(g21303) ) ;
AND2    gate13327  (.A(g996), .B(g15739), .Z(g21332) ) ;
AND2    gate13328  (.A(g1300), .B(g15740), .Z(g21333) ) ;
AND2    gate13329  (.A(g1339), .B(g15750), .Z(g21347) ) ;
AND2    gate13330  (.A(g10121), .B(g17625), .Z(g21348) ) ;
NAND2   gate13331  (.A(II12252), .B(II12253), .Z(g7869) ) ;
AND2    gate13332  (.A(g7869), .B(g16066), .Z(g21361) ) ;
NAND2   gate13333  (.A(II12278), .B(II12279), .Z(g7887) ) ;
AND2    gate13334  (.A(g7887), .B(g16090), .Z(g21378) ) ;
AND2    gate13335  (.A(g10086), .B(g17625), .Z(g21382) ) ;
NOR2    gate13336  (.A(g7851), .B(g10741), .Z(g13335) ) ;
AND2    gate13337  (.A(g13335), .B(g15799), .Z(g21394) ) ;
AND2    gate13338  (.A(g16069), .B(g13569), .Z(g21404) ) ;
NOR2    gate13339  (.A(g7873), .B(g10762), .Z(g13377) ) ;
AND2    gate13340  (.A(g13377), .B(g15811), .Z(g21405) ) ;
AND2    gate13341  (.A(g16681), .B(g13595), .Z(g21419) ) ;
AND2    gate13342  (.A(g16093), .B(g13596), .Z(g21420) ) ;
AND2    gate13343  (.A(g16119), .B(g13624), .Z(g21452) ) ;
AND2    gate13344  (.A(g16713), .B(g13625), .Z(g21453) ) ;
NAND4   gate13345  (.A(g13475), .B(g13495), .C(g13057), .D(g13459), .Z(g16181) ) ;
AND2    gate13346  (.A(g16181), .B(g10872), .Z(g21464) ) ;
AND2    gate13347  (.A(g16155), .B(g13663), .Z(g21465) ) ;
NAND3   gate13348  (.A(g13544), .B(g13528), .C(g13043), .Z(g16225) ) ;
AND2    gate13349  (.A(g16225), .B(g10881), .Z(g21512) ) ;
NAND4   gate13350  (.A(g13496), .B(g13513), .C(g13079), .D(g13476), .Z(g16196) ) ;
AND2    gate13351  (.A(g16196), .B(g10882), .Z(g21513) ) ;
NOR2    gate13352  (.A(g7909), .B(g10741), .Z(g12980) ) ;
AND2    gate13353  (.A(g12980), .B(g15674), .Z(g21557) ) ;
AND2    gate13354  (.A(g15904), .B(g13729), .Z(g21558) ) ;
NAND3   gate13355  (.A(g13573), .B(g13554), .C(g13058), .Z(g16236) ) ;
AND2    gate13356  (.A(g16236), .B(g10897), .Z(g21559) ) ;
NOR2    gate13357  (.A(g7939), .B(g10762), .Z(g13005) ) ;
AND2    gate13358  (.A(g13005), .B(g15695), .Z(g21605) ) ;
AND2    gate13359  (.A(g15959), .B(g13763), .Z(g21606) ) ;
AND2    gate13360  (.A(g142), .B(g20283), .Z(g21699) ) ;
AND2    gate13361  (.A(g150), .B(g20283), .Z(g21700) ) ;
AND2    gate13362  (.A(g153), .B(g20283), .Z(g21701) ) ;
AND2    gate13363  (.A(g157), .B(g20283), .Z(g21702) ) ;
AND2    gate13364  (.A(g146), .B(g20283), .Z(g21703) ) ;
AND2    gate13365  (.A(g164), .B(g20283), .Z(g21704) ) ;
AND2    gate13366  (.A(g209), .B(g20283), .Z(g21705) ) ;
AND2    gate13367  (.A(g222), .B(g20283), .Z(g21706) ) ;
AND2    gate13368  (.A(g191), .B(g20283), .Z(g21707) ) ;
NOR2    gate13369  (.A(g13350), .B(g6799), .Z(g15049) ) ;
AND2    gate13370  (.A(g15049), .B(g20283), .Z(g21708) ) ;
AND2    gate13371  (.A(g283), .B(g20283), .Z(g21709) ) ;
AND2    gate13372  (.A(g287), .B(g20283), .Z(g21710) ) ;
AND2    gate13373  (.A(g291), .B(g20283), .Z(g21711) ) ;
AND2    gate13374  (.A(g294), .B(g20283), .Z(g21712) ) ;
AND2    gate13375  (.A(g298), .B(g20283), .Z(g21713) ) ;
AND2    gate13376  (.A(g278), .B(g20283), .Z(g21714) ) ;
AND2    gate13377  (.A(g160), .B(g20283), .Z(g21715) ) ;
AND2    gate13378  (.A(g301), .B(g20283), .Z(g21716) ) ;
NOR2    gate13379  (.A(g6801), .B(g13350), .Z(g15051) ) ;
AND2    gate13380  (.A(g15051), .B(g21037), .Z(g21717) ) ;
AND2    gate13381  (.A(g370), .B(g21037), .Z(g21718) ) ;
AND2    gate13382  (.A(g358), .B(g21037), .Z(g21719) ) ;
AND2    gate13383  (.A(g376), .B(g21037), .Z(g21720) ) ;
AND2    gate13384  (.A(g385), .B(g21037), .Z(g21721) ) ;
AND2    gate13385  (.A(g3010), .B(g20330), .Z(g21728) ) ;
AND2    gate13386  (.A(g3021), .B(g20330), .Z(g21729) ) ;
AND2    gate13387  (.A(g3025), .B(g20330), .Z(g21730) ) ;
AND2    gate13388  (.A(g3029), .B(g20330), .Z(g21731) ) ;
AND2    gate13389  (.A(g3004), .B(g20330), .Z(g21732) ) ;
AND2    gate13390  (.A(g3034), .B(g20330), .Z(g21733) ) ;
AND2    gate13391  (.A(g3040), .B(g20330), .Z(g21734) ) ;
AND2    gate13392  (.A(g3057), .B(g20330), .Z(g21735) ) ;
AND2    gate13393  (.A(g3065), .B(g20330), .Z(g21736) ) ;
AND2    gate13394  (.A(g3068), .B(g20330), .Z(g21737) ) ;
AND2    gate13395  (.A(g3072), .B(g20330), .Z(g21738) ) ;
AND2    gate13396  (.A(g3080), .B(g20330), .Z(g21739) ) ;
AND2    gate13397  (.A(g3085), .B(g20330), .Z(g21740) ) ;
NOR2    gate13398  (.A(g13144), .B(g12859), .Z(g15086) ) ;
AND2    gate13399  (.A(g15086), .B(g20330), .Z(g21741) ) ;
AND2    gate13400  (.A(g3050), .B(g20330), .Z(g21742) ) ;
AND2    gate13401  (.A(g3100), .B(g20330), .Z(g21743) ) ;
AND2    gate13402  (.A(g3103), .B(g20330), .Z(g21744) ) ;
AND2    gate13403  (.A(g3017), .B(g20330), .Z(g21745) ) ;
AND2    gate13404  (.A(g3045), .B(g20330), .Z(g21746) ) ;
AND2    gate13405  (.A(g3061), .B(g20330), .Z(g21747) ) ;
NOR2    gate13406  (.A(g13144), .B(g12861), .Z(g15089) ) ;
AND2    gate13407  (.A(g15089), .B(g20785), .Z(g21748) ) ;
AND2    gate13408  (.A(g3155), .B(g20785), .Z(g21749) ) ;
AND2    gate13409  (.A(g3161), .B(g20785), .Z(g21750) ) ;
AND2    gate13410  (.A(g3167), .B(g20785), .Z(g21751) ) ;
AND2    gate13411  (.A(g3171), .B(g20785), .Z(g21752) ) ;
AND2    gate13412  (.A(g3179), .B(g20785), .Z(g21753) ) ;
AND2    gate13413  (.A(g3195), .B(g20785), .Z(g21754) ) ;
AND2    gate13414  (.A(g3203), .B(g20785), .Z(g21755) ) ;
AND2    gate13415  (.A(g3211), .B(g20785), .Z(g21756) ) ;
AND2    gate13416  (.A(g3187), .B(g20785), .Z(g21757) ) ;
AND2    gate13417  (.A(g3191), .B(g20785), .Z(g21758) ) ;
AND2    gate13418  (.A(g3199), .B(g20785), .Z(g21759) ) ;
AND2    gate13419  (.A(g3207), .B(g20785), .Z(g21760) ) ;
AND2    gate13420  (.A(g3215), .B(g20785), .Z(g21761) ) ;
AND2    gate13421  (.A(g3219), .B(g20785), .Z(g21762) ) ;
AND2    gate13422  (.A(g3223), .B(g20785), .Z(g21763) ) ;
AND2    gate13423  (.A(g3227), .B(g20785), .Z(g21764) ) ;
AND2    gate13424  (.A(g3231), .B(g20785), .Z(g21765) ) ;
AND2    gate13425  (.A(g3235), .B(g20785), .Z(g21766) ) ;
AND2    gate13426  (.A(g3239), .B(g20785), .Z(g21767) ) ;
AND2    gate13427  (.A(g3243), .B(g20785), .Z(g21768) ) ;
AND2    gate13428  (.A(g3247), .B(g20785), .Z(g21769) ) ;
AND2    gate13429  (.A(g3251), .B(g20785), .Z(g21770) ) ;
AND2    gate13430  (.A(g3255), .B(g20785), .Z(g21771) ) ;
AND2    gate13431  (.A(g3259), .B(g20785), .Z(g21772) ) ;
AND2    gate13432  (.A(g3263), .B(g20785), .Z(g21773) ) ;
AND2    gate13433  (.A(g3361), .B(g20391), .Z(g21774) ) ;
AND2    gate13434  (.A(g3372), .B(g20391), .Z(g21775) ) ;
AND2    gate13435  (.A(g3376), .B(g20391), .Z(g21776) ) ;
AND2    gate13436  (.A(g3380), .B(g20391), .Z(g21777) ) ;
AND2    gate13437  (.A(g3355), .B(g20391), .Z(g21778) ) ;
AND2    gate13438  (.A(g3385), .B(g20391), .Z(g21779) ) ;
AND2    gate13439  (.A(g3391), .B(g20391), .Z(g21780) ) ;
AND2    gate13440  (.A(g3408), .B(g20391), .Z(g21781) ) ;
AND2    gate13441  (.A(g3416), .B(g20391), .Z(g21782) ) ;
AND2    gate13442  (.A(g3419), .B(g20391), .Z(g21783) ) ;
AND2    gate13443  (.A(g3423), .B(g20391), .Z(g21784) ) ;
AND2    gate13444  (.A(g3431), .B(g20391), .Z(g21785) ) ;
AND2    gate13445  (.A(g3436), .B(g20391), .Z(g21786) ) ;
NOR2    gate13446  (.A(g13177), .B(g12863), .Z(g15091) ) ;
AND2    gate13447  (.A(g15091), .B(g20391), .Z(g21787) ) ;
AND2    gate13448  (.A(g3401), .B(g20391), .Z(g21788) ) ;
AND2    gate13449  (.A(g3451), .B(g20391), .Z(g21789) ) ;
AND2    gate13450  (.A(g3454), .B(g20391), .Z(g21790) ) ;
AND2    gate13451  (.A(g3368), .B(g20391), .Z(g21791) ) ;
AND2    gate13452  (.A(g3396), .B(g20391), .Z(g21792) ) ;
AND2    gate13453  (.A(g3412), .B(g20391), .Z(g21793) ) ;
NOR2    gate13454  (.A(g13177), .B(g12865), .Z(g15094) ) ;
AND2    gate13455  (.A(g15094), .B(g20924), .Z(g21794) ) ;
AND2    gate13456  (.A(g3506), .B(g20924), .Z(g21795) ) ;
AND2    gate13457  (.A(g3512), .B(g20924), .Z(g21796) ) ;
AND2    gate13458  (.A(g3518), .B(g20924), .Z(g21797) ) ;
AND2    gate13459  (.A(g3522), .B(g20924), .Z(g21798) ) ;
AND2    gate13460  (.A(g3530), .B(g20924), .Z(g21799) ) ;
AND2    gate13461  (.A(g3546), .B(g20924), .Z(g21800) ) ;
AND2    gate13462  (.A(g3554), .B(g20924), .Z(g21801) ) ;
AND2    gate13463  (.A(g3562), .B(g20924), .Z(g21802) ) ;
AND2    gate13464  (.A(g3538), .B(g20924), .Z(g21803) ) ;
AND2    gate13465  (.A(g3542), .B(g20924), .Z(g21804) ) ;
AND2    gate13466  (.A(g3550), .B(g20924), .Z(g21805) ) ;
AND2    gate13467  (.A(g3558), .B(g20924), .Z(g21806) ) ;
AND2    gate13468  (.A(g3566), .B(g20924), .Z(g21807) ) ;
AND2    gate13469  (.A(g3570), .B(g20924), .Z(g21808) ) ;
AND2    gate13470  (.A(g3574), .B(g20924), .Z(g21809) ) ;
AND2    gate13471  (.A(g3578), .B(g20924), .Z(g21810) ) ;
AND2    gate13472  (.A(g3582), .B(g20924), .Z(g21811) ) ;
AND2    gate13473  (.A(g3586), .B(g20924), .Z(g21812) ) ;
AND2    gate13474  (.A(g3590), .B(g20924), .Z(g21813) ) ;
AND2    gate13475  (.A(g3594), .B(g20924), .Z(g21814) ) ;
AND2    gate13476  (.A(g3598), .B(g20924), .Z(g21815) ) ;
AND2    gate13477  (.A(g3602), .B(g20924), .Z(g21816) ) ;
AND2    gate13478  (.A(g3606), .B(g20924), .Z(g21817) ) ;
AND2    gate13479  (.A(g3610), .B(g20924), .Z(g21818) ) ;
AND2    gate13480  (.A(g3614), .B(g20924), .Z(g21819) ) ;
AND2    gate13481  (.A(g3712), .B(g20453), .Z(g21820) ) ;
AND2    gate13482  (.A(g3723), .B(g20453), .Z(g21821) ) ;
AND2    gate13483  (.A(g3727), .B(g20453), .Z(g21822) ) ;
AND2    gate13484  (.A(g3731), .B(g20453), .Z(g21823) ) ;
AND2    gate13485  (.A(g3706), .B(g20453), .Z(g21824) ) ;
AND2    gate13486  (.A(g3736), .B(g20453), .Z(g21825) ) ;
AND2    gate13487  (.A(g3742), .B(g20453), .Z(g21826) ) ;
AND2    gate13488  (.A(g3759), .B(g20453), .Z(g21827) ) ;
AND2    gate13489  (.A(g3767), .B(g20453), .Z(g21828) ) ;
AND2    gate13490  (.A(g3770), .B(g20453), .Z(g21829) ) ;
AND2    gate13491  (.A(g3774), .B(g20453), .Z(g21830) ) ;
AND2    gate13492  (.A(g3782), .B(g20453), .Z(g21831) ) ;
AND2    gate13493  (.A(g3787), .B(g20453), .Z(g21832) ) ;
NOR2    gate13494  (.A(g13191), .B(g12867), .Z(g15096) ) ;
AND2    gate13495  (.A(g15096), .B(g20453), .Z(g21833) ) ;
AND2    gate13496  (.A(g3752), .B(g20453), .Z(g21834) ) ;
AND2    gate13497  (.A(g3802), .B(g20453), .Z(g21835) ) ;
AND2    gate13498  (.A(g3805), .B(g20453), .Z(g21836) ) ;
AND2    gate13499  (.A(g3719), .B(g20453), .Z(g21837) ) ;
AND2    gate13500  (.A(g3747), .B(g20453), .Z(g21838) ) ;
AND2    gate13501  (.A(g3763), .B(g20453), .Z(g21839) ) ;
NOR2    gate13502  (.A(g13191), .B(g12869), .Z(g15099) ) ;
AND2    gate13503  (.A(g15099), .B(g21070), .Z(g21840) ) ;
AND2    gate13504  (.A(g3857), .B(g21070), .Z(g21841) ) ;
AND2    gate13505  (.A(g3863), .B(g21070), .Z(g21842) ) ;
AND2    gate13506  (.A(g3869), .B(g21070), .Z(g21843) ) ;
AND2    gate13507  (.A(g3873), .B(g21070), .Z(g21844) ) ;
AND2    gate13508  (.A(g3881), .B(g21070), .Z(g21845) ) ;
AND2    gate13509  (.A(g3897), .B(g21070), .Z(g21846) ) ;
AND2    gate13510  (.A(g3905), .B(g21070), .Z(g21847) ) ;
AND2    gate13511  (.A(g3913), .B(g21070), .Z(g21848) ) ;
AND2    gate13512  (.A(g3889), .B(g21070), .Z(g21849) ) ;
AND2    gate13513  (.A(g3893), .B(g21070), .Z(g21850) ) ;
AND2    gate13514  (.A(g3901), .B(g21070), .Z(g21851) ) ;
AND2    gate13515  (.A(g3909), .B(g21070), .Z(g21852) ) ;
AND2    gate13516  (.A(g3917), .B(g21070), .Z(g21853) ) ;
AND2    gate13517  (.A(g3921), .B(g21070), .Z(g21854) ) ;
AND2    gate13518  (.A(g3925), .B(g21070), .Z(g21855) ) ;
AND2    gate13519  (.A(g3929), .B(g21070), .Z(g21856) ) ;
AND2    gate13520  (.A(g3933), .B(g21070), .Z(g21857) ) ;
AND2    gate13521  (.A(g3937), .B(g21070), .Z(g21858) ) ;
AND2    gate13522  (.A(g3941), .B(g21070), .Z(g21859) ) ;
AND2    gate13523  (.A(g3945), .B(g21070), .Z(g21860) ) ;
AND2    gate13524  (.A(g3949), .B(g21070), .Z(g21861) ) ;
AND2    gate13525  (.A(g3953), .B(g21070), .Z(g21862) ) ;
AND2    gate13526  (.A(g3957), .B(g21070), .Z(g21863) ) ;
AND2    gate13527  (.A(g3961), .B(g21070), .Z(g21864) ) ;
AND2    gate13528  (.A(g3965), .B(g21070), .Z(g21865) ) ;
AND2    gate13529  (.A(g4072), .B(g19801), .Z(g21866) ) ;
AND2    gate13530  (.A(g4082), .B(g19801), .Z(g21867) ) ;
AND2    gate13531  (.A(g4076), .B(g19801), .Z(g21868) ) ;
AND2    gate13532  (.A(g4087), .B(g19801), .Z(g21869) ) ;
AND2    gate13533  (.A(g4093), .B(g19801), .Z(g21870) ) ;
AND2    gate13534  (.A(g4108), .B(g19801), .Z(g21871) ) ;
AND2    gate13535  (.A(g4098), .B(g19801), .Z(g21872) ) ;
AND2    gate13536  (.A(g6946), .B(g19801), .Z(g21873) ) ;
AND2    gate13537  (.A(g4112), .B(g19801), .Z(g21874) ) ;
AND2    gate13538  (.A(g4116), .B(g19801), .Z(g21875) ) ;
AND2    gate13539  (.A(g4119), .B(g19801), .Z(g21876) ) ;
AND2    gate13540  (.A(g6888), .B(g19801), .Z(g21877) ) ;
AND2    gate13541  (.A(g4129), .B(g19801), .Z(g21878) ) ;
AND2    gate13542  (.A(g4132), .B(g19801), .Z(g21879) ) ;
AND2    gate13543  (.A(g4135), .B(g19801), .Z(g21880) ) ;
AND2    gate13544  (.A(g4064), .B(g19801), .Z(g21881) ) ;
AND2    gate13545  (.A(g4057), .B(g19801), .Z(g21882) ) ;
AND2    gate13546  (.A(g4141), .B(g19801), .Z(g21883) ) ;
AND2    gate13547  (.A(g4104), .B(g19801), .Z(g21884) ) ;
AND2    gate13548  (.A(g4122), .B(g19801), .Z(g21885) ) ;
AND2    gate13549  (.A(g4153), .B(g19801), .Z(g21886) ) ;
NOR2    gate13550  (.A(g12871), .B(g14591), .Z(g15101) ) ;
AND2    gate13551  (.A(g15101), .B(g19801), .Z(g21887) ) ;
AND2    gate13552  (.A(g4165), .B(g19801), .Z(g21888) ) ;
AND2    gate13553  (.A(g4169), .B(g19801), .Z(g21889) ) ;
AND2    gate13554  (.A(g4125), .B(g19801), .Z(g21890) ) ;
AND2    gate13555  (.A(g5022), .B(g21468), .Z(g21906) ) ;
AND2    gate13556  (.A(g5033), .B(g21468), .Z(g21907) ) ;
AND2    gate13557  (.A(g5037), .B(g21468), .Z(g21908) ) ;
AND2    gate13558  (.A(g5041), .B(g21468), .Z(g21909) ) ;
AND2    gate13559  (.A(g5016), .B(g21468), .Z(g21910) ) ;
AND2    gate13560  (.A(g5046), .B(g21468), .Z(g21911) ) ;
AND2    gate13561  (.A(g5052), .B(g21468), .Z(g21912) ) ;
AND2    gate13562  (.A(g5069), .B(g21468), .Z(g21913) ) ;
AND2    gate13563  (.A(g5077), .B(g21468), .Z(g21914) ) ;
AND2    gate13564  (.A(g5080), .B(g21468), .Z(g21915) ) ;
AND2    gate13565  (.A(g5084), .B(g21468), .Z(g21916) ) ;
AND2    gate13566  (.A(g5092), .B(g21468), .Z(g21917) ) ;
AND2    gate13567  (.A(g5097), .B(g21468), .Z(g21918) ) ;
NOR2    gate13568  (.A(g13716), .B(g12890), .Z(g15144) ) ;
AND2    gate13569  (.A(g15144), .B(g21468), .Z(g21919) ) ;
AND2    gate13570  (.A(g5062), .B(g21468), .Z(g21920) ) ;
AND2    gate13571  (.A(g5109), .B(g21468), .Z(g21921) ) ;
AND2    gate13572  (.A(g5112), .B(g21468), .Z(g21922) ) ;
AND2    gate13573  (.A(g5029), .B(g21468), .Z(g21923) ) ;
AND2    gate13574  (.A(g5057), .B(g21468), .Z(g21924) ) ;
AND2    gate13575  (.A(g5073), .B(g21468), .Z(g21925) ) ;
NOR2    gate13576  (.A(g13716), .B(g12892), .Z(g15147) ) ;
AND2    gate13577  (.A(g15147), .B(g18997), .Z(g21926) ) ;
AND2    gate13578  (.A(g5164), .B(g18997), .Z(g21927) ) ;
AND2    gate13579  (.A(g5170), .B(g18997), .Z(g21928) ) ;
AND2    gate13580  (.A(g5176), .B(g18997), .Z(g21929) ) ;
AND2    gate13581  (.A(g5180), .B(g18997), .Z(g21930) ) ;
AND2    gate13582  (.A(g5188), .B(g18997), .Z(g21931) ) ;
AND2    gate13583  (.A(g5204), .B(g18997), .Z(g21932) ) ;
AND2    gate13584  (.A(g5212), .B(g18997), .Z(g21933) ) ;
AND2    gate13585  (.A(g5220), .B(g18997), .Z(g21934) ) ;
AND2    gate13586  (.A(g5196), .B(g18997), .Z(g21935) ) ;
AND2    gate13587  (.A(g5200), .B(g18997), .Z(g21936) ) ;
AND2    gate13588  (.A(g5208), .B(g18997), .Z(g21937) ) ;
AND2    gate13589  (.A(g5216), .B(g18997), .Z(g21938) ) ;
AND2    gate13590  (.A(g5224), .B(g18997), .Z(g21939) ) ;
AND2    gate13591  (.A(g5228), .B(g18997), .Z(g21940) ) ;
AND2    gate13592  (.A(g5232), .B(g18997), .Z(g21941) ) ;
AND2    gate13593  (.A(g5236), .B(g18997), .Z(g21942) ) ;
AND2    gate13594  (.A(g5240), .B(g18997), .Z(g21943) ) ;
AND2    gate13595  (.A(g5244), .B(g18997), .Z(g21944) ) ;
AND2    gate13596  (.A(g5248), .B(g18997), .Z(g21945) ) ;
AND2    gate13597  (.A(g5252), .B(g18997), .Z(g21946) ) ;
AND2    gate13598  (.A(g5256), .B(g18997), .Z(g21947) ) ;
AND2    gate13599  (.A(g5260), .B(g18997), .Z(g21948) ) ;
AND2    gate13600  (.A(g5264), .B(g18997), .Z(g21949) ) ;
AND2    gate13601  (.A(g5268), .B(g18997), .Z(g21950) ) ;
AND2    gate13602  (.A(g5272), .B(g18997), .Z(g21951) ) ;
AND2    gate13603  (.A(g5366), .B(g21514), .Z(g21952) ) ;
AND2    gate13604  (.A(g5377), .B(g21514), .Z(g21953) ) ;
AND2    gate13605  (.A(g5381), .B(g21514), .Z(g21954) ) ;
AND2    gate13606  (.A(g5385), .B(g21514), .Z(g21955) ) ;
AND2    gate13607  (.A(g5360), .B(g21514), .Z(g21956) ) ;
AND2    gate13608  (.A(g5390), .B(g21514), .Z(g21957) ) ;
AND2    gate13609  (.A(g5396), .B(g21514), .Z(g21958) ) ;
AND2    gate13610  (.A(g5413), .B(g21514), .Z(g21959) ) ;
AND2    gate13611  (.A(g5421), .B(g21514), .Z(g21960) ) ;
AND2    gate13612  (.A(g5424), .B(g21514), .Z(g21961) ) ;
AND2    gate13613  (.A(g5428), .B(g21514), .Z(g21962) ) ;
AND2    gate13614  (.A(g5436), .B(g21514), .Z(g21963) ) ;
AND2    gate13615  (.A(g5441), .B(g21514), .Z(g21964) ) ;
NOR2    gate13616  (.A(g13745), .B(g12894), .Z(g15149) ) ;
AND2    gate13617  (.A(g15149), .B(g21514), .Z(g21965) ) ;
AND2    gate13618  (.A(g5406), .B(g21514), .Z(g21966) ) ;
AND2    gate13619  (.A(g5456), .B(g21514), .Z(g21967) ) ;
AND2    gate13620  (.A(g5459), .B(g21514), .Z(g21968) ) ;
AND2    gate13621  (.A(g5373), .B(g21514), .Z(g21969) ) ;
AND2    gate13622  (.A(g5401), .B(g21514), .Z(g21970) ) ;
AND2    gate13623  (.A(g5417), .B(g21514), .Z(g21971) ) ;
NOR2    gate13624  (.A(g13745), .B(g12896), .Z(g15152) ) ;
AND2    gate13625  (.A(g15152), .B(g19074), .Z(g21972) ) ;
AND2    gate13626  (.A(g5511), .B(g19074), .Z(g21973) ) ;
AND2    gate13627  (.A(g5517), .B(g19074), .Z(g21974) ) ;
AND2    gate13628  (.A(g5523), .B(g19074), .Z(g21975) ) ;
AND2    gate13629  (.A(g5527), .B(g19074), .Z(g21976) ) ;
AND2    gate13630  (.A(g5535), .B(g19074), .Z(g21977) ) ;
AND2    gate13631  (.A(g5551), .B(g19074), .Z(g21978) ) ;
AND2    gate13632  (.A(g5559), .B(g19074), .Z(g21979) ) ;
AND2    gate13633  (.A(g5567), .B(g19074), .Z(g21980) ) ;
AND2    gate13634  (.A(g5543), .B(g19074), .Z(g21981) ) ;
AND2    gate13635  (.A(g5547), .B(g19074), .Z(g21982) ) ;
AND2    gate13636  (.A(g5555), .B(g19074), .Z(g21983) ) ;
AND2    gate13637  (.A(g5563), .B(g19074), .Z(g21984) ) ;
AND2    gate13638  (.A(g5571), .B(g19074), .Z(g21985) ) ;
AND2    gate13639  (.A(g5575), .B(g19074), .Z(g21986) ) ;
AND2    gate13640  (.A(g5579), .B(g19074), .Z(g21987) ) ;
AND2    gate13641  (.A(g5583), .B(g19074), .Z(g21988) ) ;
AND2    gate13642  (.A(g5587), .B(g19074), .Z(g21989) ) ;
AND2    gate13643  (.A(g5591), .B(g19074), .Z(g21990) ) ;
AND2    gate13644  (.A(g5595), .B(g19074), .Z(g21991) ) ;
AND2    gate13645  (.A(g5599), .B(g19074), .Z(g21992) ) ;
AND2    gate13646  (.A(g5603), .B(g19074), .Z(g21993) ) ;
AND2    gate13647  (.A(g5607), .B(g19074), .Z(g21994) ) ;
AND2    gate13648  (.A(g5611), .B(g19074), .Z(g21995) ) ;
AND2    gate13649  (.A(g5615), .B(g19074), .Z(g21996) ) ;
AND2    gate13650  (.A(g5619), .B(g19074), .Z(g21997) ) ;
AND2    gate13651  (.A(g5712), .B(g21562), .Z(g21998) ) ;
AND2    gate13652  (.A(g5723), .B(g21562), .Z(g21999) ) ;
AND2    gate13653  (.A(g5727), .B(g21562), .Z(g22000) ) ;
AND2    gate13654  (.A(g5731), .B(g21562), .Z(g22001) ) ;
AND2    gate13655  (.A(g5706), .B(g21562), .Z(g22002) ) ;
AND2    gate13656  (.A(g5736), .B(g21562), .Z(g22003) ) ;
AND2    gate13657  (.A(g5742), .B(g21562), .Z(g22004) ) ;
AND2    gate13658  (.A(g5759), .B(g21562), .Z(g22005) ) ;
AND2    gate13659  (.A(g5767), .B(g21562), .Z(g22006) ) ;
AND2    gate13660  (.A(g5770), .B(g21562), .Z(g22007) ) ;
AND2    gate13661  (.A(g5774), .B(g21562), .Z(g22008) ) ;
AND2    gate13662  (.A(g5782), .B(g21562), .Z(g22009) ) ;
AND2    gate13663  (.A(g5787), .B(g21562), .Z(g22010) ) ;
NOR2    gate13664  (.A(g13782), .B(g12898), .Z(g15154) ) ;
AND2    gate13665  (.A(g15154), .B(g21562), .Z(g22011) ) ;
AND2    gate13666  (.A(g5752), .B(g21562), .Z(g22012) ) ;
AND2    gate13667  (.A(g5802), .B(g21562), .Z(g22013) ) ;
AND2    gate13668  (.A(g5805), .B(g21562), .Z(g22014) ) ;
AND2    gate13669  (.A(g5719), .B(g21562), .Z(g22015) ) ;
AND2    gate13670  (.A(g5747), .B(g21562), .Z(g22016) ) ;
AND2    gate13671  (.A(g5763), .B(g21562), .Z(g22017) ) ;
NOR2    gate13672  (.A(g13782), .B(g12900), .Z(g15157) ) ;
AND2    gate13673  (.A(g15157), .B(g19147), .Z(g22018) ) ;
AND2    gate13674  (.A(g5857), .B(g19147), .Z(g22019) ) ;
AND2    gate13675  (.A(g5863), .B(g19147), .Z(g22020) ) ;
AND2    gate13676  (.A(g5869), .B(g19147), .Z(g22021) ) ;
AND2    gate13677  (.A(g5873), .B(g19147), .Z(g22022) ) ;
AND2    gate13678  (.A(g5881), .B(g19147), .Z(g22023) ) ;
AND2    gate13679  (.A(g5897), .B(g19147), .Z(g22024) ) ;
AND2    gate13680  (.A(g5905), .B(g19147), .Z(g22025) ) ;
AND2    gate13681  (.A(g5913), .B(g19147), .Z(g22026) ) ;
AND2    gate13682  (.A(g5889), .B(g19147), .Z(g22027) ) ;
AND2    gate13683  (.A(g5893), .B(g19147), .Z(g22028) ) ;
AND2    gate13684  (.A(g5901), .B(g19147), .Z(g22029) ) ;
AND2    gate13685  (.A(g5909), .B(g19147), .Z(g22030) ) ;
AND2    gate13686  (.A(g5917), .B(g19147), .Z(g22031) ) ;
AND2    gate13687  (.A(g5921), .B(g19147), .Z(g22032) ) ;
AND2    gate13688  (.A(g5925), .B(g19147), .Z(g22033) ) ;
AND2    gate13689  (.A(g5929), .B(g19147), .Z(g22034) ) ;
AND2    gate13690  (.A(g5933), .B(g19147), .Z(g22035) ) ;
AND2    gate13691  (.A(g5937), .B(g19147), .Z(g22036) ) ;
AND2    gate13692  (.A(g5941), .B(g19147), .Z(g22037) ) ;
AND2    gate13693  (.A(g5945), .B(g19147), .Z(g22038) ) ;
AND2    gate13694  (.A(g5949), .B(g19147), .Z(g22039) ) ;
AND2    gate13695  (.A(g5953), .B(g19147), .Z(g22040) ) ;
AND2    gate13696  (.A(g5957), .B(g19147), .Z(g22041) ) ;
AND2    gate13697  (.A(g5961), .B(g19147), .Z(g22042) ) ;
AND2    gate13698  (.A(g5965), .B(g19147), .Z(g22043) ) ;
AND2    gate13699  (.A(g6058), .B(g21611), .Z(g22044) ) ;
AND2    gate13700  (.A(g6069), .B(g21611), .Z(g22045) ) ;
AND2    gate13701  (.A(g6073), .B(g21611), .Z(g22046) ) ;
AND2    gate13702  (.A(g6077), .B(g21611), .Z(g22047) ) ;
AND2    gate13703  (.A(g6052), .B(g21611), .Z(g22048) ) ;
AND2    gate13704  (.A(g6082), .B(g21611), .Z(g22049) ) ;
AND2    gate13705  (.A(g6088), .B(g21611), .Z(g22050) ) ;
AND2    gate13706  (.A(g6105), .B(g21611), .Z(g22051) ) ;
AND2    gate13707  (.A(g6113), .B(g21611), .Z(g22052) ) ;
AND2    gate13708  (.A(g6116), .B(g21611), .Z(g22053) ) ;
AND2    gate13709  (.A(g6120), .B(g21611), .Z(g22054) ) ;
AND2    gate13710  (.A(g6128), .B(g21611), .Z(g22055) ) ;
AND2    gate13711  (.A(g6133), .B(g21611), .Z(g22056) ) ;
NOR2    gate13712  (.A(g13809), .B(g12902), .Z(g15159) ) ;
AND2    gate13713  (.A(g15159), .B(g21611), .Z(g22057) ) ;
AND2    gate13714  (.A(g6098), .B(g21611), .Z(g22058) ) ;
AND2    gate13715  (.A(g6148), .B(g21611), .Z(g22059) ) ;
AND2    gate13716  (.A(g6151), .B(g21611), .Z(g22060) ) ;
AND2    gate13717  (.A(g6065), .B(g21611), .Z(g22061) ) ;
AND2    gate13718  (.A(g6093), .B(g21611), .Z(g22062) ) ;
AND2    gate13719  (.A(g6109), .B(g21611), .Z(g22063) ) ;
NOR2    gate13720  (.A(g13809), .B(g12904), .Z(g15162) ) ;
AND2    gate13721  (.A(g15162), .B(g19210), .Z(g22064) ) ;
AND2    gate13722  (.A(g6203), .B(g19210), .Z(g22065) ) ;
AND2    gate13723  (.A(g6209), .B(g19210), .Z(g22066) ) ;
AND2    gate13724  (.A(g6215), .B(g19210), .Z(g22067) ) ;
AND2    gate13725  (.A(g6219), .B(g19210), .Z(g22068) ) ;
AND2    gate13726  (.A(g6227), .B(g19210), .Z(g22069) ) ;
AND2    gate13727  (.A(g6243), .B(g19210), .Z(g22070) ) ;
AND2    gate13728  (.A(g6251), .B(g19210), .Z(g22071) ) ;
AND2    gate13729  (.A(g6259), .B(g19210), .Z(g22072) ) ;
AND2    gate13730  (.A(g6235), .B(g19210), .Z(g22073) ) ;
AND2    gate13731  (.A(g6239), .B(g19210), .Z(g22074) ) ;
AND2    gate13732  (.A(g6247), .B(g19210), .Z(g22075) ) ;
AND2    gate13733  (.A(g6255), .B(g19210), .Z(g22076) ) ;
AND2    gate13734  (.A(g6263), .B(g19210), .Z(g22077) ) ;
AND2    gate13735  (.A(g6267), .B(g19210), .Z(g22078) ) ;
AND2    gate13736  (.A(g6271), .B(g19210), .Z(g22079) ) ;
AND2    gate13737  (.A(g6275), .B(g19210), .Z(g22080) ) ;
AND2    gate13738  (.A(g6279), .B(g19210), .Z(g22081) ) ;
AND2    gate13739  (.A(g6283), .B(g19210), .Z(g22082) ) ;
AND2    gate13740  (.A(g6287), .B(g19210), .Z(g22083) ) ;
AND2    gate13741  (.A(g6291), .B(g19210), .Z(g22084) ) ;
AND2    gate13742  (.A(g6295), .B(g19210), .Z(g22085) ) ;
AND2    gate13743  (.A(g6299), .B(g19210), .Z(g22086) ) ;
AND2    gate13744  (.A(g6303), .B(g19210), .Z(g22087) ) ;
AND2    gate13745  (.A(g6307), .B(g19210), .Z(g22088) ) ;
AND2    gate13746  (.A(g6311), .B(g19210), .Z(g22089) ) ;
AND2    gate13747  (.A(g6404), .B(g18833), .Z(g22090) ) ;
AND2    gate13748  (.A(g6415), .B(g18833), .Z(g22091) ) ;
AND2    gate13749  (.A(g6419), .B(g18833), .Z(g22092) ) ;
AND2    gate13750  (.A(g6423), .B(g18833), .Z(g22093) ) ;
AND2    gate13751  (.A(g6398), .B(g18833), .Z(g22094) ) ;
AND2    gate13752  (.A(g6428), .B(g18833), .Z(g22095) ) ;
AND2    gate13753  (.A(g6434), .B(g18833), .Z(g22096) ) ;
AND2    gate13754  (.A(g6451), .B(g18833), .Z(g22097) ) ;
AND2    gate13755  (.A(g6459), .B(g18833), .Z(g22098) ) ;
AND2    gate13756  (.A(g6462), .B(g18833), .Z(g22099) ) ;
AND2    gate13757  (.A(g6466), .B(g18833), .Z(g22100) ) ;
AND2    gate13758  (.A(g6474), .B(g18833), .Z(g22101) ) ;
AND2    gate13759  (.A(g6479), .B(g18833), .Z(g22102) ) ;
NOR2    gate13760  (.A(g13835), .B(g12906), .Z(g15164) ) ;
AND2    gate13761  (.A(g15164), .B(g18833), .Z(g22103) ) ;
AND2    gate13762  (.A(g6444), .B(g18833), .Z(g22104) ) ;
AND2    gate13763  (.A(g6494), .B(g18833), .Z(g22105) ) ;
AND2    gate13764  (.A(g6497), .B(g18833), .Z(g22106) ) ;
AND2    gate13765  (.A(g6411), .B(g18833), .Z(g22107) ) ;
AND2    gate13766  (.A(g6439), .B(g18833), .Z(g22108) ) ;
AND2    gate13767  (.A(g6455), .B(g18833), .Z(g22109) ) ;
NOR2    gate13768  (.A(g13835), .B(g12908), .Z(g15167) ) ;
AND2    gate13769  (.A(g15167), .B(g19277), .Z(g22110) ) ;
AND2    gate13770  (.A(g6549), .B(g19277), .Z(g22111) ) ;
AND2    gate13771  (.A(g6555), .B(g19277), .Z(g22112) ) ;
AND2    gate13772  (.A(g6561), .B(g19277), .Z(g22113) ) ;
AND2    gate13773  (.A(g6565), .B(g19277), .Z(g22114) ) ;
AND2    gate13774  (.A(g6573), .B(g19277), .Z(g22115) ) ;
AND2    gate13775  (.A(g6589), .B(g19277), .Z(g22116) ) ;
AND2    gate13776  (.A(g6597), .B(g19277), .Z(g22117) ) ;
AND2    gate13777  (.A(g6605), .B(g19277), .Z(g22118) ) ;
AND2    gate13778  (.A(g6581), .B(g19277), .Z(g22119) ) ;
AND2    gate13779  (.A(g6585), .B(g19277), .Z(g22120) ) ;
AND2    gate13780  (.A(g6593), .B(g19277), .Z(g22121) ) ;
AND2    gate13781  (.A(g6601), .B(g19277), .Z(g22122) ) ;
AND2    gate13782  (.A(g6609), .B(g19277), .Z(g22123) ) ;
AND2    gate13783  (.A(g6613), .B(g19277), .Z(g22124) ) ;
AND2    gate13784  (.A(g6617), .B(g19277), .Z(g22125) ) ;
AND2    gate13785  (.A(g6621), .B(g19277), .Z(g22126) ) ;
AND2    gate13786  (.A(g6625), .B(g19277), .Z(g22127) ) ;
AND2    gate13787  (.A(g6629), .B(g19277), .Z(g22128) ) ;
AND2    gate13788  (.A(g6633), .B(g19277), .Z(g22129) ) ;
AND2    gate13789  (.A(g6637), .B(g19277), .Z(g22130) ) ;
AND2    gate13790  (.A(g6641), .B(g19277), .Z(g22131) ) ;
AND2    gate13791  (.A(g6645), .B(g19277), .Z(g22132) ) ;
AND2    gate13792  (.A(g6649), .B(g19277), .Z(g22133) ) ;
AND2    gate13793  (.A(g6653), .B(g19277), .Z(g22134) ) ;
AND2    gate13794  (.A(g6657), .B(g19277), .Z(g22135) ) ;
AND2    gate13795  (.A(g7957), .B(g19140), .Z(g22142) ) ;
AND2    gate13796  (.A(g19568), .B(g10971), .Z(g22143) ) ;
AND2    gate13797  (.A(g14555), .B(g18832), .Z(g22145) ) ;
AND2    gate13798  (.A(g14581), .B(g18880), .Z(g22149) ) ;
AND2    gate13799  (.A(g14608), .B(g18892), .Z(g22157) ) ;
NOR3    gate13800  (.A(g528), .B(g12527), .C(g11185), .Z(g13698) ) ;
AND2    gate13801  (.A(g13698), .B(g19609), .Z(g22158) ) ;
AND2    gate13802  (.A(g8005), .B(g19795), .Z(g22160) ) ;
NOR3    gate13803  (.A(g10614), .B(g13026), .C(g7285), .Z(g15594) ) ;
AND2    gate13804  (.A(g15594), .B(g18903), .Z(g22165) ) ;
AND2    gate13805  (.A(g8064), .B(g19857), .Z(g22172) ) ;
AND2    gate13806  (.A(g8119), .B(g19875), .Z(g22191) ) ;
NOR2    gate13807  (.A(g16201), .B(g13634), .Z(g19880) ) ;
AND2    gate13808  (.A(g19880), .B(g20682), .Z(g22193) ) ;
NOR2    gate13809  (.A(g16209), .B(g13672), .Z(g19906) ) ;
AND2    gate13810  (.A(g19906), .B(g20739), .Z(g22208) ) ;
NOR2    gate13811  (.A(g16210), .B(g13676), .Z(g19907) ) ;
AND2    gate13812  (.A(g19907), .B(g20751), .Z(g22209) ) ;
OR2     gate13813  (.A(g8183), .B(g12527), .Z(g13660) ) ;
AND2    gate13814  (.A(g13660), .B(g20000), .Z(g22216) ) ;
NOR2    gate13815  (.A(g16219), .B(g13709), .Z(g19951) ) ;
AND2    gate13816  (.A(g19951), .B(g20875), .Z(g22218) ) ;
NOR2    gate13817  (.A(g16220), .B(g13712), .Z(g19953) ) ;
AND2    gate13818  (.A(g19953), .B(g20887), .Z(g22219) ) ;
NOR2    gate13819  (.A(g16231), .B(g13739), .Z(g19997) ) ;
AND2    gate13820  (.A(g19997), .B(g21012), .Z(g22298) ) ;
NOR2    gate13821  (.A(g16232), .B(g13742), .Z(g19999) ) ;
AND2    gate13822  (.A(g19999), .B(g21024), .Z(g22299) ) ;
NOR2    gate13823  (.A(g16242), .B(g13779), .Z(g20027) ) ;
AND2    gate13824  (.A(g20027), .B(g21163), .Z(g22307) ) ;
AND2    gate13825  (.A(g1135), .B(g19738), .Z(g22308) ) ;
AND2    gate13826  (.A(g1478), .B(g19751), .Z(g22309) ) ;
AND2    gate13827  (.A(g19662), .B(g20235), .Z(g22310) ) ;
AND2    gate13828  (.A(g2837), .B(g20270), .Z(g22316) ) ;
NOR2    gate13829  (.A(g2712), .B(g10084), .Z(g11940) ) ;
AND2    gate13830  (.A(g11940), .B(g20329), .Z(g22329) ) ;
OR2     gate13831  (.A(g15707), .B(g13063), .Z(g19605) ) ;
AND2    gate13832  (.A(g19605), .B(g13522), .Z(g22340) ) ;
NAND2   gate13833  (.A(g14616), .B(g17571), .Z(g21287) ) ;
NAND2   gate13834  (.A(g14616), .B(g17225), .Z(g20783) ) ;
NAND2   gate13835  (.A(g14616), .B(g17595), .Z(g20784) ) ;
NAND2   gate13836  (.A(g14616), .B(g17363), .Z(g21186) ) ;
NAND2   gate13837  (.A(g14616), .B(g17364), .Z(g21187) ) ;
NAND2   gate13838  (.A(g14616), .B(g17492), .Z(g21288) ) ;
NAND2   gate13839  (.A(g14616), .B(g17493), .Z(g21289) ) ;
OR2     gate13840  (.A(g12186), .B(g9906), .Z(g12954) ) ;
AND2    gate13841  (.A(g12954), .B(g19386), .Z(g22489) ) ;
NAND2   gate13842  (.A(g14616), .B(g17596), .Z(g21334) ) ;
OR2     gate13843  (.A(g12219), .B(g9967), .Z(g12981) ) ;
AND2    gate13844  (.A(g12981), .B(g19395), .Z(g22515) ) ;
OR2     gate13845  (.A(g12220), .B(g9968), .Z(g12982) ) ;
AND2    gate13846  (.A(g12982), .B(g19398), .Z(g22518) ) ;
OR2     gate13847  (.A(g12284), .B(g10034), .Z(g13006) ) ;
AND2    gate13848  (.A(g13006), .B(g19411), .Z(g22525) ) ;
AND2    gate13849  (.A(g8766), .B(g21389), .Z(g22534) ) ;
AND2    gate13850  (.A(g14035), .B(g20248), .Z(g22538) ) ;
AND2    gate13851  (.A(g79), .B(g20078), .Z(g22588) ) ;
OR2     gate13852  (.A(g17752), .B(g17768), .Z(g19267) ) ;
AND2    gate13853  (.A(g19267), .B(g19451), .Z(g22589) ) ;
OR2     gate13854  (.A(g17753), .B(g14791), .Z(g19274) ) ;
AND2    gate13855  (.A(g19274), .B(g19452), .Z(g22590) ) ;
OR2     gate13856  (.A(g17769), .B(g14831), .Z(g19336) ) ;
AND2    gate13857  (.A(g19336), .B(g19469), .Z(g22622) ) ;
OR2     gate13858  (.A(g17770), .B(g17785), .Z(g19337) ) ;
AND2    gate13859  (.A(g19337), .B(g19470), .Z(g22623) ) ;
OR2     gate13860  (.A(g17771), .B(g14832), .Z(g19344) ) ;
AND2    gate13861  (.A(g19344), .B(g19471), .Z(g22624) ) ;
OR2     gate13862  (.A(g17784), .B(g14874), .Z(g19356) ) ;
AND2    gate13863  (.A(g19356), .B(g19476), .Z(g22632) ) ;
OR2     gate13864  (.A(g17786), .B(g14875), .Z(g19359) ) ;
AND2    gate13865  (.A(g19359), .B(g19479), .Z(g22633) ) ;
OR2     gate13866  (.A(g17810), .B(g14913), .Z(g19363) ) ;
AND2    gate13867  (.A(g19363), .B(g19489), .Z(g22637) ) ;
NOR2    gate13868  (.A(g9194), .B(g14279), .Z(g17174) ) ;
AND2    gate13869  (.A(g17174), .B(g20905), .Z(g22665) ) ;
NAND2   gate13870  (.A(g15829), .B(g10841), .Z(g19530) ) ;
NOR2    gate13871  (.A(g4064), .B(g4057), .Z(g7781) ) ;
AND2    gate13872  (.A(g19530), .B(g7781), .Z(g22680) ) ;
NOR2    gate13873  (.A(g812), .B(g9166), .Z(g11891) ) ;
AND2    gate13874  (.A(g11891), .B(g20192), .Z(g22685) ) ;
NAND2   gate13875  (.A(g15717), .B(g1056), .Z(g19335) ) ;
AND2    gate13876  (.A(g19335), .B(g19577), .Z(g22686) ) ;
NAND2   gate13877  (.A(g15723), .B(g1399), .Z(g19358) ) ;
AND2    gate13878  (.A(g19358), .B(g19600), .Z(g22710) ) ;
AND2    gate13879  (.A(g9291), .B(g20212), .Z(g22717) ) ;
AND2    gate13880  (.A(g9253), .B(g20619), .Z(g22720) ) ;
OR2     gate13881  (.A(g12920), .B(g10501), .Z(g15792) ) ;
AND2    gate13882  (.A(g15792), .B(g19612), .Z(g22752) ) ;
AND2    gate13883  (.A(g9360), .B(g20237), .Z(g22760) ) ;
AND2    gate13884  (.A(g9305), .B(g20645), .Z(g22762) ) ;
OR2     gate13885  (.A(g15507), .B(g12931), .Z(g19441) ) ;
AND2    gate13886  (.A(g19441), .B(g19629), .Z(g22831) ) ;
AND2    gate13887  (.A(g102), .B(g19630), .Z(g22834) ) ;
OR2     gate13888  (.A(g12924), .B(g10528), .Z(g15803) ) ;
AND2    gate13889  (.A(g15803), .B(g19633), .Z(g22835) ) ;
AND2    gate13890  (.A(g9429), .B(g20272), .Z(g22843) ) ;
AND2    gate13891  (.A(g9386), .B(g20676), .Z(g22846) ) ;
OR2     gate13892  (.A(g15567), .B(g12939), .Z(g19449) ) ;
AND2    gate13893  (.A(g19449), .B(g19649), .Z(g22848) ) ;
AND2    gate13894  (.A(g1227), .B(g19653), .Z(g22849) ) ;
AND2    gate13895  (.A(g496), .B(g19654), .Z(g22851) ) ;
AND2    gate13896  (.A(g9456), .B(g20734), .Z(g22859) ) ;
NAND2   gate13897  (.A(II20204), .B(II20205), .Z(g19792) ) ;
AND2    gate13898  (.A(g19792), .B(g19670), .Z(g22861) ) ;
AND2    gate13899  (.A(g1570), .B(g19673), .Z(g22862) ) ;
AND2    gate13900  (.A(g9547), .B(g20388), .Z(g22863) ) ;
AND2    gate13901  (.A(g9523), .B(g20871), .Z(g22871) ) ;
NAND2   gate13902  (.A(II20222), .B(II20223), .Z(g19854) ) ;
AND2    gate13903  (.A(g19854), .B(g19683), .Z(g22873) ) ;
OR2     gate13904  (.A(g15589), .B(g12979), .Z(g19486) ) ;
AND2    gate13905  (.A(g19486), .B(g19695), .Z(g22899) ) ;
NAND3   gate13906  (.A(g13727), .B(g13511), .C(g13527), .Z(g17137) ) ;
AND2    gate13907  (.A(g17137), .B(g19697), .Z(g22900) ) ;
NAND2   gate13908  (.A(II20166), .B(II20167), .Z(g19764) ) ;
AND2    gate13909  (.A(g19764), .B(g19719), .Z(g22920) ) ;
AND2    gate13910  (.A(g753), .B(g20540), .Z(g22937) ) ;
NAND2   gate13911  (.A(II20188), .B(II20189), .Z(g19782) ) ;
AND2    gate13912  (.A(g19782), .B(g19739), .Z(g22938) ) ;
AND2    gate13913  (.A(g9708), .B(g21062), .Z(g22939) ) ;
OR2     gate13914  (.A(g15651), .B(g13020), .Z(g19535) ) ;
AND2    gate13915  (.A(g19535), .B(g19747), .Z(g22982) ) ;
OR2     gate13916  (.A(g15672), .B(g13030), .Z(g19555) ) ;
AND2    gate13917  (.A(g19555), .B(g19760), .Z(g22990) ) ;
AND2    gate13918  (.A(g645), .B(g20248), .Z(g22991) ) ;
AND2    gate13919  (.A(g1227), .B(g19765), .Z(g22992) ) ;
OR2     gate13920  (.A(g15693), .B(g13042), .Z(g19575) ) ;
AND2    gate13921  (.A(g19575), .B(g19776), .Z(g23006) ) ;
AND2    gate13922  (.A(g681), .B(g20248), .Z(g23007) ) ;
AND2    gate13923  (.A(g1570), .B(g19783), .Z(g23008) ) ;
OR2     gate13924  (.A(g16207), .B(g13497), .Z(g20196) ) ;
AND2    gate13925  (.A(g650), .B(g20248), .Z(g23023) ) ;
OR2     gate13926  (.A(g13047), .B(g10706), .Z(g16021) ) ;
AND2    gate13927  (.A(g16021), .B(g19798), .Z(g23025) ) ;
AND2    gate13928  (.A(g655), .B(g20248), .Z(g23050) ) ;
OR2     gate13929  (.A(g13060), .B(g10724), .Z(g16052) ) ;
AND2    gate13930  (.A(g16052), .B(g19860), .Z(g23056) ) ;
AND2    gate13931  (.A(g718), .B(g20248), .Z(g23062) ) ;
OR2     gate13932  (.A(g13081), .B(g10736), .Z(g16076) ) ;
AND2    gate13933  (.A(g16076), .B(g19878), .Z(g23083) ) ;
AND2    gate13934  (.A(g10143), .B(g20765), .Z(g23103) ) ;
AND2    gate13935  (.A(g661), .B(g20248), .Z(g23104) ) ;
AND2    gate13936  (.A(g728), .B(g20248), .Z(g23130) ) ;
NOR2    gate13937  (.A(g3347), .B(g11276), .Z(g13919) ) ;
AND2    gate13938  (.A(g13919), .B(g19930), .Z(g23131) ) ;
OR2     gate13939  (.A(g16303), .B(g13632), .Z(g18994) ) ;
AND2    gate13940  (.A(g18994), .B(g7162), .Z(g23151) ) ;
NOR2    gate13941  (.A(g8663), .B(g11276), .Z(g13954) ) ;
AND2    gate13942  (.A(g13954), .B(g19964), .Z(g23165) ) ;
NOR2    gate13943  (.A(g3698), .B(g11309), .Z(g13959) ) ;
AND2    gate13944  (.A(g13959), .B(g19979), .Z(g23166) ) ;
NOR2    gate13945  (.A(g8697), .B(g11309), .Z(g13989) ) ;
AND2    gate13946  (.A(g13989), .B(g20010), .Z(g23187) ) ;
NOR2    gate13947  (.A(g4049), .B(g11363), .Z(g13994) ) ;
AND2    gate13948  (.A(g13994), .B(g20025), .Z(g23188) ) ;
NOR2    gate13949  (.A(g8734), .B(g11363), .Z(g14027) ) ;
AND2    gate13950  (.A(g14027), .B(g20040), .Z(g23201) ) ;
NAND2   gate13951  (.A(II20461), .B(II20462), .Z(g20200) ) ;
AND2    gate13952  (.A(g20200), .B(g16530), .Z(g23218) ) ;
AND2    gate13953  (.A(g19417), .B(g20067), .Z(g23220) ) ;
AND2    gate13954  (.A(g18994), .B(g4521), .Z(g23229) ) ;
AND2    gate13955  (.A(g20056), .B(g20110), .Z(g23254) ) ;
AND2    gate13956  (.A(g20069), .B(g20132), .Z(g23265) ) ;
AND2    gate13957  (.A(g19417), .B(g20146), .Z(g23280) ) ;
OR2     gate13958  (.A(g15841), .B(g13265), .Z(g19879) ) ;
AND2    gate13959  (.A(g19879), .B(g16726), .Z(g23292) ) ;
NOR2    gate13960  (.A(g822), .B(g14279), .Z(g15570) ) ;
AND2    gate13961  (.A(g15570), .B(g21393), .Z(g23348) ) ;
OR2     gate13962  (.A(g10896), .B(g10917), .Z(g13662) ) ;
AND2    gate13963  (.A(g13662), .B(g20182), .Z(g23349) ) ;
OR2     gate13964  (.A(g13287), .B(g10934), .Z(g16448) ) ;
AND2    gate13965  (.A(g16448), .B(g20194), .Z(g23372) ) ;
OR2     gate13966  (.A(g10921), .B(g10947), .Z(g13699) ) ;
AND2    gate13967  (.A(g13699), .B(g20195), .Z(g23373) ) ;
AND2    gate13968  (.A(g7239), .B(g21413), .Z(g23381) ) ;
OR2     gate13969  (.A(g15902), .B(g13299), .Z(g20034) ) ;
AND2    gate13970  (.A(g20034), .B(g20207), .Z(g23386) ) ;
OR2     gate13971  (.A(g13294), .B(g10966), .Z(g16506) ) ;
AND2    gate13972  (.A(g16506), .B(g20211), .Z(g23387) ) ;
AND2    gate13973  (.A(g9072), .B(g19757), .Z(g23389) ) ;
AND2    gate13974  (.A(g7247), .B(g21430), .Z(g23392) ) ;
OR2     gate13975  (.A(g15936), .B(g13306), .Z(g20051) ) ;
AND2    gate13976  (.A(g20051), .B(g20229), .Z(g23396) ) ;
NAND2   gate13977  (.A(II14212), .B(II14213), .Z(g11154) ) ;
AND2    gate13978  (.A(g11154), .B(g20239), .Z(g23397) ) ;
AND2    gate13979  (.A(g7262), .B(g21460), .Z(g23401) ) ;
OR2     gate13980  (.A(g15978), .B(g13313), .Z(g20063) ) ;
AND2    gate13981  (.A(g20063), .B(g20247), .Z(g23404) ) ;
NAND2   gate13982  (.A(II13066), .B(II13067), .Z(g9295) ) ;
AND2    gate13983  (.A(g9295), .B(g20273), .Z(g23407) ) ;
AND2    gate13984  (.A(g7297), .B(g21510), .Z(g23412) ) ;
OR2     gate13985  (.A(g16025), .B(g13320), .Z(g20077) ) ;
AND2    gate13986  (.A(g20077), .B(g20320), .Z(g23415) ) ;
OR2     gate13987  (.A(g16026), .B(g13321), .Z(g20082) ) ;
AND2    gate13988  (.A(g20082), .B(g20321), .Z(g23416) ) ;
AND2    gate13989  (.A(g7345), .B(g21556), .Z(g23424) ) ;
AND2    gate13990  (.A(g13771), .B(g20452), .Z(g23439) ) ;
AND2    gate13991  (.A(g13805), .B(g20510), .Z(g23451) ) ;
OR2     gate13992  (.A(g16128), .B(g13393), .Z(g20148) ) ;
AND2    gate13993  (.A(g20148), .B(g20523), .Z(g23471) ) ;
AND2    gate13994  (.A(g13830), .B(g20533), .Z(g23474) ) ;
NOR2    gate13995  (.A(g16957), .B(g11720), .Z(g19070) ) ;
AND2    gate13996  (.A(g19070), .B(g8971), .Z(g23475) ) ;
OR2     gate13997  (.A(g16163), .B(g13415), .Z(g20160) ) ;
AND2    gate13998  (.A(g20160), .B(g20541), .Z(g23484) ) ;
OR2     gate13999  (.A(g16184), .B(g13460), .Z(g20169) ) ;
AND2    gate14000  (.A(g20169), .B(g20569), .Z(g23497) ) ;
NOR2    gate14001  (.A(g17140), .B(g14207), .Z(g20234) ) ;
AND2    gate14002  (.A(g20234), .B(g12998), .Z(g23498) ) ;
NOR2    gate14003  (.A(g17150), .B(g14220), .Z(g19430) ) ;
AND2    gate14004  (.A(g19430), .B(g13007), .Z(g23513) ) ;
NOR2    gate14005  (.A(g17091), .B(g14185), .Z(g20149) ) ;
AND2    gate14006  (.A(g20149), .B(g11829), .Z(g23514) ) ;
NOR2    gate14007  (.A(g1046), .B(g7479), .Z(g10760) ) ;
AND2    gate14008  (.A(g10760), .B(g18930), .Z(g23531) ) ;
NOR2    gate14009  (.A(g17139), .B(g14206), .Z(g19400) ) ;
AND2    gate14010  (.A(g19400), .B(g11852), .Z(g23532) ) ;
NOR2    gate14011  (.A(g17176), .B(g14233), .Z(g19436) ) ;
AND2    gate14012  (.A(g19436), .B(g13015), .Z(g23533) ) ;
OR2     gate14013  (.A(g13492), .B(g11044), .Z(g16866) ) ;
AND2    gate14014  (.A(g16866), .B(g20622), .Z(g23540) ) ;
NOR2    gate14015  (.A(g1389), .B(g7503), .Z(g10793) ) ;
AND2    gate14016  (.A(g10793), .B(g18948), .Z(g23551) ) ;
NOR2    gate14017  (.A(g17151), .B(g14221), .Z(g19413) ) ;
AND2    gate14018  (.A(g19413), .B(g11875), .Z(g23553) ) ;
NOR2    gate14019  (.A(g17182), .B(g14257), .Z(g20390) ) ;
AND2    gate14020  (.A(g20390), .B(g13024), .Z(g23554) ) ;
OR2     gate14021  (.A(g13508), .B(g11114), .Z(g16882) ) ;
AND2    gate14022  (.A(g16882), .B(g20648), .Z(g23564) ) ;
AND2    gate14023  (.A(g20230), .B(g20656), .Z(g23572) ) ;
NOR2    gate14024  (.A(g17192), .B(g14295), .Z(g19444) ) ;
AND2    gate14025  (.A(g19444), .B(g13033), .Z(g23577) ) ;
NOR2    gate14026  (.A(g17152), .B(g14222), .Z(g20183) ) ;
AND2    gate14027  (.A(g20183), .B(g11900), .Z(g23581) ) ;
OR2     gate14028  (.A(g13524), .B(g11126), .Z(g16927) ) ;
AND2    gate14029  (.A(g16927), .B(g20679), .Z(g23606) ) ;
NOR2    gate14030  (.A(g17181), .B(g14256), .Z(g19388) ) ;
AND2    gate14031  (.A(g19388), .B(g11917), .Z(g23618) ) ;
NOR2    gate14032  (.A(g17199), .B(g14316), .Z(g19453) ) ;
AND2    gate14033  (.A(g19453), .B(g13045), .Z(g23619) ) ;
OR2     gate14034  (.A(g13542), .B(g11142), .Z(g16959) ) ;
AND2    gate14035  (.A(g16959), .B(g20737), .Z(g23646) ) ;
NOR2    gate14036  (.A(g17193), .B(g14296), .Z(g19401) ) ;
AND2    gate14037  (.A(g19401), .B(g11941), .Z(g23657) ) ;
NOR2    gate14038  (.A(g5352), .B(g12166), .Z(g14687) ) ;
AND2    gate14039  (.A(g14687), .B(g20852), .Z(g23658) ) ;
OR2     gate14040  (.A(g13567), .B(g11163), .Z(g16970) ) ;
AND2    gate14041  (.A(g16970), .B(g20874), .Z(g23682) ) ;
NOR2    gate14042  (.A(g10090), .B(g12166), .Z(g14726) ) ;
AND2    gate14043  (.A(g14726), .B(g20978), .Z(g23690) ) ;
NOR2    gate14044  (.A(g5698), .B(g12204), .Z(g14731) ) ;
AND2    gate14045  (.A(g14731), .B(g20993), .Z(g23691) ) ;
NOR2    gate14046  (.A(g10130), .B(g12204), .Z(g14767) ) ;
AND2    gate14047  (.A(g14767), .B(g21123), .Z(g23724) ) ;
NOR2    gate14048  (.A(g6044), .B(g12252), .Z(g14772) ) ;
AND2    gate14049  (.A(g14772), .B(g21138), .Z(g23725) ) ;
NOR2    gate14050  (.A(g10166), .B(g12252), .Z(g14816) ) ;
AND2    gate14051  (.A(g14816), .B(g21189), .Z(g23754) ) ;
NOR2    gate14052  (.A(g6390), .B(g12314), .Z(g14821) ) ;
AND2    gate14053  (.A(g14821), .B(g21204), .Z(g23755) ) ;
NOR2    gate14054  (.A(g10191), .B(g12314), .Z(g14867) ) ;
AND2    gate14055  (.A(g14867), .B(g21252), .Z(g23774) ) ;
NOR2    gate14056  (.A(g6736), .B(g12364), .Z(g14872) ) ;
AND2    gate14057  (.A(g14872), .B(g21267), .Z(g23775) ) ;
AND2    gate14058  (.A(g1105), .B(g19355), .Z(g23779) ) ;
NOR2    gate14059  (.A(g10213), .B(g12364), .Z(g14911) ) ;
AND2    gate14060  (.A(g14911), .B(g21279), .Z(g23799) ) ;
AND2    gate14061  (.A(g1448), .B(g19362), .Z(g23801) ) ;
AND2    gate14062  (.A(g4087), .B(g19364), .Z(g23811) ) ;
AND2    gate14063  (.A(g4129), .B(g19495), .Z(g23836) ) ;
AND2    gate14064  (.A(g21160), .B(g10804), .Z(g23837) ) ;
AND2    gate14065  (.A(g4093), .B(g19506), .Z(g23854) ) ;
AND2    gate14066  (.A(g4112), .B(g19455), .Z(g23855) ) ;
AND2    gate14067  (.A(g4116), .B(g19483), .Z(g23856) ) ;
AND2    gate14068  (.A(g19626), .B(g7908), .Z(g23857) ) ;
AND2    gate14069  (.A(g19389), .B(g4157), .Z(g23872) ) ;
AND2    gate14070  (.A(g21222), .B(g10815), .Z(g23873) ) ;
AND2    gate14071  (.A(g4119), .B(g19510), .Z(g23884) ) ;
AND2    gate14072  (.A(g4132), .B(g19513), .Z(g23885) ) ;
AND2    gate14073  (.A(g1129), .B(g19408), .Z(g23900) ) ;
AND2    gate14074  (.A(g19606), .B(g7963), .Z(g23901) ) ;
AND2    gate14075  (.A(g1472), .B(g19428), .Z(g23917) ) ;
AND2    gate14076  (.A(g4122), .B(g19546), .Z(g23919) ) ;
AND2    gate14077  (.A(g4135), .B(g19549), .Z(g23920) ) ;
AND2    gate14078  (.A(g19379), .B(g4146), .Z(g23921) ) ;
AND2    gate14079  (.A(g4138), .B(g19589), .Z(g23957) ) ;
AND2    gate14080  (.A(g19610), .B(g10951), .Z(g23990) ) ;
NOR3    gate14081  (.A(g12971), .B(g15614), .C(g11320), .Z(g19209) ) ;
AND2    gate14082  (.A(g19209), .B(g21428), .Z(g23991) ) ;
AND2    gate14083  (.A(g19596), .B(g10951), .Z(g23996) ) ;
AND2    gate14084  (.A(g19631), .B(g10971), .Z(g23998) ) ;
AND2    gate14085  (.A(g19651), .B(g10951), .Z(g24001) ) ;
AND2    gate14086  (.A(g19613), .B(g10971), .Z(g24002) ) ;
AND2    gate14087  (.A(g37), .B(g21225), .Z(g24004) ) ;
AND2    gate14088  (.A(g7909), .B(g19502), .Z(g24008) ) ;
AND2    gate14089  (.A(g19671), .B(g10971), .Z(g24009) ) ;
AND2    gate14090  (.A(g7939), .B(g19524), .Z(g24011) ) ;
AND2    gate14091  (.A(g14496), .B(g21561), .Z(g24012) ) ;
AND2    gate14092  (.A(g7933), .B(g19063), .Z(g24014) ) ;
AND2    gate14093  (.A(g19540), .B(g10951), .Z(g24015) ) ;
AND2    gate14094  (.A(g14528), .B(g21610), .Z(g24016) ) ;
AND2    gate14095  (.A(g17619), .B(g21653), .Z(g24139) ) ;
AND2    gate14096  (.A(g17663), .B(g21654), .Z(g24140) ) ;
AND2    gate14097  (.A(g17657), .B(g21656), .Z(g24141) ) ;
AND2    gate14098  (.A(g17700), .B(g21657), .Z(g24142) ) ;
AND2    gate14099  (.A(g17694), .B(g21659), .Z(g24143) ) ;
AND2    gate14100  (.A(g17727), .B(g21660), .Z(g24144) ) ;
AND2    gate14101  (.A(g18102), .B(g22722), .Z(g24186) ) ;
AND2    gate14102  (.A(g305), .B(g22722), .Z(g24187) ) ;
AND2    gate14103  (.A(g316), .B(g22722), .Z(g24188) ) ;
AND2    gate14104  (.A(g324), .B(g22722), .Z(g24189) ) ;
AND2    gate14105  (.A(g329), .B(g22722), .Z(g24190) ) ;
AND2    gate14106  (.A(g319), .B(g22722), .Z(g24191) ) ;
AND2    gate14107  (.A(g311), .B(g22722), .Z(g24192) ) ;
AND2    gate14108  (.A(g336), .B(g22722), .Z(g24193) ) ;
AND2    gate14109  (.A(g106), .B(g22722), .Z(g24194) ) ;
AND2    gate14110  (.A(g74), .B(g22722), .Z(g24195) ) ;
AND2    gate14111  (.A(g333), .B(g22722), .Z(g24196) ) ;
AND2    gate14112  (.A(g347), .B(g22722), .Z(g24197) ) ;
AND2    gate14113  (.A(g351), .B(g22722), .Z(g24198) ) ;
AND2    gate14114  (.A(g355), .B(g22722), .Z(g24199) ) ;
AND2    gate14115  (.A(g18200), .B(g22594), .Z(g24217) ) ;
AND2    gate14116  (.A(g872), .B(g22594), .Z(g24218) ) ;
AND2    gate14117  (.A(g225), .B(g22594), .Z(g24219) ) ;
AND2    gate14118  (.A(g255), .B(g22594), .Z(g24220) ) ;
AND2    gate14119  (.A(g232), .B(g22594), .Z(g24221) ) ;
AND2    gate14120  (.A(g262), .B(g22594), .Z(g24222) ) ;
AND2    gate14121  (.A(g239), .B(g22594), .Z(g24223) ) ;
AND2    gate14122  (.A(g269), .B(g22594), .Z(g24224) ) ;
AND2    gate14123  (.A(g246), .B(g22594), .Z(g24225) ) ;
AND2    gate14124  (.A(g446), .B(g22594), .Z(g24226) ) ;
AND2    gate14125  (.A(g890), .B(g22594), .Z(g24227) ) ;
AND2    gate14126  (.A(g862), .B(g22594), .Z(g24228) ) ;
AND2    gate14127  (.A(g901), .B(g22594), .Z(g24230) ) ;
AND2    gate14128  (.A(g4411), .B(g22550), .Z(g24283) ) ;
AND2    gate14129  (.A(g4375), .B(g22550), .Z(g24284) ) ;
AND2    gate14130  (.A(g4388), .B(g22550), .Z(g24285) ) ;
AND2    gate14131  (.A(g4405), .B(g22550), .Z(g24286) ) ;
AND2    gate14132  (.A(g4401), .B(g22550), .Z(g24287) ) ;
AND2    gate14133  (.A(g4417), .B(g22550), .Z(g24288) ) ;
AND2    gate14134  (.A(g4427), .B(g22550), .Z(g24289) ) ;
AND2    gate14135  (.A(g4430), .B(g22550), .Z(g24290) ) ;
AND2    gate14136  (.A(g18660), .B(g22550), .Z(g24291) ) ;
AND2    gate14137  (.A(g4443), .B(g22550), .Z(g24292) ) ;
AND2    gate14138  (.A(g4438), .B(g22550), .Z(g24293) ) ;
AND2    gate14139  (.A(g4452), .B(g22550), .Z(g24294) ) ;
AND2    gate14140  (.A(g4434), .B(g22550), .Z(g24295) ) ;
AND2    gate14141  (.A(g4382), .B(g22550), .Z(g24296) ) ;
AND2    gate14142  (.A(g4455), .B(g22550), .Z(g24297) ) ;
AND2    gate14143  (.A(g4456), .B(g22550), .Z(g24299) ) ;
NOR2    gate14144  (.A(g6975), .B(g13605), .Z(g15123) ) ;
AND2    gate14145  (.A(g15123), .B(g22228), .Z(g24300) ) ;
AND2    gate14146  (.A(g6961), .B(g22228), .Z(g24301) ) ;
OR2     gate14147  (.A(g13605), .B(g4581), .Z(g15124) ) ;
AND2    gate14148  (.A(g15124), .B(g22228), .Z(g24302) ) ;
AND2    gate14149  (.A(g4369), .B(g22228), .Z(g24303) ) ;
AND2    gate14150  (.A(g12875), .B(g22228), .Z(g24304) ) ;
AND2    gate14151  (.A(g4477), .B(g22228), .Z(g24305) ) ;
AND2    gate14152  (.A(g4483), .B(g22228), .Z(g24306) ) ;
AND2    gate14153  (.A(g4486), .B(g22228), .Z(g24307) ) ;
AND2    gate14154  (.A(g4489), .B(g22228), .Z(g24308) ) ;
AND2    gate14155  (.A(g4480), .B(g22228), .Z(g24309) ) ;
AND2    gate14156  (.A(g4495), .B(g22228), .Z(g24310) ) ;
AND2    gate14157  (.A(g4498), .B(g22228), .Z(g24311) ) ;
AND2    gate14158  (.A(g4501), .B(g22228), .Z(g24312) ) ;
AND2    gate14159  (.A(g4504), .B(g22228), .Z(g24313) ) ;
AND2    gate14160  (.A(g4515), .B(g22228), .Z(g24314) ) ;
AND2    gate14161  (.A(g4521), .B(g22228), .Z(g24315) ) ;
AND2    gate14162  (.A(g4527), .B(g22228), .Z(g24316) ) ;
AND2    gate14163  (.A(g4534), .B(g22228), .Z(g24317) ) ;
AND2    gate14164  (.A(g4555), .B(g22228), .Z(g24318) ) ;
AND2    gate14165  (.A(g4561), .B(g22228), .Z(g24319) ) ;
AND2    gate14166  (.A(g6973), .B(g22228), .Z(g24320) ) ;
AND2    gate14167  (.A(g4558), .B(g22228), .Z(g24321) ) ;
AND2    gate14168  (.A(g4423), .B(g22228), .Z(g24322) ) ;
AND2    gate14169  (.A(g4546), .B(g22228), .Z(g24323) ) ;
AND2    gate14170  (.A(g4540), .B(g22228), .Z(g24324) ) ;
AND2    gate14171  (.A(g4543), .B(g22228), .Z(g24325) ) ;
AND2    gate14172  (.A(g4552), .B(g22228), .Z(g24326) ) ;
AND2    gate14173  (.A(g4549), .B(g22228), .Z(g24327) ) ;
AND2    gate14174  (.A(g4567), .B(g22228), .Z(g24328) ) ;
AND2    gate14175  (.A(g4462), .B(g22228), .Z(g24329) ) ;
AND2    gate14176  (.A(g18661), .B(g22228), .Z(g24330) ) ;
AND2    gate14177  (.A(g6977), .B(g22228), .Z(g24331) ) ;
AND2    gate14178  (.A(g4459), .B(g22228), .Z(g24332) ) ;
AND2    gate14179  (.A(g4512), .B(g22228), .Z(g24333) ) ;
AND2    gate14180  (.A(g3106), .B(g22718), .Z(g24378) ) ;
AND2    gate14181  (.A(g3457), .B(g22761), .Z(g24387) ) ;
AND2    gate14182  (.A(g3115), .B(g23067), .Z(g24392) ) ;
AND2    gate14183  (.A(g3808), .B(g22844), .Z(g24393) ) ;
AND2    gate14184  (.A(g4704), .B(g22845), .Z(g24395) ) ;
AND2    gate14185  (.A(g3133), .B(g23067), .Z(g24399) ) ;
AND2    gate14186  (.A(g3466), .B(g23112), .Z(g24400) ) ;
AND2    gate14187  (.A(g4749), .B(g22857), .Z(g24402) ) ;
AND2    gate14188  (.A(g4894), .B(g22858), .Z(g24403) ) ;
OR2     gate14189  (.A(g482), .B(g12527), .Z(g13623) ) ;
AND2    gate14190  (.A(g13623), .B(g22860), .Z(g24406) ) ;
OR2     gate14191  (.A(g20581), .B(g17179), .Z(g23989) ) ;
AND2    gate14192  (.A(g23989), .B(g18946), .Z(g24408) ) ;
AND2    gate14193  (.A(g3484), .B(g23112), .Z(g24409) ) ;
AND2    gate14194  (.A(g3817), .B(g23139), .Z(g24410) ) ;
AND2    gate14195  (.A(g4760), .B(g22869), .Z(g24415) ) ;
AND2    gate14196  (.A(g4939), .B(g22870), .Z(g24416) ) ;
OR2     gate14197  (.A(g20602), .B(g17191), .Z(g23997) ) ;
AND2    gate14198  (.A(g23997), .B(g18980), .Z(g24420) ) ;
AND2    gate14199  (.A(g3835), .B(g23139), .Z(g24421) ) ;
AND2    gate14200  (.A(g4771), .B(g22896), .Z(g24422) ) ;
AND2    gate14201  (.A(g4950), .B(g22897), .Z(g24423) ) ;
AND2    gate14202  (.A(g4961), .B(g22919), .Z(g24427) ) ;
AND2    gate14203  (.A(g3125), .B(g23067), .Z(g24436) ) ;
AND2    gate14204  (.A(g3129), .B(g23067), .Z(g24450) ) ;
AND2    gate14205  (.A(g3476), .B(g23112), .Z(g24451) ) ;
AND2    gate14206  (.A(g3480), .B(g23112), .Z(g24464) ) ;
AND2    gate14207  (.A(g3827), .B(g23139), .Z(g24465) ) ;
OR2     gate14208  (.A(g490), .B(g12527), .Z(g13761) ) ;
AND2    gate14209  (.A(g13761), .B(g23047), .Z(g24467) ) ;
AND2    gate14210  (.A(g3831), .B(g23139), .Z(g24475) ) ;
OR2     gate14211  (.A(g17365), .B(g14423), .Z(g18879) ) ;
AND2    gate14212  (.A(g18879), .B(g22330), .Z(g24476) ) ;
AND2    gate14213  (.A(g6875), .B(g23055), .Z(g24482) ) ;
NOR2    gate14214  (.A(g13794), .B(g417), .Z(g16288) ) ;
NOR2    gate14215  (.A(g20035), .B(g16324), .Z(g23208) ) ;
AND2    gate14216  (.A(g6905), .B(g23082), .Z(g24488) ) ;
AND2    gate14217  (.A(g6928), .B(g23127), .Z(g24495) ) ;
NOR2    gate14218  (.A(g8725), .B(g11083), .Z(g14036) ) ;
AND2    gate14219  (.A(g14036), .B(g23850), .Z(g24498) ) ;
OR2     gate14220  (.A(g21302), .B(g17617), .Z(g22217) ) ;
AND2    gate14221  (.A(g22217), .B(g19394), .Z(g24499) ) ;
NOR2    gate14222  (.A(g8766), .B(g12259), .Z(g14000) ) ;
AND2    gate14223  (.A(g14000), .B(g23182), .Z(g24501) ) ;
NAND2   gate14224  (.A(g13945), .B(g20522), .Z(g23428) ) ;
AND2    gate14225  (.A(g23428), .B(g13223), .Z(g24502) ) ;
OR2     gate14226  (.A(g21332), .B(g17654), .Z(g22225) ) ;
AND2    gate14227  (.A(g22225), .B(g19409), .Z(g24503) ) ;
OR2     gate14228  (.A(g21333), .B(g17655), .Z(g22226) ) ;
AND2    gate14229  (.A(g22226), .B(g19410), .Z(g24504) ) ;
OR2     gate14230  (.A(g21347), .B(g17693), .Z(g22304) ) ;
AND2    gate14231  (.A(g22304), .B(g19429), .Z(g24507) ) ;
OR2     gate14232  (.A(g21394), .B(g17783), .Z(g22318) ) ;
AND2    gate14233  (.A(g22318), .B(g19468), .Z(g24523) ) ;
OR2     gate14234  (.A(g21405), .B(g17809), .Z(g22331) ) ;
AND2    gate14235  (.A(g22331), .B(g19478), .Z(g24532) ) ;
AND2    gate14236  (.A(g19516), .B(g22635), .Z(g24536) ) ;
AND2    gate14237  (.A(g3333), .B(g23285), .Z(g24545) ) ;
OR2     gate14238  (.A(g21464), .B(g12761), .Z(g22447) ) ;
AND2    gate14239  (.A(g22447), .B(g19523), .Z(g24546) ) ;
OR3     gate14240  (.A(g20184), .B(g20170), .C(II22267), .Z(g23162) ) ;
AND2    gate14241  (.A(g23162), .B(g20887), .Z(g24549) ) ;
AND2    gate14242  (.A(g3684), .B(g23308), .Z(g24550) ) ;
NOR2    gate14243  (.A(g827), .B(g14279), .Z(g17148) ) ;
AND2    gate14244  (.A(g17148), .B(g23331), .Z(g24551) ) ;
OR2     gate14245  (.A(g21512), .B(g12794), .Z(g22487) ) ;
AND2    gate14246  (.A(g22487), .B(g19538), .Z(g24552) ) ;
NOR3    gate14247  (.A(g979), .B(g16268), .C(g19853), .Z(g22983) ) ;
AND2    gate14248  (.A(g22983), .B(g19539), .Z(g24553) ) ;
OR2     gate14249  (.A(g21513), .B(g12795), .Z(g22490) ) ;
AND2    gate14250  (.A(g22490), .B(g19541), .Z(g24554) ) ;
OR3     gate14251  (.A(g20198), .B(g20185), .C(II22280), .Z(g23184) ) ;
AND2    gate14252  (.A(g23184), .B(g21024), .Z(g24555) ) ;
AND2    gate14253  (.A(g4035), .B(g23341), .Z(g24556) ) ;
OR2     gate14254  (.A(g21559), .B(g12817), .Z(g22516) ) ;
AND2    gate14255  (.A(g22516), .B(g19566), .Z(g24558) ) ;
NOR3    gate14256  (.A(g1322), .B(g16292), .C(g19873), .Z(g22993) ) ;
AND2    gate14257  (.A(g22993), .B(g19567), .Z(g24559) ) ;
OR3     gate14258  (.A(g20214), .B(g20199), .C(II22298), .Z(g23198) ) ;
AND2    gate14259  (.A(g23198), .B(g21163), .Z(g24564) ) ;
AND2    gate14260  (.A(g5115), .B(g23382), .Z(g24569) ) ;
AND2    gate14261  (.A(g5462), .B(g23393), .Z(g24572) ) ;
NOR2    gate14262  (.A(g9282), .B(g14279), .Z(g17198) ) ;
AND2    gate14263  (.A(g17198), .B(g23716), .Z(g24573) ) ;
AND2    gate14264  (.A(g5124), .B(g23590), .Z(g24581) ) ;
AND2    gate14265  (.A(g5808), .B(g23402), .Z(g24582) ) ;
AND2    gate14266  (.A(g5142), .B(g23590), .Z(g24588) ) ;
AND2    gate14267  (.A(g5471), .B(g23630), .Z(g24589) ) ;
AND2    gate14268  (.A(g6154), .B(g23413), .Z(g24590) ) ;
OR2     gate14269  (.A(g18893), .B(g18909), .Z(g22591) ) ;
AND2    gate14270  (.A(g22591), .B(g19652), .Z(g24600) ) ;
NAND2   gate14271  (.A(g13797), .B(g13764), .Z(g16507) ) ;
AND2    gate14272  (.A(g16507), .B(g22854), .Z(g24602) ) ;
AND2    gate14273  (.A(g5489), .B(g23630), .Z(g24606) ) ;
AND2    gate14274  (.A(g5817), .B(g23666), .Z(g24607) ) ;
AND2    gate14275  (.A(g6500), .B(g23425), .Z(g24608) ) ;
OR2     gate14276  (.A(g18910), .B(g18933), .Z(g22625) ) ;
AND2    gate14277  (.A(g22625), .B(g19672), .Z(g24618) ) ;
NAND3   gate14278  (.A(g13626), .B(g16278), .C(g8105), .Z(g19856) ) ;
AND2    gate14279  (.A(g19856), .B(g22866), .Z(g24622) ) ;
NAND2   gate14280  (.A(g13822), .B(g13798), .Z(g16524) ) ;
AND2    gate14281  (.A(g16524), .B(g22867), .Z(g24624) ) ;
AND2    gate14282  (.A(g22763), .B(g19679), .Z(g24627) ) ;
AND2    gate14283  (.A(g5835), .B(g23666), .Z(g24628) ) ;
AND2    gate14284  (.A(g6163), .B(g23699), .Z(g24629) ) ;
OR2     gate14285  (.A(g19655), .B(g16122), .Z(g23255) ) ;
AND2    gate14286  (.A(g23255), .B(g14149), .Z(g24630) ) ;
OR2     gate14287  (.A(g18934), .B(g15590), .Z(g22634) ) ;
AND2    gate14288  (.A(g22634), .B(g19685), .Z(g24634) ) ;
NAND3   gate14289  (.A(g13665), .B(g16299), .C(g8163), .Z(g19874) ) ;
AND2    gate14290  (.A(g19874), .B(g22883), .Z(g24635) ) ;
NAND2   gate14291  (.A(g13851), .B(g13823), .Z(g16586) ) ;
AND2    gate14292  (.A(g16586), .B(g22884), .Z(g24637) ) ;
AND2    gate14293  (.A(g22763), .B(g19690), .Z(g24638) ) ;
AND2    gate14294  (.A(g6181), .B(g23699), .Z(g24639) ) ;
AND2    gate14295  (.A(g6509), .B(g23733), .Z(g24640) ) ;
AND2    gate14296  (.A(g8290), .B(g22898), .Z(g24642) ) ;
OR2     gate14297  (.A(g18943), .B(g15611), .Z(g22636) ) ;
AND2    gate14298  (.A(g22636), .B(g19696), .Z(g24643) ) ;
AND2    gate14299  (.A(g11714), .B(g22903), .Z(g24644) ) ;
OR2     gate14300  (.A(g18950), .B(g15612), .Z(g22639) ) ;
AND2    gate14301  (.A(g22639), .B(g19709), .Z(g24645) ) ;
OR2     gate14302  (.A(g18951), .B(g15613), .Z(g22640) ) ;
AND2    gate14303  (.A(g22640), .B(g19711), .Z(g24646) ) ;
NAND3   gate14304  (.A(g13707), .B(g16319), .C(g8227), .Z(g19903) ) ;
AND2    gate14305  (.A(g19903), .B(g22907), .Z(g24647) ) ;
AND2    gate14306  (.A(g6527), .B(g23733), .Z(g24649) ) ;
OR2     gate14307  (.A(g18974), .B(g15631), .Z(g22641) ) ;
AND2    gate14308  (.A(g22641), .B(g19718), .Z(g24650) ) ;
AND2    gate14309  (.A(g2741), .B(g23472), .Z(g24651) ) ;
AND2    gate14310  (.A(g11735), .B(g22922), .Z(g24654) ) ;
AND2    gate14311  (.A(g11736), .B(g22926), .Z(g24656) ) ;
OR2     gate14312  (.A(g18981), .B(g15632), .Z(g22644) ) ;
AND2    gate14313  (.A(g22644), .B(g19730), .Z(g24657) ) ;
OR2     gate14314  (.A(g18982), .B(g15633), .Z(g22645) ) ;
AND2    gate14315  (.A(g22645), .B(g19732), .Z(g24658) ) ;
AND2    gate14316  (.A(g5134), .B(g23590), .Z(g24659) ) ;
OR2     gate14317  (.A(g18987), .B(g15652), .Z(g22648) ) ;
AND2    gate14318  (.A(g22648), .B(g19737), .Z(g24660) ) ;
AND2    gate14319  (.A(g16621), .B(g22974), .Z(g24663) ) ;
OR2     gate14320  (.A(g18992), .B(g15653), .Z(g22652) ) ;
AND2    gate14321  (.A(g22652), .B(g19741), .Z(g24664) ) ;
AND2    gate14322  (.A(g11753), .B(g22975), .Z(g24666) ) ;
AND2    gate14323  (.A(g11754), .B(g22979), .Z(g24668) ) ;
OR2     gate14324  (.A(g18993), .B(g15654), .Z(g22653) ) ;
AND2    gate14325  (.A(g22653), .B(g19742), .Z(g24669) ) ;
AND2    gate14326  (.A(g5138), .B(g23590), .Z(g24670) ) ;
AND2    gate14327  (.A(g5481), .B(g23630), .Z(g24671) ) ;
OR2     gate14328  (.A(g15650), .B(g13019), .Z(g19534) ) ;
AND2    gate14329  (.A(g19534), .B(g22981), .Z(g24672) ) ;
OR2     gate14330  (.A(g19062), .B(g15673), .Z(g22659) ) ;
AND2    gate14331  (.A(g22659), .B(g19748), .Z(g24673) ) ;
AND2    gate14332  (.A(g446), .B(g23496), .Z(g24674) ) ;
NAND2   gate14333  (.A(II18486), .B(II18487), .Z(g17568) ) ;
AND2    gate14334  (.A(g17568), .B(g22342), .Z(g24675) ) ;
AND2    gate14335  (.A(g2748), .B(g23782), .Z(g24676) ) ;
OR2     gate14336  (.A(g10619), .B(g10624), .Z(g13289) ) ;
AND2    gate14337  (.A(g13289), .B(g22985), .Z(g24679) ) ;
AND2    gate14338  (.A(g16422), .B(g22986), .Z(g24680) ) ;
AND2    gate14339  (.A(g16653), .B(g22988), .Z(g24681) ) ;
OR2     gate14340  (.A(g19069), .B(g15679), .Z(g22662) ) ;
AND2    gate14341  (.A(g22662), .B(g19754), .Z(g24682) ) ;
AND2    gate14342  (.A(g11769), .B(g22989), .Z(g24684) ) ;
AND2    gate14343  (.A(g5485), .B(g23630), .Z(g24686) ) ;
AND2    gate14344  (.A(g5827), .B(g23666), .Z(g24687) ) ;
NAND2   gate14345  (.A(II21993), .B(II21994), .Z(g22681) ) ;
NAND2   gate14346  (.A(II21977), .B(II21978), .Z(g22663) ) ;
AND2    gate14347  (.A(g22681), .B(g22663), .Z(g24688) ) ;
OR2     gate14348  (.A(g19139), .B(g15694), .Z(g22664) ) ;
AND2    gate14349  (.A(g22664), .B(g19761), .Z(g24698) ) ;
AND2    gate14350  (.A(g645), .B(g23512), .Z(g24700) ) ;
OR4     gate14351  (.A(g14334), .B(g14313), .C(g11935), .D(II18385), .Z(g17464) ) ;
AND2    gate14352  (.A(g17464), .B(g22342), .Z(g24702) ) ;
NAND2   gate14353  (.A(II18530), .B(II18531), .Z(g17592) ) ;
AND2    gate14354  (.A(g17592), .B(g22369), .Z(g24703) ) ;
NAND2   gate14355  (.A(II18537), .B(II18538), .Z(g17593) ) ;
AND2    gate14356  (.A(g17593), .B(g22384), .Z(g24704) ) ;
OR2     gate14357  (.A(g13025), .B(g10654), .Z(g15910) ) ;
AND2    gate14358  (.A(g15910), .B(g22996), .Z(g24706) ) ;
OR2     gate14359  (.A(g10625), .B(g10655), .Z(g13295) ) ;
AND2    gate14360  (.A(g13295), .B(g22997), .Z(g24707) ) ;
AND2    gate14361  (.A(g16474), .B(g22998), .Z(g24708) ) ;
AND2    gate14362  (.A(g16690), .B(g23000), .Z(g24709) ) ;
OR2     gate14363  (.A(g19145), .B(g15701), .Z(g22679) ) ;
AND2    gate14364  (.A(g22679), .B(g19771), .Z(g24710) ) ;
AND2    gate14365  (.A(g19592), .B(g23001), .Z(g24712) ) ;
AND2    gate14366  (.A(g5831), .B(g23666), .Z(g24713) ) ;
AND2    gate14367  (.A(g6173), .B(g23699), .Z(g24714) ) ;
OR2     gate14368  (.A(g13029), .B(g10665), .Z(g15935) ) ;
AND2    gate14369  (.A(g15935), .B(g23004), .Z(g24716) ) ;
OR2     gate14370  (.A(g19206), .B(g15703), .Z(g22684) ) ;
AND2    gate14371  (.A(g22684), .B(g19777), .Z(g24717) ) ;
AND2    gate14372  (.A(g681), .B(g23530), .Z(g24719) ) ;
OR4     gate14373  (.A(g14361), .B(g14335), .C(g11954), .D(II18417), .Z(g17488) ) ;
AND2    gate14374  (.A(g17488), .B(g22369), .Z(g24721) ) ;
NAND2   gate14375  (.A(II18580), .B(II18581), .Z(g17618) ) ;
AND2    gate14376  (.A(g17618), .B(g22417), .Z(g24722) ) ;
OR4     gate14377  (.A(g14364), .B(g14337), .C(g11958), .D(II18421), .Z(g17490) ) ;
AND2    gate14378  (.A(g17490), .B(g22384), .Z(g24723) ) ;
NAND2   gate14379  (.A(II18588), .B(II18589), .Z(g17624) ) ;
AND2    gate14380  (.A(g17624), .B(g22432), .Z(g24724) ) ;
OR2     gate14381  (.A(g15700), .B(g13046), .Z(g19587) ) ;
AND2    gate14382  (.A(g19587), .B(g23012), .Z(g24725) ) ;
OR2     gate14383  (.A(g13035), .B(g10675), .Z(g15965) ) ;
AND2    gate14384  (.A(g15965), .B(g23015), .Z(g24726) ) ;
OR2     gate14385  (.A(g10656), .B(g10676), .Z(g13300) ) ;
AND2    gate14386  (.A(g13300), .B(g23016), .Z(g24727) ) ;
AND2    gate14387  (.A(g16513), .B(g23017), .Z(g24728) ) ;
AND2    gate14388  (.A(g22719), .B(g23018), .Z(g24729) ) ;
AND2    gate14389  (.A(g6177), .B(g23699), .Z(g24730) ) ;
AND2    gate14390  (.A(g6519), .B(g23733), .Z(g24731) ) ;
OR2     gate14391  (.A(g19266), .B(g15711), .Z(g22708) ) ;
AND2    gate14392  (.A(g22708), .B(g19789), .Z(g24743) ) ;
AND2    gate14393  (.A(g650), .B(g23550), .Z(g24745) ) ;
OR4     gate14394  (.A(g14393), .B(g14362), .C(g11972), .D(II18449), .Z(g17510) ) ;
AND2    gate14395  (.A(g17510), .B(g22417), .Z(g24747) ) ;
NAND2   gate14396  (.A(II18626), .B(II18627), .Z(g17656) ) ;
AND2    gate14397  (.A(g17656), .B(g22457), .Z(g24748) ) ;
OR4     gate14398  (.A(g14396), .B(g14365), .C(g11976), .D(II18452), .Z(g17511) ) ;
AND2    gate14399  (.A(g17511), .B(g22432), .Z(g24749) ) ;
NAND2   gate14400  (.A(II18634), .B(II18635), .Z(g17662) ) ;
AND2    gate14401  (.A(g17662), .B(g22472), .Z(g24750) ) ;
OR2     gate14402  (.A(g15704), .B(g13059), .Z(g19604) ) ;
AND2    gate14403  (.A(g19604), .B(g23027), .Z(g24754) ) ;
OR2     gate14404  (.A(g13048), .B(g10707), .Z(g16022) ) ;
AND2    gate14405  (.A(g16022), .B(g23030), .Z(g24755) ) ;
AND2    gate14406  (.A(g7004), .B(g23563), .Z(g24757) ) ;
AND2    gate14407  (.A(g6523), .B(g23733), .Z(g24758) ) ;
OR2     gate14408  (.A(g19333), .B(g15716), .Z(g22751) ) ;
AND2    gate14409  (.A(g22751), .B(g19852), .Z(g24761) ) ;
AND2    gate14410  (.A(g655), .B(g23573), .Z(g24762) ) ;
OR4     gate14411  (.A(g14416), .B(g14394), .C(g11995), .D(II18492), .Z(g17569) ) ;
AND2    gate14412  (.A(g17569), .B(g22457), .Z(g24763) ) ;
OR4     gate14413  (.A(g14419), .B(g14397), .C(g11999), .D(II18495), .Z(g17570) ) ;
AND2    gate14414  (.A(g17570), .B(g22472), .Z(g24764) ) ;
NAND2   gate14415  (.A(II18681), .B(II18682), .Z(g17699) ) ;
AND2    gate14416  (.A(g17699), .B(g22498), .Z(g24765) ) ;
OR2     gate14417  (.A(g15712), .B(g13080), .Z(g19619) ) ;
AND2    gate14418  (.A(g19619), .B(g23058), .Z(g24769) ) ;
AND2    gate14419  (.A(g7028), .B(g23605), .Z(g24771) ) ;
NOR2    gate14420  (.A(g13622), .B(g11144), .Z(g16287) ) ;
AND2    gate14421  (.A(g16287), .B(g23061), .Z(g24772) ) ;
OR2     gate14422  (.A(g19354), .B(g15722), .Z(g22832) ) ;
AND2    gate14423  (.A(g22832), .B(g19872), .Z(g24773) ) ;
AND2    gate14424  (.A(g718), .B(g23614), .Z(g24774) ) ;
OR4     gate14425  (.A(g14450), .B(g14420), .C(g12025), .D(II18543), .Z(g17594) ) ;
AND2    gate14426  (.A(g17594), .B(g22498), .Z(g24775) ) ;
NOR2    gate14427  (.A(g8477), .B(g8479), .Z(g11345) ) ;
AND2    gate14428  (.A(g11345), .B(g23066), .Z(g24777) ) ;
AND2    gate14429  (.A(g7051), .B(g23645), .Z(g24785) ) ;
AND2    gate14430  (.A(g661), .B(g23654), .Z(g24786) ) ;
NOR2    gate14431  (.A(g8538), .B(g8540), .Z(g11384) ) ;
AND2    gate14432  (.A(g11384), .B(g23111), .Z(g24788) ) ;
AND2    gate14433  (.A(g7074), .B(g23681), .Z(g24790) ) ;
NOR2    gate14434  (.A(g8591), .B(g8593), .Z(g11414) ) ;
AND2    gate14435  (.A(g11414), .B(g23138), .Z(g24794) ) ;
AND2    gate14436  (.A(g7097), .B(g23714), .Z(g24796) ) ;
OR2     gate14437  (.A(g19372), .B(g19383), .Z(g22872) ) ;
AND2    gate14438  (.A(g22872), .B(g19960), .Z(g24797) ) ;
OR2     gate14439  (.A(g19384), .B(g15745), .Z(g22901) ) ;
AND2    gate14440  (.A(g22901), .B(g20005), .Z(g24803) ) ;
AND2    gate14441  (.A(g19662), .B(g22192), .Z(g24812) ) ;
NOR2    gate14442  (.A(g19773), .B(g12970), .Z(g22929) ) ;
AND2    gate14443  (.A(g22929), .B(g7235), .Z(g24817) ) ;
NOR2    gate14444  (.A(g10262), .B(g12259), .Z(g13944) ) ;
AND2    gate14445  (.A(g13944), .B(g23978), .Z(g24820) ) ;
AND3    gate14446  (.A(g8097), .B(g8334), .C(g3045), .Z(II24003) ) ;
AND3    gate14447  (.A(g3010), .B(g23534), .C(II24003), .Z(g24822) ) ;
NOR2    gate14448  (.A(g358), .B(g365), .Z(g8720) ) ;
AND2    gate14449  (.A(g8720), .B(g23233), .Z(g24835) ) ;
AND3    gate14450  (.A(g8334), .B(g7975), .C(g3045), .Z(II24015) ) ;
AND3    gate14451  (.A(g3010), .B(g23211), .C(II24015), .Z(g24843) ) ;
AND3    gate14452  (.A(g8155), .B(g8390), .C(g3396), .Z(II24018) ) ;
AND3    gate14453  (.A(g3361), .B(g23555), .C(II24018), .Z(g24846) ) ;
AND2    gate14454  (.A(g4165), .B(g22227), .Z(g24849) ) ;
AND3    gate14455  (.A(g3029), .B(g3034), .C(g8426), .Z(II24027) ) ;
AND3    gate14456  (.A(g3050), .B(g23534), .C(II24027), .Z(g24855) ) ;
AND3    gate14457  (.A(g8390), .B(g8016), .C(g3396), .Z(II24030) ) ;
AND3    gate14458  (.A(g3361), .B(g23223), .C(II24030), .Z(g24858) ) ;
AND3    gate14459  (.A(g8219), .B(g8443), .C(g3747), .Z(II24033) ) ;
AND3    gate14460  (.A(g3712), .B(g23582), .C(II24033), .Z(g24861) ) ;
NOR2    gate14461  (.A(g4125), .B(g7765), .Z(g11201) ) ;
AND2    gate14462  (.A(g11201), .B(g22305), .Z(g24864) ) ;
NAND2   gate14463  (.A(II14351), .B(II14352), .Z(g11323) ) ;
AND2    gate14464  (.A(g11323), .B(g23253), .Z(g24865) ) ;
AND3    gate14465  (.A(g3034), .B(g3040), .C(g8426), .Z(II24048) ) ;
AND3    gate14466  (.A(g3050), .B(g23211), .C(II24048), .Z(g24881) ) ;
AND3    gate14467  (.A(g3380), .B(g3385), .C(g8492), .Z(II24051) ) ;
AND3    gate14468  (.A(g3401), .B(g23555), .C(II24051), .Z(g24884) ) ;
AND3    gate14469  (.A(g8443), .B(g8075), .C(g3747), .Z(II24054) ) ;
AND3    gate14470  (.A(g3712), .B(g23239), .C(II24054), .Z(g24887) ) ;
NAND2   gate14471  (.A(II14509), .B(II14510), .Z(g11559) ) ;
AND2    gate14472  (.A(g11559), .B(g23264), .Z(g24892) ) ;
AND3    gate14473  (.A(g3385), .B(g3391), .C(g8492), .Z(II24064) ) ;
AND3    gate14474  (.A(g3401), .B(g23223), .C(II24064), .Z(g24897) ) ;
AND3    gate14475  (.A(g3731), .B(g3736), .C(g8553), .Z(II24067) ) ;
AND3    gate14476  (.A(g3752), .B(g23582), .C(II24067), .Z(g24900) ) ;
AND2    gate14477  (.A(g128), .B(g23889), .Z(g24903) ) ;
NAND2   gate14478  (.A(II14610), .B(II14611), .Z(g11761) ) ;
AND2    gate14479  (.A(g11761), .B(g23279), .Z(g24904) ) ;
AND3    gate14480  (.A(g3736), .B(g3742), .C(g8553), .Z(II24075) ) ;
AND3    gate14481  (.A(g3752), .B(g23239), .C(II24075), .Z(g24908) ) ;
OR3     gate14482  (.A(g21384), .B(g21363), .C(II22830), .Z(g23687) ) ;
AND2    gate14483  (.A(g23687), .B(g20682), .Z(g24912) ) ;
AND2    gate14484  (.A(g4821), .B(g23908), .Z(g24913) ) ;
AND2    gate14485  (.A(g8721), .B(g23301), .Z(g24914) ) ;
OR2     gate14486  (.A(g19487), .B(g15852), .Z(g23087) ) ;
AND2    gate14487  (.A(g23087), .B(g20158), .Z(g24915) ) ;
OR3     gate14488  (.A(g21401), .B(g21385), .C(II22852), .Z(g23721) ) ;
AND2    gate14489  (.A(g23721), .B(g20739), .Z(g24921) ) ;
AND2    gate14490  (.A(g4831), .B(g23931), .Z(g24922) ) ;
OR2     gate14491  (.A(g19500), .B(g15863), .Z(g23129) ) ;
AND2    gate14492  (.A(g23129), .B(g20167), .Z(g24923) ) ;
OR3     gate14493  (.A(g21415), .B(g21402), .C(II22880), .Z(g23751) ) ;
AND2    gate14494  (.A(g23751), .B(g20875), .Z(g24929) ) ;
AND2    gate14495  (.A(g4826), .B(g23948), .Z(g24930) ) ;
OR2     gate14496  (.A(g19521), .B(g15876), .Z(g23153) ) ;
AND2    gate14497  (.A(g23153), .B(g20178), .Z(g24931) ) ;
OR3     gate14498  (.A(g21432), .B(g21416), .C(II22912), .Z(g23771) ) ;
AND2    gate14499  (.A(g23771), .B(g21012), .Z(g24939) ) ;
AND2    gate14500  (.A(g5011), .B(g23971), .Z(g24940) ) ;
OR2     gate14501  (.A(g19536), .B(g15903), .Z(g23171) ) ;
AND2    gate14502  (.A(g23171), .B(g20190), .Z(g24941) ) ;
OR2     gate14503  (.A(g19545), .B(g15911), .Z(g23183) ) ;
AND2    gate14504  (.A(g23183), .B(g20197), .Z(g24945) ) ;
OR3     gate14505  (.A(g21462), .B(g21433), .C(II22958), .Z(g23796) ) ;
AND2    gate14506  (.A(g23796), .B(g20751), .Z(g24949) ) ;
OR2     gate14507  (.A(g19556), .B(g15937), .Z(g23193) ) ;
AND2    gate14508  (.A(g23193), .B(g20209), .Z(g24961) ) ;
OR2     gate14509  (.A(g19564), .B(g19578), .Z(g23194) ) ;
AND2    gate14510  (.A(g23194), .B(g20210), .Z(g24962) ) ;
OR2     gate14511  (.A(g19571), .B(g15966), .Z(g23197) ) ;
AND2    gate14512  (.A(g23197), .B(g20213), .Z(g24967) ) ;
OR2     gate14513  (.A(g19585), .B(g19601), .Z(g23209) ) ;
AND2    gate14514  (.A(g23209), .B(g20232), .Z(g24977) ) ;
OR2     gate14515  (.A(g19588), .B(g16023), .Z(g23217) ) ;
AND2    gate14516  (.A(g23217), .B(g20238), .Z(g24983) ) ;
AND2    gate14517  (.A(g22929), .B(g12818), .Z(g24984) ) ;
NAND2   gate14518  (.A(g14520), .B(g14489), .Z(g17412) ) ;
AND2    gate14519  (.A(g17412), .B(g23408), .Z(g24998) ) ;
NAND3   gate14520  (.A(g14342), .B(g17220), .C(g9372), .Z(g20644) ) ;
AND2    gate14521  (.A(g20644), .B(g23419), .Z(g25012) ) ;
NAND2   gate14522  (.A(g14547), .B(g14521), .Z(g17474) ) ;
AND2    gate14523  (.A(g17474), .B(g23420), .Z(g25014) ) ;
OR2     gate14524  (.A(g19637), .B(g16098), .Z(g23251) ) ;
AND2    gate14525  (.A(g23251), .B(g20432), .Z(g25030) ) ;
NAND3   gate14526  (.A(g14377), .B(g17246), .C(g9442), .Z(g20675) ) ;
AND2    gate14527  (.A(g20675), .B(g23432), .Z(g25031) ) ;
NAND2   gate14528  (.A(g14573), .B(g14548), .Z(g17500) ) ;
AND2    gate14529  (.A(g17500), .B(g23433), .Z(g25033) ) ;
AND2    gate14530  (.A(g12738), .B(g23443), .Z(g25040) ) ;
OR2     gate14531  (.A(g19660), .B(g16125), .Z(g23261) ) ;
AND2    gate14532  (.A(g23261), .B(g20494), .Z(g25041) ) ;
OR2     gate14533  (.A(g19661), .B(g16126), .Z(g23262) ) ;
AND2    gate14534  (.A(g23262), .B(g20496), .Z(g25042) ) ;
NAND3   gate14535  (.A(g14406), .B(g17290), .C(g9509), .Z(g20733) ) ;
AND2    gate14536  (.A(g20733), .B(g23447), .Z(g25043) ) ;
NAND2   gate14537  (.A(g14600), .B(g14574), .Z(g17525) ) ;
AND2    gate14538  (.A(g17525), .B(g23448), .Z(g25045) ) ;
NOR2    gate14539  (.A(g7400), .B(g10741), .Z(g13056) ) ;
AND2    gate14540  (.A(g13056), .B(g22312), .Z(g25050) ) ;
AND2    gate14541  (.A(g12778), .B(g23452), .Z(g25054) ) ;
AND2    gate14542  (.A(g12779), .B(g23456), .Z(g25056) ) ;
OR2     gate14543  (.A(g19680), .B(g16160), .Z(g23275) ) ;
AND2    gate14544  (.A(g23275), .B(g20511), .Z(g25057) ) ;
OR2     gate14545  (.A(g19681), .B(g16161), .Z(g23276) ) ;
AND2    gate14546  (.A(g23276), .B(g20513), .Z(g25058) ) ;
NAND3   gate14547  (.A(g14432), .B(g17315), .C(g9567), .Z(g20870) ) ;
AND2    gate14548  (.A(g20870), .B(g23460), .Z(g25059) ) ;
NAND2   gate14549  (.A(g14638), .B(g14601), .Z(g17586) ) ;
AND2    gate14550  (.A(g17586), .B(g23461), .Z(g25061) ) ;
NOR2    gate14551  (.A(g7446), .B(g10762), .Z(g13078) ) ;
AND2    gate14552  (.A(g13078), .B(g22325), .Z(g25063) ) ;
AND2    gate14553  (.A(g4722), .B(g22885), .Z(g25067) ) ;
AND2    gate14554  (.A(g17574), .B(g23477), .Z(g25068) ) ;
OR2     gate14555  (.A(g19691), .B(g16177), .Z(g23296) ) ;
AND2    gate14556  (.A(g23296), .B(g20535), .Z(g25069) ) ;
AND2    gate14557  (.A(g12804), .B(g23478), .Z(g25071) ) ;
AND2    gate14558  (.A(g12805), .B(g23479), .Z(g25076) ) ;
OR2     gate14559  (.A(g19692), .B(g16178), .Z(g23297) ) ;
AND2    gate14560  (.A(g23297), .B(g20536), .Z(g25077) ) ;
OR2     gate14561  (.A(g19693), .B(g16179), .Z(g23298) ) ;
AND2    gate14562  (.A(g23298), .B(g20538), .Z(g25078) ) ;
NAND3   gate14563  (.A(g14504), .B(g17399), .C(g9629), .Z(g21011) ) ;
AND2    gate14564  (.A(g21011), .B(g23483), .Z(g25079) ) ;
AND2    gate14565  (.A(g4737), .B(g22885), .Z(g25084) ) ;
AND2    gate14566  (.A(g4912), .B(g22908), .Z(g25085) ) ;
OR2     gate14567  (.A(g11019), .B(g11023), .Z(g13941) ) ;
AND2    gate14568  (.A(g13941), .B(g23488), .Z(g25086) ) ;
AND2    gate14569  (.A(g17307), .B(g23489), .Z(g25087) ) ;
AND2    gate14570  (.A(g17601), .B(g23491), .Z(g25088) ) ;
OR2     gate14571  (.A(g19715), .B(g16191), .Z(g23317) ) ;
AND2    gate14572  (.A(g23317), .B(g20553), .Z(g25089) ) ;
AND2    gate14573  (.A(g12830), .B(g23492), .Z(g25091) ) ;
AND2    gate14574  (.A(g12831), .B(g23493), .Z(g25093) ) ;
OR2     gate14575  (.A(g19716), .B(g16192), .Z(g23318) ) ;
AND2    gate14576  (.A(g23318), .B(g20554), .Z(g25094) ) ;
OR2     gate14577  (.A(g19717), .B(g16193), .Z(g23319) ) ;
AND2    gate14578  (.A(g23319), .B(g20556), .Z(g25095) ) ;
NAND2   gate14579  (.A(II22922), .B(II22923), .Z(g23778) ) ;
AND2    gate14580  (.A(g23778), .B(g20560), .Z(g25096) ) ;
AND2    gate14581  (.A(g4727), .B(g22885), .Z(g25102) ) ;
AND2    gate14582  (.A(g4927), .B(g22908), .Z(g25103) ) ;
OR2     gate14583  (.A(g13436), .B(g11027), .Z(g16800) ) ;
AND2    gate14584  (.A(g16800), .B(g23504), .Z(g25104) ) ;
OR2     gate14585  (.A(g11024), .B(g11028), .Z(g13973) ) ;
AND2    gate14586  (.A(g13973), .B(g23505), .Z(g25105) ) ;
AND2    gate14587  (.A(g17391), .B(g23506), .Z(g25106) ) ;
AND2    gate14588  (.A(g17643), .B(g23508), .Z(g25107) ) ;
OR2     gate14589  (.A(g19735), .B(g16203), .Z(g23345) ) ;
AND2    gate14590  (.A(g23345), .B(g20576), .Z(g25108) ) ;
AND2    gate14591  (.A(g10427), .B(g23509), .Z(g25110) ) ;
AND2    gate14592  (.A(g10428), .B(g23510), .Z(g25112) ) ;
OR2     gate14593  (.A(g19736), .B(g16204), .Z(g23346) ) ;
AND2    gate14594  (.A(g23346), .B(g20577), .Z(g25113) ) ;
OR2     gate14595  (.A(g19767), .B(g13514), .Z(g23374) ) ;
AND2    gate14596  (.A(g23374), .B(g20592), .Z(g25122) ) ;
AND2    gate14597  (.A(g4732), .B(g22885), .Z(g25123) ) ;
AND2    gate14598  (.A(g4917), .B(g22908), .Z(g25124) ) ;
OR2     gate14599  (.A(g16202), .B(g13491), .Z(g20187) ) ;
AND2    gate14600  (.A(g20187), .B(g23520), .Z(g25125) ) ;
OR2     gate14601  (.A(g13473), .B(g11035), .Z(g16839) ) ;
AND2    gate14602  (.A(g16839), .B(g23523), .Z(g25126) ) ;
OR2     gate14603  (.A(g11029), .B(g11036), .Z(g13997) ) ;
AND2    gate14604  (.A(g13997), .B(g23524), .Z(g25127) ) ;
AND2    gate14605  (.A(g17418), .B(g23525), .Z(g25128) ) ;
AND2    gate14606  (.A(g17682), .B(g23527), .Z(g25129) ) ;
OR2     gate14607  (.A(g19746), .B(g16212), .Z(g23358) ) ;
AND2    gate14608  (.A(g23358), .B(g20600), .Z(g25130) ) ;
AND2    gate14609  (.A(g10497), .B(g23528), .Z(g25132) ) ;
AND2    gate14610  (.A(g4717), .B(g22885), .Z(g25142) ) ;
AND2    gate14611  (.A(g4922), .B(g22908), .Z(g25143) ) ;
OR2     gate14612  (.A(g16211), .B(g13507), .Z(g20202) ) ;
AND2    gate14613  (.A(g20202), .B(g23542), .Z(g25147) ) ;
OR2     gate14614  (.A(g13493), .B(g11045), .Z(g16867) ) ;
AND2    gate14615  (.A(g16867), .B(g23545), .Z(g25148) ) ;
OR2     gate14616  (.A(g11037), .B(g11046), .Z(g14030) ) ;
AND2    gate14617  (.A(g14030), .B(g23546), .Z(g25149) ) ;
AND2    gate14618  (.A(g17480), .B(g23547), .Z(g25150) ) ;
AND2    gate14619  (.A(g17719), .B(g23549), .Z(g25151) ) ;
OR2     gate14620  (.A(g19756), .B(g16222), .Z(g23383) ) ;
AND2    gate14621  (.A(g23383), .B(g20626), .Z(g25152) ) ;
AND2    gate14622  (.A(g4907), .B(g22908), .Z(g25159) ) ;
OR2     gate14623  (.A(g16221), .B(g13523), .Z(g20217) ) ;
AND2    gate14624  (.A(g20217), .B(g23566), .Z(g25163) ) ;
OR2     gate14625  (.A(g13509), .B(g11115), .Z(g16883) ) ;
AND2    gate14626  (.A(g16883), .B(g23569), .Z(g25164) ) ;
OR2     gate14627  (.A(g11047), .B(g11116), .Z(g14062) ) ;
AND2    gate14628  (.A(g14062), .B(g23570), .Z(g25165) ) ;
AND2    gate14629  (.A(g17506), .B(g23571), .Z(g25166) ) ;
NOR2    gate14630  (.A(g9776), .B(g9778), .Z(g12234) ) ;
AND2    gate14631  (.A(g12234), .B(g23589), .Z(g25173) ) ;
OR2     gate14632  (.A(g16233), .B(g13541), .Z(g20241) ) ;
AND2    gate14633  (.A(g20241), .B(g23608), .Z(g25178) ) ;
OR2     gate14634  (.A(g13525), .B(g11127), .Z(g16928) ) ;
AND2    gate14635  (.A(g16928), .B(g23611), .Z(g25179) ) ;
OR2     gate14636  (.A(g19791), .B(g16245), .Z(g23405) ) ;
AND2    gate14637  (.A(g23405), .B(g20696), .Z(g25181) ) ;
NOR2    gate14638  (.A(g9860), .B(g9862), .Z(g12296) ) ;
AND2    gate14639  (.A(g12296), .B(g23629), .Z(g25187) ) ;
OR2     gate14640  (.A(g16243), .B(g13566), .Z(g20276) ) ;
AND2    gate14641  (.A(g20276), .B(g23648), .Z(g25192) ) ;
NOR2    gate14642  (.A(g9931), .B(g9933), .Z(g12346) ) ;
AND2    gate14643  (.A(g12346), .B(g23665), .Z(g25201) ) ;
NOR2    gate14644  (.A(g1002), .B(g19699), .Z(g22513) ) ;
AND2    gate14645  (.A(g22513), .B(g10621), .Z(g25207) ) ;
NOR2    gate14646  (.A(g9999), .B(g10001), .Z(g12418) ) ;
AND2    gate14647  (.A(g12418), .B(g23698), .Z(g25217) ) ;
NOR2    gate14648  (.A(g1345), .B(g19720), .Z(g22523) ) ;
AND2    gate14649  (.A(g22523), .B(g10652), .Z(g25223) ) ;
AND2    gate14650  (.A(g7636), .B(g22654), .Z(g25229) ) ;
NOR2    gate14651  (.A(g10057), .B(g10059), .Z(g12466) ) ;
AND2    gate14652  (.A(g12466), .B(g23732), .Z(g25238) ) ;
OR2     gate14653  (.A(g21188), .B(g17469), .Z(g22152) ) ;
AND2    gate14654  (.A(g22152), .B(g13061), .Z(g25285) ) ;
AND3    gate14655  (.A(g9364), .B(g9607), .C(g5057), .Z(II24482) ) ;
AND3    gate14656  (.A(g5022), .B(g22173), .C(II24482), .Z(g25290) ) ;
AND2    gate14657  (.A(g6888), .B(g22359), .Z(g25323) ) ;
AND3    gate14658  (.A(g9607), .B(g9229), .C(g5057), .Z(II24505) ) ;
AND3    gate14659  (.A(g5022), .B(g23764), .C(II24505), .Z(g25328) ) ;
AND3    gate14660  (.A(g9434), .B(g9672), .C(g5401), .Z(II24508) ) ;
AND3    gate14661  (.A(g5366), .B(g22194), .C(II24508), .Z(g25331) ) ;
NAND2   gate14662  (.A(II22973), .B(II22974), .Z(g23810) ) ;
NAND2   gate14663  (.A(II22945), .B(II22946), .Z(g23786) ) ;
AND2    gate14664  (.A(g23810), .B(g23786), .Z(g25357) ) ;
AND2    gate14665  (.A(g7733), .B(g22406), .Z(g25366) ) ;
AND2    gate14666  (.A(g6946), .B(g22407), .Z(g25367) ) ;
AND2    gate14667  (.A(g6946), .B(g22408), .Z(g25368) ) ;
AND3    gate14668  (.A(g5041), .B(g5046), .C(g9716), .Z(II24524) ) ;
AND3    gate14669  (.A(g5062), .B(g22173), .C(II24524), .Z(g25371) ) ;
AND3    gate14670  (.A(g9672), .B(g9264), .C(g5401), .Z(II24527) ) ;
AND3    gate14671  (.A(g5366), .B(g23789), .C(II24527), .Z(g25374) ) ;
AND3    gate14672  (.A(g9501), .B(g9733), .C(g5747), .Z(II24530) ) ;
AND3    gate14673  (.A(g5712), .B(g22210), .C(II24530), .Z(g25377) ) ;
AND2    gate14674  (.A(g22682), .B(g9772), .Z(g25408) ) ;
AND3    gate14675  (.A(g5046), .B(g5052), .C(g9716), .Z(II24546) ) ;
AND3    gate14676  (.A(g5062), .B(g23764), .C(II24546), .Z(g25411) ) ;
AND3    gate14677  (.A(g5385), .B(g5390), .C(g9792), .Z(II24549) ) ;
AND3    gate14678  (.A(g5406), .B(g22194), .C(II24549), .Z(g25414) ) ;
AND3    gate14679  (.A(g9733), .B(g9316), .C(g5747), .Z(II24552) ) ;
AND3    gate14680  (.A(g5712), .B(g23816), .C(II24552), .Z(g25417) ) ;
AND3    gate14681  (.A(g9559), .B(g9809), .C(g6093), .Z(II24555) ) ;
AND3    gate14682  (.A(g6058), .B(g22220), .C(II24555), .Z(g25420) ) ;
AND2    gate14683  (.A(g6946), .B(g22496), .Z(g25449) ) ;
AND2    gate14684  (.A(g6888), .B(g22497), .Z(g25450) ) ;
AND3    gate14685  (.A(g5390), .B(g5396), .C(g9792), .Z(II24576) ) ;
AND3    gate14686  (.A(g5406), .B(g23789), .C(II24576), .Z(g25453) ) ;
AND3    gate14687  (.A(g5731), .B(g5736), .C(g9875), .Z(II24579) ) ;
AND3    gate14688  (.A(g5752), .B(g22210), .C(II24579), .Z(g25456) ) ;
AND3    gate14689  (.A(g9809), .B(g9397), .C(g6093), .Z(II24582) ) ;
AND3    gate14690  (.A(g6058), .B(g23844), .C(II24582), .Z(g25459) ) ;
AND3    gate14691  (.A(g9621), .B(g9892), .C(g6439), .Z(II24585) ) ;
AND3    gate14692  (.A(g6404), .B(g22300), .C(II24585), .Z(g25462) ) ;
OR2     gate14693  (.A(g20093), .B(g20108), .Z(g23574) ) ;
AND2    gate14694  (.A(g23574), .B(g21346), .Z(g25466) ) ;
AND2    gate14695  (.A(g22646), .B(g9917), .Z(g25479) ) ;
AND3    gate14696  (.A(g5736), .B(g5742), .C(g9875), .Z(II24597) ) ;
AND3    gate14697  (.A(g5752), .B(g23816), .C(II24597), .Z(g25482) ) ;
AND3    gate14698  (.A(g6077), .B(g6082), .C(g9946), .Z(II24600) ) ;
AND3    gate14699  (.A(g6098), .B(g22220), .C(II24600), .Z(g25485) ) ;
AND3    gate14700  (.A(g9892), .B(g9467), .C(g6439), .Z(II24603) ) ;
AND3    gate14701  (.A(g6404), .B(g23865), .C(II24603), .Z(g25488) ) ;
OR2     gate14702  (.A(g20109), .B(g20131), .Z(g23615) ) ;
AND2    gate14703  (.A(g23615), .B(g21355), .Z(g25491) ) ;
AND2    gate14704  (.A(g6946), .B(g22527), .Z(g25502) ) ;
AND2    gate14705  (.A(g6888), .B(g22529), .Z(g25503) ) ;
AND3    gate14706  (.A(g6082), .B(g6088), .C(g9946), .Z(II24616) ) ;
AND3    gate14707  (.A(g6098), .B(g23844), .C(II24616), .Z(g25507) ) ;
AND3    gate14708  (.A(g6423), .B(g6428), .C(g10014), .Z(II24619) ) ;
AND3    gate14709  (.A(g6444), .B(g22300), .C(II24619), .Z(g25510) ) ;
AND3    gate14710  (.A(g6428), .B(g6434), .C(g10014), .Z(II24625) ) ;
AND3    gate14711  (.A(g6444), .B(g23865), .C(II24625), .Z(g25518) ) ;
AND2    gate14712  (.A(g6888), .B(g22544), .Z(g25522) ) ;
OR2     gate14713  (.A(g20165), .B(g16801), .Z(g23720) ) ;
AND2    gate14714  (.A(g23720), .B(g21400), .Z(g25526) ) ;
OR2     gate14715  (.A(g20174), .B(g16840), .Z(g23750) ) ;
AND2    gate14716  (.A(g23750), .B(g21414), .Z(g25530) ) ;
OR2     gate14717  (.A(g20188), .B(g16868), .Z(g23770) ) ;
AND2    gate14718  (.A(g23770), .B(g21431), .Z(g25536) ) ;
OR2     gate14719  (.A(g20203), .B(g16884), .Z(g23795) ) ;
AND2    gate14720  (.A(g23795), .B(g21461), .Z(g25543) ) ;
OR2     gate14721  (.A(g20218), .B(g16929), .Z(g23822) ) ;
AND2    gate14722  (.A(g23822), .B(g21511), .Z(g25551) ) ;
NOR2    gate14723  (.A(g7933), .B(g10741), .Z(g13004) ) ;
AND2    gate14724  (.A(g13004), .B(g22649), .Z(g25559) ) ;
NOR2    gate14725  (.A(g7957), .B(g10762), .Z(g13013) ) ;
AND2    gate14726  (.A(g13013), .B(g22660), .Z(g25565) ) ;
AND4    gate14727  (.A(g19919), .B(g24019), .C(g24020), .D(g24021), .Z(II24674) ) ;
AND4    gate14728  (.A(g24022), .B(g24023), .C(g24024), .D(g24025), .Z(II24675) ) ;
AND2    gate14729  (.A(II24674), .B(II24675), .Z(g25567) ) ;
AND4    gate14730  (.A(g19968), .B(g24026), .C(g24027), .D(g24028), .Z(II24679) ) ;
AND4    gate14731  (.A(g24029), .B(g24030), .C(g24031), .D(g24032), .Z(II24680) ) ;
AND2    gate14732  (.A(II24679), .B(II24680), .Z(g25568) ) ;
AND4    gate14733  (.A(g20014), .B(g24033), .C(g24034), .D(g24035), .Z(II24684) ) ;
AND4    gate14734  (.A(g24036), .B(g24037), .C(g24038), .D(g24039), .Z(II24685) ) ;
AND2    gate14735  (.A(II24684), .B(II24685), .Z(g25569) ) ;
AND4    gate14736  (.A(g20841), .B(g24040), .C(g24041), .D(g24042), .Z(II24689) ) ;
AND4    gate14737  (.A(g24043), .B(g24044), .C(g24045), .D(g24046), .Z(II24690) ) ;
AND2    gate14738  (.A(II24689), .B(II24690), .Z(g25570) ) ;
AND4    gate14739  (.A(g20982), .B(g24047), .C(g24048), .D(g24049), .Z(II24694) ) ;
AND4    gate14740  (.A(g24050), .B(g24051), .C(g24052), .D(g24053), .Z(II24695) ) ;
AND2    gate14741  (.A(II24694), .B(II24695), .Z(g25571) ) ;
AND4    gate14742  (.A(g21127), .B(g24054), .C(g24055), .D(g24056), .Z(II24699) ) ;
AND4    gate14743  (.A(g24057), .B(g24058), .C(g24059), .D(g24060), .Z(II24700) ) ;
AND2    gate14744  (.A(II24699), .B(II24700), .Z(g25572) ) ;
AND4    gate14745  (.A(g21193), .B(g24061), .C(g24062), .D(g24063), .Z(II24704) ) ;
AND4    gate14746  (.A(g24064), .B(g24065), .C(g24066), .D(g24067), .Z(II24705) ) ;
AND2    gate14747  (.A(II24704), .B(II24705), .Z(g25573) ) ;
AND4    gate14748  (.A(g21256), .B(g24068), .C(g24069), .D(g24070), .Z(II24709) ) ;
AND4    gate14749  (.A(g24071), .B(g24072), .C(g24073), .D(g24074), .Z(II24710) ) ;
AND2    gate14750  (.A(II24709), .B(II24710), .Z(g25574) ) ;
AND2    gate14751  (.A(g19402), .B(g24146), .Z(g25578) ) ;
AND2    gate14752  (.A(g19422), .B(g24147), .Z(g25579) ) ;
AND2    gate14753  (.A(g19268), .B(g24149), .Z(g25580) ) ;
AND2    gate14754  (.A(g19338), .B(g24150), .Z(g25581) ) ;
NAND2   gate14755  (.A(g21345), .B(g23363), .Z(g24989) ) ;
NAND2   gate14756  (.A(g21272), .B(g23462), .Z(g24973) ) ;
AND2    gate14757  (.A(g24989), .B(g24973), .Z(g25765) ) ;
AND2    gate14758  (.A(g2912), .B(g24560), .Z(g25768) ) ;
NAND2   gate14759  (.A(g21354), .B(g23363), .Z(g24944) ) ;
NAND2   gate14760  (.A(g21283), .B(g23462), .Z(g24934) ) ;
AND2    gate14761  (.A(g24944), .B(g24934), .Z(g25772) ) ;
AND2    gate14762  (.A(g2922), .B(g24568), .Z(g25775) ) ;
NAND2   gate14763  (.A(g21360), .B(g23363), .Z(g25532) ) ;
NAND2   gate14764  (.A(g21294), .B(g23462), .Z(g25527) ) ;
AND2    gate14765  (.A(g25532), .B(g25527), .Z(g25780) ) ;
AND2    gate14766  (.A(g2936), .B(g24571), .Z(g25782) ) ;
NAND2   gate14767  (.A(II23950), .B(II23951), .Z(g24792) ) ;
AND2    gate14768  (.A(g24792), .B(g20887), .Z(g25787) ) ;
NAND2   gate14769  (.A(II12345), .B(II12346), .Z(g8010) ) ;
AND2    gate14770  (.A(g8010), .B(g24579), .Z(g25788) ) ;
AND2    gate14771  (.A(g8097), .B(g24585), .Z(g25801) ) ;
AND2    gate14772  (.A(g8106), .B(g24586), .Z(g25802) ) ;
NAND2   gate14773  (.A(II23962), .B(II23963), .Z(g24798) ) ;
AND2    gate14774  (.A(g24798), .B(g21024), .Z(g25803) ) ;
NAND2   gate14775  (.A(II12373), .B(II12374), .Z(g8069) ) ;
AND2    gate14776  (.A(g8069), .B(g24587), .Z(g25804) ) ;
NAND2   gate14777  (.A(II23918), .B(II23919), .Z(g24760) ) ;
AND2    gate14778  (.A(g24760), .B(g13323), .Z(g25814) ) ;
AND2    gate14779  (.A(g8155), .B(g24603), .Z(g25815) ) ;
AND2    gate14780  (.A(g8164), .B(g24604), .Z(g25816) ) ;
NAND2   gate14781  (.A(II23979), .B(II23980), .Z(g24807) ) ;
AND2    gate14782  (.A(g24807), .B(g21163), .Z(g25817) ) ;
NAND2   gate14783  (.A(II12402), .B(II12403), .Z(g8124) ) ;
AND2    gate14784  (.A(g8124), .B(g24605), .Z(g25818) ) ;
AND2    gate14785  (.A(g3151), .B(g24623), .Z(g25831) ) ;
AND2    gate14786  (.A(g8219), .B(g24625), .Z(g25832) ) ;
AND2    gate14787  (.A(g8228), .B(g24626), .Z(g25833) ) ;
OR2     gate14788  (.A(g23531), .B(g20628), .Z(g25539) ) ;
AND2    gate14789  (.A(g25539), .B(g18977), .Z(g25848) ) ;
AND2    gate14790  (.A(g3502), .B(g24636), .Z(g25850) ) ;
OR2     gate14791  (.A(g23551), .B(g20658), .Z(g25545) ) ;
AND2    gate14792  (.A(g25545), .B(g18991), .Z(g25865) ) ;
AND2    gate14793  (.A(g3853), .B(g24648), .Z(g25866) ) ;
OR2     gate14794  (.A(g21419), .B(g23996), .Z(g24840) ) ;
AND2    gate14795  (.A(g24840), .B(g16182), .Z(g25870) ) ;
AND2    gate14796  (.A(g8334), .B(g24804), .Z(g25871) ) ;
AND2    gate14797  (.A(g3119), .B(g24655), .Z(g25872) ) ;
OR2     gate14798  (.A(g21453), .B(g24002), .Z(g24854) ) ;
AND2    gate14799  (.A(g24854), .B(g16197), .Z(g25873) ) ;
NAND2   gate14800  (.A(II14170), .B(II14171), .Z(g11118) ) ;
AND2    gate14801  (.A(g11118), .B(g24665), .Z(g25874) ) ;
AND2    gate14802  (.A(g8390), .B(g24809), .Z(g25875) ) ;
AND2    gate14803  (.A(g3470), .B(g24667), .Z(g25876) ) ;
NAND2   gate14804  (.A(II14186), .B(II14187), .Z(g11135) ) ;
AND2    gate14805  (.A(g11135), .B(g24683), .Z(g25879) ) ;
AND2    gate14806  (.A(g8443), .B(g24814), .Z(g25880) ) ;
AND2    gate14807  (.A(g3821), .B(g24685), .Z(g25881) ) ;
OR2     gate14808  (.A(g6804), .B(g12527), .Z(g13728) ) ;
AND2    gate14809  (.A(g13728), .B(g24699), .Z(g25883) ) ;
NAND2   gate14810  (.A(II14205), .B(II14206), .Z(g11153) ) ;
AND2    gate14811  (.A(g11153), .B(g24711), .Z(g25884) ) ;
OR2     gate14812  (.A(g23779), .B(g21285), .Z(g24390) ) ;
AND2    gate14813  (.A(g24390), .B(g19368), .Z(g25900) ) ;
OR2     gate14814  (.A(g21452), .B(g24001), .Z(g24853) ) ;
AND2    gate14815  (.A(g24853), .B(g16290), .Z(g25901) ) ;
OR2     gate14816  (.A(g23801), .B(g21296), .Z(g24398) ) ;
AND2    gate14817  (.A(g24398), .B(g19373), .Z(g25902) ) ;
NOR2    gate14818  (.A(g739), .B(g11083), .Z(g14001) ) ;
AND2    gate14819  (.A(g14001), .B(g24791), .Z(g25904) ) ;
OR2     gate14820  (.A(g21465), .B(g24009), .Z(g24879) ) ;
AND2    gate14821  (.A(g24879), .B(g16311), .Z(g25905) ) ;
OR2     gate14822  (.A(g23901), .B(g23921), .Z(g24799) ) ;
AND2    gate14823  (.A(g24799), .B(g22519), .Z(g25907) ) ;
OR2     gate14824  (.A(g23857), .B(g23872), .Z(g24782) ) ;
AND2    gate14825  (.A(g24782), .B(g22520), .Z(g25908) ) ;
AND2    gate14826  (.A(g8745), .B(g24875), .Z(g25909) ) ;
NAND4   gate14827  (.A(g20172), .B(g20163), .C(g23357), .D(g13995), .Z(g24926) ) ;
AND2    gate14828  (.A(g24926), .B(g9602), .Z(g25915) ) ;
OR2     gate14829  (.A(g23900), .B(g21361), .Z(g24432) ) ;
AND2    gate14830  (.A(g24432), .B(g19434), .Z(g25916) ) ;
NAND4   gate14831  (.A(g20186), .B(g20173), .C(g23379), .D(g14029), .Z(g24936) ) ;
AND2    gate14832  (.A(g24936), .B(g9664), .Z(g25921) ) ;
NOR2    gate14833  (.A(g8858), .B(g23324), .Z(g24959) ) ;
AND2    gate14834  (.A(g24959), .B(g20065), .Z(g25922) ) ;
OR2     gate14835  (.A(g23917), .B(g21378), .Z(g24443) ) ;
AND2    gate14836  (.A(g24443), .B(g19443), .Z(g25923) ) ;
NOR2    gate14837  (.A(g671), .B(g23324), .Z(g24976) ) ;
AND2    gate14838  (.A(g24976), .B(g16846), .Z(g25924) ) ;
NOR2    gate14839  (.A(g8898), .B(g23324), .Z(g24990) ) ;
AND2    gate14840  (.A(g24990), .B(g23234), .Z(g25925) ) ;
NOR2    gate14841  (.A(g6811), .B(g23324), .Z(g25005) ) ;
AND2    gate14842  (.A(g25005), .B(g24839), .Z(g25926) ) ;
NOR2    gate14843  (.A(g676), .B(g23324), .Z(g25004) ) ;
AND2    gate14844  (.A(g25004), .B(g20375), .Z(g25927) ) ;
NOR2    gate14845  (.A(g714), .B(g23324), .Z(g25022) ) ;
AND2    gate14846  (.A(g25022), .B(g23436), .Z(g25928) ) ;
NAND2   gate14847  (.A(g22709), .B(g22687), .Z(g24574) ) ;
AND2    gate14848  (.A(g24574), .B(g19477), .Z(g25931) ) ;
AND2    gate14849  (.A(g8997), .B(g24953), .Z(g25938) ) ;
NAND2   gate14850  (.A(g22753), .B(g22711), .Z(g24583) ) ;
AND2    gate14851  (.A(g24583), .B(g19490), .Z(g25939) ) ;
OR2     gate14852  (.A(g24008), .B(g21557), .Z(g24496) ) ;
AND2    gate14853  (.A(g24496), .B(g19537), .Z(g25946) ) ;
NOR3    gate14854  (.A(g979), .B(g23024), .C(g19778), .Z(g24701) ) ;
AND2    gate14855  (.A(g24701), .B(g19559), .Z(g25949) ) ;
OR2     gate14856  (.A(g24011), .B(g21605), .Z(g24500) ) ;
AND2    gate14857  (.A(g24500), .B(g19565), .Z(g25951) ) ;
NOR3    gate14858  (.A(g1322), .B(g23051), .C(g19793), .Z(g24720) ) ;
AND2    gate14859  (.A(g24720), .B(g19580), .Z(g25955) ) ;
NOR2    gate14860  (.A(g723), .B(g14279), .Z(g17190) ) ;
AND2    gate14861  (.A(g17190), .B(g24960), .Z(g25957) ) ;
AND2    gate14862  (.A(g1648), .B(g24963), .Z(g25959) ) ;
NAND2   gate14863  (.A(II24364), .B(II24365), .Z(g25199) ) ;
AND2    gate14864  (.A(g25199), .B(g20682), .Z(g25961) ) ;
NAND2   gate14865  (.A(II13044), .B(II13045), .Z(g9258) ) ;
AND2    gate14866  (.A(g9258), .B(g24971), .Z(g25962) ) ;
AND2    gate14867  (.A(g1657), .B(g24978), .Z(g25963) ) ;
AND2    gate14868  (.A(g1783), .B(g24979), .Z(g25964) ) ;
AND2    gate14869  (.A(g2208), .B(g24980), .Z(g25965) ) ;
AND2    gate14870  (.A(g9364), .B(g24985), .Z(g25966) ) ;
AND2    gate14871  (.A(g9373), .B(g24986), .Z(g25967) ) ;
NAND2   gate14872  (.A(II24384), .B(II24385), .Z(g25215) ) ;
AND2    gate14873  (.A(g25215), .B(g20739), .Z(g25968) ) ;
NAND2   gate14874  (.A(II13078), .B(II13079), .Z(g9310) ) ;
AND2    gate14875  (.A(g9310), .B(g24987), .Z(g25969) ) ;
AND2    gate14876  (.A(g1792), .B(g24991), .Z(g25970) ) ;
AND2    gate14877  (.A(g1917), .B(g24992), .Z(g25971) ) ;
AND2    gate14878  (.A(g2217), .B(g24993), .Z(g25972) ) ;
AND2    gate14879  (.A(g2342), .B(g24994), .Z(g25973) ) ;
AND2    gate14880  (.A(g9434), .B(g24999), .Z(g25975) ) ;
AND2    gate14881  (.A(g9443), .B(g25000), .Z(g25976) ) ;
NAND2   gate14882  (.A(II24415), .B(II24416), .Z(g25236) ) ;
AND2    gate14883  (.A(g25236), .B(g20875), .Z(g25977) ) ;
NAND2   gate14884  (.A(II13110), .B(II13111), .Z(g9391) ) ;
AND2    gate14885  (.A(g9391), .B(g25001), .Z(g25978) ) ;
OR2     gate14886  (.A(g22158), .B(g18906), .Z(g24517) ) ;
AND2    gate14887  (.A(g24517), .B(g19650), .Z(g25979) ) ;
AND2    gate14888  (.A(g1926), .B(g25006), .Z(g25980) ) ;
AND2    gate14889  (.A(g2051), .B(g25007), .Z(g25981) ) ;
AND2    gate14890  (.A(g2351), .B(g25008), .Z(g25982) ) ;
AND2    gate14891  (.A(g2476), .B(g25009), .Z(g25983) ) ;
AND2    gate14892  (.A(g5160), .B(g25013), .Z(g25986) ) ;
AND2    gate14893  (.A(g9501), .B(g25015), .Z(g25987) ) ;
AND2    gate14894  (.A(g9510), .B(g25016), .Z(g25988) ) ;
NAND2   gate14895  (.A(II24439), .B(II24440), .Z(g25258) ) ;
AND2    gate14896  (.A(g25258), .B(g21012), .Z(g25989) ) ;
NAND2   gate14897  (.A(II13140), .B(II13141), .Z(g9461) ) ;
AND2    gate14898  (.A(g9461), .B(g25017), .Z(g25990) ) ;
AND2    gate14899  (.A(g2060), .B(g25023), .Z(g25991) ) ;
AND2    gate14900  (.A(g2485), .B(g25024), .Z(g25992) ) ;
AND2    gate14901  (.A(g2610), .B(g25025), .Z(g25993) ) ;
AND2    gate14902  (.A(g5507), .B(g25032), .Z(g26019) ) ;
AND2    gate14903  (.A(g9559), .B(g25034), .Z(g26020) ) ;
AND2    gate14904  (.A(g9568), .B(g25035), .Z(g26021) ) ;
NAND2   gate14905  (.A(II24462), .B(II24463), .Z(g25271) ) ;
AND2    gate14906  (.A(g25271), .B(g20751), .Z(g26022) ) ;
NAND2   gate14907  (.A(II13183), .B(II13184), .Z(g9528) ) ;
AND2    gate14908  (.A(g9528), .B(g25036), .Z(g26023) ) ;
AND2    gate14909  (.A(g2619), .B(g25039), .Z(g26024) ) ;
AND2    gate14910  (.A(g5853), .B(g25044), .Z(g26048) ) ;
AND2    gate14911  (.A(g9621), .B(g25046), .Z(g26049) ) ;
AND2    gate14912  (.A(g9630), .B(g25047), .Z(g26050) ) ;
OR2     gate14913  (.A(g22863), .B(g19684), .Z(g24896) ) ;
AND2    gate14914  (.A(g24896), .B(g14169), .Z(g26051) ) ;
AND2    gate14915  (.A(g9607), .B(g25233), .Z(g26077) ) ;
AND2    gate14916  (.A(g5128), .B(g25055), .Z(g26078) ) ;
AND2    gate14917  (.A(g6199), .B(g25060), .Z(g26079) ) ;
AND2    gate14918  (.A(g24926), .B(g9602), .Z(g26084) ) ;
NAND2   gate14919  (.A(II14713), .B(II14714), .Z(g11906) ) ;
AND2    gate14920  (.A(g11906), .B(g25070), .Z(g26085) ) ;
AND2    gate14921  (.A(g9672), .B(g25255), .Z(g26086) ) ;
AND2    gate14922  (.A(g5475), .B(g25072), .Z(g26087) ) ;
AND2    gate14923  (.A(g6545), .B(g25080), .Z(g26088) ) ;
AND2    gate14924  (.A(g1624), .B(g25081), .Z(g26090) ) ;
AND2    gate14925  (.A(g1691), .B(g25082), .Z(g26091) ) ;
AND2    gate14926  (.A(g9766), .B(g25083), .Z(g26092) ) ;
AND2    gate14927  (.A(g24936), .B(g9664), .Z(g26094) ) ;
NAND2   gate14928  (.A(II14734), .B(II14735), .Z(g11923) ) ;
AND2    gate14929  (.A(g11923), .B(g25090), .Z(g26095) ) ;
AND2    gate14930  (.A(g9733), .B(g25268), .Z(g26096) ) ;
AND2    gate14931  (.A(g5821), .B(g25092), .Z(g26097) ) ;
AND2    gate14932  (.A(g1677), .B(g25097), .Z(g26100) ) ;
AND2    gate14933  (.A(g1760), .B(g25098), .Z(g26101) ) ;
AND2    gate14934  (.A(g1825), .B(g25099), .Z(g26102) ) ;
AND2    gate14935  (.A(g2185), .B(g25100), .Z(g26103) ) ;
AND2    gate14936  (.A(g2250), .B(g25101), .Z(g26104) ) ;
NAND2   gate14937  (.A(II14765), .B(II14766), .Z(g11944) ) ;
AND2    gate14938  (.A(g11944), .B(g25109), .Z(g26119) ) ;
AND2    gate14939  (.A(g9809), .B(g25293), .Z(g26120) ) ;
AND2    gate14940  (.A(g6167), .B(g25111), .Z(g26121) ) ;
OR2     gate14941  (.A(g22308), .B(g19207), .Z(g24557) ) ;
AND2    gate14942  (.A(g24557), .B(g19762), .Z(g26122) ) ;
AND2    gate14943  (.A(g1696), .B(g25382), .Z(g26123) ) ;
AND2    gate14944  (.A(g1811), .B(g25116), .Z(g26124) ) ;
AND2    gate14945  (.A(g1894), .B(g25117), .Z(g26125) ) ;
AND2    gate14946  (.A(g1959), .B(g25118), .Z(g26126) ) ;
AND2    gate14947  (.A(g2236), .B(g25119), .Z(g26127) ) ;
AND2    gate14948  (.A(g2319), .B(g25120), .Z(g26128) ) ;
AND2    gate14949  (.A(g2384), .B(g25121), .Z(g26129) ) ;
NAND2   gate14950  (.A(g13852), .B(g22929), .Z(g24890) ) ;
AND2    gate14951  (.A(g24890), .B(g19772), .Z(g26130) ) ;
NAND2   gate14952  (.A(II14789), .B(II14790), .Z(g11962) ) ;
AND2    gate14953  (.A(g11962), .B(g25131), .Z(g26145) ) ;
AND2    gate14954  (.A(g9892), .B(g25334), .Z(g26146) ) ;
AND2    gate14955  (.A(g6513), .B(g25133), .Z(g26147) ) ;
AND4    gate14956  (.A(g25357), .B(g11724), .C(g11709), .D(g11686), .Z(g26148) ) ;
OR2     gate14957  (.A(g22309), .B(g19275), .Z(g24565) ) ;
AND2    gate14958  (.A(g24565), .B(g19780), .Z(g26153) ) ;
AND2    gate14959  (.A(g1830), .B(g25426), .Z(g26154) ) ;
AND2    gate14960  (.A(g1945), .B(g25134), .Z(g26155) ) ;
AND2    gate14961  (.A(g2028), .B(g25135), .Z(g26156) ) ;
AND2    gate14962  (.A(g2093), .B(g25136), .Z(g26157) ) ;
AND2    gate14963  (.A(g2255), .B(g25432), .Z(g26158) ) ;
AND2    gate14964  (.A(g2370), .B(g25137), .Z(g26159) ) ;
AND2    gate14965  (.A(g2453), .B(g25138), .Z(g26160) ) ;
AND2    gate14966  (.A(g2518), .B(g25139), .Z(g26161) ) ;
NAND2   gate14967  (.A(II14817), .B(II14818), .Z(g11980) ) ;
AND2    gate14968  (.A(g11980), .B(g25153), .Z(g26165) ) ;
AND4    gate14969  (.A(g25357), .B(g11724), .C(g11709), .D(g7558), .Z(g26166) ) ;
AND4    gate14970  (.A(g25357), .B(g6856), .C(g11709), .D(g11686), .Z(g26171) ) ;
AND2    gate14971  (.A(g1964), .B(g25467), .Z(g26176) ) ;
AND2    gate14972  (.A(g2079), .B(g25154), .Z(g26177) ) ;
AND2    gate14973  (.A(g2389), .B(g25473), .Z(g26178) ) ;
AND2    gate14974  (.A(g2504), .B(g25155), .Z(g26179) ) ;
AND2    gate14975  (.A(g2587), .B(g25156), .Z(g26180) ) ;
AND2    gate14976  (.A(g2652), .B(g25157), .Z(g26181) ) ;
AND2    gate14977  (.A(g9978), .B(g25317), .Z(g26182) ) ;
OR2     gate14978  (.A(g22340), .B(g13096), .Z(g24580) ) ;
AND2    gate14979  (.A(g24580), .B(g23031), .Z(g26186) ) ;
AND4    gate14980  (.A(g25357), .B(g11724), .C(g7586), .D(g11686), .Z(g26190) ) ;
AND4    gate14981  (.A(g25357), .B(g6856), .C(g11709), .D(g7558), .Z(g26195) ) ;
AND4    gate14982  (.A(g24688), .B(g10678), .C(g10658), .D(g10627), .Z(g26200) ) ;
AND2    gate14983  (.A(g1632), .B(g25337), .Z(g26203) ) ;
AND2    gate14984  (.A(g1720), .B(g25275), .Z(g26204) ) ;
AND2    gate14985  (.A(g2098), .B(g25492), .Z(g26205) ) ;
AND2    gate14986  (.A(g2523), .B(g25495), .Z(g26206) ) ;
AND2    gate14987  (.A(g2638), .B(g25170), .Z(g26207) ) ;
AND4    gate14988  (.A(g25357), .B(g11724), .C(g7586), .D(g7558), .Z(g26213) ) ;
AND4    gate14989  (.A(g25357), .B(g6856), .C(g7586), .D(g11686), .Z(g26218) ) ;
AND4    gate14990  (.A(g24688), .B(g10678), .C(g10658), .D(g8757), .Z(g26223) ) ;
AND4    gate14991  (.A(g24688), .B(g8812), .C(g10658), .D(g10627), .Z(g26226) ) ;
AND2    gate14992  (.A(g1724), .B(g25275), .Z(g26229) ) ;
AND2    gate14993  (.A(g1768), .B(g25385), .Z(g26230) ) ;
AND2    gate14994  (.A(g1854), .B(g25300), .Z(g26231) ) ;
AND2    gate14995  (.A(g2193), .B(g25396), .Z(g26232) ) ;
AND2    gate14996  (.A(g2279), .B(g25309), .Z(g26233) ) ;
AND2    gate14997  (.A(g2657), .B(g25514), .Z(g26234) ) ;
AND4    gate14998  (.A(g25357), .B(g6856), .C(g7586), .D(g7558), .Z(g26236) ) ;
AND4    gate14999  (.A(g24688), .B(g10678), .C(g8778), .D(g10627), .Z(g26241) ) ;
AND4    gate15000  (.A(g24688), .B(g8812), .C(g10658), .D(g8757), .Z(g26244) ) ;
AND2    gate15001  (.A(g1858), .B(g25300), .Z(g26249) ) ;
AND2    gate15002  (.A(g1902), .B(g25429), .Z(g26250) ) ;
AND2    gate15003  (.A(g1988), .B(g25341), .Z(g26251) ) ;
AND2    gate15004  (.A(g2283), .B(g25309), .Z(g26252) ) ;
AND2    gate15005  (.A(g2327), .B(g25435), .Z(g26253) ) ;
AND2    gate15006  (.A(g2413), .B(g25349), .Z(g26254) ) ;
AND2    gate15007  (.A(g4253), .B(g25197), .Z(g26257) ) ;
AND2    gate15008  (.A(g12875), .B(g25231), .Z(g26258) ) ;
OR2     gate15009  (.A(g23151), .B(g8234), .Z(g24430) ) ;
AND2    gate15010  (.A(g24430), .B(g25232), .Z(g26259) ) ;
AND4    gate15011  (.A(g24688), .B(g10678), .C(g8778), .D(g8757), .Z(g26261) ) ;
AND4    gate15012  (.A(g24688), .B(g8812), .C(g8778), .D(g10627), .Z(g26264) ) ;
AND2    gate15013  (.A(g1700), .B(g25275), .Z(g26270) ) ;
AND2    gate15014  (.A(g1992), .B(g25341), .Z(g26271) ) ;
AND2    gate15015  (.A(g2036), .B(g25470), .Z(g26272) ) ;
AND2    gate15016  (.A(g2122), .B(g25389), .Z(g26273) ) ;
AND2    gate15017  (.A(g2130), .B(g25210), .Z(g26274) ) ;
AND2    gate15018  (.A(g2417), .B(g25349), .Z(g26275) ) ;
AND2    gate15019  (.A(g2461), .B(g25476), .Z(g26276) ) ;
AND2    gate15020  (.A(g2547), .B(g25400), .Z(g26277) ) ;
AND2    gate15021  (.A(g4249), .B(g25213), .Z(g26279) ) ;
AND2    gate15022  (.A(g13051), .B(g25248), .Z(g26280) ) ;
AND4    gate15023  (.A(g24688), .B(g8812), .C(g8778), .D(g8757), .Z(g26281) ) ;
AND2    gate15024  (.A(g1834), .B(g25300), .Z(g26285) ) ;
AND2    gate15025  (.A(g2126), .B(g25389), .Z(g26286) ) ;
AND2    gate15026  (.A(g2138), .B(g25225), .Z(g26287) ) ;
AND2    gate15027  (.A(g2259), .B(g25309), .Z(g26288) ) ;
AND2    gate15028  (.A(g2551), .B(g25400), .Z(g26289) ) ;
AND2    gate15029  (.A(g2595), .B(g25498), .Z(g26290) ) ;
AND2    gate15030  (.A(g2681), .B(g25439), .Z(g26291) ) ;
AND2    gate15031  (.A(g2689), .B(g25228), .Z(g26292) ) ;
AND2    gate15032  (.A(g4245), .B(g25230), .Z(g26294) ) ;
AND2    gate15033  (.A(g13070), .B(g25266), .Z(g26295) ) ;
AND2    gate15034  (.A(g1968), .B(g25341), .Z(g26300) ) ;
AND2    gate15035  (.A(g2145), .B(g25244), .Z(g26301) ) ;
AND2    gate15036  (.A(g2393), .B(g25349), .Z(g26302) ) ;
AND2    gate15037  (.A(g2685), .B(g25439), .Z(g26303) ) ;
AND2    gate15038  (.A(g2697), .B(g25246), .Z(g26304) ) ;
AND2    gate15039  (.A(g13087), .B(g25286), .Z(g26306) ) ;
AND2    gate15040  (.A(g13070), .B(g25288), .Z(g26307) ) ;
AND2    gate15041  (.A(g6961), .B(g25289), .Z(g26308) ) ;
AND2    gate15042  (.A(g2102), .B(g25389), .Z(g26310) ) ;
AND2    gate15043  (.A(g2527), .B(g25400), .Z(g26311) ) ;
AND2    gate15044  (.A(g2704), .B(g25264), .Z(g26312) ) ;
NOR2    gate15045  (.A(g4467), .B(g6961), .Z(g12645) ) ;
AND2    gate15046  (.A(g12645), .B(g25326), .Z(g26313) ) ;
AND2    gate15047  (.A(g10262), .B(g25273), .Z(g26323) ) ;
AND2    gate15048  (.A(g2661), .B(g25439), .Z(g26324) ) ;
NAND2   gate15049  (.A(g10233), .B(g4531), .Z(g12644) ) ;
AND2    gate15050  (.A(g12644), .B(g25370), .Z(g26325) ) ;
NAND2   gate15051  (.A(II13730), .B(II13731), .Z(g10307) ) ;
AND2    gate15052  (.A(g10307), .B(g25480), .Z(g26336) ) ;
AND2    gate15053  (.A(g225), .B(g24836), .Z(g26339) ) ;
OR2     gate15054  (.A(g22588), .B(g19461), .Z(g24746) ) ;
AND2    gate15055  (.A(g24746), .B(g20105), .Z(g26341) ) ;
AND2    gate15056  (.A(g13051), .B(g25505), .Z(g26345) ) ;
AND2    gate15057  (.A(g262), .B(g24850), .Z(g26347) ) ;
AND2    gate15058  (.A(g13087), .B(g25517), .Z(g26350) ) ;
AND2    gate15059  (.A(g239), .B(g24869), .Z(g26351) ) ;
NAND2   gate15060  (.A(g7232), .B(g12999), .Z(g15581) ) ;
AND2    gate15061  (.A(g15581), .B(g25523), .Z(g26356) ) ;
OR2     gate15062  (.A(g16855), .B(g20215), .Z(g22547) ) ;
AND2    gate15063  (.A(g22547), .B(g25525), .Z(g26357) ) ;
OR2     gate15064  (.A(g17057), .B(g14180), .Z(g19522) ) ;
AND2    gate15065  (.A(g19522), .B(g25528), .Z(g26358) ) ;
OR2     gate15066  (.A(g7223), .B(g7201), .Z(g10589) ) ;
AND2    gate15067  (.A(g10589), .B(g25533), .Z(g26360) ) ;
OR2     gate15068  (.A(g17123), .B(g14190), .Z(g19557) ) ;
AND2    gate15069  (.A(g19557), .B(g25538), .Z(g26362) ) ;
OR2     gate15070  (.A(g17138), .B(g14202), .Z(g19576) ) ;
AND2    gate15071  (.A(g19576), .B(g25544), .Z(g26378) ) ;
OR2     gate15072  (.A(g17636), .B(g14654), .Z(g19904) ) ;
AND2    gate15073  (.A(g19904), .B(g25546), .Z(g26379) ) ;
OR2     gate15074  (.A(g17133), .B(g14193), .Z(g19572) ) ;
AND2    gate15075  (.A(g19572), .B(g25547), .Z(g26380) ) ;
AND2    gate15076  (.A(g4456), .B(g25548), .Z(g26381) ) ;
OR2     gate15077  (.A(g22685), .B(g19594), .Z(g24813) ) ;
AND2    gate15078  (.A(g24813), .B(g20231), .Z(g26387) ) ;
OR2     gate15079  (.A(g17149), .B(g14218), .Z(g19595) ) ;
AND2    gate15080  (.A(g19595), .B(g25552), .Z(g26388) ) ;
OR2     gate15081  (.A(g17671), .B(g14681), .Z(g19949) ) ;
AND2    gate15082  (.A(g19949), .B(g25553), .Z(g26389) ) ;
AND2    gate15083  (.A(g4423), .B(g25554), .Z(g26390) ) ;
OR2     gate15084  (.A(g17145), .B(g14210), .Z(g19593) ) ;
AND2    gate15085  (.A(g19593), .B(g25555), .Z(g26391) ) ;
OR2     gate15086  (.A(g16896), .B(g14097), .Z(g19467) ) ;
AND2    gate15087  (.A(g19467), .B(g25558), .Z(g26393) ) ;
OR2     gate15088  (.A(g16751), .B(g20171), .Z(g22530) ) ;
AND2    gate15089  (.A(g22530), .B(g25560), .Z(g26394) ) ;
AND2    gate15090  (.A(g22547), .B(g25561), .Z(g26395) ) ;
OR2     gate15091  (.A(g16930), .B(g14126), .Z(g19475) ) ;
AND2    gate15092  (.A(g19475), .B(g25563), .Z(g26397) ) ;
OR3     gate15093  (.A(g22360), .B(g22409), .C(g8130), .Z(g24946) ) ;
AND2    gate15094  (.A(g24946), .B(g10474), .Z(g26398) ) ;
NAND2   gate15095  (.A(g12969), .B(g7219), .Z(g15572) ) ;
AND2    gate15096  (.A(g15572), .B(g25566), .Z(g26399) ) ;
OR2     gate15097  (.A(g16965), .B(g14148), .Z(g19488) ) ;
AND2    gate15098  (.A(g19488), .B(g24356), .Z(g26423) ) ;
AND2    gate15099  (.A(g24946), .B(g8841), .Z(g26484) ) ;
OR3     gate15100  (.A(g22360), .B(g22409), .C(g23389), .Z(g24968) ) ;
AND2    gate15101  (.A(g24968), .B(g10502), .Z(g26485) ) ;
AND2    gate15102  (.A(g4423), .B(g24358), .Z(g26486) ) ;
NAND2   gate15103  (.A(g13066), .B(g7293), .Z(g15702) ) ;
AND2    gate15104  (.A(g15702), .B(g24359), .Z(g26487) ) ;
NAND4   gate15105  (.A(g15721), .B(g15715), .C(g13091), .D(g15710), .Z(g19265) ) ;
AND2    gate15106  (.A(g19265), .B(g24364), .Z(g26511) ) ;
OR2     gate15107  (.A(g16986), .B(g14168), .Z(g19501) ) ;
AND2    gate15108  (.A(g19501), .B(g24365), .Z(g26513) ) ;
AND2    gate15109  (.A(g7400), .B(g25564), .Z(g26514) ) ;
AND2    gate15110  (.A(g24968), .B(g8876), .Z(g26516) ) ;
NAND2   gate15111  (.A(g7340), .B(g13083), .Z(g15708) ) ;
AND2    gate15112  (.A(g15708), .B(g24367), .Z(g26517) ) ;
AND2    gate15113  (.A(g319), .B(g24375), .Z(g26541) ) ;
NAND2   gate15114  (.A(g7523), .B(g10759), .Z(g13102) ) ;
AND2    gate15115  (.A(g13102), .B(g24376), .Z(g26542) ) ;
NAND2   gate15116  (.A(g11002), .B(g10601), .Z(g12910) ) ;
AND2    gate15117  (.A(g12910), .B(g24377), .Z(g26543) ) ;
AND2    gate15118  (.A(g7446), .B(g24357), .Z(g26544) ) ;
NAND3   gate15119  (.A(g12440), .B(g12399), .C(g9843), .Z(g13283) ) ;
AND2    gate15120  (.A(g13283), .B(g25027), .Z(g26547) ) ;
NAND2   gate15121  (.A(II13851), .B(II13852), .Z(g10472) ) ;
AND2    gate15122  (.A(g10472), .B(g24386), .Z(g26571) ) ;
AND2    gate15123  (.A(g7443), .B(g24439), .Z(g26572) ) ;
AND2    gate15124  (.A(g7487), .B(g24453), .Z(g26602) ) ;
NAND3   gate15125  (.A(g9985), .B(g12399), .C(g9843), .Z(g13248) ) ;
AND2    gate15126  (.A(g13248), .B(g25051), .Z(g26604) ) ;
AND2    gate15127  (.A(g1018), .B(g24510), .Z(g26606) ) ;
AND2    gate15128  (.A(g14198), .B(g24405), .Z(g26610) ) ;
OR2     gate15129  (.A(g22937), .B(g19749), .Z(g24935) ) ;
AND2    gate15130  (.A(g24935), .B(g20580), .Z(g26611) ) ;
AND2    gate15131  (.A(g901), .B(g24407), .Z(g26612) ) ;
AND2    gate15132  (.A(g1361), .B(g24518), .Z(g26613) ) ;
AND2    gate15133  (.A(g14173), .B(g24418), .Z(g26629) ) ;
AND2    gate15134  (.A(g7592), .B(g24419), .Z(g26630) ) ;
AND2    gate15135  (.A(g24964), .B(g20616), .Z(g26633) ) ;
NOR2    gate15136  (.A(g23835), .B(g14645), .Z(g25321) ) ;
AND2    gate15137  (.A(g25321), .B(g20617), .Z(g26635) ) ;
NAND2   gate15138  (.A(g7537), .B(g7523), .Z(g10796) ) ;
AND2    gate15139  (.A(g10796), .B(g24424), .Z(g26650) ) ;
OR2     gate15140  (.A(g20559), .B(g17156), .Z(g22707) ) ;
AND2    gate15141  (.A(g22707), .B(g24425), .Z(g26651) ) ;
NOR2    gate15142  (.A(g347), .B(g7541), .Z(g10799) ) ;
AND2    gate15143  (.A(g10799), .B(g24426), .Z(g26652) ) ;
AND2    gate15144  (.A(g13385), .B(g24428), .Z(g26670) ) ;
AND2    gate15145  (.A(g316), .B(g24429), .Z(g26671) ) ;
NOR2    gate15146  (.A(g23871), .B(g14645), .Z(g25407) ) ;
AND2    gate15147  (.A(g25407), .B(g20673), .Z(g26684) ) ;
NOR3    gate15148  (.A(g341), .B(g7440), .C(g13385), .Z(g15754) ) ;
AND2    gate15149  (.A(g15754), .B(g24431), .Z(g26689) ) ;
NOR2    gate15150  (.A(g23686), .B(g14645), .Z(g25446) ) ;
AND2    gate15151  (.A(g25446), .B(g20713), .Z(g26711) ) ;
NOR2    gate15152  (.A(g23577), .B(g23618), .Z(g24508) ) ;
AND2    gate15153  (.A(g24508), .B(g24463), .Z(g26712) ) ;
NOR2    gate15154  (.A(g23883), .B(g14645), .Z(g25447) ) ;
AND2    gate15155  (.A(g25447), .B(g20714), .Z(g26713) ) ;
NOR2    gate15156  (.A(g7499), .B(g351), .Z(g10709) ) ;
AND2    gate15157  (.A(g10709), .B(g24438), .Z(g26719) ) ;
NOR2    gate15158  (.A(g23513), .B(g23532), .Z(g24494) ) ;
AND2    gate15159  (.A(g24494), .B(g23578), .Z(g26749) ) ;
NOR2    gate15160  (.A(g23619), .B(g23657), .Z(g24514) ) ;
AND2    gate15161  (.A(g24514), .B(g24474), .Z(g26750) ) ;
NOR2    gate15162  (.A(g14216), .B(g11890), .Z(g16024) ) ;
AND2    gate15163  (.A(g16024), .B(g24452), .Z(g26753) ) ;
NOR2    gate15164  (.A(g23918), .B(g14645), .Z(g25501) ) ;
AND2    gate15165  (.A(g25501), .B(g20923), .Z(g26778) ) ;
NOR2    gate15166  (.A(g23533), .B(g23553), .Z(g24497) ) ;
AND2    gate15167  (.A(g24497), .B(g23620), .Z(g26779) ) ;
AND2    gate15168  (.A(g4098), .B(g24437), .Z(g26780) ) ;
OR2     gate15169  (.A(g23103), .B(g19911), .Z(g25037) ) ;
AND2    gate15170  (.A(g25037), .B(g21048), .Z(g26783) ) ;
NOR2    gate15171  (.A(g23763), .B(g14645), .Z(g25247) ) ;
AND2    gate15172  (.A(g25247), .B(g21068), .Z(g26799) ) ;
NOR2    gate15173  (.A(g23955), .B(g14645), .Z(g25521) ) ;
AND2    gate15174  (.A(g25521), .B(g21185), .Z(g26808) ) ;
AND2    gate15175  (.A(g4108), .B(g24528), .Z(g26815) ) ;
AND2    gate15176  (.A(g106), .B(g24490), .Z(g26819) ) ;
OR2     gate15177  (.A(g21404), .B(g23990), .Z(g24821) ) ;
AND2    gate15178  (.A(g24821), .B(g13103), .Z(g26821) ) ;
OR2     gate15179  (.A(g21420), .B(g23998), .Z(g24841) ) ;
AND2    gate15180  (.A(g24841), .B(g13116), .Z(g26822) ) ;
OR2     gate15181  (.A(g23811), .B(g21298), .Z(g24401) ) ;
OR2     gate15182  (.A(g21558), .B(g24015), .Z(g24907) ) ;
AND2    gate15183  (.A(g24907), .B(g15747), .Z(g26826) ) ;
OR2     gate15184  (.A(g21606), .B(g22143), .Z(g24919) ) ;
AND2    gate15185  (.A(g24919), .B(g15756), .Z(g26828) ) ;
AND2    gate15186  (.A(g2844), .B(g24505), .Z(g26829) ) ;
AND2    gate15187  (.A(g2852), .B(g24509), .Z(g26833) ) ;
AND2    gate15188  (.A(g2860), .B(g24515), .Z(g26838) ) ;
AND2    gate15189  (.A(g2988), .B(g24516), .Z(g26839) ) ;
AND2    gate15190  (.A(g2894), .B(g24522), .Z(g26842) ) ;
OR2     gate15191  (.A(g23348), .B(g20193), .Z(g25261) ) ;
AND2    gate15192  (.A(g25261), .B(g21418), .Z(g26844) ) ;
NOR2    gate15193  (.A(g22190), .B(g14645), .Z(g24391) ) ;
AND2    gate15194  (.A(g24391), .B(g21426), .Z(g26845) ) ;
AND2    gate15195  (.A(g37), .B(g24524), .Z(g26846) ) ;
AND2    gate15196  (.A(g2873), .B(g24525), .Z(g26847) ) ;
AND2    gate15197  (.A(g2950), .B(g24526), .Z(g26848) ) ;
AND2    gate15198  (.A(g2994), .B(g24527), .Z(g26849) ) ;
NAND2   gate15199  (.A(g21388), .B(g23363), .Z(g24975) ) ;
NAND2   gate15200  (.A(g21330), .B(g23462), .Z(g24958) ) ;
AND2    gate15201  (.A(g24975), .B(g24958), .Z(g26852) ) ;
AND2    gate15202  (.A(g94), .B(g24533), .Z(g26853) ) ;
AND2    gate15203  (.A(g2868), .B(g24534), .Z(g26854) ) ;
AND2    gate15204  (.A(g2960), .B(g24535), .Z(g26855) ) ;
NAND2   gate15205  (.A(g21403), .B(g23363), .Z(g25062) ) ;
NAND2   gate15206  (.A(g21344), .B(g23462), .Z(g25049) ) ;
AND2    gate15207  (.A(g25062), .B(g25049), .Z(g26857) ) ;
AND2    gate15208  (.A(g2970), .B(g24540), .Z(g26858) ) ;
NAND2   gate15209  (.A(g21417), .B(g23363), .Z(g25021) ) ;
NAND2   gate15210  (.A(g21353), .B(g23462), .Z(g25003) ) ;
AND2    gate15211  (.A(g25021), .B(g25003), .Z(g26861) ) ;
NAND2   gate15212  (.A(g21301), .B(g23363), .Z(g24974) ) ;
NAND2   gate15213  (.A(g21359), .B(g23462), .Z(g24957) ) ;
AND2    gate15214  (.A(g24974), .B(g24957), .Z(g26863) ) ;
AND2    gate15215  (.A(g2907), .B(g24548), .Z(g26864) ) ;
NAND2   gate15216  (.A(g21331), .B(g23363), .Z(g25038) ) ;
NAND2   gate15217  (.A(g21377), .B(g23462), .Z(g25020) ) ;
AND2    gate15218  (.A(g25038), .B(g25020), .Z(g26871) ) ;
AND4    gate15219  (.A(g23032), .B(g26261), .C(g26424), .D(g25550), .Z(g26977) ) ;
AND4    gate15220  (.A(g23032), .B(g26226), .C(g26424), .D(g25557), .Z(g26994) ) ;
OR2     gate15221  (.A(g1171), .B(g24591), .Z(g26334) ) ;
AND2    gate15222  (.A(g26334), .B(g7917), .Z(g27025) ) ;
OR2     gate15223  (.A(g8407), .B(g24591), .Z(g26342) ) ;
AND2    gate15224  (.A(g26342), .B(g1157), .Z(g27028) ) ;
OR2     gate15225  (.A(g8462), .B(g24591), .Z(g26327) ) ;
AND2    gate15226  (.A(g26327), .B(g11031), .Z(g27029) ) ;
OR2     gate15227  (.A(g1514), .B(g24609), .Z(g26343) ) ;
AND2    gate15228  (.A(g26343), .B(g7947), .Z(g27030) ) ;
AND4    gate15229  (.A(g7704), .B(g5180), .C(g5188), .D(g26200), .Z(g27032) ) ;
OR2     gate15230  (.A(g25207), .B(g12015), .Z(g25767) ) ;
AND2    gate15231  (.A(g25767), .B(g19273), .Z(g27033) ) ;
OR2     gate15232  (.A(g1183), .B(g24591), .Z(g26328) ) ;
AND2    gate15233  (.A(g26328), .B(g8609), .Z(g27034) ) ;
OR2     gate15234  (.A(g8466), .B(g24609), .Z(g26348) ) ;
AND2    gate15235  (.A(g26348), .B(g1500), .Z(g27035) ) ;
OR2     gate15236  (.A(g8526), .B(g24609), .Z(g26329) ) ;
AND2    gate15237  (.A(g26329), .B(g11038), .Z(g27036) ) ;
AND4    gate15238  (.A(g7738), .B(g5527), .C(g5535), .D(g26223), .Z(g27039) ) ;
AND4    gate15239  (.A(g7812), .B(g6565), .C(g6573), .D(g26226), .Z(g27040) ) ;
AND2    gate15240  (.A(g8519), .B(g26330), .Z(g27041) ) ;
OR2     gate15241  (.A(g25223), .B(g12043), .Z(g25774) ) ;
AND2    gate15242  (.A(g25774), .B(g19343), .Z(g27042) ) ;
OR2     gate15243  (.A(g1526), .B(g24609), .Z(g26335) ) ;
AND2    gate15244  (.A(g26335), .B(g8632), .Z(g27043) ) ;
AND4    gate15245  (.A(g7766), .B(g5873), .C(g5881), .D(g26241), .Z(g27044) ) ;
AND4    gate15246  (.A(g10295), .B(g3171), .C(g3179), .D(g26244), .Z(g27045) ) ;
OR2     gate15247  (.A(g25285), .B(g14543), .Z(g25789) ) ;
AND2    gate15248  (.A(g25789), .B(g22338), .Z(g27050) ) ;
AND4    gate15249  (.A(g7791), .B(g6219), .C(g6227), .D(g26261), .Z(g27057) ) ;
AND4    gate15250  (.A(g10323), .B(g3522), .C(g3530), .D(g26264), .Z(g27058) ) ;
AND4    gate15251  (.A(g7121), .B(g3873), .C(g3881), .D(g26281), .Z(g27073) ) ;
OR2     gate15252  (.A(g25323), .B(g23836), .Z(g25819) ) ;
AND2    gate15253  (.A(g25819), .B(g22456), .Z(g27083) ) ;
OR2     gate15254  (.A(g25367), .B(g23855), .Z(g25835) ) ;
AND2    gate15255  (.A(g25835), .B(g22494), .Z(g27085) ) ;
OR2     gate15256  (.A(g25368), .B(g23856), .Z(g25836) ) ;
AND2    gate15257  (.A(g25836), .B(g22495), .Z(g27086) ) ;
NOR2    gate15258  (.A(g8745), .B(g11083), .Z(g13872) ) ;
AND2    gate15259  (.A(g13872), .B(g26284), .Z(g27087) ) ;
AND2    gate15260  (.A(g25997), .B(g16423), .Z(g27090) ) ;
AND2    gate15261  (.A(g25997), .B(g16472), .Z(g27094) ) ;
AND2    gate15262  (.A(g25997), .B(g16473), .Z(g27095) ) ;
AND2    gate15263  (.A(g26026), .B(g16475), .Z(g27096) ) ;
OR2     gate15264  (.A(g25449), .B(g23884), .Z(g25867) ) ;
AND2    gate15265  (.A(g25867), .B(g22526), .Z(g27097) ) ;
OR2     gate15266  (.A(g25450), .B(g23885), .Z(g25868) ) ;
AND2    gate15267  (.A(g25868), .B(g22528), .Z(g27098) ) ;
NOR2    gate15268  (.A(g8770), .B(g11083), .Z(g14094) ) ;
AND2    gate15269  (.A(g14094), .B(g26352), .Z(g27099) ) ;
AND2    gate15270  (.A(g25997), .B(g16509), .Z(g27103) ) ;
AND2    gate15271  (.A(g25997), .B(g16510), .Z(g27104) ) ;
AND2    gate15272  (.A(g26026), .B(g16511), .Z(g27105) ) ;
AND2    gate15273  (.A(g26026), .B(g16512), .Z(g27106) ) ;
AND2    gate15274  (.A(g26055), .B(g16514), .Z(g27107) ) ;
AND2    gate15275  (.A(g25997), .B(g16522), .Z(g27113) ) ;
AND2    gate15276  (.A(g25997), .B(g16523), .Z(g27114) ) ;
AND2    gate15277  (.A(g26026), .B(g16526), .Z(g27115) ) ;
AND2    gate15278  (.A(g26026), .B(g16527), .Z(g27116) ) ;
AND2    gate15279  (.A(g26055), .B(g16528), .Z(g27117) ) ;
AND2    gate15280  (.A(g26055), .B(g16529), .Z(g27118) ) ;
OR2     gate15281  (.A(g25502), .B(g23919), .Z(g25877) ) ;
AND2    gate15282  (.A(g25877), .B(g22542), .Z(g27119) ) ;
OR2     gate15283  (.A(g25503), .B(g23920), .Z(g25878) ) ;
AND2    gate15284  (.A(g25878), .B(g22543), .Z(g27120) ) ;
AND2    gate15285  (.A(g136), .B(g26326), .Z(g27121) ) ;
AND2    gate15286  (.A(g25997), .B(g16582), .Z(g27127) ) ;
AND2    gate15287  (.A(g25997), .B(g16583), .Z(g27128) ) ;
AND2    gate15288  (.A(g26026), .B(g16584), .Z(g27129) ) ;
AND2    gate15289  (.A(g26026), .B(g16585), .Z(g27130) ) ;
AND2    gate15290  (.A(g26055), .B(g16588), .Z(g27131) ) ;
AND2    gate15291  (.A(g26055), .B(g16589), .Z(g27132) ) ;
AND2    gate15292  (.A(g25997), .B(g16602), .Z(g27134) ) ;
AND2    gate15293  (.A(g26026), .B(g16605), .Z(g27136) ) ;
AND2    gate15294  (.A(g26026), .B(g16606), .Z(g27137) ) ;
AND2    gate15295  (.A(g26055), .B(g16607), .Z(g27138) ) ;
AND2    gate15296  (.A(g26055), .B(g16608), .Z(g27139) ) ;
OR2     gate15297  (.A(g25522), .B(g23957), .Z(g25885) ) ;
AND2    gate15298  (.A(g25885), .B(g22593), .Z(g27140) ) ;
NOR2    gate15299  (.A(g8891), .B(g12259), .Z(g14121) ) ;
AND2    gate15300  (.A(g14121), .B(g26382), .Z(g27145) ) ;
AND3    gate15301  (.A(g26148), .B(g8187), .C(g1648), .Z(g27146) ) ;
AND2    gate15302  (.A(g25997), .B(g16622), .Z(g27148) ) ;
AND2    gate15303  (.A(g25997), .B(g16623), .Z(g27149) ) ;
AND2    gate15304  (.A(g26026), .B(g16626), .Z(g27151) ) ;
AND2    gate15305  (.A(g26055), .B(g16629), .Z(g27153) ) ;
AND2    gate15306  (.A(g26055), .B(g16630), .Z(g27154) ) ;
NOR2    gate15307  (.A(g146), .B(g24732), .Z(g26609) ) ;
AND2    gate15308  (.A(g26609), .B(g16645), .Z(g27158) ) ;
NOR2    gate15309  (.A(g8997), .B(g12259), .Z(g14163) ) ;
AND2    gate15310  (.A(g14163), .B(g26340), .Z(g27160) ) ;
AND3    gate15311  (.A(g26166), .B(g8241), .C(g1783), .Z(g27161) ) ;
AND3    gate15312  (.A(g26171), .B(g8259), .C(g2208), .Z(g27162) ) ;
AND2    gate15313  (.A(g25997), .B(g16651), .Z(g27177) ) ;
AND2    gate15314  (.A(g25997), .B(g16652), .Z(g27178) ) ;
AND2    gate15315  (.A(g26026), .B(g16654), .Z(g27180) ) ;
AND2    gate15316  (.A(g26026), .B(g16655), .Z(g27181) ) ;
AND2    gate15317  (.A(g26055), .B(g16658), .Z(g27183) ) ;
NOR2    gate15318  (.A(g8990), .B(g24732), .Z(g26628) ) ;
AND2    gate15319  (.A(g26628), .B(g13756), .Z(g27184) ) ;
AND3    gate15320  (.A(g26190), .B(g8302), .C(g1917), .Z(g27185) ) ;
AND3    gate15321  (.A(g26195), .B(g8316), .C(g2342), .Z(g27186) ) ;
AND2    gate15322  (.A(g25997), .B(g16685), .Z(g27201) ) ;
AND2    gate15323  (.A(g25997), .B(g13876), .Z(g27202) ) ;
AND2    gate15324  (.A(g26026), .B(g16688), .Z(g27203) ) ;
AND2    gate15325  (.A(g26026), .B(g16689), .Z(g27204) ) ;
AND2    gate15326  (.A(g26055), .B(g16691), .Z(g27206) ) ;
AND2    gate15327  (.A(g26055), .B(g16692), .Z(g27207) ) ;
AND2    gate15328  (.A(g9037), .B(g26598), .Z(g27208) ) ;
AND3    gate15329  (.A(g26213), .B(g8365), .C(g2051), .Z(g27209) ) ;
AND3    gate15330  (.A(g26218), .B(g8373), .C(g2476), .Z(g27210) ) ;
AND2    gate15331  (.A(g25997), .B(g16716), .Z(g27211) ) ;
AND2    gate15332  (.A(g25997), .B(g16717), .Z(g27212) ) ;
AND2    gate15333  (.A(g26026), .B(g16721), .Z(g27213) ) ;
AND2    gate15334  (.A(g26026), .B(g13901), .Z(g27214) ) ;
AND2    gate15335  (.A(g26055), .B(g16724), .Z(g27215) ) ;
AND2    gate15336  (.A(g26055), .B(g16725), .Z(g27216) ) ;
AND3    gate15337  (.A(g26236), .B(g8418), .C(g2610), .Z(g27217) ) ;
AND2    gate15338  (.A(g25997), .B(g16740), .Z(g27218) ) ;
AND2    gate15339  (.A(g26026), .B(g16742), .Z(g27219) ) ;
AND2    gate15340  (.A(g26026), .B(g16743), .Z(g27220) ) ;
AND2    gate15341  (.A(g26055), .B(g16747), .Z(g27221) ) ;
AND2    gate15342  (.A(g26055), .B(g13932), .Z(g27222) ) ;
AND2    gate15343  (.A(g26026), .B(g16771), .Z(g27227) ) ;
AND2    gate15344  (.A(g26055), .B(g16773), .Z(g27228) ) ;
AND2    gate15345  (.A(g26055), .B(g16774), .Z(g27229) ) ;
OR2     gate15346  (.A(g25559), .B(g24014), .Z(g25906) ) ;
AND2    gate15347  (.A(g25906), .B(g19558), .Z(g27230) ) ;
AND2    gate15348  (.A(g26055), .B(g16814), .Z(g27234) ) ;
OR2     gate15349  (.A(g25565), .B(g22142), .Z(g25910) ) ;
AND2    gate15350  (.A(g25910), .B(g19579), .Z(g27235) ) ;
OR2     gate15351  (.A(g10776), .B(g24433), .Z(g26690) ) ;
AND2    gate15352  (.A(g26690), .B(g26673), .Z(g27246) ) ;
AND2    gate15353  (.A(g2759), .B(g26745), .Z(g27247) ) ;
OR2     gate15354  (.A(g24395), .B(g22193), .Z(g25929) ) ;
AND2    gate15355  (.A(g25929), .B(g19678), .Z(g27249) ) ;
OR2     gate15356  (.A(g10776), .B(g24444), .Z(g26721) ) ;
AND2    gate15357  (.A(g26721), .B(g26694), .Z(g27251) ) ;
OR2     gate15358  (.A(g10776), .B(g24447), .Z(g26733) ) ;
AND2    gate15359  (.A(g26733), .B(g26703), .Z(g27252) ) ;
OR2     gate15360  (.A(g24402), .B(g22208), .Z(g25935) ) ;
AND2    gate15361  (.A(g25935), .B(g19688), .Z(g27254) ) ;
OR2     gate15362  (.A(g24403), .B(g22209), .Z(g25936) ) ;
AND2    gate15363  (.A(g25936), .B(g19689), .Z(g27255) ) ;
OR2     gate15364  (.A(g24406), .B(g22216), .Z(g25937) ) ;
AND2    gate15365  (.A(g25937), .B(g19698), .Z(g27256) ) ;
OR2     gate15366  (.A(g10776), .B(g24457), .Z(g26755) ) ;
AND2    gate15367  (.A(g26755), .B(g26725), .Z(g27259) ) ;
OR2     gate15368  (.A(g10776), .B(g24460), .Z(g26766) ) ;
AND2    gate15369  (.A(g26766), .B(g26737), .Z(g27260) ) ;
AND2    gate15370  (.A(g25997), .B(g17092), .Z(g27262) ) ;
OR2     gate15371  (.A(g24415), .B(g22218), .Z(g25940) ) ;
AND2    gate15372  (.A(g25940), .B(g19713), .Z(g27263) ) ;
OR2     gate15373  (.A(g24416), .B(g22219), .Z(g25941) ) ;
AND2    gate15374  (.A(g25941), .B(g19714), .Z(g27264) ) ;
OR2     gate15375  (.A(g10776), .B(g24468), .Z(g26785) ) ;
AND2    gate15376  (.A(g26785), .B(g26759), .Z(g27265) ) ;
OR2     gate15377  (.A(g10776), .B(g24471), .Z(g26789) ) ;
AND2    gate15378  (.A(g26789), .B(g26770), .Z(g27266) ) ;
AND2    gate15379  (.A(g26026), .B(g17124), .Z(g27267) ) ;
OR2     gate15380  (.A(g24422), .B(g22298), .Z(g25942) ) ;
AND2    gate15381  (.A(g25942), .B(g19733), .Z(g27268) ) ;
OR2     gate15382  (.A(g24423), .B(g22299), .Z(g25943) ) ;
AND2    gate15383  (.A(g25943), .B(g19734), .Z(g27269) ) ;
OR2     gate15384  (.A(g10776), .B(g24478), .Z(g26805) ) ;
AND2    gate15385  (.A(g26805), .B(g26793), .Z(g27270) ) ;
AND2    gate15386  (.A(g26055), .B(g17144), .Z(g27272) ) ;
OR2     gate15387  (.A(g24427), .B(g22307), .Z(g25945) ) ;
AND2    gate15388  (.A(g25945), .B(g19745), .Z(g27275) ) ;
NAND2   gate15389  (.A(II13335), .B(II13336), .Z(g9750) ) ;
AND2    gate15390  (.A(g9750), .B(g26607), .Z(g27276) ) ;
OR2     gate15391  (.A(g24651), .B(g22939), .Z(g26359) ) ;
NAND2   gate15392  (.A(II13391), .B(II13392), .Z(g9825) ) ;
AND2    gate15393  (.A(g9825), .B(g26614), .Z(g27280) ) ;
NAND2   gate15394  (.A(II13402), .B(II13403), .Z(g9830) ) ;
AND2    gate15395  (.A(g9830), .B(g26615), .Z(g27281) ) ;
NAND2   gate15396  (.A(II13453), .B(II13454), .Z(g9908) ) ;
AND2    gate15397  (.A(g9908), .B(g26631), .Z(g27284) ) ;
NAND2   gate15398  (.A(II13463), .B(II13464), .Z(g9912) ) ;
AND2    gate15399  (.A(g9912), .B(g26632), .Z(g27285) ) ;
AND2    gate15400  (.A(g6856), .B(g26634), .Z(g27286) ) ;
NOR2    gate15401  (.A(g24881), .B(g24855), .Z(g26545) ) ;
AND2    gate15402  (.A(g26545), .B(g23011), .Z(g27287) ) ;
NOR2    gate15403  (.A(g24843), .B(g24822), .Z(g26515) ) ;
AND2    gate15404  (.A(g26515), .B(g23013), .Z(g27288) ) ;
NAND2   gate15405  (.A(g7252), .B(g1636), .Z(g11969) ) ;
AND2    gate15406  (.A(g11969), .B(g26653), .Z(g27291) ) ;
AND2    gate15407  (.A(g1714), .B(g26654), .Z(g27292) ) ;
NAND2   gate15408  (.A(II13510), .B(II13511), .Z(g9972) ) ;
AND2    gate15409  (.A(g9972), .B(g26655), .Z(g27293) ) ;
NAND2   gate15410  (.A(II13519), .B(II13520), .Z(g9975) ) ;
AND2    gate15411  (.A(g9975), .B(g26656), .Z(g27294) ) ;
NOR2    gate15412  (.A(g24897), .B(g24884), .Z(g26573) ) ;
AND2    gate15413  (.A(g26573), .B(g23026), .Z(g27298) ) ;
NOR2    gate15414  (.A(g24858), .B(g24846), .Z(g26546) ) ;
AND2    gate15415  (.A(g26546), .B(g23028), .Z(g27299) ) ;
NAND2   gate15416  (.A(II15213), .B(II15214), .Z(g12370) ) ;
AND2    gate15417  (.A(g12370), .B(g26672), .Z(g27300) ) ;
NAND2   gate15418  (.A(g7275), .B(g1772), .Z(g11992) ) ;
AND2    gate15419  (.A(g11992), .B(g26679), .Z(g27301) ) ;
AND2    gate15420  (.A(g1848), .B(g26680), .Z(g27302) ) ;
NAND2   gate15421  (.A(g7280), .B(g2197), .Z(g11996) ) ;
AND2    gate15422  (.A(g11996), .B(g26681), .Z(g27303) ) ;
AND2    gate15423  (.A(g2273), .B(g26682), .Z(g27304) ) ;
NAND2   gate15424  (.A(II13565), .B(II13566), .Z(g10041) ) ;
AND2    gate15425  (.A(g10041), .B(g26683), .Z(g27305) ) ;
NOR2    gate15426  (.A(g24908), .B(g24900), .Z(g26603) ) ;
AND2    gate15427  (.A(g26603), .B(g23057), .Z(g27309) ) ;
NOR2    gate15428  (.A(g24887), .B(g24861), .Z(g26574) ) ;
AND2    gate15429  (.A(g26574), .B(g23059), .Z(g27310) ) ;
NAND2   gate15430  (.A(II15254), .B(II15255), .Z(g12431) ) ;
AND2    gate15431  (.A(g12431), .B(g26693), .Z(g27311) ) ;
NAND2   gate15432  (.A(g7322), .B(g1906), .Z(g12019) ) ;
AND2    gate15433  (.A(g12019), .B(g26700), .Z(g27312) ) ;
AND2    gate15434  (.A(g1982), .B(g26701), .Z(g27313) ) ;
NAND2   gate15435  (.A(II15263), .B(II15264), .Z(g12436) ) ;
AND2    gate15436  (.A(g12436), .B(g26702), .Z(g27314) ) ;
NAND2   gate15437  (.A(g7335), .B(g2331), .Z(g12022) ) ;
AND2    gate15438  (.A(g12022), .B(g26709), .Z(g27315) ) ;
AND2    gate15439  (.A(g2407), .B(g26710), .Z(g27316) ) ;
NOR2    gate15440  (.A(g283), .B(g24825), .Z(g26268) ) ;
AND2    gate15441  (.A(g26268), .B(g23086), .Z(g27323) ) ;
AND2    gate15442  (.A(g10150), .B(g26720), .Z(g27324) ) ;
NAND2   gate15443  (.A(II15299), .B(II15300), .Z(g12478) ) ;
AND2    gate15444  (.A(g12478), .B(g26724), .Z(g27325) ) ;
NAND2   gate15445  (.A(g7369), .B(g2040), .Z(g12048) ) ;
AND2    gate15446  (.A(g12048), .B(g26731), .Z(g27326) ) ;
AND2    gate15447  (.A(g2116), .B(g26732), .Z(g27327) ) ;
NAND2   gate15448  (.A(II15307), .B(II15308), .Z(g12482) ) ;
AND2    gate15449  (.A(g12482), .B(g26736), .Z(g27328) ) ;
NAND2   gate15450  (.A(g7387), .B(g2465), .Z(g12052) ) ;
AND2    gate15451  (.A(g12052), .B(g26743), .Z(g27329) ) ;
AND2    gate15452  (.A(g2541), .B(g26744), .Z(g27330) ) ;
AND2    gate15453  (.A(g10177), .B(g26754), .Z(g27331) ) ;
NAND2   gate15454  (.A(II15334), .B(II15335), .Z(g12538) ) ;
AND2    gate15455  (.A(g12538), .B(g26758), .Z(g27332) ) ;
AND2    gate15456  (.A(g10180), .B(g26765), .Z(g27333) ) ;
NAND2   gate15457  (.A(II15341), .B(II15342), .Z(g12539) ) ;
AND2    gate15458  (.A(g12539), .B(g26769), .Z(g27334) ) ;
NAND2   gate15459  (.A(g7431), .B(g2599), .Z(g12087) ) ;
AND2    gate15460  (.A(g12087), .B(g26776), .Z(g27335) ) ;
AND2    gate15461  (.A(g2675), .B(g26777), .Z(g27336) ) ;
AND2    gate15462  (.A(g26400), .B(g17308), .Z(g27339) ) ;
AND2    gate15463  (.A(g10199), .B(g26784), .Z(g27340) ) ;
AND2    gate15464  (.A(g10203), .B(g26788), .Z(g27341) ) ;
NAND2   gate15465  (.A(II15364), .B(II15365), .Z(g12592) ) ;
AND2    gate15466  (.A(g12592), .B(g26792), .Z(g27342) ) ;
AND2    gate15467  (.A(g26400), .B(g17389), .Z(g27346) ) ;
AND2    gate15468  (.A(g26400), .B(g17390), .Z(g27347) ) ;
AND2    gate15469  (.A(g26488), .B(g17392), .Z(g27348) ) ;
AND2    gate15470  (.A(g10217), .B(g26803), .Z(g27350) ) ;
AND2    gate15471  (.A(g10218), .B(g26804), .Z(g27351) ) ;
AND2    gate15472  (.A(g26400), .B(g17414), .Z(g27357) ) ;
AND2    gate15473  (.A(g26400), .B(g17415), .Z(g27358) ) ;
AND2    gate15474  (.A(g26488), .B(g17416), .Z(g27359) ) ;
AND2    gate15475  (.A(g26488), .B(g17417), .Z(g27360) ) ;
AND2    gate15476  (.A(g26519), .B(g17419), .Z(g27361) ) ;
OR2     gate15477  (.A(g19393), .B(g24502), .Z(g26080) ) ;
AND2    gate15478  (.A(g26080), .B(g20036), .Z(g27362) ) ;
AND2    gate15479  (.A(g10231), .B(g26812), .Z(g27363) ) ;
OR2     gate15480  (.A(g24817), .B(g23229), .Z(g25894) ) ;
AND2    gate15481  (.A(g25894), .B(g25324), .Z(g27369) ) ;
AND2    gate15482  (.A(g26400), .B(g17472), .Z(g27370) ) ;
AND2    gate15483  (.A(g26400), .B(g17473), .Z(g27371) ) ;
AND2    gate15484  (.A(g26488), .B(g17476), .Z(g27372) ) ;
AND2    gate15485  (.A(g26488), .B(g17477), .Z(g27373) ) ;
AND2    gate15486  (.A(g26519), .B(g17478), .Z(g27374) ) ;
AND2    gate15487  (.A(g26519), .B(g17479), .Z(g27375) ) ;
AND2    gate15488  (.A(g26549), .B(g17481), .Z(g27376) ) ;
OR2     gate15489  (.A(g24501), .B(g22534), .Z(g26089) ) ;
AND2    gate15490  (.A(g26089), .B(g20052), .Z(g27378) ) ;
AND2    gate15491  (.A(g26400), .B(g17496), .Z(g27384) ) ;
AND2    gate15492  (.A(g26400), .B(g17497), .Z(g27385) ) ;
AND2    gate15493  (.A(g26488), .B(g17498), .Z(g27386) ) ;
AND2    gate15494  (.A(g26488), .B(g17499), .Z(g27387) ) ;
AND2    gate15495  (.A(g26519), .B(g17502), .Z(g27388) ) ;
AND2    gate15496  (.A(g26519), .B(g17503), .Z(g27389) ) ;
AND2    gate15497  (.A(g26549), .B(g17504), .Z(g27390) ) ;
AND2    gate15498  (.A(g26549), .B(g17505), .Z(g27391) ) ;
AND2    gate15499  (.A(g26576), .B(g17507), .Z(g27392) ) ;
OR2     gate15500  (.A(g24506), .B(g22538), .Z(g26099) ) ;
AND2    gate15501  (.A(g26099), .B(g20066), .Z(g27393) ) ;
NOR2    gate15502  (.A(g24808), .B(g24802), .Z(g26314) ) ;
AND4    gate15503  (.A(g8046), .B(g26314), .C(g9187), .D(g9077), .Z(g27395) ) ;
AND2    gate15504  (.A(g26400), .B(g17518), .Z(g27404) ) ;
AND2    gate15505  (.A(g26488), .B(g17521), .Z(g27406) ) ;
AND2    gate15506  (.A(g26488), .B(g17522), .Z(g27407) ) ;
AND2    gate15507  (.A(g26519), .B(g17523), .Z(g27408) ) ;
AND2    gate15508  (.A(g26519), .B(g17524), .Z(g27409) ) ;
AND2    gate15509  (.A(g26549), .B(g17527), .Z(g27410) ) ;
AND2    gate15510  (.A(g26549), .B(g17528), .Z(g27411) ) ;
AND2    gate15511  (.A(g26576), .B(g17529), .Z(g27412) ) ;
AND2    gate15512  (.A(g26576), .B(g17530), .Z(g27413) ) ;
AND4    gate15513  (.A(g8046), .B(g26314), .C(g9187), .D(g504), .Z(g27416) ) ;
AND4    gate15514  (.A(g8038), .B(g26314), .C(g9187), .D(g9077), .Z(g27421) ) ;
AND2    gate15515  (.A(g26400), .B(g17575), .Z(g27427) ) ;
AND2    gate15516  (.A(g26400), .B(g17576), .Z(g27428) ) ;
AND2    gate15517  (.A(g26488), .B(g17579), .Z(g27430) ) ;
AND2    gate15518  (.A(g26519), .B(g17582), .Z(g27432) ) ;
AND2    gate15519  (.A(g26519), .B(g17583), .Z(g27433) ) ;
AND2    gate15520  (.A(g26549), .B(g17584), .Z(g27434) ) ;
AND2    gate15521  (.A(g26549), .B(g17585), .Z(g27435) ) ;
AND2    gate15522  (.A(g26576), .B(g17588), .Z(g27436) ) ;
AND2    gate15523  (.A(g26576), .B(g17589), .Z(g27437) ) ;
AND2    gate15524  (.A(g232), .B(g26831), .Z(g27439) ) ;
AND4    gate15525  (.A(g8046), .B(g26314), .C(g518), .D(g504), .Z(g27440) ) ;
AND4    gate15526  (.A(g8038), .B(g26314), .C(g9187), .D(g504), .Z(g27445) ) ;
AND2    gate15527  (.A(g26400), .B(g17599), .Z(g27451) ) ;
AND2    gate15528  (.A(g26400), .B(g17600), .Z(g27452) ) ;
AND2    gate15529  (.A(g26488), .B(g17602), .Z(g27454) ) ;
AND2    gate15530  (.A(g26488), .B(g17603), .Z(g27455) ) ;
AND2    gate15531  (.A(g26519), .B(g17606), .Z(g27457) ) ;
AND2    gate15532  (.A(g26549), .B(g17609), .Z(g27459) ) ;
AND2    gate15533  (.A(g26549), .B(g17610), .Z(g27460) ) ;
AND2    gate15534  (.A(g26576), .B(g17611), .Z(g27461) ) ;
AND2    gate15535  (.A(g26576), .B(g17612), .Z(g27462) ) ;
AND2    gate15536  (.A(g269), .B(g26832), .Z(g27467) ) ;
AND4    gate15537  (.A(g8046), .B(g26314), .C(g518), .D(g9077), .Z(g27469) ) ;
AND4    gate15538  (.A(g8038), .B(g26314), .C(g518), .D(g504), .Z(g27474) ) ;
AND2    gate15539  (.A(g26400), .B(g17638), .Z(g27480) ) ;
AND2    gate15540  (.A(g26400), .B(g14630), .Z(g27481) ) ;
AND2    gate15541  (.A(g26488), .B(g17641), .Z(g27482) ) ;
AND2    gate15542  (.A(g26488), .B(g17642), .Z(g27483) ) ;
AND2    gate15543  (.A(g26519), .B(g17644), .Z(g27485) ) ;
AND2    gate15544  (.A(g26519), .B(g17645), .Z(g27486) ) ;
AND2    gate15545  (.A(g26549), .B(g17648), .Z(g27488) ) ;
AND2    gate15546  (.A(g26576), .B(g17651), .Z(g27490) ) ;
AND2    gate15547  (.A(g26576), .B(g17652), .Z(g27491) ) ;
AND2    gate15548  (.A(g246), .B(g26837), .Z(g27493) ) ;
AND4    gate15549  (.A(g8038), .B(g26314), .C(g518), .D(g9077), .Z(g27494) ) ;
AND2    gate15550  (.A(g26400), .B(g17672), .Z(g27500) ) ;
AND2    gate15551  (.A(g26400), .B(g17673), .Z(g27501) ) ;
AND2    gate15552  (.A(g26488), .B(g17677), .Z(g27502) ) ;
AND2    gate15553  (.A(g26488), .B(g14668), .Z(g27503) ) ;
AND2    gate15554  (.A(g26519), .B(g17680), .Z(g27504) ) ;
AND2    gate15555  (.A(g26519), .B(g17681), .Z(g27505) ) ;
AND2    gate15556  (.A(g26549), .B(g17683), .Z(g27507) ) ;
AND2    gate15557  (.A(g26549), .B(g17684), .Z(g27508) ) ;
AND2    gate15558  (.A(g26576), .B(g17687), .Z(g27510) ) ;
AND2    gate15559  (.A(g26400), .B(g17707), .Z(g27517) ) ;
AND2    gate15560  (.A(g26488), .B(g17709), .Z(g27518) ) ;
AND2    gate15561  (.A(g26488), .B(g17710), .Z(g27519) ) ;
AND2    gate15562  (.A(g26519), .B(g17714), .Z(g27520) ) ;
AND2    gate15563  (.A(g26519), .B(g14700), .Z(g27521) ) ;
AND2    gate15564  (.A(g26549), .B(g17717), .Z(g27522) ) ;
AND2    gate15565  (.A(g26549), .B(g17718), .Z(g27523) ) ;
AND2    gate15566  (.A(g26576), .B(g17720), .Z(g27525) ) ;
AND2    gate15567  (.A(g26576), .B(g17721), .Z(g27526) ) ;
AND2    gate15568  (.A(g26488), .B(g17735), .Z(g27534) ) ;
AND2    gate15569  (.A(g26519), .B(g17737), .Z(g27535) ) ;
AND2    gate15570  (.A(g26519), .B(g17738), .Z(g27536) ) ;
AND2    gate15571  (.A(g26549), .B(g17742), .Z(g27537) ) ;
AND2    gate15572  (.A(g26549), .B(g14744), .Z(g27538) ) ;
AND2    gate15573  (.A(g26576), .B(g17745), .Z(g27539) ) ;
AND2    gate15574  (.A(g26576), .B(g17746), .Z(g27540) ) ;
OR2     gate15575  (.A(g24545), .B(g24549), .Z(g26278) ) ;
AND2    gate15576  (.A(g26278), .B(g23334), .Z(g27541) ) ;
AND2    gate15577  (.A(g26519), .B(g17756), .Z(g27545) ) ;
AND2    gate15578  (.A(g26549), .B(g17758), .Z(g27546) ) ;
AND2    gate15579  (.A(g26549), .B(g17759), .Z(g27547) ) ;
AND2    gate15580  (.A(g26576), .B(g17763), .Z(g27548) ) ;
AND2    gate15581  (.A(g26576), .B(g14785), .Z(g27549) ) ;
OR2     gate15582  (.A(g24550), .B(g24555), .Z(g26293) ) ;
AND2    gate15583  (.A(g26293), .B(g23353), .Z(g27553) ) ;
AND2    gate15584  (.A(g26549), .B(g17774), .Z(g27557) ) ;
AND2    gate15585  (.A(g26576), .B(g17776), .Z(g27558) ) ;
AND2    gate15586  (.A(g26576), .B(g17777), .Z(g27559) ) ;
OR2     gate15587  (.A(g24551), .B(g22665), .Z(g26299) ) ;
AND2    gate15588  (.A(g26299), .B(g20191), .Z(g27560) ) ;
OR2     gate15589  (.A(g24556), .B(g24564), .Z(g26305) ) ;
AND2    gate15590  (.A(g26305), .B(g23378), .Z(g27564) ) ;
AND2    gate15591  (.A(g26576), .B(g17791), .Z(g27568) ) ;
AND2    gate15592  (.A(g26690), .B(g26673), .Z(g27588) ) ;
AND2    gate15593  (.A(g26721), .B(g26694), .Z(g27594) ) ;
AND2    gate15594  (.A(g26733), .B(g26703), .Z(g27595) ) ;
AND2    gate15595  (.A(g25899), .B(g10475), .Z(g27598) ) ;
AND2    gate15596  (.A(g26755), .B(g26725), .Z(g27600) ) ;
AND2    gate15597  (.A(g26766), .B(g26737), .Z(g27601) ) ;
AND4    gate15598  (.A(g23032), .B(g26244), .C(g26424), .D(g24966), .Z(g27602) ) ;
NOR2    gate15599  (.A(g24984), .B(g11706), .Z(g25887) ) ;
AND2    gate15600  (.A(g25887), .B(g8844), .Z(g27612) ) ;
AND2    gate15601  (.A(g26785), .B(g26759), .Z(g27614) ) ;
AND2    gate15602  (.A(g26789), .B(g26770), .Z(g27615) ) ;
OR2     gate15603  (.A(g24630), .B(g13409), .Z(g26349) ) ;
AND2    gate15604  (.A(g26349), .B(g20449), .Z(g27616) ) ;
AND4    gate15605  (.A(g23032), .B(g26264), .C(g26424), .D(g24982), .Z(g27617) ) ;
NAND3   gate15606  (.A(g12440), .B(g9920), .C(g9843), .Z(g13266) ) ;
AND2    gate15607  (.A(g13266), .B(g25790), .Z(g27627) ) ;
AND2    gate15608  (.A(g26400), .B(g18061), .Z(g27628) ) ;
NOR2    gate15609  (.A(g7443), .B(g10741), .Z(g13076) ) ;
AND2    gate15610  (.A(g13076), .B(g25766), .Z(g27633) ) ;
AND2    gate15611  (.A(g26805), .B(g26793), .Z(g27634) ) ;
AND4    gate15612  (.A(g23032), .B(g26281), .C(g26424), .D(g24996), .Z(g27635) ) ;
AND2    gate15613  (.A(g26488), .B(g15344), .Z(g27645) ) ;
NOR2    gate15614  (.A(g7487), .B(g10762), .Z(g13094) ) ;
AND2    gate15615  (.A(g13094), .B(g25773), .Z(g27646) ) ;
AND2    gate15616  (.A(g25882), .B(g8974), .Z(g27648) ) ;
NAND3   gate15617  (.A(g9985), .B(g9920), .C(g9843), .Z(g10820) ) ;
AND2    gate15618  (.A(g10820), .B(g25820), .Z(g27649) ) ;
AND2    gate15619  (.A(g26519), .B(g15479), .Z(g27650) ) ;
NOR2    gate15620  (.A(g1018), .B(g19699), .Z(g22448) ) ;
AND2    gate15621  (.A(g22448), .B(g25781), .Z(g27651) ) ;
AND2    gate15622  (.A(g26549), .B(g15562), .Z(g27653) ) ;
NOR2    gate15623  (.A(g1361), .B(g19720), .Z(g22491) ) ;
AND2    gate15624  (.A(g22491), .B(g25786), .Z(g27658) ) ;
AND2    gate15625  (.A(g26576), .B(g15568), .Z(g27661) ) ;
AND2    gate15626  (.A(g1024), .B(g25911), .Z(g27664) ) ;
NOR2    gate15627  (.A(g25411), .B(g25371), .Z(g26872) ) ;
AND2    gate15628  (.A(g26872), .B(g23519), .Z(g27665) ) ;
NOR2    gate15629  (.A(g25328), .B(g25290), .Z(g26865) ) ;
AND2    gate15630  (.A(g26865), .B(g23521), .Z(g27666) ) ;
OR2     gate15631  (.A(g24674), .B(g22991), .Z(g26361) ) ;
AND2    gate15632  (.A(g26361), .B(g20601), .Z(g27667) ) ;
AND2    gate15633  (.A(g1367), .B(g25917), .Z(g27668) ) ;
AND2    gate15634  (.A(g26840), .B(g13278), .Z(g27669) ) ;
NOR2    gate15635  (.A(g25453), .B(g25414), .Z(g25769) ) ;
AND2    gate15636  (.A(g25769), .B(g23541), .Z(g27673) ) ;
NOR2    gate15637  (.A(g25374), .B(g25331), .Z(g26873) ) ;
AND2    gate15638  (.A(g26873), .B(g23543), .Z(g27674) ) ;
OR2     gate15639  (.A(g24700), .B(g23007), .Z(g26377) ) ;
AND2    gate15640  (.A(g26377), .B(g20627), .Z(g27676) ) ;
NOR2    gate15641  (.A(g7544), .B(g10741), .Z(g13021) ) ;
AND2    gate15642  (.A(g13021), .B(g25888), .Z(g27677) ) ;
AND2    gate15643  (.A(g947), .B(g25830), .Z(g27678) ) ;
NOR2    gate15644  (.A(g25482), .B(g25456), .Z(g25777) ) ;
AND2    gate15645  (.A(g25777), .B(g23565), .Z(g27682) ) ;
NOR2    gate15646  (.A(g25417), .B(g25377), .Z(g25770) ) ;
AND2    gate15647  (.A(g25770), .B(g23567), .Z(g27683) ) ;
OR2     gate15648  (.A(g24719), .B(g23023), .Z(g26386) ) ;
AND2    gate15649  (.A(g26386), .B(g20657), .Z(g27684) ) ;
NOR2    gate15650  (.A(g7577), .B(g10762), .Z(g13032) ) ;
AND2    gate15651  (.A(g13032), .B(g25895), .Z(g27685) ) ;
AND2    gate15652  (.A(g1291), .B(g25849), .Z(g27686) ) ;
NOR2    gate15653  (.A(g25507), .B(g25485), .Z(g25784) ) ;
AND2    gate15654  (.A(g25784), .B(g23607), .Z(g27690) ) ;
NOR2    gate15655  (.A(g25459), .B(g25420), .Z(g25778) ) ;
AND2    gate15656  (.A(g25778), .B(g23609), .Z(g27691) ) ;
OR2     gate15657  (.A(g24745), .B(g23050), .Z(g26392) ) ;
AND2    gate15658  (.A(g26392), .B(g20697), .Z(g27692) ) ;
NOR2    gate15659  (.A(g25518), .B(g25510), .Z(g25800) ) ;
AND2    gate15660  (.A(g25800), .B(g23647), .Z(g27696) ) ;
NOR2    gate15661  (.A(g25488), .B(g25462), .Z(g25785) ) ;
AND2    gate15662  (.A(g25785), .B(g23649), .Z(g27697) ) ;
OR2     gate15663  (.A(g24762), .B(g23062), .Z(g26396) ) ;
AND2    gate15664  (.A(g26396), .B(g20766), .Z(g27699) ) ;
OR2     gate15665  (.A(g24774), .B(g23104), .Z(g26422) ) ;
AND2    gate15666  (.A(g26422), .B(g20904), .Z(g27710) ) ;
OR2     gate15667  (.A(g24786), .B(g23130), .Z(g26512) ) ;
AND2    gate15668  (.A(g26512), .B(g21049), .Z(g27723) ) ;
AND2    gate15669  (.A(g4146), .B(g25886), .Z(g27765) ) ;
AND2    gate15670  (.A(g7670), .B(g25932), .Z(g27820) ) ;
AND2    gate15671  (.A(g7680), .B(g25892), .Z(g27821) ) ;
AND2    gate15672  (.A(g4157), .B(g25893), .Z(g27822) ) ;
NOR2    gate15673  (.A(g7716), .B(g24591), .Z(g25944) ) ;
AND2    gate15674  (.A(g25944), .B(g19369), .Z(g27932) ) ;
NOR2    gate15675  (.A(g1199), .B(g24591), .Z(g25947) ) ;
AND2    gate15676  (.A(g25947), .B(g15995), .Z(g27957) ) ;
NOR2    gate15677  (.A(g1070), .B(g24591), .Z(g25950) ) ;
AND2    gate15678  (.A(g25950), .B(g22449), .Z(g27958) ) ;
NOR2    gate15679  (.A(g7752), .B(g24609), .Z(g25948) ) ;
AND2    gate15680  (.A(g25948), .B(g19374), .Z(g27959) ) ;
NOR2    gate15681  (.A(g7750), .B(g24591), .Z(g25954) ) ;
AND2    gate15682  (.A(g25954), .B(g19597), .Z(g27962) ) ;
NOR2    gate15683  (.A(g1542), .B(g24609), .Z(g25952) ) ;
AND2    gate15684  (.A(g25952), .B(g16047), .Z(g27963) ) ;
NOR2    gate15685  (.A(g1413), .B(g24609), .Z(g25956) ) ;
AND2    gate15686  (.A(g25956), .B(g22492), .Z(g27964) ) ;
OR2     gate15687  (.A(g25366), .B(g23854), .Z(g25834) ) ;
NOR2    gate15688  (.A(g7779), .B(g24609), .Z(g25958) ) ;
AND2    gate15689  (.A(g25958), .B(g19614), .Z(g27968) ) ;
OR2     gate15690  (.A(g24903), .B(g24912), .Z(g26751) ) ;
AND2    gate15691  (.A(g26751), .B(g23924), .Z(g27981) ) ;
OR2     gate15692  (.A(g24913), .B(g24921), .Z(g26781) ) ;
AND2    gate15693  (.A(g26781), .B(g23941), .Z(g27988) ) ;
OR2     gate15694  (.A(g24922), .B(g24929), .Z(g26800) ) ;
AND2    gate15695  (.A(g26800), .B(g23964), .Z(g27992) ) ;
OR2     gate15696  (.A(g24930), .B(g24939), .Z(g26809) ) ;
AND2    gate15697  (.A(g26809), .B(g23985), .Z(g27995) ) ;
OR2     gate15698  (.A(g24940), .B(g24949), .Z(g26813) ) ;
AND2    gate15699  (.A(g26813), .B(g23995), .Z(g27997) ) ;
AND4    gate15700  (.A(g23032), .B(g26200), .C(g26424), .D(g25529), .Z(g27999) ) ;
AND4    gate15701  (.A(g23032), .B(g26223), .C(g26424), .D(g25535), .Z(g28010) ) ;
AND4    gate15702  (.A(g23032), .B(g26241), .C(g26424), .D(g25542), .Z(g28020) ) ;
AND4    gate15703  (.A(g26365), .B(g24096), .C(g24097), .D(g24098), .Z(II26530) ) ;
AND4    gate15704  (.A(g24099), .B(g24100), .C(g24101), .D(g24102), .Z(II26531) ) ;
AND3    gate15705  (.A(g24103), .B(II26530), .C(II26531), .Z(g28035) ) ;
OR2     gate15706  (.A(g26514), .B(g25050), .Z(g27970) ) ;
AND2    gate15707  (.A(g27970), .B(g18874), .Z(g28107) ) ;
AND2    gate15708  (.A(g7975), .B(g27237), .Z(g28108) ) ;
OR2     gate15709  (.A(g26544), .B(g25063), .Z(g27974) ) ;
AND2    gate15710  (.A(g27974), .B(g18886), .Z(g28110) ) ;
NOR2    gate15711  (.A(g8005), .B(g26616), .Z(g27343) ) ;
AND2    gate15712  (.A(g27343), .B(g22716), .Z(g28111) ) ;
NOR2    gate15713  (.A(g7975), .B(g26616), .Z(g27352) ) ;
AND2    gate15714  (.A(g27352), .B(g26162), .Z(g28112) ) ;
AND2    gate15715  (.A(g8016), .B(g27242), .Z(g28113) ) ;
NOR2    gate15716  (.A(g8064), .B(g26636), .Z(g27354) ) ;
AND2    gate15717  (.A(g27354), .B(g22759), .Z(g28115) ) ;
NOR2    gate15718  (.A(g8016), .B(g26636), .Z(g27366) ) ;
AND2    gate15719  (.A(g27366), .B(g26183), .Z(g28116) ) ;
AND2    gate15720  (.A(g8075), .B(g27245), .Z(g28117) ) ;
NOR2    gate15721  (.A(g8119), .B(g26657), .Z(g27368) ) ;
AND2    gate15722  (.A(g27368), .B(g22842), .Z(g28124) ) ;
NOR2    gate15723  (.A(g8075), .B(g26657), .Z(g27381) ) ;
AND2    gate15724  (.A(g27381), .B(g26209), .Z(g28125) ) ;
NOR2    gate15725  (.A(g8097), .B(g26616), .Z(g27353) ) ;
AND2    gate15726  (.A(g27353), .B(g23063), .Z(g28130) ) ;
NOR2    gate15727  (.A(g8155), .B(g26636), .Z(g27367) ) ;
AND2    gate15728  (.A(g27367), .B(g23108), .Z(g28133) ) ;
NOR2    gate15729  (.A(g8219), .B(g26657), .Z(g27382) ) ;
AND2    gate15730  (.A(g27382), .B(g23135), .Z(g28136) ) ;
NOR2    gate15731  (.A(g8334), .B(g26616), .Z(g27337) ) ;
AND2    gate15732  (.A(g27337), .B(g26054), .Z(g28139) ) ;
AND4    gate15733  (.A(g10831), .B(g11797), .C(g11261), .D(g27163), .Z(g28141) ) ;
NOR2    gate15734  (.A(g8390), .B(g26636), .Z(g27344) ) ;
AND2    gate15735  (.A(g27344), .B(g26083), .Z(g28143) ) ;
NOR2    gate15736  (.A(g8443), .B(g26657), .Z(g27355) ) ;
AND2    gate15737  (.A(g27355), .B(g26093), .Z(g28148) ) ;
AND4    gate15738  (.A(g10862), .B(g11834), .C(g11283), .D(g27187), .Z(g28150) ) ;
AND2    gate15739  (.A(g8426), .B(g27295), .Z(g28151) ) ;
NOR2    gate15740  (.A(g8519), .B(g24825), .Z(g26297) ) ;
AND2    gate15741  (.A(g26297), .B(g27279), .Z(g28152) ) ;
OR4     gate15742  (.A(g26213), .B(g26190), .C(g26166), .D(g26148), .Z(g27031) ) ;
AND2    gate15743  (.A(g8492), .B(g27306), .Z(g28154) ) ;
OR4     gate15744  (.A(g26236), .B(g26218), .C(g26195), .D(g26171), .Z(g27037) ) ;
AND2    gate15745  (.A(g8553), .B(g27317), .Z(g28159) ) ;
NOR2    gate15746  (.A(g8575), .B(g24825), .Z(g26309) ) ;
AND2    gate15747  (.A(g26309), .B(g27463), .Z(g28160) ) ;
AND2    gate15748  (.A(g8651), .B(g27528), .Z(g28164) ) ;
AND2    gate15749  (.A(g27018), .B(g22455), .Z(g28165) ) ;
OR2     gate15750  (.A(g26821), .B(g14585), .Z(g27016) ) ;
AND2    gate15751  (.A(g27016), .B(g19385), .Z(g28171) ) ;
OR2     gate15752  (.A(g26822), .B(g14610), .Z(g27019) ) ;
AND2    gate15753  (.A(g27019), .B(g19397), .Z(g28178) ) ;
AND2    gate15754  (.A(g8770), .B(g27349), .Z(g28182) ) ;
OR2     gate15755  (.A(g26826), .B(g17692), .Z(g27024) ) ;
AND2    gate15756  (.A(g27024), .B(g19421), .Z(g28183) ) ;
OR2     gate15757  (.A(g26828), .B(g17726), .Z(g27026) ) ;
AND2    gate15758  (.A(g27026), .B(g19435), .Z(g28185) ) ;
AND2    gate15759  (.A(g8891), .B(g27415), .Z(g28192) ) ;
AND2    gate15760  (.A(g8851), .B(g27629), .Z(g28193) ) ;
NOR2    gate15761  (.A(g3004), .B(g26616), .Z(g27647) ) ;
AND2    gate15762  (.A(g27647), .B(g11344), .Z(g28197) ) ;
NOR2    gate15763  (.A(g9037), .B(g24732), .Z(g26649) ) ;
AND2    gate15764  (.A(g26649), .B(g27492), .Z(g28198) ) ;
NOR2    gate15765  (.A(g9056), .B(g26616), .Z(g27479) ) ;
AND2    gate15766  (.A(g27479), .B(g16684), .Z(g28199) ) ;
NOR2    gate15767  (.A(g3355), .B(g26636), .Z(g27652) ) ;
AND2    gate15768  (.A(g27652), .B(g11383), .Z(g28200) ) ;
NOR2    gate15769  (.A(g9095), .B(g26636), .Z(g27499) ) ;
AND2    gate15770  (.A(g27499), .B(g16720), .Z(g28201) ) ;
NOR2    gate15771  (.A(g3706), .B(g26657), .Z(g27659) ) ;
AND2    gate15772  (.A(g27659), .B(g11413), .Z(g28202) ) ;
NOR2    gate15773  (.A(g9073), .B(g24732), .Z(g26098) ) ;
AND2    gate15774  (.A(g26098), .B(g27654), .Z(g28204) ) ;
NOR2    gate15775  (.A(g9180), .B(g26657), .Z(g27516) ) ;
AND2    gate15776  (.A(g27516), .B(g16746), .Z(g28205) ) ;
AND2    gate15777  (.A(g9229), .B(g27554), .Z(g28210) ) ;
NOR2    gate15778  (.A(g9253), .B(g25791), .Z(g27720) ) ;
AND2    gate15779  (.A(g27720), .B(g23380), .Z(g28213) ) ;
NOR2    gate15780  (.A(g9229), .B(g25791), .Z(g27731) ) ;
AND2    gate15781  (.A(g27731), .B(g26625), .Z(g28214) ) ;
AND2    gate15782  (.A(g9264), .B(g27565), .Z(g28215) ) ;
NOR2    gate15783  (.A(g9305), .B(g25805), .Z(g27733) ) ;
AND2    gate15784  (.A(g27733), .B(g23391), .Z(g28217) ) ;
NOR2    gate15785  (.A(g9264), .B(g25805), .Z(g27768) ) ;
AND2    gate15786  (.A(g27768), .B(g26645), .Z(g28218) ) ;
AND2    gate15787  (.A(g9316), .B(g27573), .Z(g28219) ) ;
NOR2    gate15788  (.A(g9291), .B(g26616), .Z(g27338) ) ;
AND2    gate15789  (.A(g27338), .B(g17194), .Z(g28223) ) ;
NOR2    gate15790  (.A(g9386), .B(g25821), .Z(g27770) ) ;
AND2    gate15791  (.A(g27770), .B(g23400), .Z(g28225) ) ;
NOR2    gate15792  (.A(g9316), .B(g25821), .Z(g27825) ) ;
AND2    gate15793  (.A(g27825), .B(g26667), .Z(g28226) ) ;
AND2    gate15794  (.A(g9397), .B(g27583), .Z(g28227) ) ;
OR2     gate15795  (.A(g24378), .B(g25787), .Z(g27126) ) ;
AND2    gate15796  (.A(g27126), .B(g19636), .Z(g28228) ) ;
NOR2    gate15797  (.A(g9360), .B(g26636), .Z(g27345) ) ;
AND2    gate15798  (.A(g27345), .B(g17213), .Z(g28229) ) ;
NOR2    gate15799  (.A(g9364), .B(g25791), .Z(g27732) ) ;
AND2    gate15800  (.A(g27732), .B(g23586), .Z(g28232) ) ;
NOR2    gate15801  (.A(g9456), .B(g25839), .Z(g27827) ) ;
AND2    gate15802  (.A(g27827), .B(g23411), .Z(g28233) ) ;
NOR2    gate15803  (.A(g9397), .B(g25839), .Z(g27877) ) ;
AND2    gate15804  (.A(g27877), .B(g26686), .Z(g28234) ) ;
AND2    gate15805  (.A(g9467), .B(g27592), .Z(g28235) ) ;
AND2    gate15806  (.A(g8515), .B(g27971), .Z(g28236) ) ;
AND2    gate15807  (.A(g9492), .B(g27597), .Z(g28237) ) ;
OR2     gate15808  (.A(g25788), .B(g24392), .Z(g27133) ) ;
AND2    gate15809  (.A(g27133), .B(g19658), .Z(g28238) ) ;
OR2     gate15810  (.A(g24387), .B(g25803), .Z(g27135) ) ;
AND2    gate15811  (.A(g27135), .B(g19659), .Z(g28239) ) ;
NOR2    gate15812  (.A(g9429), .B(g26657), .Z(g27356) ) ;
AND2    gate15813  (.A(g27356), .B(g17239), .Z(g28240) ) ;
NOR2    gate15814  (.A(g9434), .B(g25805), .Z(g27769) ) ;
AND2    gate15815  (.A(g27769), .B(g23626), .Z(g28242) ) ;
NOR2    gate15816  (.A(g9523), .B(g25856), .Z(g27879) ) ;
AND2    gate15817  (.A(g27879), .B(g23423), .Z(g28243) ) ;
NOR2    gate15818  (.A(g9467), .B(g25856), .Z(g27926) ) ;
AND2    gate15819  (.A(g27926), .B(g26715), .Z(g28244) ) ;
AND2    gate15820  (.A(g11367), .B(g27975), .Z(g28245) ) ;
AND2    gate15821  (.A(g8572), .B(g27976), .Z(g28246) ) ;
OR2     gate15822  (.A(g25802), .B(g24399), .Z(g27147) ) ;
AND2    gate15823  (.A(g27147), .B(g19675), .Z(g28247) ) ;
OR2     gate15824  (.A(g25804), .B(g24400), .Z(g27150) ) ;
AND2    gate15825  (.A(g27150), .B(g19676), .Z(g28248) ) ;
OR2     gate15826  (.A(g24393), .B(g25817), .Z(g27152) ) ;
AND2    gate15827  (.A(g27152), .B(g19677), .Z(g28249) ) ;
NOR2    gate15828  (.A(g9501), .B(g25821), .Z(g27826) ) ;
AND2    gate15829  (.A(g27826), .B(g23662), .Z(g28251) ) ;
OR2     gate15830  (.A(g25814), .B(g12953), .Z(g27159) ) ;
AND2    gate15831  (.A(g27159), .B(g19682), .Z(g28252) ) ;
NAND2   gate15832  (.A(II22845), .B(II22846), .Z(g23719) ) ;
AND2    gate15833  (.A(g23719), .B(g27700), .Z(g28253) ) ;
AND3    gate15834  (.A(g7268), .B(g1668), .C(g27395), .Z(g28254) ) ;
AND2    gate15835  (.A(g8515), .B(g27983), .Z(g28255) ) ;
AND2    gate15836  (.A(g11398), .B(g27984), .Z(g28256) ) ;
OR2     gate15837  (.A(g25816), .B(g24409), .Z(g27179) ) ;
AND2    gate15838  (.A(g27179), .B(g19686), .Z(g28257) ) ;
OR2     gate15839  (.A(g25818), .B(g24410), .Z(g27182) ) ;
AND2    gate15840  (.A(g27182), .B(g19687), .Z(g28258) ) ;
NOR2    gate15841  (.A(g9607), .B(g25791), .Z(g27703) ) ;
AND2    gate15842  (.A(g27703), .B(g26518), .Z(g28260) ) ;
NOR2    gate15843  (.A(g9559), .B(g25839), .Z(g27878) ) ;
AND2    gate15844  (.A(g27878), .B(g23695), .Z(g28261) ) ;
NAND2   gate15845  (.A(II22865), .B(II22866), .Z(g23747) ) ;
AND2    gate15846  (.A(g23747), .B(g27711), .Z(g28263) ) ;
AND3    gate15847  (.A(g7315), .B(g1802), .C(g27416), .Z(g28264) ) ;
AND2    gate15848  (.A(g11367), .B(g27989), .Z(g28265) ) ;
NAND2   gate15849  (.A(II22872), .B(II22873), .Z(g23748) ) ;
AND2    gate15850  (.A(g23748), .B(g27714), .Z(g28266) ) ;
AND3    gate15851  (.A(g7328), .B(g2227), .C(g27421), .Z(g28267) ) ;
AND2    gate15852  (.A(g8572), .B(g27990), .Z(g28268) ) ;
OR2     gate15853  (.A(g25833), .B(g24421), .Z(g27205) ) ;
AND2    gate15854  (.A(g27205), .B(g19712), .Z(g28269) ) ;
NOR2    gate15855  (.A(g9672), .B(g25805), .Z(g27721) ) ;
AND2    gate15856  (.A(g27721), .B(g26548), .Z(g28272) ) ;
NOR2    gate15857  (.A(g9621), .B(g25856), .Z(g27927) ) ;
AND2    gate15858  (.A(g27927), .B(g23729), .Z(g28273) ) ;
NAND2   gate15859  (.A(II22893), .B(II22894), .Z(g23761) ) ;
AND2    gate15860  (.A(g23761), .B(g27724), .Z(g28280) ) ;
AND3    gate15861  (.A(g7362), .B(g1936), .C(g27440), .Z(g28281) ) ;
NAND2   gate15862  (.A(II22900), .B(II22901), .Z(g23762) ) ;
AND2    gate15863  (.A(g23762), .B(g27727), .Z(g28282) ) ;
AND3    gate15864  (.A(g7380), .B(g2361), .C(g27445), .Z(g28283) ) ;
AND2    gate15865  (.A(g11398), .B(g27994), .Z(g28284) ) ;
AND2    gate15866  (.A(g9657), .B(g27717), .Z(g28285) ) ;
NOR2    gate15867  (.A(g9733), .B(g25821), .Z(g27734) ) ;
AND2    gate15868  (.A(g27734), .B(g26575), .Z(g28289) ) ;
NAND2   gate15869  (.A(II22930), .B(II22931), .Z(g23780) ) ;
AND2    gate15870  (.A(g23780), .B(g27759), .Z(g28290) ) ;
AND3    gate15871  (.A(g7411), .B(g2070), .C(g27469), .Z(g28291) ) ;
NAND2   gate15872  (.A(II22937), .B(II22938), .Z(g23781) ) ;
AND2    gate15873  (.A(g23781), .B(g27762), .Z(g28292) ) ;
AND3    gate15874  (.A(g7424), .B(g2495), .C(g27474), .Z(g28293) ) ;
AND2    gate15875  (.A(g9716), .B(g27670), .Z(g28299) ) ;
NOR2    gate15876  (.A(g9809), .B(g25839), .Z(g27771) ) ;
AND2    gate15877  (.A(g27771), .B(g26605), .Z(g28300) ) ;
OR2     gate15878  (.A(g25870), .B(g15678), .Z(g27224) ) ;
AND2    gate15879  (.A(g27224), .B(g19750), .Z(g28301) ) ;
NAND2   gate15880  (.A(II22966), .B(II22967), .Z(g23809) ) ;
AND2    gate15881  (.A(g23809), .B(g27817), .Z(g28302) ) ;
AND3    gate15882  (.A(g7462), .B(g2629), .C(g27494), .Z(g28303) ) ;
OR2     gate15883  (.A(g25872), .B(g24436), .Z(g27226) ) ;
AND2    gate15884  (.A(g27226), .B(g19753), .Z(g28304) ) ;
AND2    gate15885  (.A(g9792), .B(g27679), .Z(g28311) ) ;
NOR2    gate15886  (.A(g9892), .B(g25856), .Z(g27828) ) ;
AND2    gate15887  (.A(g27828), .B(g26608), .Z(g28312) ) ;
OR2     gate15888  (.A(g25873), .B(g15699), .Z(g27231) ) ;
AND2    gate15889  (.A(g27231), .B(g19766), .Z(g28313) ) ;
OR2     gate15890  (.A(g26092), .B(g24676), .Z(g27552) ) ;
OR2     gate15891  (.A(g25874), .B(g24450), .Z(g27232) ) ;
AND2    gate15892  (.A(g27232), .B(g19769), .Z(g28315) ) ;
OR2     gate15893  (.A(g25876), .B(g24451), .Z(g27233) ) ;
AND2    gate15894  (.A(g27233), .B(g19770), .Z(g28318) ) ;
AND2    gate15895  (.A(g9875), .B(g27687), .Z(g28324) ) ;
NAND2   gate15896  (.A(II26050), .B(II26051), .Z(g27365) ) ;
AND2    gate15897  (.A(g27365), .B(g19785), .Z(g28327) ) ;
OR2     gate15898  (.A(g25879), .B(g24464), .Z(g27238) ) ;
AND2    gate15899  (.A(g27238), .B(g19786), .Z(g28330) ) ;
OR2     gate15900  (.A(g25881), .B(g24465), .Z(g27239) ) ;
AND2    gate15901  (.A(g27239), .B(g19787), .Z(g28333) ) ;
AND2    gate15902  (.A(g9946), .B(g27693), .Z(g28339) ) ;
OR2     gate15903  (.A(g25883), .B(g24467), .Z(g27240) ) ;
AND2    gate15904  (.A(g27240), .B(g19790), .Z(g28341) ) ;
NAND2   gate15905  (.A(II26071), .B(II26072), .Z(g27380) ) ;
AND2    gate15906  (.A(g27380), .B(g19799), .Z(g28343) ) ;
OR2     gate15907  (.A(g25884), .B(g24475), .Z(g27243) ) ;
AND2    gate15908  (.A(g27243), .B(g19800), .Z(g28346) ) ;
AND2    gate15909  (.A(g10014), .B(g27705), .Z(g28352) ) ;
NAND2   gate15910  (.A(II26094), .B(II26095), .Z(g27401) ) ;
AND2    gate15911  (.A(g27401), .B(g19861), .Z(g28360) ) ;
OR2     gate15912  (.A(g25901), .B(g15738), .Z(g27250) ) ;
AND2    gate15913  (.A(g27250), .B(g19963), .Z(g28415) ) ;
OR2     gate15914  (.A(g25904), .B(g24498), .Z(g27257) ) ;
AND2    gate15915  (.A(g27257), .B(g20006), .Z(g28426) ) ;
OR2     gate15916  (.A(g25905), .B(g15749), .Z(g27258) ) ;
AND2    gate15917  (.A(g27258), .B(g20008), .Z(g28427) ) ;
NAND3   gate15918  (.A(g10504), .B(g26131), .C(g26105), .Z(g27273) ) ;
AND2    gate15919  (.A(g27273), .B(g10233), .Z(g28439) ) ;
OR2     gate15920  (.A(g15779), .B(g25915), .Z(g27274) ) ;
AND2    gate15921  (.A(g27274), .B(g20059), .Z(g28440) ) ;
OR2     gate15922  (.A(g15786), .B(g25921), .Z(g27278) ) ;
AND2    gate15923  (.A(g27278), .B(g20072), .Z(g28442) ) ;
OR2     gate15924  (.A(g25922), .B(g25924), .Z(g27283) ) ;
AND2    gate15925  (.A(g27283), .B(g20090), .Z(g28451) ) ;
NAND3   gate15926  (.A(g10857), .B(g26131), .C(g26105), .Z(g27582) ) ;
AND2    gate15927  (.A(g27582), .B(g10233), .Z(g28453) ) ;
NOR2    gate15928  (.A(g5016), .B(g25791), .Z(g26976) ) ;
AND2    gate15929  (.A(g26976), .B(g12233), .Z(g28454) ) ;
OR2     gate15930  (.A(g25925), .B(g25927), .Z(g27289) ) ;
AND2    gate15931  (.A(g27289), .B(g20103), .Z(g28455) ) ;
OR2     gate15932  (.A(g25926), .B(g25928), .Z(g27290) ) ;
AND2    gate15933  (.A(g27290), .B(g20104), .Z(g28456) ) ;
AND3    gate15934  (.A(g24981), .B(g26424), .C(g22698), .Z(II26948) ) ;
AND4    gate15935  (.A(g27187), .B(g12730), .C(g20887), .D(II26948), .Z(g28458) ) ;
NOR2    gate15936  (.A(g7134), .B(g25791), .Z(g27960) ) ;
AND2    gate15937  (.A(g27960), .B(g17637), .Z(g28466) ) ;
NOR2    gate15938  (.A(g5360), .B(g25805), .Z(g26993) ) ;
AND2    gate15939  (.A(g26993), .B(g12295), .Z(g28467) ) ;
AND3    gate15940  (.A(g24995), .B(g26424), .C(g22698), .Z(II26960) ) ;
AND4    gate15941  (.A(g27187), .B(g12762), .C(g21024), .D(II26960), .Z(g28471) ) ;
NOR2    gate15942  (.A(g7153), .B(g25805), .Z(g27966) ) ;
AND2    gate15943  (.A(g27966), .B(g17676), .Z(g28477) ) ;
NOR2    gate15944  (.A(g5706), .B(g25821), .Z(g27007) ) ;
AND2    gate15945  (.A(g27007), .B(g12345), .Z(g28478) ) ;
AND3    gate15946  (.A(g25011), .B(g26424), .C(g22698), .Z(II26972) ) ;
AND4    gate15947  (.A(g27187), .B(g10290), .C(g21163), .D(II26972), .Z(g28484) ) ;
NOR2    gate15948  (.A(g7170), .B(g25821), .Z(g27969) ) ;
AND2    gate15949  (.A(g27969), .B(g17713), .Z(g28488) ) ;
NOR2    gate15950  (.A(g6052), .B(g25839), .Z(g27010) ) ;
AND2    gate15951  (.A(g27010), .B(g12417), .Z(g28489) ) ;
NOR2    gate15952  (.A(g7187), .B(g25839), .Z(g27973) ) ;
AND2    gate15953  (.A(g27973), .B(g17741), .Z(g28494) ) ;
NOR2    gate15954  (.A(g6398), .B(g25856), .Z(g27012) ) ;
AND2    gate15955  (.A(g27012), .B(g12465), .Z(g28495) ) ;
NOR2    gate15956  (.A(g7212), .B(g25856), .Z(g27982) ) ;
AND2    gate15957  (.A(g27982), .B(g17762), .Z(g28499) ) ;
NOR2    gate15958  (.A(g7239), .B(g25791), .Z(g27704) ) ;
AND2    gate15959  (.A(g27704), .B(g15585), .Z(g28523) ) ;
AND2    gate15960  (.A(g6821), .B(g27084), .Z(g28524) ) ;
AND2    gate15961  (.A(g27187), .B(g12730), .Z(g28528) ) ;
OR2     gate15962  (.A(g24569), .B(g25961), .Z(g27383) ) ;
AND2    gate15963  (.A(g27383), .B(g20240), .Z(g28530) ) ;
NOR2    gate15964  (.A(g7247), .B(g25805), .Z(g27722) ) ;
AND2    gate15965  (.A(g27722), .B(g15608), .Z(g28531) ) ;
OR2     gate15966  (.A(g25957), .B(g24573), .Z(g27394) ) ;
AND2    gate15967  (.A(g27394), .B(g20265), .Z(g28532) ) ;
AND2    gate15968  (.A(g11981), .B(g27088), .Z(g28535) ) ;
AND2    gate15969  (.A(g6832), .B(g27089), .Z(g28537) ) ;
AND2    gate15970  (.A(g27187), .B(g12762), .Z(g28539) ) ;
OR2     gate15971  (.A(g25962), .B(g24581), .Z(g27403) ) ;
AND2    gate15972  (.A(g27403), .B(g20274), .Z(g28541) ) ;
OR2     gate15973  (.A(g24572), .B(g25968), .Z(g27405) ) ;
AND2    gate15974  (.A(g27405), .B(g20275), .Z(g28542) ) ;
NOR2    gate15975  (.A(g7262), .B(g25821), .Z(g27735) ) ;
AND2    gate15976  (.A(g27735), .B(g15628), .Z(g28543) ) ;
AND2    gate15977  (.A(g6821), .B(g27091), .Z(g28547) ) ;
AND2    gate15978  (.A(g12009), .B(g27092), .Z(g28550) ) ;
AND2    gate15979  (.A(g27187), .B(g10290), .Z(g28553) ) ;
OR2     gate15980  (.A(g25967), .B(g24588), .Z(g27426) ) ;
AND2    gate15981  (.A(g27426), .B(g20372), .Z(g28554) ) ;
OR2     gate15982  (.A(g25969), .B(g24589), .Z(g27429) ) ;
AND2    gate15983  (.A(g27429), .B(g20373), .Z(g28555) ) ;
OR2     gate15984  (.A(g24582), .B(g25977), .Z(g27431) ) ;
AND2    gate15985  (.A(g27431), .B(g20374), .Z(g28556) ) ;
NOR2    gate15986  (.A(g7297), .B(g25839), .Z(g27772) ) ;
AND2    gate15987  (.A(g27772), .B(g15647), .Z(g28557) ) ;
AND2    gate15988  (.A(g7301), .B(g27046), .Z(g28558) ) ;
AND2    gate15989  (.A(g11981), .B(g27100), .Z(g28563) ) ;
AND2    gate15990  (.A(g6832), .B(g27101), .Z(g28567) ) ;
OR2     gate15991  (.A(g25976), .B(g24606), .Z(g27453) ) ;
AND2    gate15992  (.A(g27453), .B(g20433), .Z(g28569) ) ;
OR2     gate15993  (.A(g25978), .B(g24607), .Z(g27456) ) ;
AND2    gate15994  (.A(g27456), .B(g20434), .Z(g28570) ) ;
OR2     gate15995  (.A(g24590), .B(g25989), .Z(g27458) ) ;
AND2    gate15996  (.A(g27458), .B(g20435), .Z(g28571) ) ;
NOR2    gate15997  (.A(g7345), .B(g25856), .Z(g27829) ) ;
AND2    gate15998  (.A(g27829), .B(g15669), .Z(g28572) ) ;
AND2    gate15999  (.A(g7349), .B(g27059), .Z(g28573) ) ;
AND2    gate16000  (.A(g12009), .B(g27112), .Z(g28583) ) ;
NOR2    gate16001  (.A(g26485), .B(g26516), .Z(g27063) ) ;
AND2    gate16002  (.A(g27063), .B(g10530), .Z(g28585) ) ;
OR2     gate16003  (.A(g25988), .B(g24628), .Z(g27484) ) ;
AND2    gate16004  (.A(g27484), .B(g20497), .Z(g28586) ) ;
OR2     gate16005  (.A(g25990), .B(g24629), .Z(g27487) ) ;
AND2    gate16006  (.A(g27487), .B(g20498), .Z(g28587) ) ;
OR2     gate16007  (.A(g24608), .B(g26022), .Z(g27489) ) ;
AND2    gate16008  (.A(g27489), .B(g20499), .Z(g28588) ) ;
OR2     gate16009  (.A(g26051), .B(g13431), .Z(g27515) ) ;
AND2    gate16010  (.A(g27515), .B(g20508), .Z(g28597) ) ;
NOR2    gate16011  (.A(g26398), .B(g26484), .Z(g27027) ) ;
AND2    gate16012  (.A(g27027), .B(g8922), .Z(g28599) ) ;
OR2     gate16013  (.A(g26021), .B(g24639), .Z(g27506) ) ;
AND2    gate16014  (.A(g27506), .B(g20514), .Z(g28601) ) ;
OR2     gate16015  (.A(g26023), .B(g24640), .Z(g27509) ) ;
AND2    gate16016  (.A(g27509), .B(g20515), .Z(g28602) ) ;
OR2     gate16017  (.A(g26050), .B(g24649), .Z(g27524) ) ;
AND2    gate16018  (.A(g27524), .B(g20539), .Z(g28612) ) ;
OR2     gate16019  (.A(g16176), .B(g26084), .Z(g27532) ) ;
AND2    gate16020  (.A(g27532), .B(g20551), .Z(g28616) ) ;
OR2     gate16021  (.A(g26078), .B(g24659), .Z(g27533) ) ;
AND2    gate16022  (.A(g27533), .B(g20552), .Z(g28617) ) ;
NOR2    gate16023  (.A(g1024), .B(g19699), .Z(g22357) ) ;
AND2    gate16024  (.A(g22357), .B(g27009), .Z(g28624) ) ;
OR2     gate16025  (.A(g16190), .B(g26094), .Z(g27542) ) ;
AND2    gate16026  (.A(g27542), .B(g20573), .Z(g28626) ) ;
OR2     gate16027  (.A(g26085), .B(g24670), .Z(g27543) ) ;
AND2    gate16028  (.A(g27543), .B(g20574), .Z(g28627) ) ;
OR2     gate16029  (.A(g26087), .B(g24671), .Z(g27544) ) ;
AND2    gate16030  (.A(g27544), .B(g20575), .Z(g28630) ) ;
NOR2    gate16031  (.A(g1367), .B(g19720), .Z(g22399) ) ;
AND2    gate16032  (.A(g22399), .B(g27011), .Z(g28637) ) ;
OR2     gate16033  (.A(g26091), .B(g24675), .Z(g27551) ) ;
AND2    gate16034  (.A(g27551), .B(g20583), .Z(g28638) ) ;
NAND2   gate16035  (.A(II26367), .B(II26368), .Z(g27767) ) ;
AND2    gate16036  (.A(g27767), .B(g20597), .Z(g28639) ) ;
OR2     gate16037  (.A(g26095), .B(g24686), .Z(g27555) ) ;
AND2    gate16038  (.A(g27555), .B(g20598), .Z(g28642) ) ;
OR2     gate16039  (.A(g26097), .B(g24687), .Z(g27556) ) ;
AND2    gate16040  (.A(g27556), .B(g20599), .Z(g28645) ) ;
NAND4   gate16041  (.A(g11192), .B(g26269), .C(g26248), .D(g479), .Z(g27282) ) ;
AND2    gate16042  (.A(g7544), .B(g27014), .Z(g28653) ) ;
AND2    gate16043  (.A(g1030), .B(g27108), .Z(g28654) ) ;
OR2     gate16044  (.A(g26100), .B(g24702), .Z(g27561) ) ;
AND2    gate16045  (.A(g27561), .B(g20603), .Z(g28655) ) ;
OR2     gate16046  (.A(g26102), .B(g24703), .Z(g27562) ) ;
AND2    gate16047  (.A(g27562), .B(g20606), .Z(g28657) ) ;
OR2     gate16048  (.A(g26104), .B(g24704), .Z(g27563) ) ;
AND2    gate16049  (.A(g27563), .B(g20611), .Z(g28658) ) ;
NAND2   gate16050  (.A(II26394), .B(II26395), .Z(g27824) ) ;
AND2    gate16051  (.A(g27824), .B(g20623), .Z(g28660) ) ;
OR2     gate16052  (.A(g26119), .B(g24713), .Z(g27566) ) ;
AND2    gate16053  (.A(g27566), .B(g20624), .Z(g28663) ) ;
OR2     gate16054  (.A(g26121), .B(g24714), .Z(g27567) ) ;
AND2    gate16055  (.A(g27567), .B(g20625), .Z(g28666) ) ;
AND2    gate16056  (.A(g7577), .B(g27017), .Z(g28672) ) ;
AND2    gate16057  (.A(g1373), .B(g27122), .Z(g28673) ) ;
OR2     gate16058  (.A(g26124), .B(g24721), .Z(g27569) ) ;
AND2    gate16059  (.A(g27569), .B(g20629), .Z(g28674) ) ;
OR2     gate16060  (.A(g26126), .B(g24722), .Z(g27570) ) ;
AND2    gate16061  (.A(g27570), .B(g20632), .Z(g28676) ) ;
OR2     gate16062  (.A(g26127), .B(g24723), .Z(g27571) ) ;
AND2    gate16063  (.A(g27571), .B(g20635), .Z(g28677) ) ;
OR2     gate16064  (.A(g26129), .B(g24724), .Z(g27572) ) ;
AND2    gate16065  (.A(g27572), .B(g20638), .Z(g28679) ) ;
NAND2   gate16066  (.A(II26418), .B(II26419), .Z(g27876) ) ;
AND2    gate16067  (.A(g27876), .B(g20649), .Z(g28683) ) ;
OR2     gate16068  (.A(g26145), .B(g24730), .Z(g27574) ) ;
AND2    gate16069  (.A(g27574), .B(g20650), .Z(g28686) ) ;
OR2     gate16070  (.A(g26147), .B(g24731), .Z(g27575) ) ;
AND2    gate16071  (.A(g27575), .B(g20651), .Z(g28689) ) ;
OR2     gate16072  (.A(g26155), .B(g24747), .Z(g27578) ) ;
AND2    gate16073  (.A(g27578), .B(g20661), .Z(g28692) ) ;
OR2     gate16074  (.A(g26157), .B(g24748), .Z(g27579) ) ;
AND2    gate16075  (.A(g27579), .B(g20664), .Z(g28694) ) ;
OR2     gate16076  (.A(g26159), .B(g24749), .Z(g27580) ) ;
AND2    gate16077  (.A(g27580), .B(g20666), .Z(g28695) ) ;
OR2     gate16078  (.A(g26161), .B(g24750), .Z(g27581) ) ;
AND2    gate16079  (.A(g27581), .B(g20669), .Z(g28697) ) ;
NAND2   gate16080  (.A(II26439), .B(II26440), .Z(g27925) ) ;
AND2    gate16081  (.A(g27925), .B(g20680), .Z(g28703) ) ;
OR2     gate16082  (.A(g26165), .B(g24758), .Z(g27584) ) ;
AND2    gate16083  (.A(g27584), .B(g20681), .Z(g28706) ) ;
OR2     gate16084  (.A(g26177), .B(g24763), .Z(g27589) ) ;
AND2    gate16085  (.A(g27589), .B(g20703), .Z(g28710) ) ;
OR2     gate16086  (.A(g26179), .B(g24764), .Z(g27590) ) ;
AND2    gate16087  (.A(g27590), .B(g20708), .Z(g28712) ) ;
OR2     gate16088  (.A(g26181), .B(g24765), .Z(g27591) ) ;
AND2    gate16089  (.A(g27591), .B(g20711), .Z(g28714) ) ;
NAND2   gate16090  (.A(II26460), .B(II26461), .Z(g27955) ) ;
AND2    gate16091  (.A(g27955), .B(g20738), .Z(g28722) ) ;
OR2     gate16092  (.A(g26207), .B(g24775), .Z(g27596) ) ;
AND2    gate16093  (.A(g27596), .B(g20779), .Z(g28725) ) ;
AND4    gate16094  (.A(g21434), .B(g26424), .C(g25274), .D(g27395), .Z(g28739) ) ;
AND4    gate16095  (.A(g21434), .B(g26424), .C(g25299), .D(g27416), .Z(g28761) ) ;
AND4    gate16096  (.A(g21434), .B(g26424), .C(g25308), .D(g27421), .Z(g28768) ) ;
AND4    gate16097  (.A(g21434), .B(g26424), .C(g25340), .D(g27440), .Z(g28789) ) ;
AND4    gate16098  (.A(g21434), .B(g26424), .C(g25348), .D(g27445), .Z(g28799) ) ;
OR2     gate16099  (.A(g26780), .B(g25229), .Z(g26972) ) ;
AND2    gate16100  (.A(g26972), .B(g13037), .Z(g28812) ) ;
AND2    gate16101  (.A(g4104), .B(g27038), .Z(g28813) ) ;
AND4    gate16102  (.A(g21434), .B(g26424), .C(g25388), .D(g27469), .Z(g28833) ) ;
AND4    gate16103  (.A(g21434), .B(g26424), .C(g25399), .D(g27474), .Z(g28846) ) ;
AND4    gate16104  (.A(g21434), .B(g26424), .C(g25438), .D(g27494), .Z(g28880) ) ;
OR2     gate16105  (.A(g26323), .B(g24820), .Z(g27663) ) ;
AND2    gate16106  (.A(g27663), .B(g21295), .Z(g28919) ) ;
AND3    gate16107  (.A(g25534), .B(g26424), .C(g22698), .Z(II27349) ) ;
AND4    gate16108  (.A(g27163), .B(g12687), .C(g20682), .D(II27349), .Z(g28982) ) ;
AND3    gate16109  (.A(g25541), .B(g26424), .C(g22698), .Z(II27364) ) ;
AND4    gate16110  (.A(g27163), .B(g12730), .C(g20739), .D(II27364), .Z(g29008) ) ;
AND3    gate16111  (.A(g25549), .B(g26424), .C(g22698), .Z(II27381) ) ;
AND4    gate16112  (.A(g27163), .B(g12762), .C(g20875), .D(II27381), .Z(g29036) ) ;
AND3    gate16113  (.A(g25556), .B(g26424), .C(g22698), .Z(II27409) ) ;
AND4    gate16114  (.A(g27163), .B(g10290), .C(g21012), .D(II27409), .Z(g29073) ) ;
AND3    gate16115  (.A(g25562), .B(g26424), .C(g22698), .Z(II27429) ) ;
AND4    gate16116  (.A(g27187), .B(g12687), .C(g20751), .D(II27429), .Z(g29110) ) ;
AND2    gate16117  (.A(g27163), .B(g12687), .Z(g29178) ) ;
AND2    gate16118  (.A(g27163), .B(g12730), .Z(g29182) ) ;
AND2    gate16119  (.A(g27163), .B(g12762), .Z(g29188) ) ;
AND2    gate16120  (.A(g27163), .B(g10290), .Z(g29192) ) ;
AND2    gate16121  (.A(g27187), .B(g12687), .Z(g29199) ) ;
AND4    gate16122  (.A(g19890), .B(g24075), .C(g24076), .D(g28032), .Z(II27503) ) ;
AND4    gate16123  (.A(g24077), .B(g24078), .C(g24079), .D(g24080), .Z(II27504) ) ;
AND3    gate16124  (.A(g24081), .B(II27503), .C(II27504), .Z(g29201) ) ;
AND4    gate16125  (.A(g19935), .B(g24082), .C(g24083), .D(g28033), .Z(II27508) ) ;
AND4    gate16126  (.A(g24084), .B(g24085), .C(g24086), .D(g24087), .Z(II27509) ) ;
AND3    gate16127  (.A(g24088), .B(II27508), .C(II27509), .Z(g29202) ) ;
AND4    gate16128  (.A(g19984), .B(g24089), .C(g24090), .D(g28034), .Z(II27513) ) ;
AND4    gate16129  (.A(g24091), .B(g24092), .C(g24093), .D(g24094), .Z(II27514) ) ;
AND3    gate16130  (.A(g24095), .B(II27513), .C(II27514), .Z(g29203) ) ;
AND4    gate16131  (.A(g20720), .B(g24104), .C(g24105), .D(g24106), .Z(II27518) ) ;
AND4    gate16132  (.A(g28036), .B(g24107), .C(g24108), .D(g24109), .Z(II27519) ) ;
AND3    gate16133  (.A(g24110), .B(II27518), .C(II27519), .Z(g29204) ) ;
AND4    gate16134  (.A(g20857), .B(g24111), .C(g24112), .D(g24113), .Z(II27523) ) ;
AND4    gate16135  (.A(g28037), .B(g24114), .C(g24115), .D(g24116), .Z(II27524) ) ;
AND3    gate16136  (.A(g24117), .B(II27523), .C(II27524), .Z(g29205) ) ;
AND4    gate16137  (.A(g20998), .B(g24118), .C(g24119), .D(g24120), .Z(II27528) ) ;
AND4    gate16138  (.A(g28038), .B(g24121), .C(g24122), .D(g24123), .Z(II27529) ) ;
AND3    gate16139  (.A(g24124), .B(II27528), .C(II27529), .Z(g29206) ) ;
AND4    gate16140  (.A(g21143), .B(g24125), .C(g24126), .D(g24127), .Z(II27533) ) ;
AND4    gate16141  (.A(g28039), .B(g24128), .C(g24129), .D(g24130), .Z(II27534) ) ;
AND3    gate16142  (.A(g24131), .B(II27533), .C(II27534), .Z(g29207) ) ;
AND4    gate16143  (.A(g21209), .B(g24132), .C(g24133), .D(g24134), .Z(II27538) ) ;
AND4    gate16144  (.A(g28040), .B(g24135), .C(g24136), .D(g24137), .Z(II27539) ) ;
AND3    gate16145  (.A(g24138), .B(II27538), .C(II27539), .Z(g29208) ) ;
NOR3    gate16146  (.A(g5164), .B(g7704), .C(g27999), .Z(g29005) ) ;
AND2    gate16147  (.A(g29005), .B(g22144), .Z(g29314) ) ;
AND3    gate16148  (.A(g29188), .B(g7051), .C(g5990), .Z(g29315) ) ;
AND3    gate16149  (.A(g28528), .B(g6875), .C(g3288), .Z(g29316) ) ;
OR2     gate16150  (.A(g27628), .B(g17119), .Z(g29068) ) ;
AND2    gate16151  (.A(g29068), .B(g22147), .Z(g29320) ) ;
NOR3    gate16152  (.A(g5511), .B(g7738), .C(g28010), .Z(g29033) ) ;
AND2    gate16153  (.A(g29033), .B(g22148), .Z(g29321) ) ;
AND3    gate16154  (.A(g29192), .B(g7074), .C(g6336), .Z(g29322) ) ;
AND3    gate16155  (.A(g28539), .B(g6905), .C(g3639), .Z(g29323) ) ;
OR2     gate16156  (.A(g27633), .B(g26572), .Z(g29078) ) ;
AND2    gate16157  (.A(g29078), .B(g18883), .Z(g29324) ) ;
OR2     gate16158  (.A(g27645), .B(g17134), .Z(g29105) ) ;
AND2    gate16159  (.A(g29105), .B(g22155), .Z(g29326) ) ;
NOR3    gate16160  (.A(g5857), .B(g7766), .C(g28020), .Z(g29070) ) ;
AND2    gate16161  (.A(g29070), .B(g22156), .Z(g29327) ) ;
AND3    gate16162  (.A(g28553), .B(g6928), .C(g3990), .Z(g29328) ) ;
AND2    gate16163  (.A(g7995), .B(g28353), .Z(g29329) ) ;
OR2     gate16164  (.A(g27646), .B(g26602), .Z(g29114) ) ;
AND2    gate16165  (.A(g29114), .B(g18894), .Z(g29330) ) ;
OR2     gate16166  (.A(g27650), .B(g17146), .Z(g29143) ) ;
AND2    gate16167  (.A(g29143), .B(g22169), .Z(g29331) ) ;
NOR3    gate16168  (.A(g6203), .B(g7791), .C(g26977), .Z(g29107) ) ;
AND2    gate16169  (.A(g29107), .B(g22170), .Z(g29332) ) ;
OR2     gate16170  (.A(g27651), .B(g26606), .Z(g29148) ) ;
AND2    gate16171  (.A(g29148), .B(g18908), .Z(g29334) ) ;
AND2    gate16172  (.A(g4704), .B(g28363), .Z(g29336) ) ;
OR2     gate16173  (.A(g27653), .B(g17153), .Z(g29166) ) ;
AND2    gate16174  (.A(g29166), .B(g22180), .Z(g29337) ) ;
NOR3    gate16175  (.A(g6549), .B(g7812), .C(g26994), .Z(g29145) ) ;
AND2    gate16176  (.A(g29145), .B(g22181), .Z(g29338) ) ;
OR2     gate16177  (.A(g27658), .B(g26613), .Z(g29168) ) ;
AND2    gate16178  (.A(g29168), .B(g18932), .Z(g29344) ) ;
AND2    gate16179  (.A(g4749), .B(g28376), .Z(g29345) ) ;
AND2    gate16180  (.A(g4894), .B(g28381), .Z(g29346) ) ;
OR2     gate16181  (.A(g27661), .B(g17177), .Z(g29176) ) ;
AND2    gate16182  (.A(g29176), .B(g22201), .Z(g29347) ) ;
AND2    gate16183  (.A(g4760), .B(g28391), .Z(g29349) ) ;
AND2    gate16184  (.A(g4939), .B(g28395), .Z(g29350) ) ;
AND2    gate16185  (.A(g4771), .B(g28406), .Z(g29351) ) ;
AND2    gate16186  (.A(g4950), .B(g28410), .Z(g29352) ) ;
AND2    gate16187  (.A(g4961), .B(g28421), .Z(g29354) ) ;
NOR2    gate16188  (.A(g8426), .B(g26616), .Z(g27364) ) ;
AND2    gate16189  (.A(g27364), .B(g28294), .Z(g29360) ) ;
NOR2    gate16190  (.A(g8492), .B(g26636), .Z(g27379) ) ;
AND2    gate16191  (.A(g27379), .B(g28307), .Z(g29362) ) ;
AND2    gate16192  (.A(g8458), .B(g28444), .Z(g29363) ) ;
NOR2    gate16193  (.A(g8553), .B(g26657), .Z(g27400) ) ;
AND2    gate16194  (.A(g27400), .B(g28321), .Z(g29364) ) ;
AND2    gate16195  (.A(g8575), .B(g28325), .Z(g29367) ) ;
OR2     gate16196  (.A(g27223), .B(g27141), .Z(g28209) ) ;
AND2    gate16197  (.A(g28209), .B(g22341), .Z(g29369) ) ;
NOR2    gate16198  (.A(g8651), .B(g11083), .Z(g13946) ) ;
AND2    gate16199  (.A(g13946), .B(g28370), .Z(g29375) ) ;
NOR2    gate16200  (.A(g8681), .B(g11083), .Z(g14002) ) ;
AND2    gate16201  (.A(g14002), .B(g28504), .Z(g29376) ) ;
OR2     gate16202  (.A(g27932), .B(g27957), .Z(g28132) ) ;
AND2    gate16203  (.A(g28132), .B(g19387), .Z(g29377) ) ;
AND2    gate16204  (.A(g28137), .B(g22493), .Z(g29378) ) ;
OR2     gate16205  (.A(g27958), .B(g27962), .Z(g28134) ) ;
AND2    gate16206  (.A(g28134), .B(g19396), .Z(g29380) ) ;
OR2     gate16207  (.A(g27959), .B(g27963), .Z(g28135) ) ;
AND2    gate16208  (.A(g28135), .B(g19399), .Z(g29381) ) ;
OR4     gate16209  (.A(g27469), .B(g27440), .C(g27416), .D(g27395), .Z(g28172) ) ;
OR2     gate16210  (.A(g27964), .B(g27968), .Z(g28138) ) ;
AND2    gate16211  (.A(g28138), .B(g19412), .Z(g29383) ) ;
OR4     gate16212  (.A(g27494), .B(g27474), .C(g27445), .D(g27421), .Z(g28179) ) ;
NOR2    gate16213  (.A(g8808), .B(g12259), .Z(g14033) ) ;
AND2    gate16214  (.A(g14033), .B(g28500), .Z(g29475) ) ;
NOR2    gate16215  (.A(g8851), .B(g12259), .Z(g14090) ) ;
AND2    gate16216  (.A(g14090), .B(g28441), .Z(g29477) ) ;
AND2    gate16217  (.A(g9073), .B(g28479), .Z(g29494) ) ;
AND2    gate16218  (.A(g1600), .B(g28755), .Z(g29509) ) ;
NAND2   gate16219  (.A(g27738), .B(g8093), .Z(g28856) ) ;
AND2    gate16220  (.A(g28856), .B(g22342), .Z(g29510) ) ;
AND2    gate16221  (.A(g1736), .B(g28783), .Z(g29511) ) ;
AND2    gate16222  (.A(g2161), .B(g28793), .Z(g29512) ) ;
NAND2   gate16223  (.A(g23975), .B(g27377), .Z(g28448) ) ;
AND2    gate16224  (.A(g28448), .B(g14095), .Z(g29513) ) ;
AND2    gate16225  (.A(g1608), .B(g28780), .Z(g29514) ) ;
NAND2   gate16226  (.A(g27738), .B(g8139), .Z(g28888) ) ;
AND2    gate16227  (.A(g28888), .B(g22342), .Z(g29515) ) ;
NAND2   gate16228  (.A(g27775), .B(g8146), .Z(g28895) ) ;
AND2    gate16229  (.A(g28895), .B(g22369), .Z(g29516) ) ;
AND2    gate16230  (.A(g1870), .B(g28827), .Z(g29517) ) ;
NAND2   gate16231  (.A(g27796), .B(g8150), .Z(g28906) ) ;
AND2    gate16232  (.A(g28906), .B(g22384), .Z(g29518) ) ;
AND2    gate16233  (.A(g2295), .B(g28840), .Z(g29519) ) ;
AND2    gate16234  (.A(g1744), .B(g28824), .Z(g29521) ) ;
NAND2   gate16235  (.A(g27775), .B(g8195), .Z(g28923) ) ;
AND2    gate16236  (.A(g28923), .B(g22369), .Z(g29522) ) ;
NAND2   gate16237  (.A(g27833), .B(g8201), .Z(g28930) ) ;
AND2    gate16238  (.A(g28930), .B(g22417), .Z(g29523) ) ;
AND2    gate16239  (.A(g2004), .B(g28864), .Z(g29524) ) ;
AND2    gate16240  (.A(g2169), .B(g28837), .Z(g29525) ) ;
NAND2   gate16241  (.A(g27796), .B(g8205), .Z(g28938) ) ;
AND2    gate16242  (.A(g28938), .B(g22384), .Z(g29526) ) ;
NAND2   gate16243  (.A(g27854), .B(g8211), .Z(g28945) ) ;
AND2    gate16244  (.A(g28945), .B(g22432), .Z(g29527) ) ;
AND2    gate16245  (.A(g2429), .B(g28874), .Z(g29528) ) ;
AND2    gate16246  (.A(g1612), .B(g28820), .Z(g29530) ) ;
AND2    gate16247  (.A(g1664), .B(g28559), .Z(g29531) ) ;
AND2    gate16248  (.A(g1878), .B(g28861), .Z(g29532) ) ;
NAND2   gate16249  (.A(g27833), .B(g8249), .Z(g28958) ) ;
AND2    gate16250  (.A(g28958), .B(g22417), .Z(g29533) ) ;
NAND2   gate16251  (.A(g27882), .B(g8255), .Z(g28965) ) ;
AND2    gate16252  (.A(g28965), .B(g22457), .Z(g29534) ) ;
AND2    gate16253  (.A(g2303), .B(g28871), .Z(g29535) ) ;
NAND2   gate16254  (.A(g27854), .B(g8267), .Z(g28969) ) ;
AND2    gate16255  (.A(g28969), .B(g22432), .Z(g29536) ) ;
NAND2   gate16256  (.A(g27903), .B(g8273), .Z(g28976) ) ;
AND2    gate16257  (.A(g28976), .B(g22472), .Z(g29537) ) ;
AND2    gate16258  (.A(g2563), .B(g28914), .Z(g29538) ) ;
AND2    gate16259  (.A(g1748), .B(g28857), .Z(g29547) ) ;
AND2    gate16260  (.A(g1798), .B(g28575), .Z(g29548) ) ;
AND2    gate16261  (.A(g2012), .B(g28900), .Z(g29549) ) ;
NAND2   gate16262  (.A(g27882), .B(g8310), .Z(g28990) ) ;
AND2    gate16263  (.A(g28990), .B(g22457), .Z(g29550) ) ;
AND2    gate16264  (.A(g2173), .B(g28867), .Z(g29551) ) ;
AND2    gate16265  (.A(g2223), .B(g28579), .Z(g29552) ) ;
AND2    gate16266  (.A(g2437), .B(g28911), .Z(g29553) ) ;
NAND2   gate16267  (.A(g27903), .B(g8324), .Z(g28997) ) ;
AND2    gate16268  (.A(g28997), .B(g22472), .Z(g29554) ) ;
NAND2   gate16269  (.A(g27933), .B(g8330), .Z(g29004) ) ;
AND2    gate16270  (.A(g29004), .B(g22498), .Z(g29555) ) ;
AND2    gate16271  (.A(g1616), .B(g28853), .Z(g29563) ) ;
AND2    gate16272  (.A(g1882), .B(g28896), .Z(g29564) ) ;
AND2    gate16273  (.A(g1932), .B(g28590), .Z(g29565) ) ;
AND2    gate16274  (.A(g2307), .B(g28907), .Z(g29566) ) ;
AND2    gate16275  (.A(g2357), .B(g28593), .Z(g29567) ) ;
AND2    gate16276  (.A(g2571), .B(g28950), .Z(g29568) ) ;
NAND2   gate16277  (.A(g27933), .B(g8381), .Z(g29028) ) ;
AND2    gate16278  (.A(g29028), .B(g22498), .Z(g29569) ) ;
AND2    gate16279  (.A(g2763), .B(g28598), .Z(g29570) ) ;
NOR2    gate16280  (.A(g3161), .B(g27602), .Z(g28452) ) ;
AND2    gate16281  (.A(g28452), .B(g11762), .Z(g29571) ) ;
AND2    gate16282  (.A(g1620), .B(g28885), .Z(g29572) ) ;
AND2    gate16283  (.A(g1752), .B(g28892), .Z(g29573) ) ;
AND2    gate16284  (.A(g2016), .B(g28931), .Z(g29574) ) ;
AND2    gate16285  (.A(g2066), .B(g28604), .Z(g29575) ) ;
AND2    gate16286  (.A(g2177), .B(g28903), .Z(g29576) ) ;
AND2    gate16287  (.A(g2441), .B(g28946), .Z(g29577) ) ;
AND2    gate16288  (.A(g2491), .B(g28606), .Z(g29578) ) ;
NOR2    gate16289  (.A(g7980), .B(g27602), .Z(g28457) ) ;
AND2    gate16290  (.A(g28457), .B(g7964), .Z(g29579) ) ;
NOR3    gate16291  (.A(g8011), .B(g27602), .C(g10295), .Z(g28519) ) ;
AND2    gate16292  (.A(g28519), .B(g14186), .Z(g29580) ) ;
NOR2    gate16293  (.A(g3512), .B(g27617), .Z(g28462) ) ;
AND2    gate16294  (.A(g28462), .B(g11796), .Z(g29581) ) ;
NOR2    gate16295  (.A(g9716), .B(g25791), .Z(g27766) ) ;
AND2    gate16296  (.A(g27766), .B(g28608), .Z(g29582) ) ;
AND2    gate16297  (.A(g1706), .B(g29018), .Z(g29584) ) ;
AND2    gate16298  (.A(g1756), .B(g28920), .Z(g29585) ) ;
AND2    gate16299  (.A(g1886), .B(g28927), .Z(g29586) ) ;
AND2    gate16300  (.A(g2181), .B(g28935), .Z(g29587) ) ;
AND2    gate16301  (.A(g2311), .B(g28942), .Z(g29588) ) ;
AND2    gate16302  (.A(g2575), .B(g28977), .Z(g29589) ) ;
AND2    gate16303  (.A(g2625), .B(g28615), .Z(g29590) ) ;
NOR2    gate16304  (.A(g10295), .B(g27602), .Z(g28552) ) ;
AND2    gate16305  (.A(g28552), .B(g11346), .Z(g29591) ) ;
NOR2    gate16306  (.A(g3171), .B(g27602), .Z(g28469) ) ;
AND2    gate16307  (.A(g28469), .B(g11832), .Z(g29592) ) ;
NOR2    gate16308  (.A(g8021), .B(g27617), .Z(g28470) ) ;
AND2    gate16309  (.A(g28470), .B(g7985), .Z(g29593) ) ;
NOR3    gate16310  (.A(g8070), .B(g27617), .C(g10323), .Z(g28529) ) ;
AND2    gate16311  (.A(g28529), .B(g14192), .Z(g29594) ) ;
NOR2    gate16312  (.A(g3863), .B(g27635), .Z(g28475) ) ;
AND2    gate16313  (.A(g28475), .B(g11833), .Z(g29595) ) ;
NOR2    gate16314  (.A(g9792), .B(g25805), .Z(g27823) ) ;
AND2    gate16315  (.A(g27823), .B(g28620), .Z(g29596) ) ;
NAND2   gate16316  (.A(g27738), .B(g14565), .Z(g28823) ) ;
AND2    gate16317  (.A(g28823), .B(g22342), .Z(g29598) ) ;
AND2    gate16318  (.A(g1710), .B(g29018), .Z(g29599) ) ;
AND2    gate16319  (.A(g1840), .B(g29049), .Z(g29600) ) ;
AND2    gate16320  (.A(g1890), .B(g28955), .Z(g29601) ) ;
AND2    gate16321  (.A(g2020), .B(g28962), .Z(g29602) ) ;
AND2    gate16322  (.A(g2265), .B(g29060), .Z(g29603) ) ;
AND2    gate16323  (.A(g2315), .B(g28966), .Z(g29604) ) ;
AND2    gate16324  (.A(g2445), .B(g28973), .Z(g29605) ) ;
NOR2    gate16325  (.A(g8059), .B(g27602), .Z(g28480) ) ;
AND2    gate16326  (.A(g28480), .B(g8011), .Z(g29606) ) ;
NOR2    gate16327  (.A(g8107), .B(g27602), .Z(g28509) ) ;
AND2    gate16328  (.A(g28509), .B(g14208), .Z(g29607) ) ;
NOR2    gate16329  (.A(g10323), .B(g27617), .Z(g28568) ) ;
AND2    gate16330  (.A(g28568), .B(g11385), .Z(g29608) ) ;
NOR2    gate16331  (.A(g3522), .B(g27617), .Z(g28482) ) ;
AND2    gate16332  (.A(g28482), .B(g11861), .Z(g29609) ) ;
NOR2    gate16333  (.A(g8080), .B(g27635), .Z(g28483) ) ;
AND2    gate16334  (.A(g28483), .B(g8026), .Z(g29610) ) ;
NOR3    gate16335  (.A(g8125), .B(g27635), .C(g7121), .Z(g28540) ) ;
AND2    gate16336  (.A(g28540), .B(g14209), .Z(g29611) ) ;
NOR2    gate16337  (.A(g9875), .B(g25821), .Z(g27875) ) ;
AND2    gate16338  (.A(g27875), .B(g28633), .Z(g29612) ) ;
OR2     gate16339  (.A(g27025), .B(g27028), .Z(g28208) ) ;
AND2    gate16340  (.A(g28208), .B(g19763), .Z(g29613) ) ;
NAND2   gate16341  (.A(g27775), .B(g14586), .Z(g28860) ) ;
AND2    gate16342  (.A(g28860), .B(g22369), .Z(g29614) ) ;
AND2    gate16343  (.A(g1844), .B(g29049), .Z(g29615) ) ;
AND2    gate16344  (.A(g1974), .B(g29085), .Z(g29616) ) ;
AND2    gate16345  (.A(g2024), .B(g28987), .Z(g29617) ) ;
NAND2   gate16346  (.A(g27796), .B(g14588), .Z(g28870) ) ;
AND2    gate16347  (.A(g28870), .B(g22384), .Z(g29618) ) ;
AND2    gate16348  (.A(g2269), .B(g29060), .Z(g29619) ) ;
AND2    gate16349  (.A(g2399), .B(g29097), .Z(g29620) ) ;
AND2    gate16350  (.A(g2449), .B(g28994), .Z(g29621) ) ;
AND2    gate16351  (.A(g2579), .B(g29001), .Z(g29622) ) ;
NOR2    gate16352  (.A(g3179), .B(g27602), .Z(g28496) ) ;
AND2    gate16353  (.A(g28496), .B(g11563), .Z(g29623) ) ;
NOR2    gate16354  (.A(g8114), .B(g27617), .Z(g28491) ) ;
AND2    gate16355  (.A(g28491), .B(g8070), .Z(g29624) ) ;
NOR2    gate16356  (.A(g8165), .B(g27617), .Z(g28514) ) ;
AND2    gate16357  (.A(g28514), .B(g14226), .Z(g29625) ) ;
NOR2    gate16358  (.A(g7121), .B(g27635), .Z(g28584) ) ;
AND2    gate16359  (.A(g28584), .B(g11415), .Z(g29626) ) ;
NOR2    gate16360  (.A(g3873), .B(g27635), .Z(g28493) ) ;
AND2    gate16361  (.A(g28493), .B(g11884), .Z(g29627) ) ;
NOR2    gate16362  (.A(g9946), .B(g25839), .Z(g27924) ) ;
AND2    gate16363  (.A(g27924), .B(g28648), .Z(g29628) ) ;
OR2     gate16364  (.A(g27029), .B(g27034), .Z(g28211) ) ;
AND2    gate16365  (.A(g28211), .B(g19779), .Z(g29629) ) ;
OR2     gate16366  (.A(g27030), .B(g27035), .Z(g28212) ) ;
AND2    gate16367  (.A(g28212), .B(g19781), .Z(g29630) ) ;
AND2    gate16368  (.A(g1682), .B(g28656), .Z(g29631) ) ;
NAND2   gate16369  (.A(g27833), .B(g14612), .Z(g28899) ) ;
AND2    gate16370  (.A(g28899), .B(g22417), .Z(g29632) ) ;
AND2    gate16371  (.A(g1978), .B(g29085), .Z(g29633) ) ;
AND2    gate16372  (.A(g2108), .B(g29121), .Z(g29634) ) ;
NAND2   gate16373  (.A(g27854), .B(g14614), .Z(g28910) ) ;
AND2    gate16374  (.A(g28910), .B(g22432), .Z(g29635) ) ;
AND2    gate16375  (.A(g2403), .B(g29097), .Z(g29636) ) ;
AND2    gate16376  (.A(g2533), .B(g29134), .Z(g29637) ) ;
AND2    gate16377  (.A(g2583), .B(g29025), .Z(g29638) ) ;
NOR2    gate16378  (.A(g3530), .B(g27617), .Z(g28510) ) ;
AND2    gate16379  (.A(g28510), .B(g11618), .Z(g29639) ) ;
NOR2    gate16380  (.A(g8172), .B(g27635), .Z(g28498) ) ;
AND2    gate16381  (.A(g28498), .B(g8125), .Z(g29640) ) ;
NOR2    gate16382  (.A(g8229), .B(g27635), .Z(g28520) ) ;
AND2    gate16383  (.A(g28520), .B(g14237), .Z(g29641) ) ;
NOR2    gate16384  (.A(g10014), .B(g25856), .Z(g27954) ) ;
AND2    gate16385  (.A(g27954), .B(g28669), .Z(g29642) ) ;
OR2     gate16386  (.A(g27036), .B(g27043), .Z(g28216) ) ;
AND2    gate16387  (.A(g28216), .B(g19794), .Z(g29644) ) ;
AND2    gate16388  (.A(g1714), .B(g29018), .Z(g29645) ) ;
AND2    gate16389  (.A(g1816), .B(g28675), .Z(g29646) ) ;
NAND2   gate16390  (.A(g27882), .B(g14641), .Z(g28934) ) ;
AND2    gate16391  (.A(g28934), .B(g22457), .Z(g29647) ) ;
AND2    gate16392  (.A(g2112), .B(g29121), .Z(g29648) ) ;
AND2    gate16393  (.A(g2241), .B(g28678), .Z(g29649) ) ;
NAND2   gate16394  (.A(g27903), .B(g14643), .Z(g28949) ) ;
AND2    gate16395  (.A(g28949), .B(g22472), .Z(g29650) ) ;
AND2    gate16396  (.A(g2537), .B(g29134), .Z(g29651) ) ;
AND2    gate16397  (.A(g2667), .B(g29157), .Z(g29652) ) ;
NOR2    gate16398  (.A(g3881), .B(g27635), .Z(g28515) ) ;
AND2    gate16399  (.A(g28515), .B(g11666), .Z(g29656) ) ;
AND2    gate16400  (.A(g1687), .B(g29015), .Z(g29661) ) ;
AND2    gate16401  (.A(g1848), .B(g29049), .Z(g29662) ) ;
AND2    gate16402  (.A(g1950), .B(g28693), .Z(g29663) ) ;
AND2    gate16403  (.A(g2273), .B(g29060), .Z(g29664) ) ;
AND2    gate16404  (.A(g2375), .B(g28696), .Z(g29665) ) ;
NAND2   gate16405  (.A(g27933), .B(g14680), .Z(g28980) ) ;
AND2    gate16406  (.A(g28980), .B(g22498), .Z(g29666) ) ;
AND2    gate16407  (.A(g2671), .B(g29157), .Z(g29667) ) ;
OR2     gate16408  (.A(g27286), .B(g26182), .Z(g28527) ) ;
AND2    gate16409  (.A(g28527), .B(g14255), .Z(g29668) ) ;
AND2    gate16410  (.A(g1821), .B(g29046), .Z(g29683) ) ;
AND2    gate16411  (.A(g1982), .B(g29085), .Z(g29684) ) ;
AND2    gate16412  (.A(g2084), .B(g28711), .Z(g29685) ) ;
AND2    gate16413  (.A(g2246), .B(g29057), .Z(g29686) ) ;
AND2    gate16414  (.A(g2407), .B(g29097), .Z(g29687) ) ;
AND2    gate16415  (.A(g2509), .B(g28713), .Z(g29688) ) ;
NAND3   gate16416  (.A(g12546), .B(g26131), .C(g27977), .Z(g28207) ) ;
AND2    gate16417  (.A(g28207), .B(g10233), .Z(g29693) ) ;
AND2    gate16418  (.A(g1955), .B(g29082), .Z(g29708) ) ;
AND2    gate16419  (.A(g2116), .B(g29121), .Z(g29709) ) ;
AND2    gate16420  (.A(g2380), .B(g29094), .Z(g29710) ) ;
AND2    gate16421  (.A(g2541), .B(g29134), .Z(g29711) ) ;
AND2    gate16422  (.A(g2643), .B(g28726), .Z(g29712) ) ;
NAND3   gate16423  (.A(g10857), .B(g27155), .C(g27142), .Z(g28512) ) ;
AND2    gate16424  (.A(g28512), .B(g11136), .Z(g29718) ) ;
AND2    gate16425  (.A(g2089), .B(g29118), .Z(g29731) ) ;
AND2    gate16426  (.A(g2514), .B(g29131), .Z(g29732) ) ;
AND2    gate16427  (.A(g2675), .B(g29157), .Z(g29733) ) ;
NAND3   gate16428  (.A(g10857), .B(g26131), .C(g27142), .Z(g28522) ) ;
AND2    gate16429  (.A(g28522), .B(g10233), .Z(g29736) ) ;
AND2    gate16430  (.A(g2648), .B(g29154), .Z(g29740) ) ;
NAND3   gate16431  (.A(g10533), .B(g26105), .C(g27004), .Z(g28288) ) ;
AND2    gate16432  (.A(g28288), .B(g10233), .Z(g29742) ) ;
NAND3   gate16433  (.A(g12546), .B(g26105), .C(g27985), .Z(g28206) ) ;
AND2    gate16434  (.A(g28206), .B(g10233), .Z(g29743) ) ;
OR2     gate16435  (.A(g27087), .B(g25909), .Z(g28279) ) ;
AND2    gate16436  (.A(g28279), .B(g20037), .Z(g29746) ) ;
OR2     gate16437  (.A(g27090), .B(g15757), .Z(g28286) ) ;
AND2    gate16438  (.A(g28286), .B(g23196), .Z(g29747) ) ;
OR2     gate16439  (.A(g27094), .B(g15783), .Z(g28295) ) ;
AND2    gate16440  (.A(g28295), .B(g23214), .Z(g29749) ) ;
OR2     gate16441  (.A(g27095), .B(g15784), .Z(g28296) ) ;
AND2    gate16442  (.A(g28296), .B(g23215), .Z(g29750) ) ;
OR2     gate16443  (.A(g27096), .B(g15785), .Z(g28297) ) ;
AND2    gate16444  (.A(g28297), .B(g23216), .Z(g29751) ) ;
NAND3   gate16445  (.A(g10857), .B(g26105), .C(g27155), .Z(g28516) ) ;
AND2    gate16446  (.A(g28516), .B(g10233), .Z(g29752) ) ;
OR2     gate16447  (.A(g27103), .B(g15793), .Z(g28305) ) ;
AND2    gate16448  (.A(g28305), .B(g23221), .Z(g29757) ) ;
OR2     gate16449  (.A(g27104), .B(g15794), .Z(g28306) ) ;
AND2    gate16450  (.A(g28306), .B(g23222), .Z(g29758) ) ;
OR2     gate16451  (.A(g27105), .B(g15795), .Z(g28308) ) ;
AND2    gate16452  (.A(g28308), .B(g23226), .Z(g29759) ) ;
OR2     gate16453  (.A(g27106), .B(g15796), .Z(g28309) ) ;
AND2    gate16454  (.A(g28309), .B(g23227), .Z(g29760) ) ;
OR2     gate16455  (.A(g27107), .B(g15797), .Z(g28310) ) ;
AND2    gate16456  (.A(g28310), .B(g23228), .Z(g29761) ) ;
NAND3   gate16457  (.A(g10533), .B(g26131), .C(g26990), .Z(g28298) ) ;
AND2    gate16458  (.A(g28298), .B(g10233), .Z(g29762) ) ;
OR2     gate16459  (.A(g27113), .B(g15804), .Z(g28316) ) ;
AND2    gate16460  (.A(g28316), .B(g23235), .Z(g29766) ) ;
OR2     gate16461  (.A(g27114), .B(g15805), .Z(g28317) ) ;
AND2    gate16462  (.A(g28317), .B(g23236), .Z(g29767) ) ;
OR2     gate16463  (.A(g27115), .B(g15807), .Z(g28319) ) ;
AND2    gate16464  (.A(g28319), .B(g23237), .Z(g29769) ) ;
OR2     gate16465  (.A(g27116), .B(g15808), .Z(g28320) ) ;
AND2    gate16466  (.A(g28320), .B(g23238), .Z(g29770) ) ;
OR2     gate16467  (.A(g27117), .B(g15809), .Z(g28322) ) ;
AND2    gate16468  (.A(g28322), .B(g23242), .Z(g29771) ) ;
OR2     gate16469  (.A(g27118), .B(g15810), .Z(g28323) ) ;
AND2    gate16470  (.A(g28323), .B(g23243), .Z(g29772) ) ;
NAND3   gate16471  (.A(g12546), .B(g27985), .C(g27977), .Z(g28203) ) ;
AND2    gate16472  (.A(g28203), .B(g10233), .Z(g29773) ) ;
NAND3   gate16473  (.A(g10504), .B(g26131), .C(g26973), .Z(g28287) ) ;
AND2    gate16474  (.A(g28287), .B(g10233), .Z(g29774) ) ;
OR2     gate16475  (.A(g27127), .B(g15812), .Z(g28328) ) ;
AND2    gate16476  (.A(g28328), .B(g23245), .Z(g29782) ) ;
OR2     gate16477  (.A(g27128), .B(g15813), .Z(g28329) ) ;
AND2    gate16478  (.A(g28329), .B(g23246), .Z(g29783) ) ;
OR2     gate16479  (.A(g27129), .B(g15814), .Z(g28331) ) ;
AND2    gate16480  (.A(g28331), .B(g23247), .Z(g29784) ) ;
OR2     gate16481  (.A(g27130), .B(g15815), .Z(g28332) ) ;
AND2    gate16482  (.A(g28332), .B(g23248), .Z(g29785) ) ;
OR2     gate16483  (.A(g27131), .B(g15817), .Z(g28334) ) ;
AND2    gate16484  (.A(g28334), .B(g23249), .Z(g29787) ) ;
OR2     gate16485  (.A(g27132), .B(g15818), .Z(g28335) ) ;
AND2    gate16486  (.A(g28335), .B(g23250), .Z(g29788) ) ;
NAND3   gate16487  (.A(g10504), .B(g26105), .C(g26987), .Z(g28270) ) ;
AND2    gate16488  (.A(g28270), .B(g10233), .Z(g29789) ) ;
OR2     gate16489  (.A(g27134), .B(g15819), .Z(g28342) ) ;
AND2    gate16490  (.A(g28342), .B(g23256), .Z(g29794) ) ;
OR2     gate16491  (.A(g27136), .B(g15820), .Z(g28344) ) ;
AND2    gate16492  (.A(g28344), .B(g23257), .Z(g29795) ) ;
OR2     gate16493  (.A(g27137), .B(g15821), .Z(g28345) ) ;
AND2    gate16494  (.A(g28345), .B(g23258), .Z(g29796) ) ;
OR2     gate16495  (.A(g27138), .B(g15822), .Z(g28347) ) ;
AND2    gate16496  (.A(g28347), .B(g23259), .Z(g29797) ) ;
OR2     gate16497  (.A(g27139), .B(g15823), .Z(g28348) ) ;
AND2    gate16498  (.A(g28348), .B(g23260), .Z(g29798) ) ;
NAND3   gate16499  (.A(g10533), .B(g27004), .C(g26990), .Z(g28271) ) ;
AND2    gate16500  (.A(g28271), .B(g10233), .Z(g29799) ) ;
NOR2    gate16501  (.A(g27467), .B(g26347), .Z(g28414) ) ;
AND2    gate16502  (.A(g28414), .B(g26836), .Z(g29803) ) ;
AND2    gate16503  (.A(g1592), .B(g29014), .Z(g29804) ) ;
OR2     gate16504  (.A(g27148), .B(g15836), .Z(g28357) ) ;
AND2    gate16505  (.A(g28357), .B(g23270), .Z(g29805) ) ;
OR2     gate16506  (.A(g27149), .B(g15837), .Z(g28358) ) ;
AND2    gate16507  (.A(g28358), .B(g23271), .Z(g29806) ) ;
OR2     gate16508  (.A(g27151), .B(g15838), .Z(g28359) ) ;
AND2    gate16509  (.A(g28359), .B(g23272), .Z(g29807) ) ;
OR2     gate16510  (.A(g27153), .B(g15839), .Z(g28361) ) ;
AND2    gate16511  (.A(g28361), .B(g23273), .Z(g29808) ) ;
OR2     gate16512  (.A(g27154), .B(g15840), .Z(g28362) ) ;
AND2    gate16513  (.A(g28362), .B(g23274), .Z(g29809) ) ;
NAND3   gate16514  (.A(g10504), .B(g26987), .C(g26973), .Z(g28259) ) ;
AND2    gate16515  (.A(g28259), .B(g11317), .Z(g29810) ) ;
OR2     gate16516  (.A(g27158), .B(g27184), .Z(g28368) ) ;
AND2    gate16517  (.A(g28368), .B(g23278), .Z(g29834) ) ;
AND2    gate16518  (.A(g28326), .B(g24866), .Z(g29835) ) ;
NOR2    gate16519  (.A(g27493), .B(g26351), .Z(g28425) ) ;
AND2    gate16520  (.A(g28425), .B(g26841), .Z(g29836) ) ;
OR2     gate16521  (.A(g27160), .B(g25938), .Z(g28369) ) ;
AND2    gate16522  (.A(g28369), .B(g20144), .Z(g29837) ) ;
AND2    gate16523  (.A(g1636), .B(g29044), .Z(g29838) ) ;
AND2    gate16524  (.A(g1728), .B(g29045), .Z(g29839) ) ;
AND2    gate16525  (.A(g2153), .B(g29056), .Z(g29840) ) ;
OR2     gate16526  (.A(g27177), .B(g15847), .Z(g28371) ) ;
AND2    gate16527  (.A(g28371), .B(g23283), .Z(g29841) ) ;
OR2     gate16528  (.A(g27178), .B(g15848), .Z(g28372) ) ;
AND2    gate16529  (.A(g28372), .B(g23284), .Z(g29842) ) ;
OR2     gate16530  (.A(g27180), .B(g15849), .Z(g28373) ) ;
AND2    gate16531  (.A(g28373), .B(g23289), .Z(g29843) ) ;
OR2     gate16532  (.A(g27181), .B(g15850), .Z(g28374) ) ;
AND2    gate16533  (.A(g28374), .B(g23290), .Z(g29844) ) ;
OR2     gate16534  (.A(g27183), .B(g15851), .Z(g28375) ) ;
AND2    gate16535  (.A(g28375), .B(g23291), .Z(g29845) ) ;
NOR2    gate16536  (.A(g27439), .B(g26339), .Z(g28340) ) ;
AND2    gate16537  (.A(g28340), .B(g24893), .Z(g29850) ) ;
AND2    gate16538  (.A(g1668), .B(g29079), .Z(g29851) ) ;
AND2    gate16539  (.A(g1772), .B(g29080), .Z(g29852) ) ;
AND2    gate16540  (.A(g1862), .B(g29081), .Z(g29853) ) ;
AND2    gate16541  (.A(g2197), .B(g29092), .Z(g29854) ) ;
AND2    gate16542  (.A(g2287), .B(g29093), .Z(g29855) ) ;
OR2     gate16543  (.A(g27201), .B(g15857), .Z(g28385) ) ;
AND2    gate16544  (.A(g28385), .B(g23303), .Z(g29856) ) ;
OR2     gate16545  (.A(g27202), .B(g13277), .Z(g28386) ) ;
AND2    gate16546  (.A(g28386), .B(g23304), .Z(g29857) ) ;
OR2     gate16547  (.A(g27203), .B(g15858), .Z(g28387) ) ;
AND2    gate16548  (.A(g28387), .B(g23306), .Z(g29858) ) ;
OR2     gate16549  (.A(g27204), .B(g15859), .Z(g28388) ) ;
AND2    gate16550  (.A(g28388), .B(g23307), .Z(g29859) ) ;
OR2     gate16551  (.A(g27206), .B(g15860), .Z(g28389) ) ;
AND2    gate16552  (.A(g28389), .B(g23312), .Z(g29860) ) ;
OR2     gate16553  (.A(g27207), .B(g15861), .Z(g28390) ) ;
AND2    gate16554  (.A(g28390), .B(g23313), .Z(g29861) ) ;
AND2    gate16555  (.A(g1802), .B(g29115), .Z(g29865) ) ;
AND2    gate16556  (.A(g1906), .B(g29116), .Z(g29866) ) ;
AND2    gate16557  (.A(g1996), .B(g29117), .Z(g29867) ) ;
AND2    gate16558  (.A(g2227), .B(g29128), .Z(g29868) ) ;
AND2    gate16559  (.A(g2331), .B(g29129), .Z(g29869) ) ;
AND2    gate16560  (.A(g2421), .B(g29130), .Z(g29870) ) ;
OR2     gate16561  (.A(g27211), .B(g15870), .Z(g28400) ) ;
AND2    gate16562  (.A(g28400), .B(g23332), .Z(g29871) ) ;
OR2     gate16563  (.A(g27212), .B(g15871), .Z(g28401) ) ;
AND2    gate16564  (.A(g28401), .B(g23333), .Z(g29872) ) ;
OR2     gate16565  (.A(g27213), .B(g15873), .Z(g28402) ) ;
AND2    gate16566  (.A(g28402), .B(g23336), .Z(g29874) ) ;
OR2     gate16567  (.A(g27214), .B(g13282), .Z(g28403) ) ;
AND2    gate16568  (.A(g28403), .B(g23337), .Z(g29875) ) ;
OR2     gate16569  (.A(g27215), .B(g15874), .Z(g28404) ) ;
AND2    gate16570  (.A(g28404), .B(g23339), .Z(g29876) ) ;
OR2     gate16571  (.A(g27216), .B(g15875), .Z(g28405) ) ;
AND2    gate16572  (.A(g28405), .B(g23340), .Z(g29877) ) ;
AND2    gate16573  (.A(g1936), .B(g29149), .Z(g29880) ) ;
AND2    gate16574  (.A(g2040), .B(g29150), .Z(g29881) ) ;
AND2    gate16575  (.A(g2361), .B(g29151), .Z(g29882) ) ;
AND2    gate16576  (.A(g2465), .B(g29152), .Z(g29883) ) ;
AND2    gate16577  (.A(g2555), .B(g29153), .Z(g29884) ) ;
OR2     gate16578  (.A(g27218), .B(g15880), .Z(g28416) ) ;
AND2    gate16579  (.A(g28416), .B(g23350), .Z(g29885) ) ;
OR2     gate16580  (.A(g27219), .B(g15881), .Z(g28417) ) ;
AND2    gate16581  (.A(g28417), .B(g23351), .Z(g29887) ) ;
OR2     gate16582  (.A(g27220), .B(g15882), .Z(g28418) ) ;
AND2    gate16583  (.A(g28418), .B(g23352), .Z(g29888) ) ;
OR2     gate16584  (.A(g27221), .B(g15884), .Z(g28419) ) ;
AND2    gate16585  (.A(g28419), .B(g23355), .Z(g29890) ) ;
OR2     gate16586  (.A(g27222), .B(g13290), .Z(g28420) ) ;
AND2    gate16587  (.A(g28420), .B(g23356), .Z(g29891) ) ;
AND2    gate16588  (.A(g2070), .B(g29169), .Z(g29894) ) ;
AND2    gate16589  (.A(g2495), .B(g29170), .Z(g29895) ) ;
AND2    gate16590  (.A(g2599), .B(g29171), .Z(g29896) ) ;
OR2     gate16591  (.A(g27227), .B(g15912), .Z(g28428) ) ;
AND2    gate16592  (.A(g28428), .B(g23375), .Z(g29899) ) ;
OR2     gate16593  (.A(g27228), .B(g15913), .Z(g28429) ) ;
AND2    gate16594  (.A(g28429), .B(g23376), .Z(g29901) ) ;
OR2     gate16595  (.A(g27229), .B(g15914), .Z(g28430) ) ;
AND2    gate16596  (.A(g28430), .B(g23377), .Z(g29902) ) ;
AND2    gate16597  (.A(g2629), .B(g29177), .Z(g29907) ) ;
OR2     gate16598  (.A(g27234), .B(g15967), .Z(g28435) ) ;
AND2    gate16599  (.A(g28435), .B(g23388), .Z(g29909) ) ;
NOR2    gate16600  (.A(g7301), .B(g10741), .Z(g13031) ) ;
AND2    gate16601  (.A(g13031), .B(g29190), .Z(g29924) ) ;
AND2    gate16602  (.A(g1604), .B(g28736), .Z(g29926) ) ;
NOR2    gate16603  (.A(g7349), .B(g10762), .Z(g13044) ) ;
AND2    gate16604  (.A(g13044), .B(g29196), .Z(g29937) ) ;
NAND2   gate16605  (.A(II22684), .B(II22685), .Z(g23552) ) ;
AND2    gate16606  (.A(g23552), .B(g28889), .Z(g29938) ) ;
AND2    gate16607  (.A(g1740), .B(g28758), .Z(g29940) ) ;
AND2    gate16608  (.A(g2165), .B(g28765), .Z(g29943) ) ;
NAND2   gate16609  (.A(II22711), .B(II22712), .Z(g23575) ) ;
AND2    gate16610  (.A(g23575), .B(g28924), .Z(g29949) ) ;
AND2    gate16611  (.A(g1874), .B(g28786), .Z(g29951) ) ;
NAND2   gate16612  (.A(II22718), .B(II22719), .Z(g23576) ) ;
AND2    gate16613  (.A(g23576), .B(g28939), .Z(g29952) ) ;
AND2    gate16614  (.A(g2299), .B(g28796), .Z(g29954) ) ;
NOR2    gate16615  (.A(g5170), .B(g27999), .Z(g28953) ) ;
AND2    gate16616  (.A(g28953), .B(g12823), .Z(g29959) ) ;
NAND2   gate16617  (.A(II22754), .B(II22755), .Z(g23616) ) ;
AND2    gate16618  (.A(g23616), .B(g28959), .Z(g29962) ) ;
AND2    gate16619  (.A(g2008), .B(g28830), .Z(g29964) ) ;
NAND2   gate16620  (.A(II22761), .B(II22762), .Z(g23617) ) ;
AND2    gate16621  (.A(g23617), .B(g28970), .Z(g29966) ) ;
AND2    gate16622  (.A(g2433), .B(g28843), .Z(g29968) ) ;
AND2    gate16623  (.A(g28121), .B(g20509), .Z(g29969) ) ;
NOR2    gate16624  (.A(g9234), .B(g27999), .Z(g28981) ) ;
AND2    gate16625  (.A(g28981), .B(g9206), .Z(g29973) ) ;
NOR3    gate16626  (.A(g9259), .B(g27999), .C(g7704), .Z(g29173) ) ;
AND2    gate16627  (.A(g29173), .B(g12914), .Z(g29974) ) ;
NOR2    gate16628  (.A(g5517), .B(g28010), .Z(g28986) ) ;
AND2    gate16629  (.A(g28986), .B(g10420), .Z(g29975) ) ;
NAND2   gate16630  (.A(II22793), .B(II22794), .Z(g23655) ) ;
AND2    gate16631  (.A(g23655), .B(g28991), .Z(g29979) ) ;
NAND2   gate16632  (.A(II22800), .B(II22801), .Z(g23656) ) ;
AND2    gate16633  (.A(g23656), .B(g28998), .Z(g29982) ) ;
AND2    gate16634  (.A(g2567), .B(g28877), .Z(g29984) ) ;
AND2    gate16635  (.A(g28127), .B(g20532), .Z(g29985) ) ;
NOR3    gate16636  (.A(g3155), .B(g10295), .C(g27602), .Z(g28468) ) ;
AND2    gate16637  (.A(g28468), .B(g23473), .Z(g29986) ) ;
OR2     gate16638  (.A(g27187), .B(g27163), .Z(g29197) ) ;
NOR2    gate16639  (.A(g7704), .B(g27999), .Z(g29187) ) ;
AND2    gate16640  (.A(g29187), .B(g12235), .Z(g29988) ) ;
NOR2    gate16641  (.A(g5180), .B(g27999), .Z(g29006) ) ;
AND2    gate16642  (.A(g29006), .B(g10489), .Z(g29989) ) ;
NOR2    gate16643  (.A(g9269), .B(g28010), .Z(g29007) ) ;
AND2    gate16644  (.A(g29007), .B(g9239), .Z(g29990) ) ;
NOR3    gate16645  (.A(g9311), .B(g28010), .C(g7738), .Z(g29179) ) ;
AND2    gate16646  (.A(g29179), .B(g12922), .Z(g29991) ) ;
NOR2    gate16647  (.A(g5863), .B(g28020), .Z(g29012) ) ;
AND2    gate16648  (.A(g29012), .B(g10490), .Z(g29992) ) ;
NAND2   gate16649  (.A(II22823), .B(II22824), .Z(g23685) ) ;
AND2    gate16650  (.A(g23685), .B(g29029), .Z(g30000) ) ;
OR2     gate16651  (.A(g27262), .B(g16185), .Z(g28490) ) ;
AND2    gate16652  (.A(g28490), .B(g23486), .Z(g30001) ) ;
NOR3    gate16653  (.A(g3506), .B(g10323), .C(g27617), .Z(g28481) ) ;
AND2    gate16654  (.A(g28481), .B(g23487), .Z(g30002) ) ;
NOR2    gate16655  (.A(g27598), .B(g27612), .Z(g28149) ) ;
AND2    gate16656  (.A(g28149), .B(g9021), .Z(g30003) ) ;
NOR2    gate16657  (.A(g27649), .B(g26604), .Z(g28521) ) ;
AND2    gate16658  (.A(g28521), .B(g25837), .Z(g30004) ) ;
OR2     gate16659  (.A(g27669), .B(g14261), .Z(g28230) ) ;
AND2    gate16660  (.A(g28230), .B(g24394), .Z(g30005) ) ;
NOR2    gate16661  (.A(g9300), .B(g27999), .Z(g29032) ) ;
AND2    gate16662  (.A(g29032), .B(g9259), .Z(g30006) ) ;
NOR2    gate16663  (.A(g9374), .B(g27999), .Z(g29141) ) ;
AND2    gate16664  (.A(g29141), .B(g12929), .Z(g30007) ) ;
NOR2    gate16665  (.A(g7738), .B(g28010), .Z(g29191) ) ;
AND2    gate16666  (.A(g29191), .B(g12297), .Z(g30008) ) ;
NOR2    gate16667  (.A(g5527), .B(g28010), .Z(g29034) ) ;
AND2    gate16668  (.A(g29034), .B(g10518), .Z(g30009) ) ;
NOR2    gate16669  (.A(g9321), .B(g28020), .Z(g29035) ) ;
AND2    gate16670  (.A(g29035), .B(g9274), .Z(g30010) ) ;
NOR3    gate16671  (.A(g9392), .B(g28020), .C(g7766), .Z(g29183) ) ;
AND2    gate16672  (.A(g29183), .B(g12930), .Z(g30011) ) ;
NOR2    gate16673  (.A(g6209), .B(g26977), .Z(g29040) ) ;
AND2    gate16674  (.A(g29040), .B(g10519), .Z(g30015) ) ;
AND2    gate16675  (.A(g28508), .B(g20570), .Z(g30023) ) ;
OR2     gate16676  (.A(g27267), .B(g16199), .Z(g28497) ) ;
AND2    gate16677  (.A(g28497), .B(g23501), .Z(g30024) ) ;
NOR3    gate16678  (.A(g3857), .B(g7121), .C(g27635), .Z(g28492) ) ;
AND2    gate16679  (.A(g28492), .B(g23502), .Z(g30025) ) ;
NOR2    gate16680  (.A(g27627), .B(g26547), .Z(g28476) ) ;
AND2    gate16681  (.A(g28476), .B(g25064), .Z(g30026) ) ;
NOR2    gate16682  (.A(g5188), .B(g27999), .Z(g29104) ) ;
AND2    gate16683  (.A(g29104), .B(g12550), .Z(g30027) ) ;
NOR2    gate16684  (.A(g9381), .B(g28010), .Z(g29069) ) ;
AND2    gate16685  (.A(g29069), .B(g9311), .Z(g30028) ) ;
NOR2    gate16686  (.A(g9444), .B(g28010), .Z(g29164) ) ;
AND2    gate16687  (.A(g29164), .B(g12936), .Z(g30029) ) ;
NOR2    gate16688  (.A(g7766), .B(g28020), .Z(g29198) ) ;
AND2    gate16689  (.A(g29198), .B(g12347), .Z(g30030) ) ;
NOR2    gate16690  (.A(g5873), .B(g28020), .Z(g29071) ) ;
AND2    gate16691  (.A(g29071), .B(g10540), .Z(g30031) ) ;
NOR2    gate16692  (.A(g9402), .B(g26977), .Z(g29072) ) ;
AND2    gate16693  (.A(g29072), .B(g9326), .Z(g30032) ) ;
NOR3    gate16694  (.A(g9462), .B(g26977), .C(g7791), .Z(g29189) ) ;
AND2    gate16695  (.A(g29189), .B(g12937), .Z(g30033) ) ;
NOR2    gate16696  (.A(g6555), .B(g26994), .Z(g29077) ) ;
AND2    gate16697  (.A(g29077), .B(g10541), .Z(g30034) ) ;
NOR2    gate16698  (.A(g1030), .B(g19699), .Z(g22539) ) ;
AND2    gate16699  (.A(g22539), .B(g28120), .Z(g30035) ) ;
OR2     gate16700  (.A(g27272), .B(g16208), .Z(g28511) ) ;
AND2    gate16701  (.A(g28511), .B(g23518), .Z(g30041) ) ;
NOR2    gate16702  (.A(g5535), .B(g28010), .Z(g29142) ) ;
AND2    gate16703  (.A(g29142), .B(g12601), .Z(g30042) ) ;
NOR2    gate16704  (.A(g9451), .B(g28020), .Z(g29106) ) ;
AND2    gate16705  (.A(g29106), .B(g9392), .Z(g30043) ) ;
NOR2    gate16706  (.A(g9511), .B(g28020), .Z(g29174) ) ;
AND2    gate16707  (.A(g29174), .B(g12944), .Z(g30044) ) ;
NOR2    gate16708  (.A(g7791), .B(g26977), .Z(g29200) ) ;
AND2    gate16709  (.A(g29200), .B(g12419), .Z(g30045) ) ;
NOR2    gate16710  (.A(g6219), .B(g26977), .Z(g29108) ) ;
AND2    gate16711  (.A(g29108), .B(g10564), .Z(g30046) ) ;
NOR2    gate16712  (.A(g9472), .B(g26994), .Z(g29109) ) ;
AND2    gate16713  (.A(g29109), .B(g9407), .Z(g30047) ) ;
NOR3    gate16714  (.A(g9529), .B(g26994), .C(g7812), .Z(g29193) ) ;
AND2    gate16715  (.A(g29193), .B(g12945), .Z(g30048) ) ;
NOR2    gate16716  (.A(g7528), .B(g10741), .Z(g13114) ) ;
AND2    gate16717  (.A(g13114), .B(g28167), .Z(g30049) ) ;
NOR2    gate16718  (.A(g1373), .B(g19720), .Z(g22545) ) ;
AND2    gate16719  (.A(g22545), .B(g28126), .Z(g30050) ) ;
OR2     gate16720  (.A(g27276), .B(g26123), .Z(g28513) ) ;
AND2    gate16721  (.A(g28513), .B(g20604), .Z(g30051) ) ;
NOR2    gate16722  (.A(g5881), .B(g28020), .Z(g29165) ) ;
AND2    gate16723  (.A(g29165), .B(g12659), .Z(g30056) ) ;
NOR2    gate16724  (.A(g9518), .B(g26977), .Z(g29144) ) ;
AND2    gate16725  (.A(g29144), .B(g9462), .Z(g30057) ) ;
NOR2    gate16726  (.A(g9569), .B(g26977), .Z(g29180) ) ;
AND2    gate16727  (.A(g29180), .B(g12950), .Z(g30058) ) ;
NOR2    gate16728  (.A(g7812), .B(g26994), .Z(g28106) ) ;
AND2    gate16729  (.A(g28106), .B(g12467), .Z(g30059) ) ;
NOR2    gate16730  (.A(g6565), .B(g26994), .Z(g29146) ) ;
AND2    gate16731  (.A(g29146), .B(g10581), .Z(g30060) ) ;
AND2    gate16732  (.A(g1036), .B(g28188), .Z(g30061) ) ;
NOR2    gate16733  (.A(g7553), .B(g10762), .Z(g13129) ) ;
AND2    gate16734  (.A(g13129), .B(g28174), .Z(g30062) ) ;
OR2     gate16735  (.A(g27280), .B(g26154), .Z(g28517) ) ;
AND2    gate16736  (.A(g28517), .B(g20630), .Z(g30064) ) ;
OR2     gate16737  (.A(g27281), .B(g26158), .Z(g28518) ) ;
AND2    gate16738  (.A(g28518), .B(g20636), .Z(g30066) ) ;
NOR2    gate16739  (.A(g6227), .B(g26977), .Z(g29175) ) ;
AND2    gate16740  (.A(g29175), .B(g12708), .Z(g30069) ) ;
NOR2    gate16741  (.A(g9576), .B(g26994), .Z(g29167) ) ;
AND2    gate16742  (.A(g29167), .B(g9529), .Z(g30070) ) ;
NOR2    gate16743  (.A(g9631), .B(g26994), .Z(g29184) ) ;
AND2    gate16744  (.A(g29184), .B(g12975), .Z(g30071) ) ;
AND2    gate16745  (.A(g1379), .B(g28194), .Z(g30073) ) ;
OR2     gate16746  (.A(g27284), .B(g26176), .Z(g28525) ) ;
AND2    gate16747  (.A(g28525), .B(g20662), .Z(g30075) ) ;
OR2     gate16748  (.A(g27285), .B(g26178), .Z(g28526) ) ;
AND2    gate16749  (.A(g28526), .B(g20667), .Z(g30078) ) ;
AND2    gate16750  (.A(g28121), .B(g20674), .Z(g30080) ) ;
NOR2    gate16751  (.A(g6573), .B(g26994), .Z(g29181) ) ;
AND2    gate16752  (.A(g29181), .B(g12752), .Z(g30082) ) ;
OR2     gate16753  (.A(g27291), .B(g26203), .Z(g28533) ) ;
AND2    gate16754  (.A(g28533), .B(g20698), .Z(g30083) ) ;
OR2     gate16755  (.A(g27292), .B(g26204), .Z(g28534) ) ;
AND2    gate16756  (.A(g28534), .B(g20700), .Z(g30084) ) ;
OR2     gate16757  (.A(g27293), .B(g26205), .Z(g28536) ) ;
AND2    gate16758  (.A(g28536), .B(g20704), .Z(g30086) ) ;
OR2     gate16759  (.A(g27294), .B(g26206), .Z(g28538) ) ;
AND2    gate16760  (.A(g28538), .B(g20709), .Z(g30089) ) ;
AND2    gate16761  (.A(g28127), .B(g20716), .Z(g30091) ) ;
OR2     gate16762  (.A(g27300), .B(g26229), .Z(g28544) ) ;
AND2    gate16763  (.A(g28544), .B(g20767), .Z(g30094) ) ;
OR2     gate16764  (.A(g27301), .B(g26230), .Z(g28545) ) ;
AND2    gate16765  (.A(g28545), .B(g20768), .Z(g30095) ) ;
OR2     gate16766  (.A(g27302), .B(g26231), .Z(g28546) ) ;
AND2    gate16767  (.A(g28546), .B(g20770), .Z(g30096) ) ;
OR2     gate16768  (.A(g27303), .B(g26232), .Z(g28548) ) ;
AND2    gate16769  (.A(g28548), .B(g20774), .Z(g30098) ) ;
OR2     gate16770  (.A(g27304), .B(g26233), .Z(g28549) ) ;
AND2    gate16771  (.A(g28549), .B(g20776), .Z(g30099) ) ;
OR2     gate16772  (.A(g27305), .B(g26234), .Z(g28551) ) ;
AND2    gate16773  (.A(g28551), .B(g20780), .Z(g30101) ) ;
OR2     gate16774  (.A(g27311), .B(g26249), .Z(g28560) ) ;
AND2    gate16775  (.A(g28560), .B(g20909), .Z(g30107) ) ;
OR2     gate16776  (.A(g27312), .B(g26250), .Z(g28561) ) ;
AND2    gate16777  (.A(g28561), .B(g20910), .Z(g30108) ) ;
OR2     gate16778  (.A(g27313), .B(g26251), .Z(g28562) ) ;
AND2    gate16779  (.A(g28562), .B(g20912), .Z(g30109) ) ;
OR2     gate16780  (.A(g27314), .B(g26252), .Z(g28564) ) ;
AND2    gate16781  (.A(g28564), .B(g20916), .Z(g30110) ) ;
OR2     gate16782  (.A(g27315), .B(g26253), .Z(g28565) ) ;
AND2    gate16783  (.A(g28565), .B(g20917), .Z(g30111) ) ;
OR2     gate16784  (.A(g27316), .B(g26254), .Z(g28566) ) ;
AND2    gate16785  (.A(g28566), .B(g20919), .Z(g30112) ) ;
OR2     gate16786  (.A(g27324), .B(g26270), .Z(g28574) ) ;
AND2    gate16787  (.A(g28574), .B(g21050), .Z(g30118) ) ;
OR2     gate16788  (.A(g27325), .B(g26271), .Z(g28576) ) ;
AND2    gate16789  (.A(g28576), .B(g21051), .Z(g30120) ) ;
OR2     gate16790  (.A(g27326), .B(g26272), .Z(g28577) ) ;
AND2    gate16791  (.A(g28577), .B(g21052), .Z(g30121) ) ;
OR2     gate16792  (.A(g27327), .B(g26273), .Z(g28578) ) ;
AND2    gate16793  (.A(g28578), .B(g21054), .Z(g30122) ) ;
OR2     gate16794  (.A(g27328), .B(g26275), .Z(g28580) ) ;
AND2    gate16795  (.A(g28580), .B(g21055), .Z(g30124) ) ;
OR2     gate16796  (.A(g27329), .B(g26276), .Z(g28581) ) ;
AND2    gate16797  (.A(g28581), .B(g21056), .Z(g30125) ) ;
OR2     gate16798  (.A(g27330), .B(g26277), .Z(g28582) ) ;
AND2    gate16799  (.A(g28582), .B(g21058), .Z(g30126) ) ;
OR2     gate16800  (.A(g27331), .B(g26285), .Z(g28589) ) ;
AND2    gate16801  (.A(g28589), .B(g21178), .Z(g30131) ) ;
OR2     gate16802  (.A(g27332), .B(g26286), .Z(g28591) ) ;
AND2    gate16803  (.A(g28591), .B(g21179), .Z(g30133) ) ;
OR2     gate16804  (.A(g27333), .B(g26288), .Z(g28592) ) ;
AND2    gate16805  (.A(g28592), .B(g21180), .Z(g30135) ) ;
OR2     gate16806  (.A(g27334), .B(g26289), .Z(g28594) ) ;
AND2    gate16807  (.A(g28594), .B(g21181), .Z(g30137) ) ;
OR2     gate16808  (.A(g27335), .B(g26290), .Z(g28595) ) ;
AND2    gate16809  (.A(g28595), .B(g21182), .Z(g30138) ) ;
OR2     gate16810  (.A(g27336), .B(g26291), .Z(g28596) ) ;
AND2    gate16811  (.A(g28596), .B(g21184), .Z(g30139) ) ;
OR2     gate16812  (.A(g27339), .B(g16427), .Z(g28600) ) ;
AND2    gate16813  (.A(g28600), .B(g23749), .Z(g30140) ) ;
OR2     gate16814  (.A(g27340), .B(g26300), .Z(g28603) ) ;
AND2    gate16815  (.A(g28603), .B(g21247), .Z(g30145) ) ;
OR2     gate16816  (.A(g27341), .B(g26302), .Z(g28605) ) ;
AND2    gate16817  (.A(g28605), .B(g21248), .Z(g30149) ) ;
OR2     gate16818  (.A(g27342), .B(g26303), .Z(g28607) ) ;
AND2    gate16819  (.A(g28607), .B(g21249), .Z(g30151) ) ;
OR2     gate16820  (.A(g27346), .B(g16483), .Z(g28609) ) ;
AND2    gate16821  (.A(g28609), .B(g23767), .Z(g30152) ) ;
OR2     gate16822  (.A(g27347), .B(g16484), .Z(g28610) ) ;
AND2    gate16823  (.A(g28610), .B(g23768), .Z(g30153) ) ;
OR2     gate16824  (.A(g27348), .B(g16485), .Z(g28611) ) ;
AND2    gate16825  (.A(g28611), .B(g23769), .Z(g30154) ) ;
OR2     gate16826  (.A(g27350), .B(g26310), .Z(g28613) ) ;
AND2    gate16827  (.A(g28613), .B(g21274), .Z(g30158) ) ;
OR2     gate16828  (.A(g27351), .B(g26311), .Z(g28614) ) ;
AND2    gate16829  (.A(g28614), .B(g21275), .Z(g30161) ) ;
OR2     gate16830  (.A(g27357), .B(g16516), .Z(g28618) ) ;
AND2    gate16831  (.A(g28618), .B(g23787), .Z(g30164) ) ;
OR2     gate16832  (.A(g27358), .B(g16517), .Z(g28619) ) ;
AND2    gate16833  (.A(g28619), .B(g23788), .Z(g30165) ) ;
OR2     gate16834  (.A(g27359), .B(g16518), .Z(g28621) ) ;
AND2    gate16835  (.A(g28621), .B(g23792), .Z(g30166) ) ;
OR2     gate16836  (.A(g27360), .B(g16519), .Z(g28622) ) ;
AND2    gate16837  (.A(g28622), .B(g23793), .Z(g30167) ) ;
OR2     gate16838  (.A(g27361), .B(g16520), .Z(g28623) ) ;
AND2    gate16839  (.A(g28623), .B(g23794), .Z(g30168) ) ;
OR2     gate16840  (.A(g27363), .B(g26324), .Z(g28625) ) ;
AND2    gate16841  (.A(g28625), .B(g21286), .Z(g30172) ) ;
OR2     gate16842  (.A(g27821), .B(g26815), .Z(g28118) ) ;
AND2    gate16843  (.A(g28118), .B(g13082), .Z(g30173) ) ;
OR2     gate16844  (.A(g27370), .B(g16531), .Z(g28628) ) ;
AND2    gate16845  (.A(g28628), .B(g23812), .Z(g30174) ) ;
OR2     gate16846  (.A(g27371), .B(g16532), .Z(g28629) ) ;
AND2    gate16847  (.A(g28629), .B(g23813), .Z(g30175) ) ;
OR2     gate16848  (.A(g27372), .B(g16534), .Z(g28631) ) ;
AND2    gate16849  (.A(g28631), .B(g23814), .Z(g30177) ) ;
OR2     gate16850  (.A(g27373), .B(g16535), .Z(g28632) ) ;
AND2    gate16851  (.A(g28632), .B(g23815), .Z(g30178) ) ;
OR2     gate16852  (.A(g27374), .B(g16536), .Z(g28634) ) ;
AND2    gate16853  (.A(g28634), .B(g23819), .Z(g30179) ) ;
OR2     gate16854  (.A(g27375), .B(g16537), .Z(g28635) ) ;
AND2    gate16855  (.A(g28635), .B(g23820), .Z(g30180) ) ;
OR2     gate16856  (.A(g27376), .B(g16538), .Z(g28636) ) ;
AND2    gate16857  (.A(g28636), .B(g23821), .Z(g30181) ) ;
OR2     gate16858  (.A(g27384), .B(g16590), .Z(g28640) ) ;
AND2    gate16859  (.A(g28640), .B(g23838), .Z(g30185) ) ;
OR2     gate16860  (.A(g27385), .B(g16591), .Z(g28641) ) ;
AND2    gate16861  (.A(g28641), .B(g23839), .Z(g30186) ) ;
OR2     gate16862  (.A(g27386), .B(g16592), .Z(g28643) ) ;
AND2    gate16863  (.A(g28643), .B(g23840), .Z(g30187) ) ;
OR2     gate16864  (.A(g27387), .B(g16593), .Z(g28644) ) ;
AND2    gate16865  (.A(g28644), .B(g23841), .Z(g30188) ) ;
OR2     gate16866  (.A(g27388), .B(g16595), .Z(g28646) ) ;
AND2    gate16867  (.A(g28646), .B(g23842), .Z(g30190) ) ;
OR2     gate16868  (.A(g27389), .B(g16596), .Z(g28647) ) ;
AND2    gate16869  (.A(g28647), .B(g23843), .Z(g30191) ) ;
OR2     gate16870  (.A(g27390), .B(g16597), .Z(g28649) ) ;
AND2    gate16871  (.A(g28649), .B(g23847), .Z(g30192) ) ;
OR2     gate16872  (.A(g27391), .B(g16598), .Z(g28650) ) ;
AND2    gate16873  (.A(g28650), .B(g23848), .Z(g30193) ) ;
OR2     gate16874  (.A(g27392), .B(g16599), .Z(g28651) ) ;
AND2    gate16875  (.A(g28651), .B(g23849), .Z(g30194) ) ;
OR2     gate16876  (.A(g27404), .B(g16610), .Z(g28659) ) ;
AND2    gate16877  (.A(g28659), .B(g23858), .Z(g30196) ) ;
OR2     gate16878  (.A(g27406), .B(g16611), .Z(g28661) ) ;
AND2    gate16879  (.A(g28661), .B(g23859), .Z(g30197) ) ;
OR2     gate16880  (.A(g27407), .B(g16612), .Z(g28662) ) ;
AND2    gate16881  (.A(g28662), .B(g23860), .Z(g30198) ) ;
OR2     gate16882  (.A(g27408), .B(g16613), .Z(g28664) ) ;
AND2    gate16883  (.A(g28664), .B(g23861), .Z(g30199) ) ;
OR2     gate16884  (.A(g27409), .B(g16614), .Z(g28665) ) ;
AND2    gate16885  (.A(g28665), .B(g23862), .Z(g30200) ) ;
OR2     gate16886  (.A(g27410), .B(g16616), .Z(g28667) ) ;
AND2    gate16887  (.A(g28667), .B(g23863), .Z(g30202) ) ;
OR2     gate16888  (.A(g27411), .B(g16617), .Z(g28668) ) ;
AND2    gate16889  (.A(g28668), .B(g23864), .Z(g30203) ) ;
OR2     gate16890  (.A(g27412), .B(g16618), .Z(g28670) ) ;
AND2    gate16891  (.A(g28670), .B(g23868), .Z(g30204) ) ;
OR2     gate16892  (.A(g27413), .B(g16619), .Z(g28671) ) ;
AND2    gate16893  (.A(g28671), .B(g23869), .Z(g30205) ) ;
OR2     gate16894  (.A(g27427), .B(g16633), .Z(g28680) ) ;
AND2    gate16895  (.A(g28680), .B(g23874), .Z(g30207) ) ;
OR2     gate16896  (.A(g27428), .B(g16634), .Z(g28681) ) ;
AND2    gate16897  (.A(g28681), .B(g23875), .Z(g30208) ) ;
OR2     gate16898  (.A(g27430), .B(g16635), .Z(g28682) ) ;
AND2    gate16899  (.A(g28682), .B(g23876), .Z(g30209) ) ;
OR2     gate16900  (.A(g27432), .B(g16636), .Z(g28684) ) ;
AND2    gate16901  (.A(g28684), .B(g23877), .Z(g30210) ) ;
OR2     gate16902  (.A(g27433), .B(g16637), .Z(g28685) ) ;
AND2    gate16903  (.A(g28685), .B(g23878), .Z(g30211) ) ;
OR2     gate16904  (.A(g27434), .B(g16638), .Z(g28687) ) ;
AND2    gate16905  (.A(g28687), .B(g23879), .Z(g30212) ) ;
OR2     gate16906  (.A(g27435), .B(g16639), .Z(g28688) ) ;
AND2    gate16907  (.A(g28688), .B(g23880), .Z(g30213) ) ;
OR2     gate16908  (.A(g27436), .B(g16641), .Z(g28690) ) ;
AND2    gate16909  (.A(g28690), .B(g23881), .Z(g30215) ) ;
OR2     gate16910  (.A(g27437), .B(g16642), .Z(g28691) ) ;
AND2    gate16911  (.A(g28691), .B(g23882), .Z(g30216) ) ;
OR2     gate16912  (.A(g27451), .B(g16666), .Z(g28698) ) ;
AND2    gate16913  (.A(g28698), .B(g23887), .Z(g30219) ) ;
OR2     gate16914  (.A(g27452), .B(g16667), .Z(g28699) ) ;
AND2    gate16915  (.A(g28699), .B(g23888), .Z(g30220) ) ;
OR2     gate16916  (.A(g27454), .B(g16668), .Z(g28700) ) ;
AND2    gate16917  (.A(g28700), .B(g23893), .Z(g30221) ) ;
OR2     gate16918  (.A(g27455), .B(g16669), .Z(g28701) ) ;
AND2    gate16919  (.A(g28701), .B(g23894), .Z(g30222) ) ;
OR2     gate16920  (.A(g27457), .B(g16670), .Z(g28702) ) ;
AND2    gate16921  (.A(g28702), .B(g23895), .Z(g30223) ) ;
OR2     gate16922  (.A(g27459), .B(g16671), .Z(g28704) ) ;
AND2    gate16923  (.A(g28704), .B(g23896), .Z(g30224) ) ;
OR2     gate16924  (.A(g27460), .B(g16672), .Z(g28705) ) ;
AND2    gate16925  (.A(g28705), .B(g23897), .Z(g30225) ) ;
OR2     gate16926  (.A(g27461), .B(g16673), .Z(g28707) ) ;
AND2    gate16927  (.A(g28707), .B(g23898), .Z(g30226) ) ;
OR2     gate16928  (.A(g27462), .B(g16674), .Z(g28708) ) ;
AND2    gate16929  (.A(g28708), .B(g23899), .Z(g30227) ) ;
OR2     gate16930  (.A(g27480), .B(g16700), .Z(g28715) ) ;
AND2    gate16931  (.A(g28715), .B(g23903), .Z(g30228) ) ;
OR2     gate16932  (.A(g27481), .B(g13887), .Z(g28716) ) ;
AND2    gate16933  (.A(g28716), .B(g23904), .Z(g30229) ) ;
OR2     gate16934  (.A(g27482), .B(g16701), .Z(g28717) ) ;
AND2    gate16935  (.A(g28717), .B(g23906), .Z(g30230) ) ;
OR2     gate16936  (.A(g27483), .B(g16702), .Z(g28718) ) ;
AND2    gate16937  (.A(g28718), .B(g23907), .Z(g30231) ) ;
OR2     gate16938  (.A(g27485), .B(g16703), .Z(g28719) ) ;
AND2    gate16939  (.A(g28719), .B(g23912), .Z(g30232) ) ;
OR2     gate16940  (.A(g27486), .B(g16704), .Z(g28720) ) ;
AND2    gate16941  (.A(g28720), .B(g23913), .Z(g30233) ) ;
OR2     gate16942  (.A(g27488), .B(g16705), .Z(g28721) ) ;
AND2    gate16943  (.A(g28721), .B(g23914), .Z(g30234) ) ;
OR2     gate16944  (.A(g27490), .B(g16706), .Z(g28723) ) ;
AND2    gate16945  (.A(g28723), .B(g23915), .Z(g30235) ) ;
OR2     gate16946  (.A(g27491), .B(g16707), .Z(g28724) ) ;
AND2    gate16947  (.A(g28724), .B(g23916), .Z(g30236) ) ;
OR2     gate16948  (.A(g27500), .B(g16729), .Z(g28727) ) ;
AND2    gate16949  (.A(g28727), .B(g23922), .Z(g30238) ) ;
OR2     gate16950  (.A(g27501), .B(g16730), .Z(g28728) ) ;
AND2    gate16951  (.A(g28728), .B(g23923), .Z(g30239) ) ;
OR2     gate16952  (.A(g27502), .B(g16732), .Z(g28729) ) ;
AND2    gate16953  (.A(g28729), .B(g23926), .Z(g30241) ) ;
OR2     gate16954  (.A(g27503), .B(g13912), .Z(g28730) ) ;
AND2    gate16955  (.A(g28730), .B(g23927), .Z(g30242) ) ;
OR2     gate16956  (.A(g27504), .B(g16733), .Z(g28731) ) ;
AND2    gate16957  (.A(g28731), .B(g23929), .Z(g30243) ) ;
OR2     gate16958  (.A(g27505), .B(g16734), .Z(g28732) ) ;
AND2    gate16959  (.A(g28732), .B(g23930), .Z(g30244) ) ;
OR2     gate16960  (.A(g27507), .B(g16735), .Z(g28733) ) ;
AND2    gate16961  (.A(g28733), .B(g23935), .Z(g30245) ) ;
OR2     gate16962  (.A(g27508), .B(g16736), .Z(g28734) ) ;
AND2    gate16963  (.A(g28734), .B(g23936), .Z(g30246) ) ;
OR2     gate16964  (.A(g27510), .B(g16737), .Z(g28735) ) ;
AND2    gate16965  (.A(g28735), .B(g23937), .Z(g30247) ) ;
OR2     gate16966  (.A(g27517), .B(g16758), .Z(g28743) ) ;
AND2    gate16967  (.A(g28743), .B(g23938), .Z(g30248) ) ;
OR2     gate16968  (.A(g27518), .B(g16759), .Z(g28744) ) ;
AND2    gate16969  (.A(g28744), .B(g23939), .Z(g30250) ) ;
OR2     gate16970  (.A(g27519), .B(g16760), .Z(g28745) ) ;
AND2    gate16971  (.A(g28745), .B(g23940), .Z(g30251) ) ;
OR2     gate16972  (.A(g27520), .B(g16762), .Z(g28746) ) ;
AND2    gate16973  (.A(g28746), .B(g23943), .Z(g30253) ) ;
OR2     gate16974  (.A(g27521), .B(g13942), .Z(g28747) ) ;
AND2    gate16975  (.A(g28747), .B(g23944), .Z(g30254) ) ;
OR2     gate16976  (.A(g27522), .B(g16763), .Z(g28748) ) ;
AND2    gate16977  (.A(g28748), .B(g23946), .Z(g30255) ) ;
OR2     gate16978  (.A(g27523), .B(g16764), .Z(g28749) ) ;
AND2    gate16979  (.A(g28749), .B(g23947), .Z(g30256) ) ;
OR2     gate16980  (.A(g27525), .B(g16765), .Z(g28750) ) ;
AND2    gate16981  (.A(g28750), .B(g23952), .Z(g30257) ) ;
OR2     gate16982  (.A(g27526), .B(g16766), .Z(g28751) ) ;
AND2    gate16983  (.A(g28751), .B(g23953), .Z(g30258) ) ;
OR2     gate16984  (.A(g27534), .B(g16802), .Z(g28772) ) ;
AND2    gate16985  (.A(g28772), .B(g23961), .Z(g30261) ) ;
OR2     gate16986  (.A(g27535), .B(g16803), .Z(g28773) ) ;
AND2    gate16987  (.A(g28773), .B(g23962), .Z(g30263) ) ;
OR2     gate16988  (.A(g27536), .B(g16804), .Z(g28774) ) ;
AND2    gate16989  (.A(g28774), .B(g23963), .Z(g30264) ) ;
OR2     gate16990  (.A(g27537), .B(g16806), .Z(g28775) ) ;
AND2    gate16991  (.A(g28775), .B(g23966), .Z(g30266) ) ;
OR2     gate16992  (.A(g27538), .B(g13974), .Z(g28776) ) ;
AND2    gate16993  (.A(g28776), .B(g23967), .Z(g30267) ) ;
OR2     gate16994  (.A(g27539), .B(g16807), .Z(g28777) ) ;
AND2    gate16995  (.A(g28777), .B(g23969), .Z(g30268) ) ;
OR2     gate16996  (.A(g27540), .B(g16808), .Z(g28778) ) ;
AND2    gate16997  (.A(g28778), .B(g23970), .Z(g30269) ) ;
OR2     gate16998  (.A(g27545), .B(g16841), .Z(g28814) ) ;
AND2    gate16999  (.A(g28814), .B(g23982), .Z(g30272) ) ;
OR2     gate17000  (.A(g27546), .B(g16842), .Z(g28815) ) ;
AND2    gate17001  (.A(g28815), .B(g23983), .Z(g30274) ) ;
OR2     gate17002  (.A(g27547), .B(g16843), .Z(g28816) ) ;
AND2    gate17003  (.A(g28816), .B(g23984), .Z(g30275) ) ;
OR2     gate17004  (.A(g27548), .B(g16845), .Z(g28817) ) ;
AND2    gate17005  (.A(g28817), .B(g23987), .Z(g30277) ) ;
OR2     gate17006  (.A(g27549), .B(g13998), .Z(g28818) ) ;
AND2    gate17007  (.A(g28818), .B(g23988), .Z(g30278) ) ;
OR2     gate17008  (.A(g27557), .B(g16869), .Z(g28850) ) ;
AND2    gate17009  (.A(g28850), .B(g23992), .Z(g30281) ) ;
OR2     gate17010  (.A(g27558), .B(g16870), .Z(g28851) ) ;
AND2    gate17011  (.A(g28851), .B(g23993), .Z(g30283) ) ;
OR2     gate17012  (.A(g27559), .B(g16871), .Z(g28852) ) ;
AND2    gate17013  (.A(g28852), .B(g23994), .Z(g30284) ) ;
OR2     gate17014  (.A(g27568), .B(g16885), .Z(g28884) ) ;
AND2    gate17015  (.A(g28884), .B(g24000), .Z(g30289) ) ;
AND3    gate17016  (.A(g29178), .B(g7004), .C(g5297), .Z(g30308) ) ;
AND3    gate17017  (.A(g29182), .B(g7028), .C(g5644), .Z(g30315) ) ;
AND3    gate17018  (.A(g29199), .B(g7097), .C(g6682), .Z(g30316) ) ;
AND2    gate17019  (.A(g21358), .B(g29385), .Z(g30564) ) ;
NOR2    gate17020  (.A(g7995), .B(g24732), .Z(g26247) ) ;
AND2    gate17021  (.A(g26247), .B(g29507), .Z(g30566) ) ;
AND2    gate17022  (.A(g18898), .B(g29800), .Z(g30576) ) ;
NOR2    gate17023  (.A(g8033), .B(g24732), .Z(g26267) ) ;
AND2    gate17024  (.A(g26267), .B(g29679), .Z(g30577) ) ;
NAND2   gate17025  (.A(g24383), .B(g28109), .Z(g29355) ) ;
AND2    gate17026  (.A(g19666), .B(g29355), .Z(g30583) ) ;
AND2    gate17027  (.A(g18898), .B(g29811), .Z(g30589) ) ;
AND2    gate17028  (.A(g18911), .B(g29812), .Z(g30590) ) ;
OR2     gate17029  (.A(g28624), .B(g27664), .Z(g30270) ) ;
AND2    gate17030  (.A(g30270), .B(g18929), .Z(g30592) ) ;
AND2    gate17031  (.A(g18898), .B(g29846), .Z(g30594) ) ;
AND2    gate17032  (.A(g18911), .B(g29847), .Z(g30595) ) ;
OR2     gate17033  (.A(g28637), .B(g27668), .Z(g30279) ) ;
AND2    gate17034  (.A(g30279), .B(g18947), .Z(g30596) ) ;
AND2    gate17035  (.A(g18898), .B(g29862), .Z(g30598) ) ;
AND2    gate17036  (.A(g18911), .B(g29863), .Z(g30599) ) ;
OR2     gate17037  (.A(g28653), .B(g27677), .Z(g30287) ) ;
AND2    gate17038  (.A(g30287), .B(g18975), .Z(g30600) ) ;
AND2    gate17039  (.A(g18911), .B(g29878), .Z(g30604) ) ;
OR2     gate17040  (.A(g28672), .B(g27685), .Z(g30291) ) ;
AND2    gate17041  (.A(g30291), .B(g18989), .Z(g30607) ) ;
NOR2    gate17042  (.A(g8458), .B(g24825), .Z(g26338) ) ;
AND2    gate17043  (.A(g26338), .B(g29597), .Z(g30612) ) ;
NOR2    gate17044  (.A(g7528), .B(g28167), .Z(g29359) ) ;
AND2    gate17045  (.A(g11330), .B(g29359), .Z(g30670) ) ;
OR2     gate17046  (.A(g28812), .B(g14453), .Z(g29319) ) ;
AND2    gate17047  (.A(g29319), .B(g22317), .Z(g30671) ) ;
NOR2    gate17048  (.A(g8522), .B(g24825), .Z(g26346) ) ;
AND2    gate17049  (.A(g26346), .B(g29778), .Z(g30730) ) ;
NOR2    gate17050  (.A(g7553), .B(g28174), .Z(g29361) ) ;
AND2    gate17051  (.A(g11374), .B(g29361), .Z(g30731) ) ;
NOR2    gate17052  (.A(g6875), .B(g28458), .Z(g29873) ) ;
AND2    gate17053  (.A(g29873), .B(g20887), .Z(g30914) ) ;
NOR2    gate17054  (.A(g3288), .B(g28458), .Z(g29886) ) ;
AND2    gate17055  (.A(g29886), .B(g24778), .Z(g30915) ) ;
AND2    gate17056  (.A(g8681), .B(g29707), .Z(g30918) ) ;
NOR2    gate17057  (.A(g6895), .B(g28458), .Z(g29898) ) ;
AND2    gate17058  (.A(g29898), .B(g23286), .Z(g30919) ) ;
NOR2    gate17059  (.A(g6905), .B(g28471), .Z(g29889) ) ;
AND2    gate17060  (.A(g29889), .B(g21024), .Z(g30920) ) ;
NOR2    gate17061  (.A(g3639), .B(g28471), .Z(g29900) ) ;
AND2    gate17062  (.A(g29900), .B(g24789), .Z(g30921) ) ;
NOR2    gate17063  (.A(g6918), .B(g28471), .Z(g29908) ) ;
AND2    gate17064  (.A(g29908), .B(g23309), .Z(g30925) ) ;
NOR2    gate17065  (.A(g6928), .B(g28484), .Z(g29903) ) ;
AND2    gate17066  (.A(g29903), .B(g21163), .Z(g30926) ) ;
NOR2    gate17067  (.A(g3990), .B(g28484), .Z(g29910) ) ;
AND2    gate17068  (.A(g29910), .B(g24795), .Z(g30927) ) ;
NOR2    gate17069  (.A(g6941), .B(g28484), .Z(g29915) ) ;
AND2    gate17070  (.A(g29915), .B(g23342), .Z(g30930) ) ;
AND2    gate17071  (.A(g8808), .B(g29745), .Z(g30935) ) ;
AND2    gate17072  (.A(g8830), .B(g29916), .Z(g30936) ) ;
AND2    gate17073  (.A(g8895), .B(g29933), .Z(g30982) ) ;
OR2     gate17074  (.A(g28108), .B(g28112), .Z(g29476) ) ;
AND2    gate17075  (.A(g29476), .B(g22758), .Z(g31015) ) ;
OR2     gate17076  (.A(g28111), .B(g22160), .Z(g29478) ) ;
AND2    gate17077  (.A(g29478), .B(g22840), .Z(g31016) ) ;
OR2     gate17078  (.A(g28113), .B(g28116), .Z(g29479) ) ;
AND2    gate17079  (.A(g29479), .B(g22841), .Z(g31017) ) ;
OR2     gate17080  (.A(g28115), .B(g22172), .Z(g29480) ) ;
AND2    gate17081  (.A(g29480), .B(g22855), .Z(g31018) ) ;
OR2     gate17082  (.A(g28117), .B(g28125), .Z(g29481) ) ;
AND2    gate17083  (.A(g29481), .B(g22856), .Z(g31019) ) ;
NAND2   gate17084  (.A(g22405), .B(g24631), .Z(g26025) ) ;
OR2     gate17085  (.A(g25801), .B(g28130), .Z(g29483) ) ;
AND2    gate17086  (.A(g29483), .B(g22865), .Z(g31066) ) ;
OR2     gate17087  (.A(g28124), .B(g22191), .Z(g29484) ) ;
AND2    gate17088  (.A(g29484), .B(g22868), .Z(g31067) ) ;
OR2     gate17089  (.A(g28237), .B(g27247), .Z(g29793) ) ;
AND2    gate17090  (.A(g29793), .B(g14150), .Z(g31069) ) ;
NAND2   gate17091  (.A(g24631), .B(g23956), .Z(g25985) ) ;
OR2     gate17092  (.A(g25815), .B(g28133), .Z(g29487) ) ;
AND2    gate17093  (.A(g29487), .B(g22882), .Z(g31115) ) ;
OR2     gate17094  (.A(g25832), .B(g28136), .Z(g29490) ) ;
AND2    gate17095  (.A(g29490), .B(g22906), .Z(g31118) ) ;
AND2    gate17096  (.A(g1700), .B(g29976), .Z(g31120) ) ;
NAND2   gate17097  (.A(II15003), .B(II15004), .Z(g12144) ) ;
AND2    gate17098  (.A(g12144), .B(g29993), .Z(g31122) ) ;
AND2    gate17099  (.A(g1834), .B(g29994), .Z(g31123) ) ;
AND2    gate17100  (.A(g2259), .B(g29997), .Z(g31124) ) ;
OR2     gate17101  (.A(g28139), .B(g25871), .Z(g29502) ) ;
AND2    gate17102  (.A(g29502), .B(g22973), .Z(g31125) ) ;
NAND2   gate17103  (.A(II15042), .B(II15043), .Z(g12187) ) ;
AND2    gate17104  (.A(g12187), .B(g30016), .Z(g31128) ) ;
AND2    gate17105  (.A(g1968), .B(g30017), .Z(g31129) ) ;
NAND2   gate17106  (.A(II15052), .B(II15053), .Z(g12191) ) ;
AND2    gate17107  (.A(g12191), .B(g30019), .Z(g31130) ) ;
AND2    gate17108  (.A(g2393), .B(g30020), .Z(g31131) ) ;
OR2     gate17109  (.A(g28143), .B(g25875), .Z(g29504) ) ;
AND2    gate17110  (.A(g29504), .B(g22987), .Z(g31132) ) ;
NAND2   gate17111  (.A(II15079), .B(II15080), .Z(g12221) ) ;
AND2    gate17112  (.A(g12221), .B(g30036), .Z(g31139) ) ;
AND2    gate17113  (.A(g2102), .B(g30037), .Z(g31140) ) ;
NAND2   gate17114  (.A(II15088), .B(II15089), .Z(g12224) ) ;
AND2    gate17115  (.A(g12224), .B(g30038), .Z(g31141) ) ;
AND2    gate17116  (.A(g2527), .B(g30039), .Z(g31142) ) ;
OR2     gate17117  (.A(g28148), .B(g25880), .Z(g29506) ) ;
AND2    gate17118  (.A(g29506), .B(g22999), .Z(g31143) ) ;
AND2    gate17119  (.A(g9970), .B(g30052), .Z(g31145) ) ;
NAND2   gate17120  (.A(II15122), .B(II15123), .Z(g12285) ) ;
AND2    gate17121  (.A(g12285), .B(g30053), .Z(g31146) ) ;
NAND2   gate17122  (.A(II15129), .B(II15130), .Z(g12286) ) ;
AND2    gate17123  (.A(g12286), .B(g30054), .Z(g31147) ) ;
AND2    gate17124  (.A(g2661), .B(g30055), .Z(g31148) ) ;
OR2     gate17125  (.A(g28152), .B(g27041), .Z(g29508) ) ;
AND2    gate17126  (.A(g29508), .B(g23021), .Z(g31149) ) ;
AND2    gate17127  (.A(g1682), .B(g30063), .Z(g31150) ) ;
AND2    gate17128  (.A(g10037), .B(g30065), .Z(g31151) ) ;
AND2    gate17129  (.A(g10039), .B(g30067), .Z(g31152) ) ;
NAND2   gate17130  (.A(II15175), .B(II15176), .Z(g12336) ) ;
AND2    gate17131  (.A(g12336), .B(g30068), .Z(g31153) ) ;
AND2    gate17132  (.A(g1816), .B(g30074), .Z(g31166) ) ;
AND2    gate17133  (.A(g10080), .B(g30076), .Z(g31167) ) ;
AND2    gate17134  (.A(g2241), .B(g30077), .Z(g31168) ) ;
AND2    gate17135  (.A(g10083), .B(g30079), .Z(g31169) ) ;
NOR2    gate17136  (.A(g7004), .B(g28982), .Z(g30240) ) ;
AND2    gate17137  (.A(g30240), .B(g20682), .Z(g31182) ) ;
NOR2    gate17138  (.A(g5297), .B(g28982), .Z(g30249) ) ;
AND2    gate17139  (.A(g30249), .B(g25174), .Z(g31183) ) ;
AND2    gate17140  (.A(g1950), .B(g30085), .Z(g31184) ) ;
AND2    gate17141  (.A(g10114), .B(g30087), .Z(g31185) ) ;
AND2    gate17142  (.A(g2375), .B(g30088), .Z(g31186) ) ;
AND2    gate17143  (.A(g10118), .B(g30090), .Z(g31187) ) ;
AND2    gate17144  (.A(g20028), .B(g29653), .Z(g31188) ) ;
NOR2    gate17145  (.A(g7018), .B(g28982), .Z(g30260) ) ;
AND2    gate17146  (.A(g30260), .B(g23890), .Z(g31206) ) ;
NOR2    gate17147  (.A(g7028), .B(g29008), .Z(g30252) ) ;
AND2    gate17148  (.A(g30252), .B(g20739), .Z(g31207) ) ;
NOR2    gate17149  (.A(g5644), .B(g29008), .Z(g30262) ) ;
AND2    gate17150  (.A(g30262), .B(g25188), .Z(g31208) ) ;
AND2    gate17151  (.A(g2084), .B(g30097), .Z(g31209) ) ;
AND2    gate17152  (.A(g2509), .B(g30100), .Z(g31210) ) ;
AND2    gate17153  (.A(g10156), .B(g30102), .Z(g31211) ) ;
AND2    gate17154  (.A(g20028), .B(g29669), .Z(g31212) ) ;
NOR2    gate17155  (.A(g7041), .B(g29008), .Z(g30271) ) ;
AND2    gate17156  (.A(g30271), .B(g23909), .Z(g31218) ) ;
NOR2    gate17157  (.A(g7051), .B(g29036), .Z(g30265) ) ;
AND2    gate17158  (.A(g30265), .B(g20875), .Z(g31219) ) ;
NOR2    gate17159  (.A(g5990), .B(g29036), .Z(g30273) ) ;
AND2    gate17160  (.A(g30273), .B(g25202), .Z(g31220) ) ;
AND2    gate17161  (.A(g2643), .B(g30113), .Z(g31222) ) ;
AND2    gate17162  (.A(g20028), .B(g29689), .Z(g31223) ) ;
NOR2    gate17163  (.A(g7064), .B(g29036), .Z(g30280) ) ;
AND2    gate17164  (.A(g30280), .B(g23932), .Z(g31224) ) ;
NOR2    gate17165  (.A(g7074), .B(g29073), .Z(g30276) ) ;
AND2    gate17166  (.A(g30276), .B(g21012), .Z(g31225) ) ;
NOR2    gate17167  (.A(g6336), .B(g29073), .Z(g30282) ) ;
AND2    gate17168  (.A(g30282), .B(g25218), .Z(g31226) ) ;
AND2    gate17169  (.A(g20028), .B(g29713), .Z(g31228) ) ;
NOR2    gate17170  (.A(g7087), .B(g29073), .Z(g30288) ) ;
AND2    gate17171  (.A(g30288), .B(g23949), .Z(g31229) ) ;
NOR2    gate17172  (.A(g7097), .B(g29110), .Z(g30285) ) ;
AND2    gate17173  (.A(g30285), .B(g20751), .Z(g31230) ) ;
NOR2    gate17174  (.A(g6682), .B(g29110), .Z(g30290) ) ;
AND2    gate17175  (.A(g30290), .B(g25239), .Z(g31231) ) ;
NOR2    gate17176  (.A(g7110), .B(g29110), .Z(g30294) ) ;
AND2    gate17177  (.A(g30294), .B(g23972), .Z(g31232) ) ;
OR2     gate17178  (.A(g13738), .B(g28439), .Z(g29366) ) ;
AND2    gate17179  (.A(g29366), .B(g25325), .Z(g31237) ) ;
OR2     gate17180  (.A(g28182), .B(g27099), .Z(g29583) ) ;
AND2    gate17181  (.A(g29583), .B(g20053), .Z(g31238) ) ;
NOR2    gate17182  (.A(g2988), .B(g12228), .Z(g14793) ) ;
AND2    gate17183  (.A(g14793), .B(g30206), .Z(g31240) ) ;
OR2     gate17184  (.A(g13832), .B(g28453), .Z(g29373) ) ;
AND2    gate17185  (.A(g29373), .B(g25409), .Z(g31242) ) ;
OR2     gate17186  (.A(g28192), .B(g27145), .Z(g29643) ) ;
AND2    gate17187  (.A(g29643), .B(g20101), .Z(g31252) ) ;
NOR2    gate17188  (.A(g12821), .B(g2988), .Z(g14754) ) ;
AND2    gate17189  (.A(g14754), .B(g30259), .Z(g31261) ) ;
NOR2    gate17190  (.A(g28739), .B(g14537), .Z(g30129) ) ;
AND2    gate17191  (.A(g30129), .B(g27742), .Z(g31266) ) ;
OR2     gate17192  (.A(g28197), .B(g10873), .Z(g29692) ) ;
AND2    gate17193  (.A(g29692), .B(g23282), .Z(g31270) ) ;
OR2     gate17194  (.A(g28198), .B(g27208), .Z(g29706) ) ;
AND2    gate17195  (.A(g29706), .B(g23300), .Z(g31271) ) ;
NOR2    gate17196  (.A(g28739), .B(g7252), .Z(g30117) ) ;
AND2    gate17197  (.A(g30117), .B(g27742), .Z(g31272) ) ;
NOR2    gate17198  (.A(g28761), .B(g14566), .Z(g30143) ) ;
AND2    gate17199  (.A(g30143), .B(g27779), .Z(g31273) ) ;
NOR2    gate17200  (.A(g28768), .B(g14567), .Z(g30147) ) ;
AND2    gate17201  (.A(g30147), .B(g27800), .Z(g31275) ) ;
OR2     gate17202  (.A(g28199), .B(g15856), .Z(g29716) ) ;
AND2    gate17203  (.A(g29716), .B(g23302), .Z(g31278) ) ;
OR2     gate17204  (.A(g28200), .B(g10883), .Z(g29717) ) ;
AND2    gate17205  (.A(g29717), .B(g23305), .Z(g31280) ) ;
NOR2    gate17206  (.A(g28739), .B(g7268), .Z(g30106) ) ;
AND2    gate17207  (.A(g30106), .B(g27742), .Z(g31281) ) ;
NOR2    gate17208  (.A(g28761), .B(g7275), .Z(g30130) ) ;
AND2    gate17209  (.A(g30130), .B(g27779), .Z(g31282) ) ;
NOR2    gate17210  (.A(g28789), .B(g14587), .Z(g30156) ) ;
AND2    gate17211  (.A(g30156), .B(g27837), .Z(g31283) ) ;
NOR2    gate17212  (.A(g28768), .B(g7280), .Z(g30134) ) ;
AND2    gate17213  (.A(g30134), .B(g27800), .Z(g31285) ) ;
NOR2    gate17214  (.A(g28799), .B(g14589), .Z(g30159) ) ;
AND2    gate17215  (.A(g30159), .B(g27858), .Z(g31286) ) ;
OR2     gate17216  (.A(g28201), .B(g15872), .Z(g29734) ) ;
AND2    gate17217  (.A(g29734), .B(g23335), .Z(g31290) ) ;
OR2     gate17218  (.A(g28202), .B(g10898), .Z(g29735) ) ;
AND2    gate17219  (.A(g29735), .B(g23338), .Z(g31292) ) ;
NOR2    gate17220  (.A(g28761), .B(g7315), .Z(g30119) ) ;
AND2    gate17221  (.A(g30119), .B(g27779), .Z(g31296) ) ;
NOR2    gate17222  (.A(g28789), .B(g7322), .Z(g30144) ) ;
AND2    gate17223  (.A(g30144), .B(g27837), .Z(g31297) ) ;
NOR2    gate17224  (.A(g28833), .B(g14613), .Z(g30169) ) ;
AND2    gate17225  (.A(g30169), .B(g27886), .Z(g31298) ) ;
NOR2    gate17226  (.A(g28768), .B(g7328), .Z(g30123) ) ;
AND2    gate17227  (.A(g30123), .B(g27800), .Z(g31299) ) ;
NOR2    gate17228  (.A(g28799), .B(g7335), .Z(g30148) ) ;
AND2    gate17229  (.A(g30148), .B(g27858), .Z(g31300) ) ;
NOR2    gate17230  (.A(g28846), .B(g14615), .Z(g30170) ) ;
AND2    gate17231  (.A(g30170), .B(g27907), .Z(g31301) ) ;
OR2     gate17232  (.A(g28205), .B(g15883), .Z(g29741) ) ;
AND2    gate17233  (.A(g29741), .B(g23354), .Z(g31305) ) ;
NOR2    gate17234  (.A(g28789), .B(g7362), .Z(g30132) ) ;
AND2    gate17235  (.A(g30132), .B(g27837), .Z(g31309) ) ;
NOR2    gate17236  (.A(g28833), .B(g7369), .Z(g30157) ) ;
AND2    gate17237  (.A(g30157), .B(g27886), .Z(g31310) ) ;
NOR2    gate17238  (.A(g28799), .B(g7380), .Z(g30136) ) ;
AND2    gate17239  (.A(g30136), .B(g27858), .Z(g31312) ) ;
NOR2    gate17240  (.A(g28846), .B(g7387), .Z(g30160) ) ;
AND2    gate17241  (.A(g30160), .B(g27907), .Z(g31313) ) ;
NOR2    gate17242  (.A(g28880), .B(g14644), .Z(g30183) ) ;
AND2    gate17243  (.A(g30183), .B(g27937), .Z(g31314) ) ;
NOR2    gate17244  (.A(g28833), .B(g7411), .Z(g30146) ) ;
AND2    gate17245  (.A(g30146), .B(g27886), .Z(g31321) ) ;
NOR2    gate17246  (.A(g28846), .B(g7424), .Z(g30150) ) ;
AND2    gate17247  (.A(g30150), .B(g27907), .Z(g31323) ) ;
NOR2    gate17248  (.A(g28880), .B(g7431), .Z(g30171) ) ;
AND2    gate17249  (.A(g30171), .B(g27937), .Z(g31324) ) ;
OR2     gate17250  (.A(g28210), .B(g28214), .Z(g29748) ) ;
AND2    gate17251  (.A(g29748), .B(g23390), .Z(g31374) ) ;
OR3     gate17252  (.A(g21326), .B(g21340), .C(II24117), .Z(g24952) ) ;
NOR2    gate17253  (.A(g28880), .B(g7462), .Z(g30162) ) ;
AND2    gate17254  (.A(g30162), .B(g27937), .Z(g31467) ) ;
OR2     gate17255  (.A(g28213), .B(g22720), .Z(g29753) ) ;
AND2    gate17256  (.A(g29753), .B(g23398), .Z(g31470) ) ;
OR2     gate17257  (.A(g28215), .B(g28218), .Z(g29754) ) ;
AND2    gate17258  (.A(g29754), .B(g23399), .Z(g31471) ) ;
OR2     gate17259  (.A(g22717), .B(g28223), .Z(g29756) ) ;
AND2    gate17260  (.A(g29756), .B(g23406), .Z(g31475) ) ;
OR2     gate17261  (.A(g28217), .B(g22762), .Z(g29763) ) ;
AND2    gate17262  (.A(g29763), .B(g23409), .Z(g31477) ) ;
OR2     gate17263  (.A(g28219), .B(g28226), .Z(g29764) ) ;
AND2    gate17264  (.A(g29764), .B(g23410), .Z(g31478) ) ;
AND2    gate17265  (.A(g1644), .B(g30296), .Z(g31480) ) ;
OR2     gate17266  (.A(g22760), .B(g28229), .Z(g29768) ) ;
AND2    gate17267  (.A(g29768), .B(g23417), .Z(g31481) ) ;
OR2     gate17268  (.A(g25966), .B(g28232), .Z(g29775) ) ;
AND2    gate17269  (.A(g29775), .B(g23418), .Z(g31484) ) ;
OR2     gate17270  (.A(g28225), .B(g22846), .Z(g29776) ) ;
AND2    gate17271  (.A(g29776), .B(g23421), .Z(g31485) ) ;
OR2     gate17272  (.A(g28227), .B(g28234), .Z(g29777) ) ;
AND2    gate17273  (.A(g29777), .B(g23422), .Z(g31486) ) ;
AND2    gate17274  (.A(g1779), .B(g30302), .Z(g31488) ) ;
AND2    gate17275  (.A(g2204), .B(g30305), .Z(g31489) ) ;
OR2     gate17276  (.A(g22843), .B(g28240), .Z(g29786) ) ;
AND2    gate17277  (.A(g29786), .B(g23429), .Z(g31490) ) ;
OR2     gate17278  (.A(g25975), .B(g28242), .Z(g29790) ) ;
AND2    gate17279  (.A(g29790), .B(g23431), .Z(g31492) ) ;
OR2     gate17280  (.A(g28233), .B(g22859), .Z(g29791) ) ;
AND2    gate17281  (.A(g29791), .B(g23434), .Z(g31493) ) ;
OR2     gate17282  (.A(g28235), .B(g28244), .Z(g29792) ) ;
AND2    gate17283  (.A(g29792), .B(g23435), .Z(g31494) ) ;
AND2    gate17284  (.A(g1913), .B(g30309), .Z(g31495) ) ;
AND2    gate17285  (.A(g2338), .B(g30312), .Z(g31496) ) ;
AND2    gate17286  (.A(g20041), .B(g29930), .Z(g31497) ) ;
OR2     gate17287  (.A(g25987), .B(g28251), .Z(g29801) ) ;
AND2    gate17288  (.A(g29801), .B(g23446), .Z(g31499) ) ;
OR2     gate17289  (.A(g28243), .B(g22871), .Z(g29802) ) ;
AND2    gate17290  (.A(g29802), .B(g23449), .Z(g31500) ) ;
AND2    gate17291  (.A(g2047), .B(g29310), .Z(g31501) ) ;
AND2    gate17292  (.A(g2472), .B(g29311), .Z(g31502) ) ;
AND2    gate17293  (.A(g20041), .B(g29945), .Z(g31503) ) ;
NOR2    gate17294  (.A(g28585), .B(g28599), .Z(g29370) ) ;
AND2    gate17295  (.A(g29370), .B(g10553), .Z(g31504) ) ;
AND2    gate17296  (.A(g30195), .B(g24379), .Z(g31505) ) ;
OR2     gate17297  (.A(g26020), .B(g28261), .Z(g29813) ) ;
AND2    gate17298  (.A(g29813), .B(g23459), .Z(g31508) ) ;
AND2    gate17299  (.A(g2606), .B(g29318), .Z(g31513) ) ;
AND2    gate17300  (.A(g20041), .B(g29956), .Z(g31514) ) ;
OR2     gate17301  (.A(g28260), .B(g26077), .Z(g29848) ) ;
AND2    gate17302  (.A(g29848), .B(g23476), .Z(g31516) ) ;
OR2     gate17303  (.A(g26049), .B(g28273), .Z(g29849) ) ;
AND2    gate17304  (.A(g29849), .B(g23482), .Z(g31517) ) ;
AND2    gate17305  (.A(g20041), .B(g29970), .Z(g31518) ) ;
OR2     gate17306  (.A(g28272), .B(g26086), .Z(g29864) ) ;
AND2    gate17307  (.A(g29864), .B(g23490), .Z(g31519) ) ;
OR2     gate17308  (.A(g28289), .B(g26096), .Z(g29879) ) ;
AND2    gate17309  (.A(g29879), .B(g23507), .Z(g31520) ) ;
AND2    gate17310  (.A(g7528), .B(g29333), .Z(g31523) ) ;
AND2    gate17311  (.A(g29897), .B(g20593), .Z(g31524) ) ;
OR2     gate17312  (.A(g28300), .B(g26120), .Z(g29892) ) ;
AND2    gate17313  (.A(g29892), .B(g23526), .Z(g31525) ) ;
NOR2    gate17314  (.A(g1036), .B(g19699), .Z(g22521) ) ;
AND2    gate17315  (.A(g22521), .B(g29342), .Z(g31526) ) ;
AND2    gate17316  (.A(g7553), .B(g29343), .Z(g31527) ) ;
OR2     gate17317  (.A(g28312), .B(g26146), .Z(g29904) ) ;
AND2    gate17318  (.A(g29904), .B(g23548), .Z(g31540) ) ;
NOR2    gate17319  (.A(g1379), .B(g19720), .Z(g22536) ) ;
AND2    gate17320  (.A(g22536), .B(g29348), .Z(g31541) ) ;
OR2     gate17321  (.A(g28813), .B(g27820), .Z(g29325) ) ;
AND2    gate17322  (.A(g29325), .B(g13062), .Z(g31654) ) ;
OR2     gate17323  (.A(g28454), .B(g11366), .Z(g30081) ) ;
AND2    gate17324  (.A(g30081), .B(g23886), .Z(g31707) ) ;
OR2     gate17325  (.A(g28466), .B(g16699), .Z(g30092) ) ;
AND2    gate17326  (.A(g30092), .B(g23902), .Z(g31744) ) ;
OR2     gate17327  (.A(g28467), .B(g11397), .Z(g30093) ) ;
AND2    gate17328  (.A(g30093), .B(g23905), .Z(g31746) ) ;
OR2     gate17329  (.A(g28477), .B(g16731), .Z(g30103) ) ;
AND2    gate17330  (.A(g30103), .B(g23925), .Z(g31750) ) ;
OR2     gate17331  (.A(g28478), .B(g11427), .Z(g30104) ) ;
AND2    gate17332  (.A(g30104), .B(g23928), .Z(g31752) ) ;
OR2     gate17333  (.A(g28488), .B(g16761), .Z(g30114) ) ;
AND2    gate17334  (.A(g30114), .B(g23942), .Z(g31756) ) ;
OR2     gate17335  (.A(g28489), .B(g11449), .Z(g30115) ) ;
AND2    gate17336  (.A(g30115), .B(g23945), .Z(g31758) ) ;
AND2    gate17337  (.A(g21291), .B(g29385), .Z(g31759) ) ;
OR2     gate17338  (.A(g28494), .B(g16805), .Z(g30127) ) ;
AND2    gate17339  (.A(g30127), .B(g23965), .Z(g31763) ) ;
OR2     gate17340  (.A(g28495), .B(g11497), .Z(g30128) ) ;
AND2    gate17341  (.A(g30128), .B(g23968), .Z(g31765) ) ;
OR2     gate17342  (.A(g28499), .B(g16844), .Z(g30141) ) ;
AND2    gate17343  (.A(g30141), .B(g23986), .Z(g31769) ) ;
AND2    gate17344  (.A(g21329), .B(g29385), .Z(g31776) ) ;
AND2    gate17345  (.A(g21343), .B(g29385), .Z(g31777) ) ;
AND2    gate17346  (.A(g21369), .B(g29385), .Z(g31778) ) ;
OR2     gate17347  (.A(g23381), .B(g28523), .Z(g30163) ) ;
AND2    gate17348  (.A(g30163), .B(g23999), .Z(g31780) ) ;
OR2     gate17349  (.A(g23392), .B(g28531), .Z(g30176) ) ;
AND2    gate17350  (.A(g30176), .B(g24003), .Z(g31784) ) ;
OR2     gate17351  (.A(g23401), .B(g28543), .Z(g30189) ) ;
AND2    gate17352  (.A(g30189), .B(g24010), .Z(g31786) ) ;
AND2    gate17353  (.A(g21281), .B(g29385), .Z(g31787) ) ;
AND2    gate17354  (.A(g21352), .B(g29385), .Z(g31788) ) ;
OR2     gate17355  (.A(g23412), .B(g28557), .Z(g30201) ) ;
AND2    gate17356  (.A(g30201), .B(g24013), .Z(g31789) ) ;
AND2    gate17357  (.A(g21299), .B(g29385), .Z(g31790) ) ;
OR2     gate17358  (.A(g23424), .B(g28572), .Z(g30214) ) ;
AND2    gate17359  (.A(g30214), .B(g24017), .Z(g31792) ) ;
AND2    gate17360  (.A(g939), .B(g30735), .Z(g31933) ) ;
OR2     gate17361  (.A(g29937), .B(g28573), .Z(g31670) ) ;
AND2    gate17362  (.A(g31670), .B(g18827), .Z(g31934) ) ;
AND2    gate17363  (.A(g31213), .B(g24005), .Z(g31936) ) ;
AND2    gate17364  (.A(g943), .B(g30735), .Z(g31940) ) ;
AND2    gate17365  (.A(g1283), .B(g30825), .Z(g31941) ) ;
AND2    gate17366  (.A(g4717), .B(g30614), .Z(g31943) ) ;
OR2     gate17367  (.A(g29959), .B(g29973), .Z(g31745) ) ;
AND2    gate17368  (.A(g31745), .B(g22146), .Z(g31944) ) ;
AND2    gate17369  (.A(g30670), .B(g18884), .Z(g31948) ) ;
AND2    gate17370  (.A(g1287), .B(g30825), .Z(g31949) ) ;
AND2    gate17371  (.A(g4907), .B(g30673), .Z(g31959) ) ;
OR2     gate17372  (.A(g29974), .B(g29988), .Z(g31749) ) ;
AND2    gate17373  (.A(g31749), .B(g22153), .Z(g31960) ) ;
OR2     gate17374  (.A(g29975), .B(g29990), .Z(g31751) ) ;
AND2    gate17375  (.A(g31751), .B(g22154), .Z(g31961) ) ;
AND2    gate17376  (.A(g8033), .B(g31013), .Z(g31962) ) ;
AND2    gate17377  (.A(g30731), .B(g18895), .Z(g31963) ) ;
OR2     gate17378  (.A(g29989), .B(g30006), .Z(g31754) ) ;
AND2    gate17379  (.A(g31754), .B(g22166), .Z(g31966) ) ;
OR2     gate17380  (.A(g29991), .B(g30008), .Z(g31755) ) ;
AND2    gate17381  (.A(g31755), .B(g22167), .Z(g31967) ) ;
OR2     gate17382  (.A(g29992), .B(g30010), .Z(g31757) ) ;
AND2    gate17383  (.A(g31757), .B(g22168), .Z(g31968) ) ;
AND2    gate17384  (.A(g31189), .B(g22139), .Z(g31969) ) ;
OR2     gate17385  (.A(g30007), .B(g30027), .Z(g31760) ) ;
AND2    gate17386  (.A(g31760), .B(g22176), .Z(g31974) ) ;
OR2     gate17387  (.A(g30009), .B(g30028), .Z(g31761) ) ;
AND2    gate17388  (.A(g31761), .B(g22177), .Z(g31975) ) ;
OR2     gate17389  (.A(g30011), .B(g30030), .Z(g31762) ) ;
AND2    gate17390  (.A(g31762), .B(g22178), .Z(g31976) ) ;
OR2     gate17391  (.A(g30015), .B(g30032), .Z(g31764) ) ;
AND2    gate17392  (.A(g31764), .B(g22179), .Z(g31977) ) ;
AND2    gate17393  (.A(g4722), .B(g30614), .Z(g31985) ) ;
OR2     gate17394  (.A(g30029), .B(g30042), .Z(g31766) ) ;
AND2    gate17395  (.A(g31766), .B(g22197), .Z(g31986) ) ;
OR2     gate17396  (.A(g30031), .B(g30043), .Z(g31767) ) ;
AND2    gate17397  (.A(g31767), .B(g22198), .Z(g31987) ) ;
OR2     gate17398  (.A(g30033), .B(g30045), .Z(g31768) ) ;
AND2    gate17399  (.A(g31768), .B(g22199), .Z(g31988) ) ;
OR2     gate17400  (.A(g30034), .B(g30047), .Z(g31770) ) ;
AND2    gate17401  (.A(g31770), .B(g22200), .Z(g31989) ) ;
OR2     gate17402  (.A(g30035), .B(g28654), .Z(g31772) ) ;
AND2    gate17403  (.A(g31772), .B(g18945), .Z(g31990) ) ;
AND2    gate17404  (.A(g4912), .B(g30673), .Z(g31991) ) ;
OR2     gate17405  (.A(g30044), .B(g30056), .Z(g31773) ) ;
AND2    gate17406  (.A(g31773), .B(g22213), .Z(g31992) ) ;
OR2     gate17407  (.A(g30046), .B(g30057), .Z(g31774) ) ;
AND2    gate17408  (.A(g31774), .B(g22214), .Z(g31993) ) ;
OR2     gate17409  (.A(g30048), .B(g30059), .Z(g31775) ) ;
AND2    gate17410  (.A(g31775), .B(g22215), .Z(g31994) ) ;
AND2    gate17411  (.A(g28274), .B(g30569), .Z(g31995) ) ;
OR2     gate17412  (.A(g30050), .B(g28673), .Z(g31779) ) ;
AND2    gate17413  (.A(g31779), .B(g18979), .Z(g31996) ) ;
OR2     gate17414  (.A(g30058), .B(g30069), .Z(g31781) ) ;
AND2    gate17415  (.A(g31781), .B(g22223), .Z(g32008) ) ;
OR2     gate17416  (.A(g30060), .B(g30070), .Z(g31782) ) ;
AND2    gate17417  (.A(g31782), .B(g22224), .Z(g32009) ) ;
OR2     gate17418  (.A(g30071), .B(g30082), .Z(g31785) ) ;
AND2    gate17419  (.A(g31785), .B(g22303), .Z(g32010) ) ;
AND2    gate17420  (.A(g8287), .B(g31134), .Z(g32011) ) ;
AND2    gate17421  (.A(g8297), .B(g31233), .Z(g32012) ) ;
AND2    gate17422  (.A(g8673), .B(g30614), .Z(g32013) ) ;
AND2    gate17423  (.A(g8715), .B(g30673), .Z(g32014) ) ;
AND2    gate17424  (.A(g8522), .B(g31138), .Z(g32016) ) ;
AND2    gate17425  (.A(g4146), .B(g30937), .Z(g32018) ) ;
OR2     gate17426  (.A(g30173), .B(g14571), .Z(g30579) ) ;
AND2    gate17427  (.A(g30579), .B(g22358), .Z(g32019) ) ;
AND2    gate17428  (.A(g4157), .B(g30937), .Z(g32020) ) ;
AND2    gate17429  (.A(g30569), .B(g29339), .Z(g32028) ) ;
NOR2    gate17430  (.A(g4785), .B(g29697), .Z(g31318) ) ;
AND2    gate17431  (.A(g31318), .B(g16482), .Z(g32029) ) ;
AND2    gate17432  (.A(g4172), .B(g30937), .Z(g32030) ) ;
NOR2    gate17433  (.A(g8796), .B(g29697), .Z(g31372) ) ;
AND2    gate17434  (.A(g31372), .B(g13464), .Z(g32031) ) ;
NOR2    gate17435  (.A(g4975), .B(g29725), .Z(g31373) ) ;
AND2    gate17436  (.A(g31373), .B(g16515), .Z(g32032) ) ;
NOR2    gate17437  (.A(g8830), .B(g11083), .Z(g14124) ) ;
AND2    gate17438  (.A(g14124), .B(g31239), .Z(g32034) ) ;
AND2    gate17439  (.A(g4176), .B(g30937), .Z(g32035) ) ;
NOR2    gate17440  (.A(g8822), .B(g29725), .Z(g31469) ) ;
AND2    gate17441  (.A(g31469), .B(g13486), .Z(g32036) ) ;
NOR2    gate17442  (.A(g4709), .B(g29697), .Z(g31476) ) ;
AND2    gate17443  (.A(g31476), .B(g20070), .Z(g32039) ) ;
NOR2    gate17444  (.A(g8895), .B(g12259), .Z(g14122) ) ;
AND2    gate17445  (.A(g14122), .B(g31243), .Z(g32040) ) ;
NOR2    gate17446  (.A(g8859), .B(g11083), .Z(g13913) ) ;
AND2    gate17447  (.A(g13913), .B(g31262), .Z(g32041) ) ;
OR2     gate17448  (.A(g24652), .B(g25995), .Z(g27244) ) ;
AND2    gate17449  (.A(g27244), .B(g31070), .Z(g32042) ) ;
NOR2    gate17450  (.A(g8883), .B(g29697), .Z(g31482) ) ;
AND2    gate17451  (.A(g31482), .B(g16173), .Z(g32043) ) ;
NOR2    gate17452  (.A(g4899), .B(g29725), .Z(g31483) ) ;
AND2    gate17453  (.A(g31483), .B(g20085), .Z(g32044) ) ;
NOR2    gate17454  (.A(g8938), .B(g29725), .Z(g31491) ) ;
AND2    gate17455  (.A(g31491), .B(g16187), .Z(g32045) ) ;
AND2    gate17456  (.A(g10925), .B(g30735), .Z(g32046) ) ;
OR2     gate17457  (.A(g24880), .B(g25953), .Z(g27248) ) ;
AND2    gate17458  (.A(g27248), .B(g31070), .Z(g32047) ) ;
NOR2    gate17459  (.A(g9030), .B(g29540), .Z(g31498) ) ;
AND2    gate17460  (.A(g31498), .B(g13869), .Z(g32048) ) ;
AND2    gate17461  (.A(g10902), .B(g30735), .Z(g32049) ) ;
AND2    gate17462  (.A(g11003), .B(g30825), .Z(g32050) ) ;
NOR2    gate17463  (.A(g4793), .B(g29540), .Z(g31506) ) ;
AND2    gate17464  (.A(g31506), .B(g10831), .Z(g32051) ) ;
NOR2    gate17465  (.A(g9064), .B(g29556), .Z(g31507) ) ;
AND2    gate17466  (.A(g31507), .B(g13885), .Z(g32052) ) ;
NOR2    gate17467  (.A(g9044), .B(g12259), .Z(g14176) ) ;
AND2    gate17468  (.A(g14176), .B(g31509), .Z(g32053) ) ;
AND2    gate17469  (.A(g10890), .B(g30735), .Z(g32054) ) ;
AND2    gate17470  (.A(g10999), .B(g30825), .Z(g32055) ) ;
OR2     gate17471  (.A(g24547), .B(g26053), .Z(g27271) ) ;
AND2    gate17472  (.A(g27271), .B(g31021), .Z(g32056) ) ;
AND2    gate17473  (.A(g4727), .B(g30614), .Z(g32067) ) ;
NOR2    gate17474  (.A(g4983), .B(g29556), .Z(g31515) ) ;
AND2    gate17475  (.A(g31515), .B(g10862), .Z(g32068) ) ;
AND2    gate17476  (.A(g10878), .B(g30735), .Z(g32069) ) ;
AND2    gate17477  (.A(g10967), .B(g30825), .Z(g32070) ) ;
OR2     gate17478  (.A(g24620), .B(g25974), .Z(g27236) ) ;
AND2    gate17479  (.A(g27236), .B(g31070), .Z(g32071) ) ;
AND2    gate17480  (.A(g4917), .B(g30673), .Z(g32082) ) ;
AND2    gate17481  (.A(g947), .B(g30735), .Z(g32083) ) ;
AND2    gate17482  (.A(g10948), .B(g30825), .Z(g32084) ) ;
OR2     gate17483  (.A(g24661), .B(g26052), .Z(g27253) ) ;
AND2    gate17484  (.A(g27253), .B(g31021), .Z(g32085) ) ;
AND2    gate17485  (.A(g7597), .B(g30735), .Z(g32086) ) ;
AND2    gate17486  (.A(g1291), .B(g30825), .Z(g32087) ) ;
OR2     gate17487  (.A(g24584), .B(g25984), .Z(g27241) ) ;
AND2    gate17488  (.A(g27241), .B(g31070), .Z(g32088) ) ;
OR2     gate17489  (.A(g24544), .B(g25996), .Z(g27261) ) ;
AND2    gate17490  (.A(g27261), .B(g31021), .Z(g32089) ) ;
AND2    gate17491  (.A(g7619), .B(g30825), .Z(g32095) ) ;
AND2    gate17492  (.A(g31601), .B(g29893), .Z(g32096) ) ;
OR2     gate17493  (.A(g24566), .B(g24678), .Z(g25960) ) ;
AND2    gate17494  (.A(g25960), .B(g31021), .Z(g32097) ) ;
AND2    gate17495  (.A(g4732), .B(g30614), .Z(g32098) ) ;
AND2    gate17496  (.A(g31609), .B(g29905), .Z(g32103) ) ;
AND2    gate17497  (.A(g31616), .B(g29906), .Z(g32104) ) ;
AND2    gate17498  (.A(g4922), .B(g30673), .Z(g32105) ) ;
AND2    gate17499  (.A(g31601), .B(g29911), .Z(g32106) ) ;
AND2    gate17500  (.A(g31624), .B(g29912), .Z(g32107) ) ;
AND2    gate17501  (.A(g31631), .B(g29913), .Z(g32108) ) ;
AND2    gate17502  (.A(g31609), .B(g29920), .Z(g32109) ) ;
AND2    gate17503  (.A(g31639), .B(g29921), .Z(g32110) ) ;
AND2    gate17504  (.A(g31616), .B(g29922), .Z(g32111) ) ;
AND2    gate17505  (.A(g31646), .B(g29923), .Z(g32112) ) ;
AND2    gate17506  (.A(g31601), .B(g29925), .Z(g32113) ) ;
AND2    gate17507  (.A(g31624), .B(g29927), .Z(g32114) ) ;
AND2    gate17508  (.A(g31631), .B(g29928), .Z(g32115) ) ;
AND2    gate17509  (.A(g31658), .B(g29929), .Z(g32116) ) ;
AND2    gate17510  (.A(g31609), .B(g29939), .Z(g32119) ) ;
AND2    gate17511  (.A(g31639), .B(g29941), .Z(g32120) ) ;
AND2    gate17512  (.A(g31616), .B(g29942), .Z(g32121) ) ;
AND2    gate17513  (.A(g31646), .B(g29944), .Z(g32122) ) ;
AND2    gate17514  (.A(g31601), .B(g29948), .Z(g32126) ) ;
AND2    gate17515  (.A(g31624), .B(g29950), .Z(g32127) ) ;
AND2    gate17516  (.A(g31631), .B(g29953), .Z(g32128) ) ;
AND2    gate17517  (.A(g31658), .B(g29955), .Z(g32129) ) ;
AND2    gate17518  (.A(g31601), .B(g29960), .Z(g32139) ) ;
AND2    gate17519  (.A(g31609), .B(g29961), .Z(g32140) ) ;
AND2    gate17520  (.A(g31639), .B(g29963), .Z(g32141) ) ;
AND2    gate17521  (.A(g31616), .B(g29965), .Z(g32142) ) ;
AND2    gate17522  (.A(g31646), .B(g29967), .Z(g32143) ) ;
AND2    gate17523  (.A(g31609), .B(g29977), .Z(g32145) ) ;
AND2    gate17524  (.A(g31624), .B(g29978), .Z(g32146) ) ;
AND2    gate17525  (.A(g31616), .B(g29980), .Z(g32147) ) ;
AND2    gate17526  (.A(g31631), .B(g29981), .Z(g32148) ) ;
AND2    gate17527  (.A(g31658), .B(g29983), .Z(g32149) ) ;
AND2    gate17528  (.A(g31624), .B(g29995), .Z(g32150) ) ;
AND2    gate17529  (.A(g31639), .B(g29996), .Z(g32151) ) ;
AND2    gate17530  (.A(g31631), .B(g29998), .Z(g32152) ) ;
AND2    gate17531  (.A(g31646), .B(g29999), .Z(g32153) ) ;
OR2     gate17532  (.A(g29570), .B(g28285), .Z(g31277) ) ;
AND2    gate17533  (.A(g31277), .B(g14184), .Z(g32154) ) ;
AND2    gate17534  (.A(g31639), .B(g30018), .Z(g32156) ) ;
AND2    gate17535  (.A(g31646), .B(g30021), .Z(g32157) ) ;
AND2    gate17536  (.A(g31658), .B(g30022), .Z(g32158) ) ;
AND2    gate17537  (.A(g31658), .B(g30040), .Z(g32159) ) ;
OR2     gate17538  (.A(g29360), .B(g28151), .Z(g31001) ) ;
AND2    gate17539  (.A(g31001), .B(g22995), .Z(g32160) ) ;
AND2    gate17540  (.A(g3151), .B(g31154), .Z(g32161) ) ;
OR2     gate17541  (.A(g29362), .B(g28154), .Z(g31002) ) ;
AND2    gate17542  (.A(g31002), .B(g23014), .Z(g32162) ) ;
AND2    gate17543  (.A(g3502), .B(g31170), .Z(g32163) ) ;
OR2     gate17544  (.A(g13807), .B(g29773), .Z(g30733) ) ;
AND2    gate17545  (.A(g30733), .B(g25171), .Z(g32164) ) ;
NAND2   gate17546  (.A(II29254), .B(II29255), .Z(g31669) ) ;
AND2    gate17547  (.A(g31669), .B(g27742), .Z(g32165) ) ;
OR2     gate17548  (.A(g29364), .B(g28159), .Z(g31007) ) ;
AND2    gate17549  (.A(g31007), .B(g23029), .Z(g32166) ) ;
AND2    gate17550  (.A(g3853), .B(g31194), .Z(g32167) ) ;
OR2     gate17551  (.A(g13564), .B(g29693), .Z(g30597) ) ;
AND2    gate17552  (.A(g30597), .B(g25185), .Z(g32168) ) ;
OR2     gate17553  (.A(g29367), .B(g28160), .Z(g31014) ) ;
AND2    gate17554  (.A(g31014), .B(g23046), .Z(g32169) ) ;
NAND2   gate17555  (.A(II29262), .B(II29263), .Z(g31671) ) ;
AND2    gate17556  (.A(g31671), .B(g27779), .Z(g32170) ) ;
NAND2   gate17557  (.A(II29270), .B(II29271), .Z(g31706) ) ;
AND2    gate17558  (.A(g31706), .B(g27800), .Z(g32171) ) ;
AND2    gate17559  (.A(g2767), .B(g31608), .Z(g32172) ) ;
AND2    gate17560  (.A(g160), .B(g31134), .Z(g32173) ) ;
NAND2   gate17561  (.A(II29278), .B(II29279), .Z(g31708) ) ;
AND2    gate17562  (.A(g31708), .B(g27837), .Z(g32174) ) ;
NAND2   gate17563  (.A(II29285), .B(II29286), .Z(g31709) ) ;
AND2    gate17564  (.A(g31709), .B(g27858), .Z(g32175) ) ;
AND2    gate17565  (.A(g2779), .B(g31623), .Z(g32176) ) ;
OR2     gate17566  (.A(g13604), .B(g29736), .Z(g30608) ) ;
AND2    gate17567  (.A(g30608), .B(g25214), .Z(g32177) ) ;
NAND2   gate17568  (.A(II29296), .B(II29297), .Z(g31747) ) ;
AND2    gate17569  (.A(g31747), .B(g27886), .Z(g32178) ) ;
NAND2   gate17570  (.A(II29303), .B(II29304), .Z(g31748) ) ;
AND2    gate17571  (.A(g31748), .B(g27907), .Z(g32179) ) ;
AND2    gate17572  (.A(g2791), .B(g31638), .Z(g32180) ) ;
OR2     gate17573  (.A(g29375), .B(g28164), .Z(g31020) ) ;
AND2    gate17574  (.A(g31020), .B(g19912), .Z(g32181) ) ;
NAND2   gate17575  (.A(II29314), .B(II29315), .Z(g31753) ) ;
AND2    gate17576  (.A(g31753), .B(g27937), .Z(g32182) ) ;
AND2    gate17577  (.A(g2795), .B(g31653), .Z(g32183) ) ;
OR2     gate17578  (.A(g13671), .B(g29743), .Z(g30611) ) ;
AND2    gate17579  (.A(g30611), .B(g25249), .Z(g32184) ) ;
OR2     gate17580  (.A(g13737), .B(g29752), .Z(g30672) ) ;
AND2    gate17581  (.A(g30672), .B(g25287), .Z(g32187) ) ;
NAND4   gate17582  (.A(g24924), .B(g24916), .C(g24905), .D(g26863), .Z(g27586) ) ;
AND2    gate17583  (.A(g27586), .B(g31376), .Z(g32188) ) ;
OR2     gate17584  (.A(g13833), .B(g29789), .Z(g30824) ) ;
AND2    gate17585  (.A(g30824), .B(g25369), .Z(g32189) ) ;
AND2    gate17586  (.A(g142), .B(g31233), .Z(g32190) ) ;
NAND4   gate17587  (.A(g24972), .B(g24950), .C(g24906), .D(g26861), .Z(g27593) ) ;
AND2    gate17588  (.A(g27593), .B(g31376), .Z(g32191) ) ;
OR2     gate17589  (.A(g13778), .B(g29762), .Z(g30732) ) ;
AND2    gate17590  (.A(g30732), .B(g25410), .Z(g32193) ) ;
AND2    gate17591  (.A(g30601), .B(g28436), .Z(g32194) ) ;
OR2     gate17592  (.A(g13808), .B(g29774), .Z(g30734) ) ;
AND2    gate17593  (.A(g30734), .B(g25451), .Z(g32195) ) ;
NAND4   gate17594  (.A(g24917), .B(g25018), .C(g24918), .D(g26857), .Z(g27587) ) ;
AND2    gate17595  (.A(g27587), .B(g31376), .Z(g32196) ) ;
OR2     gate17596  (.A(g29477), .B(g28193), .Z(g31144) ) ;
AND2    gate17597  (.A(g31144), .B(g20088), .Z(g32197) ) ;
AND2    gate17598  (.A(g4253), .B(g31327), .Z(g32198) ) ;
OR2     gate17599  (.A(g13853), .B(g29799), .Z(g30916) ) ;
AND2    gate17600  (.A(g30916), .B(g25506), .Z(g32199) ) ;
NAND4   gate17601  (.A(g24951), .B(g24932), .C(g24925), .D(g26852), .Z(g27468) ) ;
AND2    gate17602  (.A(g27468), .B(g31376), .Z(g32200) ) ;
AND2    gate17603  (.A(g4249), .B(g31327), .Z(g32203) ) ;
AND2    gate17604  (.A(g4245), .B(g31327), .Z(g32204) ) ;
AND2    gate17605  (.A(g30922), .B(g28463), .Z(g32205) ) ;
OR2     gate17606  (.A(g13633), .B(g29742), .Z(g30609) ) ;
AND2    gate17607  (.A(g30609), .B(g25524), .Z(g32206) ) ;
OR2     gate17608  (.A(g29494), .B(g28204), .Z(g31221) ) ;
AND2    gate17609  (.A(g31221), .B(g23323), .Z(g32207) ) ;
AND2    gate17610  (.A(g4300), .B(g31327), .Z(g32224) ) ;
OR2     gate17611  (.A(g25959), .B(g29510), .Z(g31241) ) ;
AND2    gate17612  (.A(g31241), .B(g20266), .Z(g32232) ) ;
AND2    gate17613  (.A(g31601), .B(g30292), .Z(g32234) ) ;
OR2     gate17614  (.A(g25963), .B(g29515), .Z(g31244) ) ;
AND2    gate17615  (.A(g31244), .B(g20323), .Z(g32241) ) ;
OR2     gate17616  (.A(g25964), .B(g29516), .Z(g31245) ) ;
AND2    gate17617  (.A(g31245), .B(g20324), .Z(g32242) ) ;
AND2    gate17618  (.A(g31609), .B(g30297), .Z(g32244) ) ;
OR2     gate17619  (.A(g25965), .B(g29518), .Z(g31246) ) ;
AND2    gate17620  (.A(g31246), .B(g20326), .Z(g32246) ) ;
AND2    gate17621  (.A(g31616), .B(g30299), .Z(g32248) ) ;
OR2     gate17622  (.A(g29513), .B(g13324), .Z(g31247) ) ;
AND2    gate17623  (.A(g31247), .B(g20379), .Z(g32254) ) ;
OR2     gate17624  (.A(g25970), .B(g29522), .Z(g31248) ) ;
AND2    gate17625  (.A(g31248), .B(g20381), .Z(g32255) ) ;
OR2     gate17626  (.A(g25971), .B(g29523), .Z(g31249) ) ;
AND2    gate17627  (.A(g31249), .B(g20382), .Z(g32256) ) ;
AND2    gate17628  (.A(g31624), .B(g30303), .Z(g32258) ) ;
OR2     gate17629  (.A(g25972), .B(g29526), .Z(g31250) ) ;
AND2    gate17630  (.A(g31250), .B(g20385), .Z(g32260) ) ;
OR2     gate17631  (.A(g25973), .B(g29527), .Z(g31251) ) ;
AND2    gate17632  (.A(g31251), .B(g20386), .Z(g32261) ) ;
AND2    gate17633  (.A(g31631), .B(g30306), .Z(g32263) ) ;
AND2    gate17634  (.A(g2799), .B(g30567), .Z(g32265) ) ;
OR2     gate17635  (.A(g25980), .B(g29533), .Z(g31253) ) ;
AND2    gate17636  (.A(g31253), .B(g20443), .Z(g32269) ) ;
OR2     gate17637  (.A(g25981), .B(g29534), .Z(g31254) ) ;
AND2    gate17638  (.A(g31254), .B(g20444), .Z(g32270) ) ;
AND2    gate17639  (.A(g31639), .B(g30310), .Z(g32272) ) ;
OR2     gate17640  (.A(g25982), .B(g29536), .Z(g31255) ) ;
AND2    gate17641  (.A(g31255), .B(g20446), .Z(g32273) ) ;
OR2     gate17642  (.A(g25983), .B(g29537), .Z(g31256) ) ;
AND2    gate17643  (.A(g31256), .B(g20447), .Z(g32274) ) ;
AND2    gate17644  (.A(g31646), .B(g30313), .Z(g32276) ) ;
AND2    gate17645  (.A(g2811), .B(g30572), .Z(g32278) ) ;
OR2     gate17646  (.A(g29531), .B(g28253), .Z(g31257) ) ;
AND2    gate17647  (.A(g31257), .B(g20500), .Z(g32281) ) ;
OR2     gate17648  (.A(g25991), .B(g29550), .Z(g31258) ) ;
AND2    gate17649  (.A(g31258), .B(g20503), .Z(g32282) ) ;
OR2     gate17650  (.A(g25992), .B(g29554), .Z(g31259) ) ;
AND2    gate17651  (.A(g31259), .B(g20506), .Z(g32283) ) ;
OR2     gate17652  (.A(g25993), .B(g29555), .Z(g31260) ) ;
AND2    gate17653  (.A(g31260), .B(g20507), .Z(g32284) ) ;
AND2    gate17654  (.A(g31658), .B(g29312), .Z(g32286) ) ;
AND2    gate17655  (.A(g2823), .B(g30578), .Z(g32287) ) ;
OR2     gate17656  (.A(g29548), .B(g28263), .Z(g31267) ) ;
AND2    gate17657  (.A(g31267), .B(g20525), .Z(g32290) ) ;
OR2     gate17658  (.A(g29552), .B(g28266), .Z(g31268) ) ;
AND2    gate17659  (.A(g31268), .B(g20527), .Z(g32291) ) ;
OR2     gate17660  (.A(g26024), .B(g29569), .Z(g31269) ) ;
AND2    gate17661  (.A(g31269), .B(g20530), .Z(g32292) ) ;
AND2    gate17662  (.A(g2827), .B(g30593), .Z(g32293) ) ;
NAND3   gate17663  (.A(g25425), .B(g25381), .C(g25780), .Z(g27931) ) ;
AND2    gate17664  (.A(g27931), .B(g31376), .Z(g32295) ) ;
OR2     gate17665  (.A(g29565), .B(g28280), .Z(g31274) ) ;
AND2    gate17666  (.A(g31274), .B(g20544), .Z(g32300) ) ;
OR2     gate17667  (.A(g29567), .B(g28282), .Z(g31276) ) ;
AND2    gate17668  (.A(g31276), .B(g20547), .Z(g32301) ) ;
OR2     gate17669  (.A(g29571), .B(g29579), .Z(g31279) ) ;
AND2    gate17670  (.A(g31279), .B(g23485), .Z(g32302) ) ;
NAND2   gate17671  (.A(g24943), .B(g25772), .Z(g27550) ) ;
AND2    gate17672  (.A(g27550), .B(g31376), .Z(g32303) ) ;
OR2     gate17673  (.A(g29575), .B(g28290), .Z(g31284) ) ;
AND2    gate17674  (.A(g31284), .B(g20564), .Z(g32304) ) ;
OR2     gate17675  (.A(g29578), .B(g28292), .Z(g31287) ) ;
AND2    gate17676  (.A(g31287), .B(g20567), .Z(g32305) ) ;
OR2     gate17677  (.A(g29580), .B(g29591), .Z(g31289) ) ;
AND2    gate17678  (.A(g31289), .B(g23499), .Z(g32306) ) ;
OR2     gate17679  (.A(g29581), .B(g29593), .Z(g31291) ) ;
AND2    gate17680  (.A(g31291), .B(g23500), .Z(g32307) ) ;
OR2     gate17681  (.A(g29582), .B(g28299), .Z(g31293) ) ;
AND2    gate17682  (.A(g31293), .B(g23503), .Z(g32308) ) ;
AND2    gate17683  (.A(g5160), .B(g31528), .Z(g32309) ) ;
NAND4   gate17684  (.A(g25019), .B(g25002), .C(g24988), .D(g25765), .Z(g27577) ) ;
AND2    gate17685  (.A(g27577), .B(g31376), .Z(g32310) ) ;
OR2     gate17686  (.A(g26090), .B(g29598), .Z(g31295) ) ;
AND2    gate17687  (.A(g31295), .B(g20582), .Z(g32311) ) ;
OR2     gate17688  (.A(g29590), .B(g28302), .Z(g31302) ) ;
AND2    gate17689  (.A(g31302), .B(g20591), .Z(g32312) ) ;
OR2     gate17690  (.A(g29592), .B(g29606), .Z(g31303) ) ;
AND2    gate17691  (.A(g31303), .B(g23515), .Z(g32313) ) ;
OR2     gate17692  (.A(g29594), .B(g29608), .Z(g31304) ) ;
AND2    gate17693  (.A(g31304), .B(g23516), .Z(g32314) ) ;
OR2     gate17694  (.A(g29595), .B(g29610), .Z(g31306) ) ;
AND2    gate17695  (.A(g31306), .B(g23517), .Z(g32315) ) ;
OR2     gate17696  (.A(g29596), .B(g28311), .Z(g31307) ) ;
AND2    gate17697  (.A(g31307), .B(g23522), .Z(g32316) ) ;
AND2    gate17698  (.A(g5507), .B(g31542), .Z(g32317) ) ;
NAND4   gate17699  (.A(g24942), .B(g24933), .C(g25048), .D(g26871), .Z(g27613) ) ;
AND2    gate17700  (.A(g27613), .B(g31376), .Z(g32321) ) ;
OR2     gate17701  (.A(g26101), .B(g29614), .Z(g31308) ) ;
AND2    gate17702  (.A(g31308), .B(g20605), .Z(g32322) ) ;
OR2     gate17703  (.A(g26103), .B(g29618), .Z(g31311) ) ;
AND2    gate17704  (.A(g31311), .B(g20610), .Z(g32323) ) ;
OR2     gate17705  (.A(g29607), .B(g29623), .Z(g31315) ) ;
AND2    gate17706  (.A(g31315), .B(g23537), .Z(g32324) ) ;
OR2     gate17707  (.A(g29609), .B(g29624), .Z(g31316) ) ;
AND2    gate17708  (.A(g31316), .B(g23538), .Z(g32325) ) ;
OR2     gate17709  (.A(g29611), .B(g29626), .Z(g31317) ) ;
AND2    gate17710  (.A(g31317), .B(g23539), .Z(g32326) ) ;
OR2     gate17711  (.A(g29612), .B(g28324), .Z(g31319) ) ;
AND2    gate17712  (.A(g31319), .B(g23544), .Z(g32327) ) ;
AND2    gate17713  (.A(g5853), .B(g31554), .Z(g32328) ) ;
OR2     gate17714  (.A(g26125), .B(g29632), .Z(g31320) ) ;
AND2    gate17715  (.A(g31320), .B(g20631), .Z(g32330) ) ;
OR2     gate17716  (.A(g26128), .B(g29635), .Z(g31322) ) ;
AND2    gate17717  (.A(g31322), .B(g20637), .Z(g32331) ) ;
OR2     gate17718  (.A(g29625), .B(g29639), .Z(g31325) ) ;
AND2    gate17719  (.A(g31325), .B(g23558), .Z(g32332) ) ;
OR2     gate17720  (.A(g29627), .B(g29640), .Z(g31326) ) ;
AND2    gate17721  (.A(g31326), .B(g23559), .Z(g32333) ) ;
OR2     gate17722  (.A(g29628), .B(g28339), .Z(g31375) ) ;
AND2    gate17723  (.A(g31375), .B(g23568), .Z(g32334) ) ;
AND2    gate17724  (.A(g6199), .B(g31566), .Z(g32335) ) ;
AND2    gate17725  (.A(g31596), .B(g11842), .Z(g32336) ) ;
OR2     gate17726  (.A(g26156), .B(g29647), .Z(g31465) ) ;
AND2    gate17727  (.A(g31465), .B(g20663), .Z(g32337) ) ;
OR2     gate17728  (.A(g26160), .B(g29650), .Z(g31466) ) ;
AND2    gate17729  (.A(g31466), .B(g20668), .Z(g32338) ) ;
OR2     gate17730  (.A(g29668), .B(g13583), .Z(g31474) ) ;
AND2    gate17731  (.A(g31474), .B(g20672), .Z(g32339) ) ;
OR2     gate17732  (.A(g29641), .B(g29656), .Z(g31468) ) ;
AND2    gate17733  (.A(g31468), .B(g23585), .Z(g32340) ) ;
OR2     gate17734  (.A(g29642), .B(g28352), .Z(g31472) ) ;
AND2    gate17735  (.A(g31472), .B(g23610), .Z(g32341) ) ;
AND2    gate17736  (.A(g6545), .B(g31579), .Z(g32342) ) ;
OR2     gate17737  (.A(g26180), .B(g29666), .Z(g31473) ) ;
AND2    gate17738  (.A(g31473), .B(g20710), .Z(g32343) ) ;
AND2    gate17739  (.A(g2138), .B(g31672), .Z(g32345) ) ;
AND2    gate17740  (.A(g2145), .B(g31672), .Z(g32348) ) ;
AND2    gate17741  (.A(g2697), .B(g31710), .Z(g32350) ) ;
AND2    gate17742  (.A(g2704), .B(g31710), .Z(g32356) ) ;
AND2    gate17743  (.A(g2130), .B(g31672), .Z(g32369) ) ;
AND2    gate17744  (.A(g2689), .B(g31710), .Z(g32376) ) ;
AND2    gate17745  (.A(g4698), .B(g30983), .Z(g32396) ) ;
NOR2    gate17746  (.A(g4801), .B(g29540), .Z(g31068) ) ;
AND2    gate17747  (.A(g31068), .B(g15830), .Z(g32397) ) ;
AND2    gate17748  (.A(g4743), .B(g30989), .Z(g32400) ) ;
NOR2    gate17749  (.A(g7892), .B(g29540), .Z(g31116) ) ;
AND2    gate17750  (.A(g31116), .B(g13432), .Z(g32401) ) ;
AND2    gate17751  (.A(g4888), .B(g30990), .Z(g32402) ) ;
NOR2    gate17752  (.A(g4991), .B(g29556), .Z(g31117) ) ;
AND2    gate17753  (.A(g31117), .B(g15842), .Z(g32403) ) ;
AND2    gate17754  (.A(g4754), .B(g30996), .Z(g32409) ) ;
AND2    gate17755  (.A(g4933), .B(g30997), .Z(g32410) ) ;
NOR2    gate17756  (.A(g7898), .B(g29556), .Z(g31119) ) ;
AND2    gate17757  (.A(g31119), .B(g13469), .Z(g32411) ) ;
AND2    gate17758  (.A(g4765), .B(g30998), .Z(g32412) ) ;
NOR2    gate17759  (.A(g4776), .B(g29540), .Z(g31121) ) ;
AND2    gate17760  (.A(g31121), .B(g19518), .Z(g32413) ) ;
AND2    gate17761  (.A(g4944), .B(g30999), .Z(g32414) ) ;
NOR2    gate17762  (.A(g7928), .B(g29540), .Z(g31126) ) ;
AND2    gate17763  (.A(g31126), .B(g16239), .Z(g32418) ) ;
AND2    gate17764  (.A(g4955), .B(g31000), .Z(g32419) ) ;
NOR2    gate17765  (.A(g4966), .B(g29556), .Z(g31127) ) ;
AND2    gate17766  (.A(g31127), .B(g19533), .Z(g32420) ) ;
OR2     gate17767  (.A(g29924), .B(g28558), .Z(g31668) ) ;
AND2    gate17768  (.A(g31668), .B(g21604), .Z(g32425) ) ;
NOR2    gate17769  (.A(g7953), .B(g29556), .Z(g31133) ) ;
AND2    gate17770  (.A(g31133), .B(g16261), .Z(g32428) ) ;
AND2    gate17771  (.A(g31591), .B(g32404), .Z(g33071) ) ;
OR2     gate17772  (.A(g31488), .B(g29949), .Z(g32386) ) ;
AND2    gate17773  (.A(g32386), .B(g18828), .Z(g33073) ) ;
OR2     gate17774  (.A(g31489), .B(g29952), .Z(g32387) ) ;
AND2    gate17775  (.A(g32387), .B(g18830), .Z(g33074) ) ;
OR2     gate17776  (.A(g31495), .B(g29962), .Z(g32388) ) ;
AND2    gate17777  (.A(g32388), .B(g18875), .Z(g33081) ) ;
OR2     gate17778  (.A(g31496), .B(g29966), .Z(g32389) ) ;
AND2    gate17779  (.A(g32389), .B(g18877), .Z(g33082) ) ;
OR2     gate17780  (.A(g31501), .B(g29979), .Z(g32390) ) ;
AND2    gate17781  (.A(g32390), .B(g18887), .Z(g33086) ) ;
OR2     gate17782  (.A(g31502), .B(g29982), .Z(g32391) ) ;
AND2    gate17783  (.A(g32391), .B(g18888), .Z(g33087) ) ;
OR2     gate17784  (.A(g31513), .B(g30000), .Z(g32392) ) ;
AND2    gate17785  (.A(g32392), .B(g18897), .Z(g33091) ) ;
OR2     gate17786  (.A(g31523), .B(g30049), .Z(g32395) ) ;
AND2    gate17787  (.A(g32395), .B(g18944), .Z(g33099) ) ;
OR2     gate17788  (.A(g31526), .B(g30061), .Z(g32398) ) ;
AND2    gate17789  (.A(g32398), .B(g18976), .Z(g33101) ) ;
OR2     gate17790  (.A(g31527), .B(g30062), .Z(g32399) ) ;
AND2    gate17791  (.A(g32399), .B(g18978), .Z(g33102) ) ;
NOR2    gate17792  (.A(g8287), .B(g24732), .Z(g26296) ) ;
AND2    gate17793  (.A(g26296), .B(g32137), .Z(g33104) ) ;
NOR2    gate17794  (.A(g8297), .B(g24825), .Z(g26298) ) ;
AND2    gate17795  (.A(g26298), .B(g32138), .Z(g33105) ) ;
OR2     gate17796  (.A(g31541), .B(g30073), .Z(g32408) ) ;
AND2    gate17797  (.A(g32408), .B(g18990), .Z(g33106) ) ;
AND2    gate17798  (.A(g32404), .B(g32415), .Z(g33110) ) ;
AND2    gate17799  (.A(g24005), .B(g32421), .Z(g33111) ) ;
OR2     gate17800  (.A(g31654), .B(g14544), .Z(g31964) ) ;
AND2    gate17801  (.A(g31964), .B(g22339), .Z(g33113) ) ;
AND2    gate17802  (.A(g22139), .B(g31945), .Z(g33114) ) ;
AND2    gate17803  (.A(g8748), .B(g32212), .Z(g33121) ) ;
AND2    gate17804  (.A(g8859), .B(g32192), .Z(g33122) ) ;
AND2    gate17805  (.A(g8945), .B(g32296), .Z(g33124) ) ;
AND2    gate17806  (.A(g9044), .B(g32201), .Z(g33126) ) ;
OR2     gate17807  (.A(g30566), .B(g29329), .Z(g32037) ) ;
AND2    gate17808  (.A(g32037), .B(g22830), .Z(g33186) ) ;
OR2     gate17809  (.A(g30612), .B(g29363), .Z(g32094) ) ;
AND2    gate17810  (.A(g32094), .B(g23005), .Z(g33233) ) ;
AND2    gate17811  (.A(g32394), .B(g25198), .Z(g33237) ) ;
OR2     gate17812  (.A(g24482), .B(g30914), .Z(g32117) ) ;
AND2    gate17813  (.A(g32117), .B(g19902), .Z(g33239) ) ;
AND2    gate17814  (.A(g32173), .B(g23128), .Z(g33241) ) ;
OR2     gate17815  (.A(g30915), .B(g30919), .Z(g32123) ) ;
AND2    gate17816  (.A(g32123), .B(g19931), .Z(g33242) ) ;
OR2     gate17817  (.A(g24488), .B(g30920), .Z(g32124) ) ;
AND2    gate17818  (.A(g32124), .B(g19947), .Z(g33243) ) ;
AND2    gate17819  (.A(g32190), .B(g23152), .Z(g33244) ) ;
OR2     gate17820  (.A(g30918), .B(g29376), .Z(g32125) ) ;
AND2    gate17821  (.A(g32125), .B(g19961), .Z(g33245) ) ;
OR2     gate17822  (.A(g30921), .B(g30925), .Z(g32130) ) ;
AND2    gate17823  (.A(g32130), .B(g19980), .Z(g33247) ) ;
OR2     gate17824  (.A(g24495), .B(g30926), .Z(g32131) ) ;
AND2    gate17825  (.A(g32131), .B(g19996), .Z(g33248) ) ;
OR2     gate17826  (.A(g30927), .B(g30930), .Z(g32144) ) ;
AND2    gate17827  (.A(g32144), .B(g20026), .Z(g33249) ) ;
OR2     gate17828  (.A(g30935), .B(g29475), .Z(g32155) ) ;
AND2    gate17829  (.A(g32155), .B(g20064), .Z(g33252) ) ;
AND2    gate17830  (.A(g32393), .B(g25481), .Z(g33263) ) ;
NOR2    gate17831  (.A(g30583), .B(g4358), .Z(g31965) ) ;
AND2    gate17832  (.A(g31965), .B(g21306), .Z(g33264) ) ;
NOR2    gate17833  (.A(g9024), .B(g30583), .Z(g31970) ) ;
AND2    gate17834  (.A(g31970), .B(g15582), .Z(g33269) ) ;
OR2     gate17835  (.A(g8928), .B(g30583), .Z(g32427) ) ;
AND2    gate17836  (.A(g32427), .B(g31971), .Z(g33304) ) ;
NOR2    gate17837  (.A(g30583), .B(g4349), .Z(g31935) ) ;
AND2    gate17838  (.A(g31935), .B(g17811), .Z(g33305) ) ;
NOR2    gate17839  (.A(g8977), .B(g30583), .Z(g31942) ) ;
AND2    gate17840  (.A(g31942), .B(g12925), .Z(g33311) ) ;
OR2     gate17841  (.A(g31069), .B(g13410), .Z(g32202) ) ;
AND2    gate17842  (.A(g32202), .B(g20450), .Z(g33322) ) ;
OR2     gate17843  (.A(g31120), .B(g29584), .Z(g32208) ) ;
AND2    gate17844  (.A(g32208), .B(g20561), .Z(g33327) ) ;
OR2     gate17845  (.A(g31122), .B(g29599), .Z(g32209) ) ;
AND2    gate17846  (.A(g32209), .B(g20584), .Z(g33328) ) ;
OR2     gate17847  (.A(g31123), .B(g29600), .Z(g32210) ) ;
AND2    gate17848  (.A(g32210), .B(g20585), .Z(g33329) ) ;
OR2     gate17849  (.A(g31124), .B(g29603), .Z(g32211) ) ;
AND2    gate17850  (.A(g32211), .B(g20588), .Z(g33330) ) ;
OR2     gate17851  (.A(g31128), .B(g29615), .Z(g32216) ) ;
AND2    gate17852  (.A(g32216), .B(g20607), .Z(g33331) ) ;
OR2     gate17853  (.A(g31129), .B(g29616), .Z(g32217) ) ;
AND2    gate17854  (.A(g32217), .B(g20608), .Z(g33332) ) ;
OR2     gate17855  (.A(g31130), .B(g29619), .Z(g32218) ) ;
AND2    gate17856  (.A(g32218), .B(g20612), .Z(g33333) ) ;
OR2     gate17857  (.A(g31131), .B(g29620), .Z(g32219) ) ;
AND2    gate17858  (.A(g32219), .B(g20613), .Z(g33334) ) ;
OR2     gate17859  (.A(g31139), .B(g29633), .Z(g32220) ) ;
AND2    gate17860  (.A(g32220), .B(g20633), .Z(g33338) ) ;
OR2     gate17861  (.A(g31140), .B(g29634), .Z(g32221) ) ;
AND2    gate17862  (.A(g32221), .B(g20634), .Z(g33339) ) ;
OR2     gate17863  (.A(g31141), .B(g29636), .Z(g32222) ) ;
AND2    gate17864  (.A(g32222), .B(g20639), .Z(g33340) ) ;
OR2     gate17865  (.A(g31142), .B(g29637), .Z(g32223) ) ;
AND2    gate17866  (.A(g32223), .B(g20640), .Z(g33341) ) ;
OR2     gate17867  (.A(g31145), .B(g29645), .Z(g32226) ) ;
AND2    gate17868  (.A(g32226), .B(g20660), .Z(g33342) ) ;
OR2     gate17869  (.A(g31146), .B(g29648), .Z(g32227) ) ;
AND2    gate17870  (.A(g32227), .B(g20665), .Z(g33343) ) ;
OR2     gate17871  (.A(g31147), .B(g29651), .Z(g32228) ) ;
AND2    gate17872  (.A(g32228), .B(g20670), .Z(g33344) ) ;
OR2     gate17873  (.A(g31148), .B(g29652), .Z(g32229) ) ;
AND2    gate17874  (.A(g32229), .B(g20671), .Z(g33345) ) ;
OR2     gate17875  (.A(g31150), .B(g29661), .Z(g32233) ) ;
AND2    gate17876  (.A(g32233), .B(g20699), .Z(g33349) ) ;
OR2     gate17877  (.A(g31151), .B(g29662), .Z(g32235) ) ;
AND2    gate17878  (.A(g32235), .B(g20702), .Z(g33350) ) ;
OR2     gate17879  (.A(g31152), .B(g29664), .Z(g32236) ) ;
AND2    gate17880  (.A(g32236), .B(g20707), .Z(g33351) ) ;
OR2     gate17881  (.A(g31153), .B(g29667), .Z(g32237) ) ;
AND2    gate17882  (.A(g32237), .B(g20712), .Z(g33352) ) ;
OR2     gate17883  (.A(g24757), .B(g31182), .Z(g32240) ) ;
AND2    gate17884  (.A(g32240), .B(g20732), .Z(g33353) ) ;
OR2     gate17885  (.A(g31166), .B(g29683), .Z(g32243) ) ;
AND2    gate17886  (.A(g32243), .B(g20769), .Z(g33355) ) ;
OR2     gate17887  (.A(g31167), .B(g29684), .Z(g32245) ) ;
AND2    gate17888  (.A(g32245), .B(g20772), .Z(g33356) ) ;
OR2     gate17889  (.A(g31168), .B(g29686), .Z(g32247) ) ;
AND2    gate17890  (.A(g32247), .B(g20775), .Z(g33357) ) ;
OR2     gate17891  (.A(g31169), .B(g29687), .Z(g32249) ) ;
AND2    gate17892  (.A(g32249), .B(g20778), .Z(g33358) ) ;
OR2     gate17893  (.A(g31183), .B(g31206), .Z(g32252) ) ;
AND2    gate17894  (.A(g32252), .B(g20853), .Z(g33359) ) ;
OR2     gate17895  (.A(g24771), .B(g31207), .Z(g32253) ) ;
AND2    gate17896  (.A(g32253), .B(g20869), .Z(g33360) ) ;
OR2     gate17897  (.A(g31184), .B(g29708), .Z(g32257) ) ;
AND2    gate17898  (.A(g32257), .B(g20911), .Z(g33361) ) ;
OR2     gate17899  (.A(g31185), .B(g29709), .Z(g32259) ) ;
AND2    gate17900  (.A(g32259), .B(g20914), .Z(g33362) ) ;
OR2     gate17901  (.A(g31186), .B(g29710), .Z(g32262) ) ;
AND2    gate17902  (.A(g32262), .B(g20918), .Z(g33363) ) ;
OR2     gate17903  (.A(g31187), .B(g29711), .Z(g32264) ) ;
AND2    gate17904  (.A(g32264), .B(g20921), .Z(g33364) ) ;
OR2     gate17905  (.A(g31208), .B(g31218), .Z(g32267) ) ;
AND2    gate17906  (.A(g32267), .B(g20994), .Z(g33365) ) ;
OR2     gate17907  (.A(g24785), .B(g31219), .Z(g32268) ) ;
AND2    gate17908  (.A(g32268), .B(g21010), .Z(g33366) ) ;
OR2     gate17909  (.A(g31209), .B(g29731), .Z(g32271) ) ;
AND2    gate17910  (.A(g32271), .B(g21053), .Z(g33367) ) ;
OR2     gate17911  (.A(g31210), .B(g29732), .Z(g32275) ) ;
AND2    gate17912  (.A(g32275), .B(g21057), .Z(g33368) ) ;
OR2     gate17913  (.A(g31211), .B(g29733), .Z(g32277) ) ;
AND2    gate17914  (.A(g32277), .B(g21060), .Z(g33369) ) ;
OR2     gate17915  (.A(g31220), .B(g31224), .Z(g32279) ) ;
AND2    gate17916  (.A(g32279), .B(g21139), .Z(g33370) ) ;
OR2     gate17917  (.A(g24790), .B(g31225), .Z(g32280) ) ;
AND2    gate17918  (.A(g32280), .B(g21155), .Z(g33371) ) ;
OR2     gate17919  (.A(g31222), .B(g29740), .Z(g32285) ) ;
AND2    gate17920  (.A(g32285), .B(g21183), .Z(g33372) ) ;
OR2     gate17921  (.A(g31226), .B(g31229), .Z(g32288) ) ;
AND2    gate17922  (.A(g32288), .B(g21205), .Z(g33373) ) ;
OR2     gate17923  (.A(g24796), .B(g31230), .Z(g32289) ) ;
AND2    gate17924  (.A(g32289), .B(g21221), .Z(g33374) ) ;
OR2     gate17925  (.A(g31231), .B(g31232), .Z(g32294) ) ;
AND2    gate17926  (.A(g32294), .B(g21268), .Z(g33376) ) ;
AND2    gate17927  (.A(g30984), .B(g32364), .Z(g33379) ) ;
AND2    gate17928  (.A(g11842), .B(g32318), .Z(g33381) ) ;
OR2     gate17929  (.A(g29804), .B(g31266), .Z(g32344) ) ;
AND2    gate17930  (.A(g32344), .B(g21362), .Z(g33392) ) ;
OR2     gate17931  (.A(g29838), .B(g31272), .Z(g32346) ) ;
AND2    gate17932  (.A(g32346), .B(g21379), .Z(g33399) ) ;
OR2     gate17933  (.A(g29839), .B(g31273), .Z(g32347) ) ;
AND2    gate17934  (.A(g32347), .B(g21380), .Z(g33400) ) ;
OR2     gate17935  (.A(g29840), .B(g31275), .Z(g32349) ) ;
AND2    gate17936  (.A(g32349), .B(g21381), .Z(g33401) ) ;
OR2     gate17937  (.A(g29851), .B(g31281), .Z(g32351) ) ;
AND2    gate17938  (.A(g32351), .B(g21395), .Z(g33402) ) ;
OR2     gate17939  (.A(g29852), .B(g31282), .Z(g32352) ) ;
AND2    gate17940  (.A(g32352), .B(g21396), .Z(g33403) ) ;
OR2     gate17941  (.A(g29853), .B(g31283), .Z(g32353) ) ;
AND2    gate17942  (.A(g32353), .B(g21397), .Z(g33404) ) ;
OR2     gate17943  (.A(g29854), .B(g31285), .Z(g32354) ) ;
AND2    gate17944  (.A(g32354), .B(g21398), .Z(g33405) ) ;
OR2     gate17945  (.A(g29855), .B(g31286), .Z(g32355) ) ;
AND2    gate17946  (.A(g32355), .B(g21399), .Z(g33406) ) ;
OR2     gate17947  (.A(g29865), .B(g31296), .Z(g32357) ) ;
AND2    gate17948  (.A(g32357), .B(g21406), .Z(g33407) ) ;
OR2     gate17949  (.A(g29866), .B(g31297), .Z(g32358) ) ;
AND2    gate17950  (.A(g32358), .B(g21407), .Z(g33408) ) ;
OR2     gate17951  (.A(g29867), .B(g31298), .Z(g32359) ) ;
AND2    gate17952  (.A(g32359), .B(g21408), .Z(g33409) ) ;
OR2     gate17953  (.A(g29868), .B(g31299), .Z(g32360) ) ;
AND2    gate17954  (.A(g32360), .B(g21409), .Z(g33410) ) ;
OR2     gate17955  (.A(g29869), .B(g31300), .Z(g32361) ) ;
AND2    gate17956  (.A(g32361), .B(g21410), .Z(g33411) ) ;
OR2     gate17957  (.A(g29870), .B(g31301), .Z(g32362) ) ;
AND2    gate17958  (.A(g32362), .B(g21411), .Z(g33412) ) ;
OR2     gate17959  (.A(g29880), .B(g31309), .Z(g32367) ) ;
AND2    gate17960  (.A(g32367), .B(g21421), .Z(g33414) ) ;
OR2     gate17961  (.A(g29881), .B(g31310), .Z(g32368) ) ;
AND2    gate17962  (.A(g32368), .B(g21422), .Z(g33415) ) ;
OR2     gate17963  (.A(g29882), .B(g31312), .Z(g32370) ) ;
AND2    gate17964  (.A(g32370), .B(g21423), .Z(g33416) ) ;
OR2     gate17965  (.A(g29883), .B(g31313), .Z(g32371) ) ;
AND2    gate17966  (.A(g32371), .B(g21424), .Z(g33417) ) ;
OR2     gate17967  (.A(g29884), .B(g31314), .Z(g32372) ) ;
AND2    gate17968  (.A(g32372), .B(g21425), .Z(g33418) ) ;
OR2     gate17969  (.A(g29894), .B(g31321), .Z(g32373) ) ;
AND2    gate17970  (.A(g32373), .B(g21454), .Z(g33420) ) ;
OR2     gate17971  (.A(g29895), .B(g31323), .Z(g32374) ) ;
AND2    gate17972  (.A(g32374), .B(g21455), .Z(g33421) ) ;
OR2     gate17973  (.A(g29896), .B(g31324), .Z(g32375) ) ;
AND2    gate17974  (.A(g32375), .B(g21456), .Z(g33422) ) ;
OR2     gate17975  (.A(g30576), .B(g29336), .Z(g32225) ) ;
AND2    gate17976  (.A(g32225), .B(g29657), .Z(g33423) ) ;
OR2     gate17977  (.A(g29907), .B(g31467), .Z(g32380) ) ;
AND2    gate17978  (.A(g32380), .B(g21466), .Z(g33425) ) ;
OR2     gate17979  (.A(g30589), .B(g29345), .Z(g32230) ) ;
AND2    gate17980  (.A(g32230), .B(g29672), .Z(g33428) ) ;
OR2     gate17981  (.A(g30590), .B(g29346), .Z(g32231) ) ;
AND2    gate17982  (.A(g32231), .B(g29676), .Z(g33429) ) ;
AND2    gate17983  (.A(g32364), .B(g32377), .Z(g33431) ) ;
OR2     gate17984  (.A(g30594), .B(g29349), .Z(g32238) ) ;
AND2    gate17985  (.A(g32238), .B(g29694), .Z(g33433) ) ;
OR2     gate17986  (.A(g30595), .B(g29350), .Z(g32239) ) ;
AND2    gate17987  (.A(g32239), .B(g29702), .Z(g33434) ) ;
OR2     gate17988  (.A(g30598), .B(g29351), .Z(g32250) ) ;
AND2    gate17989  (.A(g32250), .B(g29719), .Z(g33440) ) ;
OR2     gate17990  (.A(g30599), .B(g29352), .Z(g32251) ) ;
AND2    gate17991  (.A(g32251), .B(g29722), .Z(g33441) ) ;
OR2     gate17992  (.A(g31480), .B(g29938), .Z(g32385) ) ;
AND2    gate17993  (.A(g32385), .B(g21607), .Z(g33446) ) ;
OR2     gate17994  (.A(g30604), .B(g29354), .Z(g32266) ) ;
AND2    gate17995  (.A(g32266), .B(g29737), .Z(g33450) ) ;
AND4    gate17996  (.A(g29385), .B(g32456), .C(g32457), .D(g32458), .Z(II31001) ) ;
AND4    gate17997  (.A(g32459), .B(g32460), .C(g32461), .D(g32462), .Z(II31002) ) ;
AND3    gate17998  (.A(g32463), .B(II31001), .C(II31002), .Z(g33461) ) ;
AND4    gate17999  (.A(g31376), .B(g31796), .C(g32464), .D(g32465), .Z(II31006) ) ;
AND4    gate18000  (.A(g32466), .B(g32467), .C(g32468), .D(g32469), .Z(II31007) ) ;
AND3    gate18001  (.A(g32470), .B(II31006), .C(II31007), .Z(g33462) ) ;
AND4    gate18002  (.A(g30735), .B(g31797), .C(g32471), .D(g32472), .Z(II31011) ) ;
AND4    gate18003  (.A(g32473), .B(g32474), .C(g32475), .D(g32476), .Z(II31012) ) ;
AND3    gate18004  (.A(g32477), .B(II31011), .C(II31012), .Z(g33463) ) ;
AND4    gate18005  (.A(g30825), .B(g31798), .C(g32478), .D(g32479), .Z(II31016) ) ;
AND4    gate18006  (.A(g32480), .B(g32481), .C(g32482), .D(g32483), .Z(II31017) ) ;
AND3    gate18007  (.A(g32484), .B(II31016), .C(II31017), .Z(g33464) ) ;
AND4    gate18008  (.A(g31070), .B(g31799), .C(g32485), .D(g32486), .Z(II31021) ) ;
AND4    gate18009  (.A(g32487), .B(g32488), .C(g32489), .D(g32490), .Z(II31022) ) ;
AND3    gate18010  (.A(g32491), .B(II31021), .C(II31022), .Z(g33465) ) ;
AND4    gate18011  (.A(g31194), .B(g31800), .C(g32492), .D(g32493), .Z(II31026) ) ;
AND4    gate18012  (.A(g32494), .B(g32495), .C(g32496), .D(g32497), .Z(II31027) ) ;
AND3    gate18013  (.A(g32498), .B(II31026), .C(II31027), .Z(g33466) ) ;
AND4    gate18014  (.A(g30614), .B(g31801), .C(g32499), .D(g32500), .Z(II31031) ) ;
AND4    gate18015  (.A(g32501), .B(g32502), .C(g32503), .D(g32504), .Z(II31032) ) ;
AND3    gate18016  (.A(g32505), .B(II31031), .C(II31032), .Z(g33467) ) ;
AND4    gate18017  (.A(g30673), .B(g31802), .C(g32506), .D(g32507), .Z(II31036) ) ;
AND4    gate18018  (.A(g32508), .B(g32509), .C(g32510), .D(g32511), .Z(II31037) ) ;
AND3    gate18019  (.A(g32512), .B(II31036), .C(II31037), .Z(g33468) ) ;
AND4    gate18020  (.A(g31566), .B(g31803), .C(g32513), .D(g32514), .Z(II31041) ) ;
AND4    gate18021  (.A(g32515), .B(g32516), .C(g32517), .D(g32518), .Z(II31042) ) ;
AND3    gate18022  (.A(g32519), .B(II31041), .C(II31042), .Z(g33469) ) ;
AND4    gate18023  (.A(g29385), .B(g32521), .C(g32522), .D(g32523), .Z(II31046) ) ;
AND4    gate18024  (.A(g32524), .B(g32525), .C(g32526), .D(g32527), .Z(II31047) ) ;
AND3    gate18025  (.A(g32528), .B(II31046), .C(II31047), .Z(g33470) ) ;
AND4    gate18026  (.A(g31376), .B(g31804), .C(g32529), .D(g32530), .Z(II31051) ) ;
AND4    gate18027  (.A(g32531), .B(g32532), .C(g32533), .D(g32534), .Z(II31052) ) ;
AND3    gate18028  (.A(g32535), .B(II31051), .C(II31052), .Z(g33471) ) ;
AND4    gate18029  (.A(g30735), .B(g31805), .C(g32536), .D(g32537), .Z(II31056) ) ;
AND4    gate18030  (.A(g32538), .B(g32539), .C(g32540), .D(g32541), .Z(II31057) ) ;
AND3    gate18031  (.A(g32542), .B(II31056), .C(II31057), .Z(g33472) ) ;
AND4    gate18032  (.A(g30825), .B(g31806), .C(g32543), .D(g32544), .Z(II31061) ) ;
AND4    gate18033  (.A(g32545), .B(g32546), .C(g32547), .D(g32548), .Z(II31062) ) ;
AND3    gate18034  (.A(g32549), .B(II31061), .C(II31062), .Z(g33473) ) ;
AND4    gate18035  (.A(g31070), .B(g31807), .C(g32550), .D(g32551), .Z(II31066) ) ;
AND4    gate18036  (.A(g32552), .B(g32553), .C(g32554), .D(g32555), .Z(II31067) ) ;
AND3    gate18037  (.A(g32556), .B(II31066), .C(II31067), .Z(g33474) ) ;
AND4    gate18038  (.A(g31170), .B(g31808), .C(g32557), .D(g32558), .Z(II31071) ) ;
AND4    gate18039  (.A(g32559), .B(g32560), .C(g32561), .D(g32562), .Z(II31072) ) ;
AND3    gate18040  (.A(g32563), .B(II31071), .C(II31072), .Z(g33475) ) ;
AND4    gate18041  (.A(g30614), .B(g31809), .C(g32564), .D(g32565), .Z(II31076) ) ;
AND4    gate18042  (.A(g32566), .B(g32567), .C(g32568), .D(g32569), .Z(II31077) ) ;
AND3    gate18043  (.A(g32570), .B(II31076), .C(II31077), .Z(g33476) ) ;
AND4    gate18044  (.A(g30673), .B(g31810), .C(g32571), .D(g32572), .Z(II31081) ) ;
AND4    gate18045  (.A(g32573), .B(g32574), .C(g32575), .D(g32576), .Z(II31082) ) ;
AND3    gate18046  (.A(g32577), .B(II31081), .C(II31082), .Z(g33477) ) ;
AND4    gate18047  (.A(g31554), .B(g31811), .C(g32578), .D(g32579), .Z(II31086) ) ;
AND4    gate18048  (.A(g32580), .B(g32581), .C(g32582), .D(g32583), .Z(II31087) ) ;
AND3    gate18049  (.A(g32584), .B(II31086), .C(II31087), .Z(g33478) ) ;
AND4    gate18050  (.A(g29385), .B(g32586), .C(g32587), .D(g32588), .Z(II31091) ) ;
AND4    gate18051  (.A(g32589), .B(g32590), .C(g32591), .D(g32592), .Z(II31092) ) ;
AND3    gate18052  (.A(g32593), .B(II31091), .C(II31092), .Z(g33479) ) ;
AND4    gate18053  (.A(g31376), .B(g31812), .C(g32594), .D(g32595), .Z(II31096) ) ;
AND4    gate18054  (.A(g32596), .B(g32597), .C(g32598), .D(g32599), .Z(II31097) ) ;
AND3    gate18055  (.A(g32600), .B(II31096), .C(II31097), .Z(g33480) ) ;
AND4    gate18056  (.A(g30735), .B(g31813), .C(g32601), .D(g32602), .Z(II31101) ) ;
AND4    gate18057  (.A(g32603), .B(g32604), .C(g32605), .D(g32606), .Z(II31102) ) ;
AND3    gate18058  (.A(g32607), .B(II31101), .C(II31102), .Z(g33481) ) ;
AND4    gate18059  (.A(g30825), .B(g31814), .C(g32608), .D(g32609), .Z(II31106) ) ;
AND4    gate18060  (.A(g32610), .B(g32611), .C(g32612), .D(g32613), .Z(II31107) ) ;
AND3    gate18061  (.A(g32614), .B(II31106), .C(II31107), .Z(g33482) ) ;
AND4    gate18062  (.A(g31070), .B(g31815), .C(g32615), .D(g32616), .Z(II31111) ) ;
AND4    gate18063  (.A(g32617), .B(g32618), .C(g32619), .D(g32620), .Z(II31112) ) ;
AND3    gate18064  (.A(g32621), .B(II31111), .C(II31112), .Z(g33483) ) ;
AND4    gate18065  (.A(g31154), .B(g31816), .C(g32622), .D(g32623), .Z(II31116) ) ;
AND4    gate18066  (.A(g32624), .B(g32625), .C(g32626), .D(g32627), .Z(II31117) ) ;
AND3    gate18067  (.A(g32628), .B(II31116), .C(II31117), .Z(g33484) ) ;
AND4    gate18068  (.A(g30614), .B(g31817), .C(g32629), .D(g32630), .Z(II31121) ) ;
AND4    gate18069  (.A(g32631), .B(g32632), .C(g32633), .D(g32634), .Z(II31122) ) ;
AND3    gate18070  (.A(g32635), .B(II31121), .C(II31122), .Z(g33485) ) ;
AND4    gate18071  (.A(g30673), .B(g31818), .C(g32636), .D(g32637), .Z(II31126) ) ;
AND4    gate18072  (.A(g32638), .B(g32639), .C(g32640), .D(g32641), .Z(II31127) ) ;
AND3    gate18073  (.A(g32642), .B(II31126), .C(II31127), .Z(g33486) ) ;
AND4    gate18074  (.A(g31542), .B(g31819), .C(g32643), .D(g32644), .Z(II31131) ) ;
AND4    gate18075  (.A(g32645), .B(g32646), .C(g32647), .D(g32648), .Z(II31132) ) ;
AND3    gate18076  (.A(g32649), .B(II31131), .C(II31132), .Z(g33487) ) ;
AND4    gate18077  (.A(g29385), .B(g32651), .C(g32652), .D(g32653), .Z(II31136) ) ;
AND4    gate18078  (.A(g32654), .B(g32655), .C(g32656), .D(g32657), .Z(II31137) ) ;
AND3    gate18079  (.A(g32658), .B(II31136), .C(II31137), .Z(g33488) ) ;
AND4    gate18080  (.A(g31376), .B(g31820), .C(g32659), .D(g32660), .Z(II31141) ) ;
AND4    gate18081  (.A(g32661), .B(g32662), .C(g32663), .D(g32664), .Z(II31142) ) ;
AND3    gate18082  (.A(g32665), .B(II31141), .C(II31142), .Z(g33489) ) ;
AND4    gate18083  (.A(g30735), .B(g31821), .C(g32666), .D(g32667), .Z(II31146) ) ;
AND4    gate18084  (.A(g32668), .B(g32669), .C(g32670), .D(g32671), .Z(II31147) ) ;
AND3    gate18085  (.A(g32672), .B(II31146), .C(II31147), .Z(g33490) ) ;
AND4    gate18086  (.A(g30825), .B(g31822), .C(g32673), .D(g32674), .Z(II31151) ) ;
AND4    gate18087  (.A(g32675), .B(g32676), .C(g32677), .D(g32678), .Z(II31152) ) ;
AND3    gate18088  (.A(g32679), .B(II31151), .C(II31152), .Z(g33491) ) ;
AND4    gate18089  (.A(g31070), .B(g31823), .C(g32680), .D(g32681), .Z(II31156) ) ;
AND4    gate18090  (.A(g32682), .B(g32683), .C(g32684), .D(g32685), .Z(II31157) ) ;
AND3    gate18091  (.A(g32686), .B(II31156), .C(II31157), .Z(g33492) ) ;
AND4    gate18092  (.A(g30614), .B(g31824), .C(g32687), .D(g32688), .Z(II31161) ) ;
AND4    gate18093  (.A(g32689), .B(g32690), .C(g32691), .D(g32692), .Z(II31162) ) ;
AND3    gate18094  (.A(g32693), .B(II31161), .C(II31162), .Z(g33493) ) ;
AND4    gate18095  (.A(g30673), .B(g31825), .C(g32694), .D(g32695), .Z(II31166) ) ;
AND4    gate18096  (.A(g32696), .B(g32697), .C(g32698), .D(g32699), .Z(II31167) ) ;
AND3    gate18097  (.A(g32700), .B(II31166), .C(II31167), .Z(g33494) ) ;
AND4    gate18098  (.A(g31528), .B(g31826), .C(g32701), .D(g32702), .Z(II31171) ) ;
AND4    gate18099  (.A(g32703), .B(g32704), .C(g32705), .D(g32706), .Z(II31172) ) ;
AND3    gate18100  (.A(g32707), .B(II31171), .C(II31172), .Z(g33495) ) ;
AND4    gate18101  (.A(g31579), .B(g31827), .C(g32708), .D(g32709), .Z(II31176) ) ;
AND4    gate18102  (.A(g32710), .B(g32711), .C(g32712), .D(g32713), .Z(II31177) ) ;
AND3    gate18103  (.A(g32714), .B(II31176), .C(II31177), .Z(g33496) ) ;
AND4    gate18104  (.A(g29385), .B(g32716), .C(g32717), .D(g32718), .Z(II31181) ) ;
AND4    gate18105  (.A(g32719), .B(g32720), .C(g32721), .D(g32722), .Z(II31182) ) ;
AND3    gate18106  (.A(g32723), .B(II31181), .C(II31182), .Z(g33497) ) ;
AND4    gate18107  (.A(g31376), .B(g31828), .C(g32724), .D(g32725), .Z(II31186) ) ;
AND4    gate18108  (.A(g32726), .B(g32727), .C(g32728), .D(g32729), .Z(II31187) ) ;
AND3    gate18109  (.A(g32730), .B(II31186), .C(II31187), .Z(g33498) ) ;
AND4    gate18110  (.A(g30735), .B(g31829), .C(g32731), .D(g32732), .Z(II31191) ) ;
AND4    gate18111  (.A(g32733), .B(g32734), .C(g32735), .D(g32736), .Z(II31192) ) ;
AND3    gate18112  (.A(g32737), .B(II31191), .C(II31192), .Z(g33499) ) ;
AND4    gate18113  (.A(g30825), .B(g31830), .C(g32738), .D(g32739), .Z(II31196) ) ;
AND4    gate18114  (.A(g32740), .B(g32741), .C(g32742), .D(g32743), .Z(II31197) ) ;
AND3    gate18115  (.A(g32744), .B(II31196), .C(II31197), .Z(g33500) ) ;
AND4    gate18116  (.A(g31672), .B(g31831), .C(g32745), .D(g32746), .Z(II31201) ) ;
AND4    gate18117  (.A(g32747), .B(g32748), .C(g32749), .D(g32750), .Z(II31202) ) ;
AND3    gate18118  (.A(g32751), .B(II31201), .C(II31202), .Z(g33501) ) ;
AND4    gate18119  (.A(g31710), .B(g31832), .C(g32752), .D(g32753), .Z(II31206) ) ;
AND4    gate18120  (.A(g32754), .B(g32755), .C(g32756), .D(g32757), .Z(II31207) ) ;
AND3    gate18121  (.A(g32758), .B(II31206), .C(II31207), .Z(g33502) ) ;
AND4    gate18122  (.A(g31021), .B(g31833), .C(g32759), .D(g32760), .Z(II31211) ) ;
AND4    gate18123  (.A(g32761), .B(g32762), .C(g32763), .D(g32764), .Z(II31212) ) ;
AND3    gate18124  (.A(g32765), .B(II31211), .C(II31212), .Z(g33503) ) ;
AND4    gate18125  (.A(g30937), .B(g31834), .C(g32766), .D(g32767), .Z(II31216) ) ;
AND4    gate18126  (.A(g32768), .B(g32769), .C(g32770), .D(g32771), .Z(II31217) ) ;
AND3    gate18127  (.A(g32772), .B(II31216), .C(II31217), .Z(g33504) ) ;
AND4    gate18128  (.A(g31327), .B(g31835), .C(g32773), .D(g32774), .Z(II31221) ) ;
AND4    gate18129  (.A(g32775), .B(g32776), .C(g32777), .D(g32778), .Z(II31222) ) ;
AND3    gate18130  (.A(g32779), .B(II31221), .C(II31222), .Z(g33505) ) ;
AND4    gate18131  (.A(g29385), .B(g32781), .C(g32782), .D(g32783), .Z(II31226) ) ;
AND4    gate18132  (.A(g32784), .B(g32785), .C(g32786), .D(g32787), .Z(II31227) ) ;
AND3    gate18133  (.A(g32788), .B(II31226), .C(II31227), .Z(g33506) ) ;
AND4    gate18134  (.A(g31376), .B(g31836), .C(g32789), .D(g32790), .Z(II31231) ) ;
AND4    gate18135  (.A(g32791), .B(g32792), .C(g32793), .D(g32794), .Z(II31232) ) ;
AND3    gate18136  (.A(g32795), .B(II31231), .C(II31232), .Z(g33507) ) ;
AND4    gate18137  (.A(g30735), .B(g31837), .C(g32796), .D(g32797), .Z(II31236) ) ;
AND4    gate18138  (.A(g32798), .B(g32799), .C(g32800), .D(g32801), .Z(II31237) ) ;
AND3    gate18139  (.A(g32802), .B(II31236), .C(II31237), .Z(g33508) ) ;
AND4    gate18140  (.A(g30825), .B(g31838), .C(g32803), .D(g32804), .Z(II31241) ) ;
AND4    gate18141  (.A(g32805), .B(g32806), .C(g32807), .D(g32808), .Z(II31242) ) ;
AND3    gate18142  (.A(g32809), .B(II31241), .C(II31242), .Z(g33509) ) ;
AND4    gate18143  (.A(g31672), .B(g31839), .C(g32810), .D(g32811), .Z(II31246) ) ;
AND4    gate18144  (.A(g32812), .B(g32813), .C(g32814), .D(g32815), .Z(II31247) ) ;
AND3    gate18145  (.A(g32816), .B(II31246), .C(II31247), .Z(g33510) ) ;
AND4    gate18146  (.A(g31710), .B(g31840), .C(g32817), .D(g32818), .Z(II31251) ) ;
AND4    gate18147  (.A(g32819), .B(g32820), .C(g32821), .D(g32822), .Z(II31252) ) ;
AND3    gate18148  (.A(g32823), .B(II31251), .C(II31252), .Z(g33511) ) ;
AND4    gate18149  (.A(g31021), .B(g31841), .C(g32824), .D(g32825), .Z(II31256) ) ;
AND4    gate18150  (.A(g32826), .B(g32827), .C(g32828), .D(g32829), .Z(II31257) ) ;
AND3    gate18151  (.A(g32830), .B(II31256), .C(II31257), .Z(g33512) ) ;
AND4    gate18152  (.A(g30937), .B(g31842), .C(g32831), .D(g32832), .Z(II31261) ) ;
AND4    gate18153  (.A(g32833), .B(g32834), .C(g32835), .D(g32836), .Z(II31262) ) ;
AND3    gate18154  (.A(g32837), .B(II31261), .C(II31262), .Z(g33513) ) ;
AND4    gate18155  (.A(g31327), .B(g31843), .C(g32838), .D(g32839), .Z(II31266) ) ;
AND4    gate18156  (.A(g32840), .B(g32841), .C(g32842), .D(g32843), .Z(II31267) ) ;
AND3    gate18157  (.A(g32844), .B(II31266), .C(II31267), .Z(g33514) ) ;
AND4    gate18158  (.A(g29385), .B(g32846), .C(g32847), .D(g32848), .Z(II31271) ) ;
AND4    gate18159  (.A(g32849), .B(g32850), .C(g32851), .D(g32852), .Z(II31272) ) ;
AND3    gate18160  (.A(g32853), .B(II31271), .C(II31272), .Z(g33515) ) ;
AND4    gate18161  (.A(g31376), .B(g31844), .C(g32854), .D(g32855), .Z(II31276) ) ;
AND4    gate18162  (.A(g32856), .B(g32857), .C(g32858), .D(g32859), .Z(II31277) ) ;
AND3    gate18163  (.A(g32860), .B(II31276), .C(II31277), .Z(g33516) ) ;
AND4    gate18164  (.A(g30735), .B(g31845), .C(g32861), .D(g32862), .Z(II31281) ) ;
AND4    gate18165  (.A(g32863), .B(g32864), .C(g32865), .D(g32866), .Z(II31282) ) ;
AND3    gate18166  (.A(g32867), .B(II31281), .C(II31282), .Z(g33517) ) ;
AND4    gate18167  (.A(g30825), .B(g31846), .C(g32868), .D(g32869), .Z(II31286) ) ;
AND4    gate18168  (.A(g32870), .B(g32871), .C(g32872), .D(g32873), .Z(II31287) ) ;
AND3    gate18169  (.A(g32874), .B(II31286), .C(II31287), .Z(g33518) ) ;
AND4    gate18170  (.A(g31021), .B(g31847), .C(g32875), .D(g32876), .Z(II31291) ) ;
AND4    gate18171  (.A(g32877), .B(g32878), .C(g32879), .D(g32880), .Z(II31292) ) ;
AND3    gate18172  (.A(g32881), .B(II31291), .C(II31292), .Z(g33519) ) ;
AND4    gate18173  (.A(g30937), .B(g31848), .C(g32882), .D(g32883), .Z(II31296) ) ;
AND4    gate18174  (.A(g32884), .B(g32885), .C(g32886), .D(g32887), .Z(II31297) ) ;
AND3    gate18175  (.A(g32888), .B(II31296), .C(II31297), .Z(g33520) ) ;
AND4    gate18176  (.A(g31327), .B(g31849), .C(g32889), .D(g32890), .Z(II31301) ) ;
AND4    gate18177  (.A(g32891), .B(g32892), .C(g32893), .D(g32894), .Z(II31302) ) ;
AND3    gate18178  (.A(g32895), .B(II31301), .C(II31302), .Z(g33521) ) ;
AND4    gate18179  (.A(g30614), .B(g31850), .C(g32896), .D(g32897), .Z(II31306) ) ;
AND4    gate18180  (.A(g32898), .B(g32899), .C(g32900), .D(g32901), .Z(II31307) ) ;
AND3    gate18181  (.A(g32902), .B(II31306), .C(II31307), .Z(g33522) ) ;
AND4    gate18182  (.A(g30673), .B(g31851), .C(g32903), .D(g32904), .Z(II31311) ) ;
AND4    gate18183  (.A(g32905), .B(g32906), .C(g32907), .D(g32908), .Z(II31312) ) ;
AND3    gate18184  (.A(g32909), .B(II31311), .C(II31312), .Z(g33523) ) ;
AND4    gate18185  (.A(g29385), .B(g32911), .C(g32912), .D(g32913), .Z(II31316) ) ;
AND4    gate18186  (.A(g32914), .B(g32915), .C(g32916), .D(g32917), .Z(II31317) ) ;
AND3    gate18187  (.A(g32918), .B(II31316), .C(II31317), .Z(g33524) ) ;
AND4    gate18188  (.A(g31376), .B(g31852), .C(g32919), .D(g32920), .Z(II31321) ) ;
AND4    gate18189  (.A(g32921), .B(g32922), .C(g32923), .D(g32924), .Z(II31322) ) ;
AND3    gate18190  (.A(g32925), .B(II31321), .C(II31322), .Z(g33525) ) ;
AND4    gate18191  (.A(g30735), .B(g31853), .C(g32926), .D(g32927), .Z(II31326) ) ;
AND4    gate18192  (.A(g32928), .B(g32929), .C(g32930), .D(g32931), .Z(II31327) ) ;
AND3    gate18193  (.A(g32932), .B(II31326), .C(II31327), .Z(g33526) ) ;
AND4    gate18194  (.A(g30825), .B(g31854), .C(g32933), .D(g32934), .Z(II31331) ) ;
AND4    gate18195  (.A(g32935), .B(g32936), .C(g32937), .D(g32938), .Z(II31332) ) ;
AND3    gate18196  (.A(g32939), .B(II31331), .C(II31332), .Z(g33527) ) ;
AND4    gate18197  (.A(g31672), .B(g31855), .C(g32940), .D(g32941), .Z(II31336) ) ;
AND4    gate18198  (.A(g32942), .B(g32943), .C(g32944), .D(g32945), .Z(II31337) ) ;
AND3    gate18199  (.A(g32946), .B(II31336), .C(II31337), .Z(g33528) ) ;
AND4    gate18200  (.A(g31710), .B(g31856), .C(g32947), .D(g32948), .Z(II31341) ) ;
AND4    gate18201  (.A(g32949), .B(g32950), .C(g32951), .D(g32952), .Z(II31342) ) ;
AND3    gate18202  (.A(g32953), .B(II31341), .C(II31342), .Z(g33529) ) ;
AND4    gate18203  (.A(g31021), .B(g31857), .C(g32954), .D(g32955), .Z(II31346) ) ;
AND4    gate18204  (.A(g32956), .B(g32957), .C(g32958), .D(g32959), .Z(II31347) ) ;
AND3    gate18205  (.A(g32960), .B(II31346), .C(II31347), .Z(g33530) ) ;
AND4    gate18206  (.A(g30937), .B(g31858), .C(g32961), .D(g32962), .Z(II31351) ) ;
AND4    gate18207  (.A(g32963), .B(g32964), .C(g32965), .D(g32966), .Z(II31352) ) ;
AND3    gate18208  (.A(g32967), .B(II31351), .C(II31352), .Z(g33531) ) ;
AND4    gate18209  (.A(g31327), .B(g31859), .C(g32968), .D(g32969), .Z(II31356) ) ;
AND4    gate18210  (.A(g32970), .B(g32971), .C(g32972), .D(g32973), .Z(II31357) ) ;
AND3    gate18211  (.A(g32974), .B(II31356), .C(II31357), .Z(g33532) ) ;
OR2     gate18212  (.A(g32258), .B(g29951), .Z(g33386) ) ;
AND2    gate18213  (.A(g33386), .B(g18829), .Z(g33639) ) ;
OR2     gate18214  (.A(g32263), .B(g29954), .Z(g33387) ) ;
AND2    gate18215  (.A(g33387), .B(g18831), .Z(g33640) ) ;
OR2     gate18216  (.A(g32272), .B(g29964), .Z(g33389) ) ;
AND2    gate18217  (.A(g33389), .B(g18876), .Z(g33646) ) ;
OR2     gate18218  (.A(g32276), .B(g29968), .Z(g33390) ) ;
AND2    gate18219  (.A(g33390), .B(g18878), .Z(g33647) ) ;
OR2     gate18220  (.A(g32286), .B(g29984), .Z(g33393) ) ;
AND2    gate18221  (.A(g33393), .B(g18889), .Z(g33652) ) ;
AND2    gate18222  (.A(g30991), .B(g33443), .Z(g33657) ) ;
NOR2    gate18223  (.A(g8606), .B(g32057), .Z(g33125) ) ;
AND2    gate18224  (.A(g33125), .B(g7970), .Z(g33676) ) ;
AND2    gate18225  (.A(g33443), .B(g31937), .Z(g33677) ) ;
NOR2    gate18226  (.A(g4653), .B(g32057), .Z(g33128) ) ;
AND2    gate18227  (.A(g33128), .B(g4688), .Z(g33680) ) ;
NOR2    gate18228  (.A(g8630), .B(g32072), .Z(g33129) ) ;
AND2    gate18229  (.A(g33129), .B(g7991), .Z(g33681) ) ;
NOR2    gate18230  (.A(g8650), .B(g32057), .Z(g33139) ) ;
AND2    gate18231  (.A(g33139), .B(g13565), .Z(g33684) ) ;
NOR2    gate18232  (.A(g4843), .B(g32072), .Z(g33132) ) ;
AND2    gate18233  (.A(g33132), .B(g4878), .Z(g33687) ) ;
NOR2    gate18234  (.A(g4664), .B(g32057), .Z(g33144) ) ;
AND2    gate18235  (.A(g33144), .B(g11006), .Z(g33689) ) ;
NOR2    gate18236  (.A(g4669), .B(g32057), .Z(g33146) ) ;
AND2    gate18237  (.A(g33146), .B(g16280), .Z(g33690) ) ;
NOR2    gate18238  (.A(g8677), .B(g32072), .Z(g33145) ) ;
AND2    gate18239  (.A(g33145), .B(g13594), .Z(g33693) ) ;
NOR2    gate18240  (.A(g8672), .B(g32057), .Z(g33160) ) ;
AND2    gate18241  (.A(g33160), .B(g13330), .Z(g33697) ) ;
NOR2    gate18242  (.A(g4854), .B(g32072), .Z(g33148) ) ;
AND2    gate18243  (.A(g33148), .B(g11012), .Z(g33700) ) ;
NOR2    gate18244  (.A(g4859), .B(g32072), .Z(g33162) ) ;
AND2    gate18245  (.A(g33162), .B(g16305), .Z(g33701) ) ;
NOR2    gate18246  (.A(g8714), .B(g32072), .Z(g33174) ) ;
AND2    gate18247  (.A(g33174), .B(g13346), .Z(g33707) ) ;
NOR2    gate18248  (.A(g8748), .B(g11083), .Z(g14037) ) ;
AND2    gate18249  (.A(g14037), .B(g33246), .Z(g33710) ) ;
NOR2    gate18250  (.A(g32090), .B(g8350), .Z(g33135) ) ;
AND2    gate18251  (.A(g33135), .B(g19416), .Z(g33715) ) ;
NOR2    gate18252  (.A(g8774), .B(g11083), .Z(g14092) ) ;
AND2    gate18253  (.A(g14092), .B(g33306), .Z(g33717) ) ;
NOR2    gate18254  (.A(g32090), .B(g7788), .Z(g33147) ) ;
AND2    gate18255  (.A(g33147), .B(g19432), .Z(g33718) ) ;
NOR2    gate18256  (.A(g32099), .B(g8400), .Z(g33141) ) ;
AND2    gate18257  (.A(g33141), .B(g19433), .Z(g33719) ) ;
NOR2    gate18258  (.A(g32090), .B(g7806), .Z(g33161) ) ;
AND2    gate18259  (.A(g33161), .B(g19439), .Z(g33720) ) ;
NOR2    gate18260  (.A(g32099), .B(g7809), .Z(g33163) ) ;
AND2    gate18261  (.A(g33163), .B(g19440), .Z(g33721) ) ;
NOR2    gate18262  (.A(g32099), .B(g7828), .Z(g33175) ) ;
AND2    gate18263  (.A(g33175), .B(g19445), .Z(g33722) ) ;
NOR2    gate18264  (.A(g8854), .B(g12259), .Z(g14091) ) ;
AND2    gate18265  (.A(g14091), .B(g33299), .Z(g33723) ) ;
NOR2    gate18266  (.A(g8945), .B(g12259), .Z(g14145) ) ;
AND2    gate18267  (.A(g14145), .B(g33258), .Z(g33724) ) ;
OR2     gate18268  (.A(g32397), .B(g32401), .Z(g33115) ) ;
AND2    gate18269  (.A(g33115), .B(g19499), .Z(g33727) ) ;
AND4    gate18270  (.A(g7202), .B(g4621), .C(g33127), .D(g4633), .Z(g33730) ) ;
OR2     gate18271  (.A(g32403), .B(g32411), .Z(g33116) ) ;
AND2    gate18272  (.A(g33116), .B(g19520), .Z(g33731) ) ;
AND3    gate18273  (.A(g31003), .B(g8350), .C(g7788), .Z(II31593) ) ;
AND3    gate18274  (.A(g7806), .B(g33136), .C(II31593), .Z(g33734) ) ;
OR2     gate18275  (.A(g32413), .B(g32418), .Z(g33118) ) ;
AND2    gate18276  (.A(g33118), .B(g19553), .Z(g33735) ) ;
AND3    gate18277  (.A(g31009), .B(g8400), .C(g7809), .Z(II31600) ) ;
AND3    gate18278  (.A(g7828), .B(g33142), .C(II31600), .Z(g33742) ) ;
OR2     gate18279  (.A(g32420), .B(g32428), .Z(g33119) ) ;
AND2    gate18280  (.A(g33119), .B(g19574), .Z(g33743) ) ;
NOR2    gate18281  (.A(g32278), .B(g31503), .Z(g33133) ) ;
AND2    gate18282  (.A(g33133), .B(g20269), .Z(g33758) ) ;
OR2     gate18283  (.A(g31962), .B(g30577), .Z(g33123) ) ;
AND2    gate18284  (.A(g33123), .B(g22847), .Z(g33759) ) ;
NOR2    gate18285  (.A(g32293), .B(g31518), .Z(g33143) ) ;
AND2    gate18286  (.A(g33143), .B(g20328), .Z(g33760) ) ;
NOR2    gate18287  (.A(g32180), .B(g31223), .Z(g33107) ) ;
AND2    gate18288  (.A(g33107), .B(g20531), .Z(g33784) ) ;
NOR2    gate18289  (.A(g32172), .B(g31188), .Z(g33100) ) ;
AND2    gate18290  (.A(g33100), .B(g20550), .Z(g33785) ) ;
NOR2    gate18291  (.A(g32265), .B(g31497), .Z(g33130) ) ;
AND2    gate18292  (.A(g33130), .B(g20572), .Z(g33786) ) ;
NOR2    gate18293  (.A(g32176), .B(g31212), .Z(g33103) ) ;
AND2    gate18294  (.A(g33103), .B(g20595), .Z(g33787) ) ;
OR2     gate18295  (.A(g32016), .B(g30730), .Z(g33159) ) ;
AND2    gate18296  (.A(g33159), .B(g23022), .Z(g33789) ) ;
NOR2    gate18297  (.A(g32183), .B(g31228), .Z(g33108) ) ;
AND2    gate18298  (.A(g33108), .B(g20643), .Z(g33790) ) ;
NOR2    gate18299  (.A(g32287), .B(g31514), .Z(g33138) ) ;
AND2    gate18300  (.A(g33138), .B(g20782), .Z(g33795) ) ;
NOR2    gate18301  (.A(g31261), .B(g32205), .Z(g33117) ) ;
AND2    gate18302  (.A(g33117), .B(g25267), .Z(g33796) ) ;
OR2     gate18303  (.A(g32029), .B(g32031), .Z(g33227) ) ;
AND2    gate18304  (.A(g33227), .B(g20058), .Z(g33798) ) ;
NOR2    gate18305  (.A(g31997), .B(g10275), .Z(g33437) ) ;
AND2    gate18306  (.A(g33437), .B(g25327), .Z(g33801) ) ;
NOR2    gate18307  (.A(g31950), .B(g4628), .Z(g33097) ) ;
AND2    gate18308  (.A(g33097), .B(g14545), .Z(g33802) ) ;
OR2     gate18309  (.A(g32032), .B(g32036), .Z(g33231) ) ;
AND2    gate18310  (.A(g33231), .B(g20071), .Z(g33803) ) ;
OR2     gate18311  (.A(g32034), .B(g30936), .Z(g33232) ) ;
AND2    gate18312  (.A(g33232), .B(g20079), .Z(g33805) ) ;
NOR2    gate18313  (.A(g31240), .B(g32194), .Z(g33112) ) ;
AND2    gate18314  (.A(g33112), .B(g25452), .Z(g33807) ) ;
NOR2    gate18315  (.A(g31997), .B(g4584), .Z(g33109) ) ;
AND2    gate18316  (.A(g33109), .B(g22161), .Z(g33808) ) ;
NOR2    gate18317  (.A(g31997), .B(g6978), .Z(g33432) ) ;
AND2    gate18318  (.A(g33432), .B(g30184), .Z(g33809) ) ;
NOR2    gate18319  (.A(g10278), .B(g31950), .Z(g33427) ) ;
AND2    gate18320  (.A(g33427), .B(g12768), .Z(g33810) ) ;
NOR2    gate18321  (.A(g31950), .B(g4633), .Z(g33439) ) ;
AND2    gate18322  (.A(g33439), .B(g17573), .Z(g33811) ) ;
NOR2    gate18323  (.A(g31997), .B(g4616), .Z(g33098) ) ;
AND2    gate18324  (.A(g33098), .B(g28144), .Z(g33814) ) ;
NOR2    gate18325  (.A(g10311), .B(g31950), .Z(g33449) ) ;
AND2    gate18326  (.A(g33449), .B(g12911), .Z(g33815) ) ;
OR2     gate18327  (.A(g32039), .B(g32043), .Z(g33234) ) ;
AND2    gate18328  (.A(g33234), .B(g20096), .Z(g33816) ) ;
OR2     gate18329  (.A(g32040), .B(g30982), .Z(g33235) ) ;
AND2    gate18330  (.A(g33235), .B(g20102), .Z(g33817) ) ;
OR2     gate18331  (.A(g32044), .B(g32045), .Z(g33236) ) ;
AND2    gate18332  (.A(g33236), .B(g20113), .Z(g33818) ) ;
NOR2    gate18333  (.A(g31997), .B(g7163), .Z(g33075) ) ;
AND2    gate18334  (.A(g33075), .B(g26830), .Z(g33820) ) ;
OR2     gate18335  (.A(g32048), .B(g32051), .Z(g33238) ) ;
AND2    gate18336  (.A(g33238), .B(g20153), .Z(g33821) ) ;
AND2    gate18337  (.A(g33385), .B(g20157), .Z(g33822) ) ;
NOR2    gate18338  (.A(g31997), .B(g4593), .Z(g33090) ) ;
AND2    gate18339  (.A(g33090), .B(g24411), .Z(g33828) ) ;
OR2     gate18340  (.A(g32052), .B(g32068), .Z(g33240) ) ;
AND2    gate18341  (.A(g33240), .B(g20164), .Z(g33829) ) ;
AND2    gate18342  (.A(g33382), .B(g20166), .Z(g33830) ) ;
NOR2    gate18343  (.A(g31997), .B(g7224), .Z(g33088) ) ;
AND2    gate18344  (.A(g33088), .B(g27991), .Z(g33832) ) ;
NOR2    gate18345  (.A(g31997), .B(g4601), .Z(g33093) ) ;
AND2    gate18346  (.A(g33093), .B(g25852), .Z(g33833) ) ;
NOR2    gate18347  (.A(g31997), .B(g7236), .Z(g33095) ) ;
AND2    gate18348  (.A(g33095), .B(g29172), .Z(g33834) ) ;
AND2    gate18349  (.A(g4340), .B(g33413), .Z(g33835) ) ;
NOR2    gate18350  (.A(g31997), .B(g4608), .Z(g33096) ) ;
AND2    gate18351  (.A(g33096), .B(g27020), .Z(g33836) ) ;
OR2     gate18352  (.A(g32096), .B(g29509), .Z(g33251) ) ;
AND2    gate18353  (.A(g33251), .B(g20233), .Z(g33837) ) ;
OR2     gate18354  (.A(g32103), .B(g29511), .Z(g33253) ) ;
AND2    gate18355  (.A(g33253), .B(g20267), .Z(g33840) ) ;
OR2     gate18356  (.A(g32104), .B(g29512), .Z(g33254) ) ;
AND2    gate18357  (.A(g33254), .B(g20268), .Z(g33841) ) ;
OR2     gate18358  (.A(g32106), .B(g29514), .Z(g33255) ) ;
AND2    gate18359  (.A(g33255), .B(g20322), .Z(g33842) ) ;
OR2     gate18360  (.A(g32107), .B(g29517), .Z(g33256) ) ;
AND2    gate18361  (.A(g33256), .B(g20325), .Z(g33843) ) ;
OR2     gate18362  (.A(g32108), .B(g29519), .Z(g33257) ) ;
AND2    gate18363  (.A(g33257), .B(g20327), .Z(g33844) ) ;
OR2     gate18364  (.A(g32109), .B(g29521), .Z(g33259) ) ;
AND2    gate18365  (.A(g33259), .B(g20380), .Z(g33846) ) ;
OR2     gate18366  (.A(g32110), .B(g29524), .Z(g33260) ) ;
AND2    gate18367  (.A(g33260), .B(g20383), .Z(g33847) ) ;
OR2     gate18368  (.A(g32111), .B(g29525), .Z(g33261) ) ;
AND2    gate18369  (.A(g33261), .B(g20384), .Z(g33848) ) ;
OR2     gate18370  (.A(g32112), .B(g29528), .Z(g33262) ) ;
AND2    gate18371  (.A(g33262), .B(g20387), .Z(g33849) ) ;
OR2     gate18372  (.A(g32113), .B(g29530), .Z(g33265) ) ;
AND2    gate18373  (.A(g33265), .B(g20441), .Z(g33855) ) ;
OR2     gate18374  (.A(g32114), .B(g29532), .Z(g33266) ) ;
AND2    gate18375  (.A(g33266), .B(g20442), .Z(g33856) ) ;
OR2     gate18376  (.A(g32115), .B(g29535), .Z(g33267) ) ;
AND2    gate18377  (.A(g33267), .B(g20445), .Z(g33857) ) ;
OR2     gate18378  (.A(g32116), .B(g29538), .Z(g33268) ) ;
AND2    gate18379  (.A(g33268), .B(g20448), .Z(g33858) ) ;
AND2    gate18380  (.A(g33426), .B(g10531), .Z(g33859) ) ;
OR2     gate18381  (.A(g32119), .B(g29547), .Z(g33270) ) ;
AND2    gate18382  (.A(g33270), .B(g20501), .Z(g33860) ) ;
OR2     gate18383  (.A(g32120), .B(g29549), .Z(g33271) ) ;
AND2    gate18384  (.A(g33271), .B(g20502), .Z(g33861) ) ;
OR2     gate18385  (.A(g32121), .B(g29551), .Z(g33272) ) ;
AND2    gate18386  (.A(g33272), .B(g20504), .Z(g33862) ) ;
OR2     gate18387  (.A(g32122), .B(g29553), .Z(g33273) ) ;
AND2    gate18388  (.A(g33273), .B(g20505), .Z(g33863) ) ;
OR2     gate18389  (.A(g32126), .B(g29563), .Z(g33274) ) ;
AND2    gate18390  (.A(g33274), .B(g20524), .Z(g33864) ) ;
OR2     gate18391  (.A(g32127), .B(g29564), .Z(g33275) ) ;
AND2    gate18392  (.A(g33275), .B(g20526), .Z(g33865) ) ;
OR2     gate18393  (.A(g32128), .B(g29566), .Z(g33276) ) ;
AND2    gate18394  (.A(g33276), .B(g20528), .Z(g33866) ) ;
OR2     gate18395  (.A(g32129), .B(g29568), .Z(g33277) ) ;
AND2    gate18396  (.A(g33277), .B(g20529), .Z(g33867) ) ;
OR2     gate18397  (.A(g32139), .B(g29572), .Z(g33278) ) ;
AND2    gate18398  (.A(g33278), .B(g20542), .Z(g33868) ) ;
OR2     gate18399  (.A(g32140), .B(g29573), .Z(g33279) ) ;
AND2    gate18400  (.A(g33279), .B(g20543), .Z(g33869) ) ;
OR2     gate18401  (.A(g32141), .B(g29574), .Z(g33280) ) ;
AND2    gate18402  (.A(g33280), .B(g20545), .Z(g33870) ) ;
OR2     gate18403  (.A(g32142), .B(g29576), .Z(g33281) ) ;
AND2    gate18404  (.A(g33281), .B(g20546), .Z(g33871) ) ;
OR2     gate18405  (.A(g32143), .B(g29577), .Z(g33282) ) ;
AND2    gate18406  (.A(g33282), .B(g20548), .Z(g33872) ) ;
OR2     gate18407  (.A(g32154), .B(g13477), .Z(g33291) ) ;
AND2    gate18408  (.A(g33291), .B(g20549), .Z(g33873) ) ;
OR2     gate18409  (.A(g32145), .B(g29585), .Z(g33286) ) ;
AND2    gate18410  (.A(g33286), .B(g20562), .Z(g33876) ) ;
OR2     gate18411  (.A(g32146), .B(g29586), .Z(g33287) ) ;
AND2    gate18412  (.A(g33287), .B(g20563), .Z(g33877) ) ;
OR2     gate18413  (.A(g32147), .B(g29587), .Z(g33288) ) ;
AND2    gate18414  (.A(g33288), .B(g20565), .Z(g33878) ) ;
OR2     gate18415  (.A(g32148), .B(g29588), .Z(g33289) ) ;
AND2    gate18416  (.A(g33289), .B(g20566), .Z(g33879) ) ;
OR2     gate18417  (.A(g32149), .B(g29589), .Z(g33290) ) ;
AND2    gate18418  (.A(g33290), .B(g20568), .Z(g33880) ) ;
OR2     gate18419  (.A(g32150), .B(g29601), .Z(g33292) ) ;
AND2    gate18420  (.A(g33292), .B(g20586), .Z(g33881) ) ;
OR2     gate18421  (.A(g32151), .B(g29602), .Z(g33293) ) ;
AND2    gate18422  (.A(g33293), .B(g20587), .Z(g33882) ) ;
OR2     gate18423  (.A(g32152), .B(g29604), .Z(g33294) ) ;
AND2    gate18424  (.A(g33294), .B(g20589), .Z(g33883) ) ;
OR2     gate18425  (.A(g32153), .B(g29605), .Z(g33295) ) ;
AND2    gate18426  (.A(g33295), .B(g20590), .Z(g33884) ) ;
OR2     gate18427  (.A(g32156), .B(g29617), .Z(g33296) ) ;
AND2    gate18428  (.A(g33296), .B(g20609), .Z(g33885) ) ;
OR2     gate18429  (.A(g32157), .B(g29621), .Z(g33297) ) ;
AND2    gate18430  (.A(g33297), .B(g20614), .Z(g33886) ) ;
OR2     gate18431  (.A(g32158), .B(g29622), .Z(g33298) ) ;
AND2    gate18432  (.A(g33298), .B(g20615), .Z(g33887) ) ;
OR2     gate18433  (.A(g32159), .B(g29638), .Z(g33303) ) ;
AND2    gate18434  (.A(g33303), .B(g20641), .Z(g33889) ) ;
OR2     gate18435  (.A(g29631), .B(g32165), .Z(g33310) ) ;
AND2    gate18436  (.A(g33310), .B(g20659), .Z(g33890) ) ;
OR2     gate18437  (.A(g29646), .B(g32170), .Z(g33312) ) ;
AND2    gate18438  (.A(g33312), .B(g20701), .Z(g33892) ) ;
OR2     gate18439  (.A(g29649), .B(g32171), .Z(g33313) ) ;
AND2    gate18440  (.A(g33313), .B(g20706), .Z(g33893) ) ;
OR2     gate18441  (.A(g29663), .B(g32174), .Z(g33314) ) ;
AND2    gate18442  (.A(g33314), .B(g20771), .Z(g33896) ) ;
OR2     gate18443  (.A(g29665), .B(g32175), .Z(g33315) ) ;
AND2    gate18444  (.A(g33315), .B(g20777), .Z(g33897) ) ;
NOR2    gate18445  (.A(g31978), .B(g7627), .Z(g33419) ) ;
AND2    gate18446  (.A(g33419), .B(g15655), .Z(g33898) ) ;
AND2    gate18447  (.A(g32132), .B(g33335), .Z(g33899) ) ;
OR2     gate18448  (.A(g29685), .B(g32178), .Z(g33316) ) ;
AND2    gate18449  (.A(g33316), .B(g20913), .Z(g33900) ) ;
OR2     gate18450  (.A(g29688), .B(g32179), .Z(g33317) ) ;
AND2    gate18451  (.A(g33317), .B(g20920), .Z(g33901) ) ;
NOR2    gate18452  (.A(g31978), .B(g4311), .Z(g33085) ) ;
AND2    gate18453  (.A(g33085), .B(g13202), .Z(g33902) ) ;
NOR2    gate18454  (.A(g31978), .B(g7643), .Z(g33447) ) ;
AND2    gate18455  (.A(g33447), .B(g19146), .Z(g33903) ) ;
OR2     gate18456  (.A(g29712), .B(g32182), .Z(g33321) ) ;
AND2    gate18457  (.A(g33321), .B(g21059), .Z(g33904) ) ;
NOR2    gate18458  (.A(g31978), .B(g4322), .Z(g33089) ) ;
AND2    gate18459  (.A(g33089), .B(g15574), .Z(g33905) ) ;
NOR2    gate18460  (.A(g31978), .B(g7655), .Z(g33084) ) ;
AND2    gate18461  (.A(g33084), .B(g22311), .Z(g33906) ) ;
NOR2    gate18462  (.A(g31978), .B(g4332), .Z(g33092) ) ;
AND2    gate18463  (.A(g33092), .B(g18935), .Z(g33908) ) ;
NOR2    gate18464  (.A(g4659), .B(g32057), .Z(g33131) ) ;
AND2    gate18465  (.A(g33131), .B(g10708), .Z(g33909) ) ;
NOR2    gate18466  (.A(g7686), .B(g32057), .Z(g33134) ) ;
AND2    gate18467  (.A(g33134), .B(g7836), .Z(g33910) ) ;
NOR2    gate18468  (.A(g4849), .B(g32072), .Z(g33137) ) ;
AND2    gate18469  (.A(g33137), .B(g10725), .Z(g33911) ) ;
NOR2    gate18470  (.A(g7693), .B(g32072), .Z(g33140) ) ;
AND2    gate18471  (.A(g33140), .B(g7846), .Z(g33915) ) ;
NOR2    gate18472  (.A(g31950), .B(g4621), .Z(g33438) ) ;
AND2    gate18473  (.A(g33438), .B(g10795), .Z(g33919) ) ;
NOR2    gate18474  (.A(g7785), .B(g31950), .Z(g33448) ) ;
AND2    gate18475  (.A(g33448), .B(g7202), .Z(g33922) ) ;
AND2    gate18476  (.A(g33335), .B(g33346), .Z(g33924) ) ;
NOR2    gate18477  (.A(g31950), .B(g4639), .Z(g33094) ) ;
AND2    gate18478  (.A(g33094), .B(g21412), .Z(g33927) ) ;
OR2     gate18479  (.A(g32234), .B(g29926), .Z(g33380) ) ;
AND2    gate18480  (.A(g33380), .B(g21560), .Z(g33941) ) ;
OR2     gate18481  (.A(g32244), .B(g29940), .Z(g33383) ) ;
AND2    gate18482  (.A(g33383), .B(g21608), .Z(g33942) ) ;
OR2     gate18483  (.A(g32248), .B(g29943), .Z(g33384) ) ;
AND2    gate18484  (.A(g33384), .B(g21609), .Z(g33943) ) ;
AND2    gate18485  (.A(g33766), .B(g22942), .Z(g34045) ) ;
AND2    gate18486  (.A(g33772), .B(g22942), .Z(g34050) ) ;
AND2    gate18487  (.A(g33778), .B(g22942), .Z(g34054) ) ;
AND2    gate18488  (.A(g33800), .B(g23076), .Z(g34061) ) ;
AND2    gate18489  (.A(g33806), .B(g23121), .Z(g34063) ) ;
AND2    gate18490  (.A(g33813), .B(g23148), .Z(g34065) ) ;
AND2    gate18491  (.A(g33730), .B(g19352), .Z(g34066) ) ;
AND2    gate18492  (.A(g8774), .B(g33797), .Z(g34069) ) ;
AND2    gate18493  (.A(g8854), .B(g33799), .Z(g34071) ) ;
AND2    gate18494  (.A(g33839), .B(g24872), .Z(g34072) ) ;
AND2    gate18495  (.A(g8948), .B(g33823), .Z(g34073) ) ;
OR2     gate18496  (.A(g32396), .B(g33423), .Z(g33685) ) ;
AND2    gate18497  (.A(g33685), .B(g19498), .Z(g34074) ) ;
OR2     gate18498  (.A(g32400), .B(g33428), .Z(g33692) ) ;
AND2    gate18499  (.A(g33692), .B(g19517), .Z(g34075) ) ;
OR2     gate18500  (.A(g32402), .B(g33429), .Z(g33694) ) ;
AND2    gate18501  (.A(g33694), .B(g19519), .Z(g34076) ) ;
OR2     gate18502  (.A(g32409), .B(g33433), .Z(g33699) ) ;
AND2    gate18503  (.A(g33699), .B(g19531), .Z(g34078) ) ;
OR2     gate18504  (.A(g32410), .B(g33434), .Z(g33703) ) ;
AND2    gate18505  (.A(g33703), .B(g19532), .Z(g34079) ) ;
OR2     gate18506  (.A(g32412), .B(g33440), .Z(g33706) ) ;
AND2    gate18507  (.A(g33706), .B(g19552), .Z(g34081) ) ;
OR2     gate18508  (.A(g32414), .B(g33441), .Z(g33709) ) ;
AND2    gate18509  (.A(g33709), .B(g19554), .Z(g34082) ) ;
OR2     gate18510  (.A(g32419), .B(g33450), .Z(g33714) ) ;
AND2    gate18511  (.A(g33714), .B(g19573), .Z(g34083) ) ;
AND2    gate18512  (.A(g9214), .B(g33851), .Z(g34084) ) ;
AND2    gate18513  (.A(g33912), .B(g23599), .Z(g34102) ) ;
AND2    gate18514  (.A(g33916), .B(g23639), .Z(g34104) ) ;
AND2    gate18515  (.A(g33917), .B(g23675), .Z(g34106) ) ;
AND2    gate18516  (.A(g33918), .B(g23708), .Z(g34109) ) ;
OR2     gate18517  (.A(g33104), .B(g32011), .Z(g33732) ) ;
AND2    gate18518  (.A(g33732), .B(g22935), .Z(g34110) ) ;
OR2     gate18519  (.A(g33105), .B(g32012), .Z(g33733) ) ;
AND2    gate18520  (.A(g33733), .B(g22936), .Z(g34111) ) ;
AND2    gate18521  (.A(g33734), .B(g19744), .Z(g34113) ) ;
AND2    gate18522  (.A(g33920), .B(g23742), .Z(g34114) ) ;
NAND4   gate18523  (.A(g33394), .B(g12491), .C(g12819), .D(g12796), .Z(g33933) ) ;
AND2    gate18524  (.A(g33933), .B(g25140), .Z(g34116) ) ;
AND2    gate18525  (.A(g33742), .B(g19755), .Z(g34117) ) ;
NAND3   gate18526  (.A(g33394), .B(g12767), .C(g9848), .Z(g33930) ) ;
AND2    gate18527  (.A(g33930), .B(g25158), .Z(g34120) ) ;
AND2    gate18528  (.A(g33845), .B(g23958), .Z(g34133) ) ;
AND2    gate18529  (.A(g33926), .B(g23802), .Z(g34135) ) ;
AND2    gate18530  (.A(g33850), .B(g23293), .Z(g34136) ) ;
AND2    gate18531  (.A(g33928), .B(g23802), .Z(g34137) ) ;
AND2    gate18532  (.A(g33929), .B(g23828), .Z(g34138) ) ;
AND2    gate18533  (.A(g33827), .B(g23314), .Z(g34139) ) ;
AND2    gate18534  (.A(g33931), .B(g23802), .Z(g34140) ) ;
AND2    gate18535  (.A(g33932), .B(g23828), .Z(g34141) ) ;
AND2    gate18536  (.A(g33934), .B(g23828), .Z(g34143) ) ;
OR2     gate18537  (.A(g33122), .B(g32041), .Z(g33788) ) ;
AND2    gate18538  (.A(g33788), .B(g20091), .Z(g34146) ) ;
OR2     gate18539  (.A(g33126), .B(g32053), .Z(g33794) ) ;
AND2    gate18540  (.A(g33794), .B(g20159), .Z(g34157) ) ;
NAND3   gate18541  (.A(g33394), .B(g4462), .C(g4467), .Z(g33925) ) ;
AND2    gate18542  (.A(g33925), .B(g24360), .Z(g34171) ) ;
NAND3   gate18543  (.A(g33394), .B(g10737), .C(g10308), .Z(g33679) ) ;
AND2    gate18544  (.A(g33679), .B(g24368), .Z(g34173) ) ;
AND2    gate18545  (.A(g33712), .B(g24361), .Z(g34178) ) ;
AND2    gate18546  (.A(g33686), .B(g24372), .Z(g34179) ) ;
AND2    gate18547  (.A(g33716), .B(g24373), .Z(g34180) ) ;
AND2    gate18548  (.A(g33691), .B(g24384), .Z(g34182) ) ;
AND2    gate18549  (.A(g33695), .B(g24385), .Z(g34183) ) ;
AND2    gate18550  (.A(g33698), .B(g24388), .Z(g34184) ) ;
AND2    gate18551  (.A(g33702), .B(g24389), .Z(g34185) ) ;
AND2    gate18552  (.A(g33705), .B(g24396), .Z(g34186) ) ;
AND2    gate18553  (.A(g33708), .B(g24397), .Z(g34187) ) ;
AND2    gate18554  (.A(g33713), .B(g24404), .Z(g34191) ) ;
AND2    gate18555  (.A(g33682), .B(g24485), .Z(g34196) ) ;
AND2    gate18556  (.A(g33688), .B(g24491), .Z(g34198) ) ;
AND2    gate18557  (.A(g33726), .B(g24537), .Z(g34203) ) ;
AND2    gate18558  (.A(g33729), .B(g24541), .Z(g34205) ) ;
OR2     gate18559  (.A(g33264), .B(g33269), .Z(g33891) ) ;
AND2    gate18560  (.A(g33891), .B(g21349), .Z(g34211) ) ;
AND2    gate18561  (.A(g33761), .B(g22689), .Z(g34212) ) ;
AND2    gate18562  (.A(g33766), .B(g22689), .Z(g34213) ) ;
AND2    gate18563  (.A(g33772), .B(g22689), .Z(g34214) ) ;
AND2    gate18564  (.A(g33778), .B(g22670), .Z(g34215) ) ;
AND2    gate18565  (.A(g33778), .B(g22689), .Z(g34216) ) ;
AND2    gate18566  (.A(g33736), .B(g22876), .Z(g34217) ) ;
AND2    gate18567  (.A(g33744), .B(g22670), .Z(g34218) ) ;
AND2    gate18568  (.A(g33736), .B(g22942), .Z(g34219) ) ;
AND2    gate18569  (.A(g33744), .B(g22876), .Z(g34223) ) ;
AND2    gate18570  (.A(g33736), .B(g22670), .Z(g34224) ) ;
AND2    gate18571  (.A(g33744), .B(g22942), .Z(g34225) ) ;
OR2     gate18572  (.A(g33305), .B(g33311), .Z(g33914) ) ;
AND2    gate18573  (.A(g33914), .B(g21467), .Z(g34226) ) ;
AND2    gate18574  (.A(g33750), .B(g22942), .Z(g34228) ) ;
AND2    gate18575  (.A(g33761), .B(g22942), .Z(g34230) ) ;
OR2     gate18576  (.A(g33898), .B(g33902), .Z(g34231) ) ;
AND2    gate18577  (.A(g34231), .B(g19208), .Z(g34279) ) ;
OR2     gate18578  (.A(g33903), .B(g33905), .Z(g34043) ) ;
AND2    gate18579  (.A(g34043), .B(g19276), .Z(g34281) ) ;
OR2     gate18580  (.A(g33906), .B(g33908), .Z(g34046) ) ;
AND2    gate18581  (.A(g34046), .B(g19351), .Z(g34284) ) ;
OR2     gate18582  (.A(g8807), .B(g550), .Z(g11370) ) ;
OR2     gate18583  (.A(g33909), .B(g33910), .Z(g34055) ) ;
AND2    gate18584  (.A(g34055), .B(g19366), .Z(g34291) ) ;
OR2     gate18585  (.A(g33911), .B(g33915), .Z(g34057) ) ;
AND2    gate18586  (.A(g34057), .B(g19370), .Z(g34295) ) ;
OR2     gate18587  (.A(g222), .B(g199), .Z(g8679) ) ;
OR2     gate18588  (.A(g33919), .B(g33922), .Z(g34064) ) ;
AND2    gate18589  (.A(g34064), .B(g19415), .Z(g34301) ) ;
NOR2    gate18590  (.A(g8948), .B(g11083), .Z(g13947) ) ;
AND2    gate18591  (.A(g13947), .B(g34147), .Z(g34309) ) ;
NOR2    gate18592  (.A(g9003), .B(g11083), .Z(g14003) ) ;
AND2    gate18593  (.A(g14003), .B(g34162), .Z(g34310) ) ;
OR2     gate18594  (.A(g209), .B(g538), .Z(g9535) ) ;
NOR2    gate18595  (.A(g9162), .B(g12259), .Z(g14188) ) ;
AND2    gate18596  (.A(g14188), .B(g34174), .Z(g34322) ) ;
NOR2    gate18597  (.A(g9214), .B(g12259), .Z(g14064) ) ;
AND2    gate18598  (.A(g14064), .B(g34161), .Z(g34324) ) ;
OR2     gate18599  (.A(g10685), .B(g546), .Z(g14511) ) ;
OR2     gate18600  (.A(g4300), .B(g4242), .Z(g9984) ) ;
OR2     gate18601  (.A(g33676), .B(g33680), .Z(g34090) ) ;
AND2    gate18602  (.A(g34090), .B(g19865), .Z(g34334) ) ;
OR2     gate18603  (.A(g301), .B(g534), .Z(g8461) ) ;
OR2     gate18604  (.A(g33681), .B(g33687), .Z(g34095) ) ;
AND2    gate18605  (.A(g34095), .B(g19881), .Z(g34337) ) ;
OR2     gate18606  (.A(g33684), .B(g33689), .Z(g34099) ) ;
AND2    gate18607  (.A(g34099), .B(g19905), .Z(g34338) ) ;
OR2     gate18608  (.A(g33690), .B(g33697), .Z(g34100) ) ;
AND2    gate18609  (.A(g34100), .B(g19950), .Z(g34340) ) ;
OR2     gate18610  (.A(g33693), .B(g33700), .Z(g34101) ) ;
AND2    gate18611  (.A(g34101), .B(g19952), .Z(g34341) ) ;
OR2     gate18612  (.A(g33701), .B(g33707), .Z(g34103) ) ;
AND2    gate18613  (.A(g34103), .B(g19998), .Z(g34342) ) ;
OR2     gate18614  (.A(g33710), .B(g33121), .Z(g34107) ) ;
AND2    gate18615  (.A(g34107), .B(g20038), .Z(g34344) ) ;
OR2     gate18616  (.A(g33724), .B(g33124), .Z(g34125) ) ;
AND2    gate18617  (.A(g34125), .B(g20128), .Z(g34348) ) ;
OR2     gate18618  (.A(g33758), .B(g19656), .Z(g34148) ) ;
AND2    gate18619  (.A(g34148), .B(g20389), .Z(g34363) ) ;
NAND3   gate18620  (.A(g33669), .B(g10583), .C(g7442), .Z(g34048) ) ;
AND2    gate18621  (.A(g34048), .B(g24366), .Z(g34364) ) ;
OR2     gate18622  (.A(g33760), .B(g19674), .Z(g34149) ) ;
AND2    gate18623  (.A(g34149), .B(g20451), .Z(g34365) ) ;
OR2     gate18624  (.A(g933), .B(g939), .Z(g7404) ) ;
NOR2    gate18625  (.A(g33859), .B(g11772), .Z(g34067) ) ;
AND2    gate18626  (.A(g34067), .B(g10554), .Z(g34370) ) ;
OR2     gate18627  (.A(g1277), .B(g1283), .Z(g7450) ) ;
OR2     gate18628  (.A(g11330), .B(g943), .Z(g13077) ) ;
OR2     gate18629  (.A(g11374), .B(g1287), .Z(g13095) ) ;
OR2     gate18630  (.A(g33784), .B(g19740), .Z(g34158) ) ;
AND2    gate18631  (.A(g34158), .B(g20571), .Z(g34380) ) ;
OR2     gate18632  (.A(g33785), .B(g19752), .Z(g34166) ) ;
AND2    gate18633  (.A(g34166), .B(g20594), .Z(g34381) ) ;
OR2     gate18634  (.A(g33786), .B(g19768), .Z(g34167) ) ;
AND2    gate18635  (.A(g34167), .B(g20618), .Z(g34382) ) ;
OR2     gate18636  (.A(g33787), .B(g19784), .Z(g34168) ) ;
AND2    gate18637  (.A(g34168), .B(g20642), .Z(g34385) ) ;
OR2     gate18638  (.A(g7517), .B(g952), .Z(g10800) ) ;
OR2     gate18639  (.A(g7533), .B(g1296), .Z(g10802) ) ;
OR2     gate18640  (.A(g33790), .B(g19855), .Z(g34170) ) ;
AND2    gate18641  (.A(g34170), .B(g20715), .Z(g34389) ) ;
OR2     gate18642  (.A(g33795), .B(g19914), .Z(g34172) ) ;
AND2    gate18643  (.A(g34172), .B(g21069), .Z(g34390) ) ;
OR2     gate18644  (.A(g33801), .B(g33808), .Z(g34189) ) ;
AND2    gate18645  (.A(g34189), .B(g21304), .Z(g34393) ) ;
OR2     gate18646  (.A(g33802), .B(g33810), .Z(g34190) ) ;
AND2    gate18647  (.A(g34190), .B(g21305), .Z(g34394) ) ;
OR2     gate18648  (.A(g33809), .B(g33814), .Z(g34193) ) ;
AND2    gate18649  (.A(g34193), .B(g21336), .Z(g34395) ) ;
OR2     gate18650  (.A(g33811), .B(g33815), .Z(g34194) ) ;
AND2    gate18651  (.A(g34194), .B(g21337), .Z(g34396) ) ;
OR2     gate18652  (.A(g4153), .B(g4172), .Z(g7673) ) ;
OR2     gate18653  (.A(g4072), .B(g4176), .Z(g7684) ) ;
OR2     gate18654  (.A(g33820), .B(g33828), .Z(g34199) ) ;
AND2    gate18655  (.A(g34199), .B(g21383), .Z(g34401) ) ;
OR2     gate18656  (.A(g33832), .B(g33833), .Z(g34204) ) ;
AND2    gate18657  (.A(g34204), .B(g21427), .Z(g34410) ) ;
AND2    gate18658  (.A(g34094), .B(g22670), .Z(g34413) ) ;
OR2     gate18659  (.A(g33834), .B(g33836), .Z(g34206) ) ;
AND2    gate18660  (.A(g34206), .B(g21457), .Z(g34414) ) ;
OR2     gate18661  (.A(g33835), .B(g33304), .Z(g34207) ) ;
AND2    gate18662  (.A(g34207), .B(g21458), .Z(g34415) ) ;
OR2     gate18663  (.A(g2886), .B(g2946), .Z(g7834) ) ;
OR2     gate18664  (.A(g2902), .B(g17058), .Z(g20083) ) ;
OR2     gate18665  (.A(g2917), .B(g26483), .Z(g27450) ) ;
OR2     gate18666  (.A(g34178), .B(g25067), .Z(g34399) ) ;
AND2    gate18667  (.A(g34399), .B(g18891), .Z(g34476) ) ;
OR2     gate18668  (.A(g2927), .B(g25010), .Z(g26344) ) ;
OR2     gate18669  (.A(g34179), .B(g25084), .Z(g34402) ) ;
AND2    gate18670  (.A(g34402), .B(g18904), .Z(g34478) ) ;
OR2     gate18671  (.A(g34180), .B(g25085), .Z(g34403) ) ;
AND2    gate18672  (.A(g34403), .B(g18905), .Z(g34479) ) ;
OR2     gate18673  (.A(g34182), .B(g25102), .Z(g34404) ) ;
AND2    gate18674  (.A(g34404), .B(g18916), .Z(g34481) ) ;
OR2     gate18675  (.A(g34183), .B(g25103), .Z(g34405) ) ;
AND2    gate18676  (.A(g34405), .B(g18917), .Z(g34482) ) ;
OR2     gate18677  (.A(g34184), .B(g25123), .Z(g34406) ) ;
AND2    gate18678  (.A(g34406), .B(g18938), .Z(g34483) ) ;
OR2     gate18679  (.A(g34185), .B(g25124), .Z(g34407) ) ;
AND2    gate18680  (.A(g34407), .B(g18939), .Z(g34484) ) ;
OR2     gate18681  (.A(g34186), .B(g25142), .Z(g34411) ) ;
AND2    gate18682  (.A(g34411), .B(g18952), .Z(g34485) ) ;
OR2     gate18683  (.A(g34187), .B(g25143), .Z(g34412) ) ;
AND2    gate18684  (.A(g34412), .B(g18953), .Z(g34486) ) ;
OR2     gate18685  (.A(g34191), .B(g25159), .Z(g34416) ) ;
AND2    gate18686  (.A(g34416), .B(g18983), .Z(g34487) ) ;
OR2     gate18687  (.A(g27678), .B(g34196), .Z(g34417) ) ;
AND2    gate18688  (.A(g34417), .B(g18988), .Z(g34488) ) ;
OR2     gate18689  (.A(g27686), .B(g34198), .Z(g34421) ) ;
AND2    gate18690  (.A(g34421), .B(g19068), .Z(g34489) ) ;
AND2    gate18691  (.A(g34272), .B(g33430), .Z(g34492) ) ;
OR2     gate18692  (.A(g27765), .B(g34203), .Z(g34273) ) ;
AND2    gate18693  (.A(g34273), .B(g19360), .Z(g34493) ) ;
OR2     gate18694  (.A(g27822), .B(g34205), .Z(g34274) ) ;
AND2    gate18695  (.A(g34274), .B(g19365), .Z(g34495) ) ;
AND2    gate18696  (.A(g34275), .B(g33072), .Z(g34497) ) ;
OR2     gate18697  (.A(g2941), .B(g11691), .Z(g13888) ) ;
OR2     gate18698  (.A(g2955), .B(g29914), .Z(g31288) ) ;
AND2    gate18699  (.A(g34276), .B(g30568), .Z(g34500) ) ;
OR2     gate18700  (.A(g2965), .B(g24965), .Z(g26363) ) ;
OR2     gate18701  (.A(g26829), .B(g34212), .Z(g34278) ) ;
AND2    gate18702  (.A(g34278), .B(g19437), .Z(g34503) ) ;
AND2    gate18703  (.A(g8833), .B(g34354), .Z(g34506) ) ;
OR2     gate18704  (.A(g26833), .B(g34213), .Z(g34280) ) ;
AND2    gate18705  (.A(g34280), .B(g19454), .Z(g34507) ) ;
OR2     gate18706  (.A(g26838), .B(g34214), .Z(g34282) ) ;
AND2    gate18707  (.A(g34282), .B(g19472), .Z(g34508) ) ;
OR2     gate18708  (.A(g26839), .B(g34215), .Z(g34283) ) ;
AND2    gate18709  (.A(g34283), .B(g19473), .Z(g34509) ) ;
AND2    gate18710  (.A(g9003), .B(g34346), .Z(g34513) ) ;
OR2     gate18711  (.A(g26842), .B(g34216), .Z(g34286) ) ;
AND2    gate18712  (.A(g34286), .B(g19480), .Z(g34514) ) ;
OR2     gate18713  (.A(g26846), .B(g34217), .Z(g34288) ) ;
AND2    gate18714  (.A(g34288), .B(g19491), .Z(g34515) ) ;
OR2     gate18715  (.A(g26847), .B(g34218), .Z(g34289) ) ;
AND2    gate18716  (.A(g34289), .B(g19492), .Z(g34516) ) ;
OR2     gate18717  (.A(g26848), .B(g34219), .Z(g34290) ) ;
AND2    gate18718  (.A(g34290), .B(g19493), .Z(g34517) ) ;
OR2     gate18719  (.A(g26853), .B(g34223), .Z(g34292) ) ;
AND2    gate18720  (.A(g34292), .B(g19503), .Z(g34518) ) ;
OR2     gate18721  (.A(g26854), .B(g34224), .Z(g34293) ) ;
AND2    gate18722  (.A(g34293), .B(g19504), .Z(g34519) ) ;
OR2     gate18723  (.A(g26855), .B(g34225), .Z(g34294) ) ;
AND2    gate18724  (.A(g34294), .B(g19505), .Z(g34520) ) ;
AND2    gate18725  (.A(g9162), .B(g34351), .Z(g34523) ) ;
AND2    gate18726  (.A(g9083), .B(g34359), .Z(g34524) ) ;
OR2     gate18727  (.A(g26858), .B(g34228), .Z(g34297) ) ;
AND2    gate18728  (.A(g34297), .B(g19528), .Z(g34525) ) ;
OR2     gate18729  (.A(g26864), .B(g34230), .Z(g34300) ) ;
AND2    gate18730  (.A(g34300), .B(g19569), .Z(g34526) ) ;
OR2     gate18731  (.A(g25768), .B(g34045), .Z(g34303) ) ;
AND2    gate18732  (.A(g34303), .B(g19603), .Z(g34527) ) ;
OR2     gate18733  (.A(g25775), .B(g34050), .Z(g34305) ) ;
AND2    gate18734  (.A(g34305), .B(g19617), .Z(g34528) ) ;
OR2     gate18735  (.A(g25782), .B(g34054), .Z(g34306) ) ;
AND2    gate18736  (.A(g34306), .B(g19634), .Z(g34529) ) ;
OR2     gate18737  (.A(g25831), .B(g34061), .Z(g34314) ) ;
AND2    gate18738  (.A(g34314), .B(g19710), .Z(g34532) ) ;
OR2     gate18739  (.A(g25850), .B(g34063), .Z(g34318) ) ;
AND2    gate18740  (.A(g34318), .B(g19731), .Z(g34533) ) ;
OR2     gate18741  (.A(g25866), .B(g34065), .Z(g34321) ) ;
AND2    gate18742  (.A(g34321), .B(g19743), .Z(g34534) ) ;
OR2     gate18743  (.A(g34069), .B(g33717), .Z(g34330) ) ;
AND2    gate18744  (.A(g34330), .B(g20054), .Z(g34538) ) ;
OR2     gate18745  (.A(g27121), .B(g34072), .Z(g34331) ) ;
AND2    gate18746  (.A(g34331), .B(g20087), .Z(g34541) ) ;
OR2     gate18747  (.A(g34071), .B(g33723), .Z(g34332) ) ;
AND2    gate18748  (.A(g34332), .B(g20089), .Z(g34542) ) ;
OR2     gate18749  (.A(g25986), .B(g34102), .Z(g34347) ) ;
AND2    gate18750  (.A(g34347), .B(g20495), .Z(g34554) ) ;
OR2     gate18751  (.A(g26019), .B(g34104), .Z(g34349) ) ;
AND2    gate18752  (.A(g34349), .B(g20512), .Z(g34555) ) ;
OR2     gate18753  (.A(g26048), .B(g34106), .Z(g34350) ) ;
AND2    gate18754  (.A(g34350), .B(g20537), .Z(g34556) ) ;
OR2     gate18755  (.A(g26079), .B(g34109), .Z(g34352) ) ;
AND2    gate18756  (.A(g34352), .B(g20555), .Z(g34557) ) ;
OR2     gate18757  (.A(g26088), .B(g34114), .Z(g34353) ) ;
AND2    gate18758  (.A(g34353), .B(g20578), .Z(g34558) ) ;
OR2     gate18759  (.A(g26257), .B(g34133), .Z(g34366) ) ;
AND2    gate18760  (.A(g34366), .B(g17366), .Z(g34560) ) ;
OR2     gate18761  (.A(g26274), .B(g34135), .Z(g34368) ) ;
AND2    gate18762  (.A(g34368), .B(g17410), .Z(g34561) ) ;
OR2     gate18763  (.A(g26279), .B(g34136), .Z(g34369) ) ;
AND2    gate18764  (.A(g34369), .B(g17411), .Z(g34562) ) ;
OR2     gate18765  (.A(g26287), .B(g34137), .Z(g34372) ) ;
AND2    gate18766  (.A(g34372), .B(g17465), .Z(g34563) ) ;
OR2     gate18767  (.A(g26292), .B(g34138), .Z(g34373) ) ;
AND2    gate18768  (.A(g34373), .B(g17466), .Z(g34564) ) ;
OR2     gate18769  (.A(g26294), .B(g34139), .Z(g34374) ) ;
AND2    gate18770  (.A(g34374), .B(g17471), .Z(g34565) ) ;
OR2     gate18771  (.A(g26301), .B(g34140), .Z(g34376) ) ;
AND2    gate18772  (.A(g34376), .B(g17489), .Z(g34566) ) ;
OR2     gate18773  (.A(g26304), .B(g34141), .Z(g34377) ) ;
AND2    gate18774  (.A(g34377), .B(g17491), .Z(g34567) ) ;
OR2     gate18775  (.A(g26312), .B(g34143), .Z(g34379) ) ;
AND2    gate18776  (.A(g34379), .B(g17512), .Z(g34568) ) ;
OR2     gate18777  (.A(g2975), .B(g26364), .Z(g27225) ) ;
AND2    gate18778  (.A(g34387), .B(g33326), .Z(g34572) ) ;
OR2     gate18779  (.A(g2856), .B(g22531), .Z(g24577) ) ;
OR2     gate18780  (.A(g2882), .B(g23825), .Z(g24578) ) ;
OR2     gate18781  (.A(g2864), .B(g28220), .Z(g29539) ) ;
NAND2   gate18782  (.A(g7780), .B(g21156), .Z(g22864) ) ;
OR2     gate18783  (.A(g2999), .B(g2932), .Z(g7764) ) ;
OR2     gate18784  (.A(g2848), .B(g22585), .Z(g24653) ) ;
OR2     gate18785  (.A(g2890), .B(g23267), .Z(g24705) ) ;
OR2     gate18786  (.A(g2980), .B(g7831), .Z(g11025) ) ;
OR2     gate18787  (.A(g2898), .B(g24561), .Z(g26082) ) ;
AND2    gate18788  (.A(g34573), .B(g18885), .Z(g34655) ) ;
AND2    gate18789  (.A(g34574), .B(g18896), .Z(g34658) ) ;
AND2    gate18790  (.A(g34575), .B(g18907), .Z(g34661) ) ;
AND2    gate18791  (.A(g34576), .B(g18931), .Z(g34662) ) ;
AND2    gate18792  (.A(g34583), .B(g19067), .Z(g34665) ) ;
AND2    gate18793  (.A(g34587), .B(g19144), .Z(g34666) ) ;
AND2    gate18794  (.A(g34471), .B(g33424), .Z(g34667) ) ;
AND2    gate18795  (.A(g34490), .B(g19431), .Z(g34678) ) ;
NOR2    gate18796  (.A(g8833), .B(g11083), .Z(g14093) ) ;
AND2    gate18797  (.A(g14093), .B(g34539), .Z(g34679) ) ;
AND2    gate18798  (.A(g34491), .B(g19438), .Z(g34681) ) ;
NOR2    gate18799  (.A(g8899), .B(g11083), .Z(g14178) ) ;
AND2    gate18800  (.A(g14178), .B(g34545), .Z(g34684) ) ;
NOR2    gate18801  (.A(g9000), .B(g12259), .Z(g14164) ) ;
AND2    gate18802  (.A(g14164), .B(g34550), .Z(g34685) ) ;
OR2     gate18803  (.A(g26849), .B(g34413), .Z(g34494) ) ;
AND2    gate18804  (.A(g34494), .B(g19494), .Z(g34686) ) ;
NOR2    gate18805  (.A(g9083), .B(g12259), .Z(g14181) ) ;
AND2    gate18806  (.A(g14181), .B(g34543), .Z(g34687) ) ;
AND2    gate18807  (.A(g34530), .B(g19885), .Z(g34694) ) ;
AND2    gate18808  (.A(g34531), .B(g20004), .Z(g34696) ) ;
OR2     gate18809  (.A(g34309), .B(g34073), .Z(g34535) ) ;
AND2    gate18810  (.A(g34535), .B(g20129), .Z(g34700) ) ;
AND2    gate18811  (.A(g34536), .B(g20179), .Z(g34701) ) ;
OR2     gate18812  (.A(g34324), .B(g34084), .Z(g34537) ) ;
AND2    gate18813  (.A(g34537), .B(g20208), .Z(g34702) ) ;
NOR2    gate18814  (.A(g34370), .B(g27648), .Z(g34496) ) ;
AND2    gate18815  (.A(g34496), .B(g10570), .Z(g34706) ) ;
AND2    gate18816  (.A(g34544), .B(g20579), .Z(g34707) ) ;
AND2    gate18817  (.A(g34549), .B(g17242), .Z(g34709) ) ;
AND2    gate18818  (.A(g34553), .B(g20903), .Z(g34710) ) ;
AND2    gate18819  (.A(g34570), .B(g33375), .Z(g34715) ) ;
AND2    gate18820  (.A(g34660), .B(g33442), .Z(g34738) ) ;
AND2    gate18821  (.A(g34664), .B(g19414), .Z(g34740) ) ;
AND2    gate18822  (.A(g8899), .B(g34697), .Z(g34741) ) ;
AND2    gate18823  (.A(g9000), .B(g34698), .Z(g34742) ) ;
AND2    gate18824  (.A(g8951), .B(g34703), .Z(g34743) ) ;
AND2    gate18825  (.A(g34668), .B(g19481), .Z(g34744) ) ;
AND2    gate18826  (.A(g34669), .B(g19482), .Z(g34745) ) ;
AND2    gate18827  (.A(g34670), .B(g19526), .Z(g34746) ) ;
AND2    gate18828  (.A(g34671), .B(g19527), .Z(g34747) ) ;
AND2    gate18829  (.A(g34672), .B(g19529), .Z(g34748) ) ;
AND2    gate18830  (.A(g34673), .B(g19542), .Z(g34750) ) ;
AND2    gate18831  (.A(g34674), .B(g19543), .Z(g34751) ) ;
AND2    gate18832  (.A(g34675), .B(g19544), .Z(g34752) ) ;
AND2    gate18833  (.A(g34676), .B(g19586), .Z(g34753) ) ;
AND2    gate18834  (.A(g34677), .B(g19602), .Z(g34754) ) ;
AND2    gate18835  (.A(g34680), .B(g19618), .Z(g34756) ) ;
AND2    gate18836  (.A(g34682), .B(g19635), .Z(g34757) ) ;
AND2    gate18837  (.A(g34683), .B(g19657), .Z(g34758) ) ;
AND2    gate18838  (.A(g34689), .B(g19915), .Z(g34763) ) ;
AND2    gate18839  (.A(g34691), .B(g20009), .Z(g34764) ) ;
AND2    gate18840  (.A(g34692), .B(g20057), .Z(g34765) ) ;
OR2     gate18841  (.A(g34513), .B(g34310), .Z(g34693) ) ;
AND2    gate18842  (.A(g34693), .B(g20147), .Z(g34771) ) ;
OR2     gate18843  (.A(g34523), .B(g34322), .Z(g34695) ) ;
AND2    gate18844  (.A(g34695), .B(g20180), .Z(g34774) ) ;
AND2    gate18845  (.A(g34711), .B(g33888), .Z(g34782) ) ;
NOR2    gate18846  (.A(g8951), .B(g11083), .Z(g14165) ) ;
AND2    gate18847  (.A(g14165), .B(g34766), .Z(g34811) ) ;
OR2     gate18848  (.A(g34679), .B(g34506), .Z(g34761) ) ;
AND2    gate18849  (.A(g34761), .B(g20080), .Z(g34841) ) ;
OR2     gate18850  (.A(g34687), .B(g34524), .Z(g34762) ) ;
AND2    gate18851  (.A(g34762), .B(g20168), .Z(g34842) ) ;
AND2    gate18852  (.A(g16540), .B(g34813), .Z(g34857) ) ;
AND2    gate18853  (.A(g16540), .B(g34816), .Z(g34858) ) ;
AND2    gate18854  (.A(g16540), .B(g34820), .Z(g34859) ) ;
AND2    gate18855  (.A(g16540), .B(g34823), .Z(g34860) ) ;
AND2    gate18856  (.A(g16540), .B(g34827), .Z(g34861) ) ;
AND2    gate18857  (.A(g16540), .B(g34830), .Z(g34862) ) ;
AND2    gate18858  (.A(g16540), .B(g34833), .Z(g34863) ) ;
AND2    gate18859  (.A(g16540), .B(g34836), .Z(g34865) ) ;
OR2     gate18860  (.A(g34741), .B(g34684), .Z(g34819) ) ;
AND2    gate18861  (.A(g34819), .B(g20106), .Z(g34866) ) ;
OR2     gate18862  (.A(g34742), .B(g34685), .Z(g34826) ) ;
AND2    gate18863  (.A(g34826), .B(g20145), .Z(g34867) ) ;
AND2    gate18864  (.A(g34813), .B(g19866), .Z(g34868) ) ;
AND2    gate18865  (.A(g34816), .B(g19869), .Z(g34869) ) ;
AND2    gate18866  (.A(g34820), .B(g19882), .Z(g34870) ) ;
AND2    gate18867  (.A(g34823), .B(g19908), .Z(g34871) ) ;
AND2    gate18868  (.A(g34827), .B(g19954), .Z(g34872) ) ;
AND2    gate18869  (.A(g34830), .B(g20046), .Z(g34873) ) ;
AND2    gate18870  (.A(g34833), .B(g20060), .Z(g34874) ) ;
AND2    gate18871  (.A(g34836), .B(g20073), .Z(g34875) ) ;
AND2    gate18872  (.A(g34844), .B(g20534), .Z(g34876) ) ;
OR2     gate18873  (.A(g34811), .B(g34743), .Z(g34856) ) ;
AND2    gate18874  (.A(g34856), .B(g20130), .Z(g34909) ) ;
AND2    gate18875  (.A(g16540), .B(g34935), .Z(g34948) ) ;
AND2    gate18876  (.A(g34935), .B(g19957), .Z(g34953) ) ;
OR2     gate18877  (.A(g2984), .B(g34912), .Z(g34931) ) ;
AND2    gate18878  (.A(g34944), .B(g23019), .Z(g34961) ) ;
AND2    gate18879  (.A(g34945), .B(g23020), .Z(g34962) ) ;
AND2    gate18880  (.A(g34946), .B(g23041), .Z(g34963) ) ;
AND2    gate18881  (.A(g34947), .B(g23060), .Z(g34964) ) ;
AND2    gate18882  (.A(g34949), .B(g23084), .Z(g34965) ) ;
AND2    gate18883  (.A(g34950), .B(g23170), .Z(g34966) ) ;
AND2    gate18884  (.A(g34951), .B(g23189), .Z(g34967) ) ;
AND2    gate18885  (.A(g34952), .B(g23203), .Z(g34968) ) ;
AND2    gate18886  (.A(g34960), .B(g19570), .Z(g34969) ) ;
AND2    gate18887  (.A(g34998), .B(g23085), .Z(g34999) ) ;
OR3     gate18888  (.A(g1157), .B(g1239), .C(g990), .Z(II12583) ) ;
OR3     gate18889  (.A(g1500), .B(g1582), .C(g1333), .Z(II12611) ) ;
OR4     gate18890  (.A(g4188), .B(g4194), .C(g4197), .D(g4200), .Z(II12782) ) ;
OR4     gate18891  (.A(g4204), .B(g4207), .C(g4210), .D(g4180), .Z(II12783) ) ;
OR2     gate18892  (.A(II12782), .B(II12783), .Z(g8790) ) ;
OR2     gate18893  (.A(g1644), .B(g1664), .Z(g8863) ) ;
OR2     gate18894  (.A(g1779), .B(g1798), .Z(g8904) ) ;
OR2     gate18895  (.A(g2204), .B(g2223), .Z(g8905) ) ;
OR4     gate18896  (.A(g4235), .B(g4232), .C(g4229), .D(g4226), .Z(II12902) ) ;
OR4     gate18897  (.A(g4222), .B(g4219), .C(g4216), .D(g4213), .Z(II12903) ) ;
OR2     gate18898  (.A(II12902), .B(II12903), .Z(g8921) ) ;
OR2     gate18899  (.A(g1913), .B(g1932), .Z(g8956) ) ;
OR2     gate18900  (.A(g2338), .B(g2357), .Z(g8957) ) ;
OR2     gate18901  (.A(g2047), .B(g2066), .Z(g9012) ) ;
OR2     gate18902  (.A(g2472), .B(g2491), .Z(g9013) ) ;
OR2     gate18903  (.A(g2606), .B(g2625), .Z(g9055) ) ;
OR2     gate18904  (.A(g1008), .B(g969), .Z(g9483) ) ;
OR2     gate18905  (.A(g1351), .B(g1312), .Z(g9536) ) ;
NAND2   gate18906  (.A(II11878), .B(II11879), .Z(g7223) ) ;
NAND2   gate18907  (.A(II11865), .B(II11866), .Z(g7201) ) ;
OR3     gate18908  (.A(g490), .B(g482), .C(g8038), .Z(g11372) ) ;
OR2     gate18909  (.A(g8583), .B(g8530), .Z(g11380) ) ;
NAND3   gate18910  (.A(g4628), .B(g7202), .C(g4621), .Z(g10511) ) ;
OR3     gate18911  (.A(g329), .B(g319), .C(g10796), .Z(g13091) ) ;
OR2     gate18912  (.A(g7396), .B(g10684), .Z(g13794) ) ;
NOR2    gate18913  (.A(g513), .B(g9040), .Z(g11184) ) ;
OR2     gate18914  (.A(g209), .B(g10685), .Z(g13858) ) ;
OR2     gate18915  (.A(g8643), .B(g11380), .Z(g13914) ) ;
NOR3    gate18916  (.A(g4776), .B(g7892), .C(g9030), .Z(g11213) ) ;
NOR3    gate18917  (.A(g4776), .B(g4801), .C(g9030), .Z(g11191) ) ;
OR2     gate18918  (.A(g11213), .B(g11191), .Z(g13938) ) ;
NOR2    gate18919  (.A(g4191), .B(g8790), .Z(g11448) ) ;
NAND2   gate18920  (.A(II12877), .B(II12878), .Z(g8913) ) ;
NOR3    gate18921  (.A(g4966), .B(g7898), .C(g9064), .Z(g11232) ) ;
NOR3    gate18922  (.A(g4966), .B(g4991), .C(g9064), .Z(g11203) ) ;
OR2     gate18923  (.A(g11232), .B(g11203), .Z(g13972) ) ;
NAND2   gate18924  (.A(II12841), .B(II12842), .Z(g8871) ) ;
NOR2    gate18925  (.A(g8921), .B(g4185), .Z(g11771) ) ;
OR2     gate18926  (.A(g8871), .B(g11771), .Z(g14187) ) ;
NOR2    gate18927  (.A(g7479), .B(g1041), .Z(g10819) ) ;
NOR2    gate18928  (.A(g7503), .B(g1384), .Z(g10821) ) ;
OR2     gate18929  (.A(g8690), .B(g13914), .Z(g16811) ) ;
OR3     gate18930  (.A(g14028), .B(g11773), .C(g11755), .Z(g16876) ) ;
OR3     gate18931  (.A(g14061), .B(g11804), .C(g11780), .Z(g16926) ) ;
NOR2    gate18932  (.A(g11914), .B(g9638), .Z(g14413) ) ;
NOR2    gate18933  (.A(g12112), .B(g9585), .Z(g14391) ) ;
NOR2    gate18934  (.A(g12078), .B(g9484), .Z(g14360) ) ;
OR3     gate18935  (.A(g14413), .B(g14391), .C(g14360), .Z(II18385) ) ;
NOR2    gate18936  (.A(g12044), .B(g9337), .Z(g14334) ) ;
NOR2    gate18937  (.A(g12016), .B(g9250), .Z(g14313) ) ;
NOR2    gate18938  (.A(g9485), .B(g7267), .Z(g11935) ) ;
NOR2    gate18939  (.A(g11936), .B(g9692), .Z(g14444) ) ;
NOR2    gate18940  (.A(g12145), .B(g9639), .Z(g14414) ) ;
NOR2    gate18941  (.A(g12114), .B(g9537), .Z(g14392) ) ;
OR3     gate18942  (.A(g14444), .B(g14414), .C(g14392), .Z(II18417) ) ;
NOR2    gate18943  (.A(g12079), .B(g9413), .Z(g14361) ) ;
NOR2    gate18944  (.A(g12045), .B(g9283), .Z(g14335) ) ;
NOR2    gate18945  (.A(g9538), .B(g7314), .Z(g11954) ) ;
NOR2    gate18946  (.A(g11938), .B(g9698), .Z(g14447) ) ;
NOR2    gate18947  (.A(g12149), .B(g9648), .Z(g14417) ) ;
NOR2    gate18948  (.A(g12118), .B(g9542), .Z(g14395) ) ;
OR3     gate18949  (.A(g14447), .B(g14417), .C(g14395), .Z(II18421) ) ;
NOR2    gate18950  (.A(g12083), .B(g9415), .Z(g14364) ) ;
NOR2    gate18951  (.A(g12049), .B(g9284), .Z(g14337) ) ;
NOR2    gate18952  (.A(g9543), .B(g7327), .Z(g11958) ) ;
NOR2    gate18953  (.A(g11955), .B(g9753), .Z(g14512) ) ;
NOR2    gate18954  (.A(g12188), .B(g9693), .Z(g14445) ) ;
NOR2    gate18955  (.A(g12147), .B(g9590), .Z(g14415) ) ;
OR3     gate18956  (.A(g14512), .B(g14445), .C(g14415), .Z(II18449) ) ;
NOR2    gate18957  (.A(g12115), .B(g9488), .Z(g14393) ) ;
NOR2    gate18958  (.A(g12080), .B(g9338), .Z(g14362) ) ;
NOR2    gate18959  (.A(g9591), .B(g7361), .Z(g11972) ) ;
NOR2    gate18960  (.A(g11959), .B(g9760), .Z(g14514) ) ;
NOR2    gate18961  (.A(g12192), .B(g9699), .Z(g14448) ) ;
NOR2    gate18962  (.A(g12151), .B(g9594), .Z(g14418) ) ;
OR3     gate18963  (.A(g14514), .B(g14448), .C(g14418), .Z(II18452) ) ;
NOR2    gate18964  (.A(g12119), .B(g9489), .Z(g14396) ) ;
NOR2    gate18965  (.A(g12084), .B(g9339), .Z(g14365) ) ;
NOR2    gate18966  (.A(g9595), .B(g7379), .Z(g11976) ) ;
NOR2    gate18967  (.A(g11973), .B(g9828), .Z(g14538) ) ;
NOR2    gate18968  (.A(g12222), .B(g9754), .Z(g14513) ) ;
NOR2    gate18969  (.A(g12190), .B(g9644), .Z(g14446) ) ;
OR3     gate18970  (.A(g14538), .B(g14513), .C(g14446), .Z(II18492) ) ;
NOR2    gate18971  (.A(g12148), .B(g9541), .Z(g14416) ) ;
NOR2    gate18972  (.A(g12116), .B(g9414), .Z(g14394) ) ;
NOR2    gate18973  (.A(g9645), .B(g7410), .Z(g11995) ) ;
NOR2    gate18974  (.A(g11977), .B(g9833), .Z(g14539) ) ;
NOR2    gate18975  (.A(g12225), .B(g9761), .Z(g14515) ) ;
NOR2    gate18976  (.A(g12194), .B(g9653), .Z(g14449) ) ;
OR3     gate18977  (.A(g14539), .B(g14515), .C(g14449), .Z(II18495) ) ;
NOR2    gate18978  (.A(g12152), .B(g9546), .Z(g14419) ) ;
NOR2    gate18979  (.A(g12120), .B(g9416), .Z(g14397) ) ;
NOR2    gate18980  (.A(g9654), .B(g7423), .Z(g11999) ) ;
NOR2    gate18981  (.A(g12000), .B(g9915), .Z(g14568) ) ;
NOR2    gate18982  (.A(g12287), .B(g9834), .Z(g14540) ) ;
NOR2    gate18983  (.A(g12227), .B(g9704), .Z(g14516) ) ;
OR3     gate18984  (.A(g14568), .B(g14540), .C(g14516), .Z(II18543) ) ;
NOR2    gate18985  (.A(g12195), .B(g9598), .Z(g14450) ) ;
NOR2    gate18986  (.A(g12153), .B(g9490), .Z(g14420) ) ;
NOR2    gate18987  (.A(g9705), .B(g7461), .Z(g12025) ) ;
OR2     gate18988  (.A(g7696), .B(g16811), .Z(g19525) ) ;
OR2     gate18989  (.A(g691), .B(g16893), .Z(g20522) ) ;
OR2     gate18990  (.A(g20773), .B(g20922), .Z(g22531) ) ;
OR2     gate18991  (.A(g20915), .B(g21061), .Z(g22585) ) ;
OR2     gate18992  (.A(g7763), .B(g19525), .Z(g22669) ) ;
NAND4   gate18993  (.A(g16875), .B(g14014), .C(g16625), .D(g16604), .Z(g20236) ) ;
NAND4   gate18994  (.A(g17668), .B(g17634), .C(g17597), .D(g14569), .Z(g20133) ) ;
NAND4   gate18995  (.A(g17513), .B(g14517), .C(g17468), .D(g14422), .Z(g20111) ) ;
OR3     gate18996  (.A(g20236), .B(g20133), .C(g20111), .Z(II22267) ) ;
NAND4   gate18997  (.A(g16770), .B(g13918), .C(g16719), .D(g13896), .Z(g20184) ) ;
NAND4   gate18998  (.A(g16741), .B(g13897), .C(g16687), .D(g13866), .Z(g20170) ) ;
NAND4   gate18999  (.A(g16925), .B(g14054), .C(g16657), .D(g16628), .Z(g20271) ) ;
NAND4   gate19000  (.A(g17705), .B(g17669), .C(g17635), .D(g14590), .Z(g20150) ) ;
NAND4   gate19001  (.A(g17572), .B(g14542), .C(g17495), .D(g14452), .Z(g20134) ) ;
OR3     gate19002  (.A(g20271), .B(g20150), .C(g20134), .Z(II22280) ) ;
NAND4   gate19003  (.A(g16813), .B(g13958), .C(g16745), .D(g13927), .Z(g20198) ) ;
NAND4   gate19004  (.A(g16772), .B(g13928), .C(g16723), .D(g13882), .Z(g20185) ) ;
NAND4   gate19005  (.A(g16956), .B(g14088), .C(g16694), .D(g16660), .Z(g20371) ) ;
NAND4   gate19006  (.A(g17732), .B(g17706), .C(g17670), .D(g14625), .Z(g20161) ) ;
NAND4   gate19007  (.A(g17598), .B(g14570), .C(g17514), .D(g14519), .Z(g20151) ) ;
OR3     gate19008  (.A(g20371), .B(g20161), .C(g20151), .Z(II22298) ) ;
NAND4   gate19009  (.A(g16854), .B(g13993), .C(g16776), .D(g13967), .Z(g20214) ) ;
NAND4   gate19010  (.A(g16815), .B(g13968), .C(g16749), .D(g13907), .Z(g20199) ) ;
NAND4   gate19011  (.A(g17788), .B(g14803), .C(g17578), .D(g17520), .Z(g21429) ) ;
NAND4   gate19012  (.A(g15741), .B(g15734), .C(g15728), .D(g13097), .Z(g21338) ) ;
NAND4   gate19013  (.A(g15719), .B(g13067), .C(g15709), .D(g13040), .Z(g21307) ) ;
OR3     gate19014  (.A(g21429), .B(g21338), .C(g21307), .Z(II22830) ) ;
NAND4   gate19015  (.A(g17734), .B(g14686), .C(g17675), .D(g14663), .Z(g21384) ) ;
NAND4   gate19016  (.A(g17708), .B(g14664), .C(g17640), .D(g14598), .Z(g21363) ) ;
NAND4   gate19017  (.A(g17814), .B(g14854), .C(g17605), .D(g17581), .Z(g21459) ) ;
NAND4   gate19018  (.A(g15751), .B(g15742), .C(g15735), .D(g13108), .Z(g21350) ) ;
NAND4   gate19019  (.A(g15725), .B(g13084), .C(g15713), .D(g13050), .Z(g21339) ) ;
OR3     gate19020  (.A(g21459), .B(g21350), .C(g21339), .Z(II22852) ) ;
NAND4   gate19021  (.A(g17755), .B(g14730), .C(g17712), .D(g14695), .Z(g21401) ) ;
NAND4   gate19022  (.A(g17736), .B(g14696), .C(g17679), .D(g14636), .Z(g21385) ) ;
NAND4   gate19023  (.A(g17820), .B(g14898), .C(g17647), .D(g17608), .Z(g21509) ) ;
NAND4   gate19024  (.A(g15780), .B(g15752), .C(g15743), .D(g13118), .Z(g21356) ) ;
NAND4   gate19025  (.A(g15729), .B(g13098), .C(g15720), .D(g13069), .Z(g21351) ) ;
OR3     gate19026  (.A(g21509), .B(g21356), .C(g21351), .Z(II22880) ) ;
NAND4   gate19027  (.A(g17773), .B(g14771), .C(g17740), .D(g14739), .Z(g21415) ) ;
NAND4   gate19028  (.A(g17757), .B(g14740), .C(g17716), .D(g14674), .Z(g21402) ) ;
NAND4   gate19029  (.A(g17846), .B(g14946), .C(g17686), .D(g17650), .Z(g21555) ) ;
NAND4   gate19030  (.A(g15787), .B(g15781), .C(g15753), .D(g13131), .Z(g21364) ) ;
NAND4   gate19031  (.A(g15736), .B(g13109), .C(g15726), .D(g13086), .Z(g21357) ) ;
OR3     gate19032  (.A(g21555), .B(g21364), .C(g21357), .Z(II22912) ) ;
NAND4   gate19033  (.A(g17790), .B(g14820), .C(g17761), .D(g14780), .Z(g21432) ) ;
NAND4   gate19034  (.A(g17775), .B(g14781), .C(g17744), .D(g14706), .Z(g21416) ) ;
NAND4   gate19035  (.A(g17872), .B(g14987), .C(g17723), .D(g17689), .Z(g21603) ) ;
NAND4   gate19036  (.A(g15798), .B(g15788), .C(g15782), .D(g13139), .Z(g21386) ) ;
NAND4   gate19037  (.A(g15744), .B(g13119), .C(g15730), .D(g13100), .Z(g21365) ) ;
OR3     gate19038  (.A(g21603), .B(g21386), .C(g21365), .Z(II22958) ) ;
NAND4   gate19039  (.A(g17816), .B(g14871), .C(g17779), .D(g14829), .Z(g21462) ) ;
NAND4   gate19040  (.A(g17792), .B(g14830), .C(g17765), .D(g14750), .Z(g21433) ) ;
OR2     gate19041  (.A(g20705), .B(g20781), .Z(g23825) ) ;
OR4     gate19042  (.A(g19919), .B(g19968), .C(g20014), .D(g20841), .Z(II23162) ) ;
OR4     gate19043  (.A(g20982), .B(g21127), .C(g21193), .D(g21256), .Z(II23163) ) ;
OR2     gate19044  (.A(g7831), .B(g22138), .Z(g24363) ) ;
NOR2    gate19045  (.A(g19345), .B(g15718), .Z(g22400) ) ;
OR2     gate19046  (.A(g10878), .B(g22400), .Z(g24433) ) ;
OR2     gate19047  (.A(g10890), .B(g22400), .Z(g24444) ) ;
NOR2    gate19048  (.A(g19345), .B(g15724), .Z(g22450) ) ;
OR2     gate19049  (.A(g10948), .B(g22450), .Z(g24447) ) ;
OR2     gate19050  (.A(g10902), .B(g22400), .Z(g24457) ) ;
OR2     gate19051  (.A(g10967), .B(g22450), .Z(g24460) ) ;
OR2     gate19052  (.A(g10925), .B(g22400), .Z(g24468) ) ;
OR2     gate19053  (.A(g10999), .B(g22450), .Z(g24471) ) ;
OR2     gate19054  (.A(g11003), .B(g22450), .Z(g24478) ) ;
NOR2    gate19055  (.A(g19699), .B(g1002), .Z(g22488) ) ;
NOR2    gate19056  (.A(g19720), .B(g1345), .Z(g22517) ) ;
OR4     gate19057  (.A(g22904), .B(g22927), .C(g22980), .D(g23444), .Z(II23755) ) ;
OR4     gate19058  (.A(g23457), .B(g23480), .C(g23494), .D(g23511), .Z(II23756) ) ;
OR2     gate19059  (.A(II23755), .B(II23756), .Z(g24561) ) ;
OR3     gate19060  (.A(g23088), .B(g23154), .C(g23172), .Z(II24117) ) ;
OR2     gate19061  (.A(g22667), .B(g23825), .Z(g24965) ) ;
OR2     gate19062  (.A(g23267), .B(g2932), .Z(g25010) ) ;
OR2     gate19063  (.A(g24139), .B(g24140), .Z(g25575) ) ;
OR2     gate19064  (.A(g24141), .B(g24142), .Z(g25576) ) ;
OR2     gate19065  (.A(g24143), .B(g24144), .Z(g25577) ) ;
OR4     gate19066  (.A(g25411), .B(g25371), .C(g25328), .D(g25290), .Z(g25791) ) ;
OR4     gate19067  (.A(g25453), .B(g25414), .C(g25374), .D(g25331), .Z(g25805) ) ;
OR4     gate19068  (.A(g25482), .B(g25456), .C(g25417), .D(g25377), .Z(g25821) ) ;
OR4     gate19069  (.A(g25507), .B(g25485), .C(g25459), .D(g25420), .Z(g25839) ) ;
OR4     gate19070  (.A(g25518), .B(g25510), .C(g25488), .D(g25462), .Z(g25856) ) ;
NOR2    gate19071  (.A(g19699), .B(g1018), .Z(g22514) ) ;
NOR2    gate19072  (.A(g19720), .B(g1361), .Z(g22524) ) ;
NAND2   gate19073  (.A(g22755), .B(g22713), .Z(g24566) ) ;
NAND2   gate19074  (.A(g22994), .B(g23010), .Z(g24678) ) ;
NAND2   gate19075  (.A(g22833), .B(g22642), .Z(g24591) ) ;
NAND2   gate19076  (.A(g22850), .B(g22650), .Z(g24609) ) ;
NOR2    gate19077  (.A(g22550), .B(g7222), .Z(g25504) ) ;
NOR2    gate19078  (.A(g22228), .B(g10334), .Z(g25141) ) ;
OR4     gate19079  (.A(g24881), .B(g24855), .C(g24843), .D(g24822), .Z(g26616) ) ;
OR4     gate19080  (.A(g24897), .B(g24884), .C(g24858), .D(g24846), .Z(g26636) ) ;
OR4     gate19081  (.A(g24908), .B(g24900), .C(g24887), .D(g24861), .Z(g26657) ) ;
OR3     gate19082  (.A(g20204), .B(g20242), .C(g24363), .Z(g26866) ) ;
OR4     gate19083  (.A(g25567), .B(g25568), .C(g25569), .D(g25570), .Z(II25612) ) ;
OR4     gate19084  (.A(g25571), .B(g25572), .C(g25573), .D(g25574), .Z(II25613) ) ;
OR2     gate19085  (.A(II25612), .B(II25613), .Z(g26874) ) ;
NOR2    gate19086  (.A(g17619), .B(g17663), .Z(g21652) ) ;
NOR2    gate19087  (.A(g17657), .B(g17700), .Z(g21655) ) ;
NOR2    gate19088  (.A(g17694), .B(g17727), .Z(g21658) ) ;
OR2     gate19089  (.A(g25578), .B(g25579), .Z(g26878) ) ;
OR2     gate19090  (.A(g25580), .B(g25581), .Z(g26879) ) ;
OR3     gate19091  (.A(g12), .B(g22150), .C(g20277), .Z(II25736) ) ;
NOR2    gate19092  (.A(g19699), .B(g1024), .Z(g22522) ) ;
NOR2    gate19093  (.A(g19720), .B(g1367), .Z(g22537) ) ;
NAND2   gate19094  (.A(g22902), .B(g22874), .Z(g24620) ) ;
NAND2   gate19095  (.A(g24576), .B(g22837), .Z(g25974) ) ;
NAND3   gate19096  (.A(g22852), .B(g22836), .C(g22715), .Z(g24584) ) ;
NAND2   gate19097  (.A(g24567), .B(g22668), .Z(g25984) ) ;
NAND3   gate19098  (.A(g22712), .B(g22940), .C(g22757), .Z(g24652) ) ;
NAND2   gate19099  (.A(g24621), .B(g22853), .Z(g25995) ) ;
NAND3   gate19100  (.A(g23281), .B(g23266), .C(g22839), .Z(g24880) ) ;
NAND3   gate19101  (.A(g22756), .B(g24570), .C(g22688), .Z(g25953) ) ;
NAND3   gate19102  (.A(g23210), .B(g23195), .C(g22984), .Z(g24661) ) ;
NAND3   gate19103  (.A(g22714), .B(g24662), .C(g22921), .Z(g26052) ) ;
NAND3   gate19104  (.A(g22666), .B(g22661), .C(g22651), .Z(g24544) ) ;
NAND2   gate19105  (.A(g24601), .B(g22838), .Z(g25996) ) ;
NAND3   gate19106  (.A(g22638), .B(g22643), .C(g22754), .Z(g24547) ) ;
NAND3   gate19107  (.A(g22875), .B(g24677), .C(g22941), .Z(g26053) ) ;
NOR2    gate19108  (.A(II23162), .B(II23163), .Z(g24018) ) ;
OR4     gate19109  (.A(g19890), .B(g19935), .C(g19984), .D(g26365), .Z(II26522) ) ;
OR4     gate19110  (.A(g20720), .B(g20857), .C(g20998), .D(g21143), .Z(II26523) ) ;
NOR2    gate19111  (.A(g19402), .B(g19422), .Z(g24145) ) ;
NOR2    gate19112  (.A(g19268), .B(g19338), .Z(g24148) ) ;
OR4     gate19113  (.A(g27073), .B(g27058), .C(g27045), .D(g27040), .Z(II26643) ) ;
OR4     gate19114  (.A(g27057), .B(g27044), .C(g27039), .D(g27032), .Z(II26644) ) ;
OR4     gate19115  (.A(g27209), .B(g27185), .C(g27161), .D(g27146), .Z(g28186) ) ;
NOR2    gate19116  (.A(g19699), .B(g1030), .Z(g22535) ) ;
OR4     gate19117  (.A(g27217), .B(g27210), .C(g27186), .D(g27162), .Z(g28191) ) ;
NOR2    gate19118  (.A(g19720), .B(g1373), .Z(g22540) ) ;
NAND2   gate19119  (.A(II25908), .B(II25909), .Z(g27223) ) ;
NAND2   gate19120  (.A(II25846), .B(II25847), .Z(g27141) ) ;
OR4     gate19121  (.A(g22881), .B(g22905), .C(g22928), .D(g27402), .Z(II26741) ) ;
OR4     gate19122  (.A(g23430), .B(g23445), .C(g23458), .D(g23481), .Z(II26742) ) ;
OR3     gate19123  (.A(g23495), .B(II26741), .C(II26742), .Z(g28220) ) ;
OR2     gate19124  (.A(g28524), .B(g27588), .Z(g29482) ) ;
OR2     gate19125  (.A(g28535), .B(g27594), .Z(g29485) ) ;
OR2     gate19126  (.A(g28537), .B(g27595), .Z(g29486) ) ;
OR2     gate19127  (.A(g28547), .B(g27600), .Z(g29488) ) ;
OR2     gate19128  (.A(g28550), .B(g27601), .Z(g29489) ) ;
OR2     gate19129  (.A(g28563), .B(g27614), .Z(g29495) ) ;
OR2     gate19130  (.A(g28567), .B(g27615), .Z(g29496) ) ;
OR2     gate19131  (.A(g28583), .B(g27634), .Z(g29501) ) ;
OR4     gate19132  (.A(g28291), .B(g28281), .C(g28264), .D(g28254), .Z(g29520) ) ;
OR4     gate19133  (.A(g28303), .B(g28293), .C(g28283), .D(g28267), .Z(g29529) ) ;
OR3     gate19134  (.A(g2946), .B(g24561), .C(g28220), .Z(II28147) ) ;
OR3     gate19135  (.A(g22531), .B(g22585), .C(II28147), .Z(g29914) ) ;
OR4     gate19136  (.A(g29201), .B(g29202), .C(g29203), .D(g28035), .Z(II28566) ) ;
OR4     gate19137  (.A(g29204), .B(g29205), .C(g29206), .D(g29207), .Z(II28567) ) ;
OR3     gate19138  (.A(g29208), .B(II28566), .C(II28567), .Z(g30317) ) ;
OR4     gate19139  (.A(g29328), .B(g29323), .C(g29316), .D(g30316), .Z(II29351) ) ;
OR4     gate19140  (.A(g29322), .B(g29315), .C(g30315), .D(g30308), .Z(II29352) ) ;
NOR3    gate19141  (.A(g21209), .B(II26522), .C(II26523), .Z(g28031) ) ;
NOR2    gate19142  (.A(g4507), .B(g29365), .Z(g30613) ) ;
OR3     gate19143  (.A(g26105), .B(g26131), .C(g30613), .Z(g32426) ) ;
OR4     gate19144  (.A(g29385), .B(g31376), .C(g30735), .D(g30825), .Z(II29985) ) ;
OR4     gate19145  (.A(g31070), .B(g31194), .C(g30614), .D(g30673), .Z(II29986) ) ;
OR4     gate19146  (.A(g29385), .B(g31376), .C(g30735), .D(g30825), .Z(II30054) ) ;
OR4     gate19147  (.A(g31070), .B(g31170), .C(g30614), .D(g30673), .Z(II30055) ) ;
OR4     gate19148  (.A(g29385), .B(g31376), .C(g30735), .D(g30825), .Z(II30123) ) ;
OR4     gate19149  (.A(g31070), .B(g31154), .C(g30614), .D(g30673), .Z(II30124) ) ;
OR4     gate19150  (.A(g29385), .B(g31376), .C(g30735), .D(g30825), .Z(II30192) ) ;
OR4     gate19151  (.A(g31070), .B(g30614), .C(g30673), .D(g31528), .Z(II30193) ) ;
OR4     gate19152  (.A(g29385), .B(g31376), .C(g30735), .D(g30825), .Z(II30261) ) ;
OR4     gate19153  (.A(g31672), .B(g31710), .C(g31021), .D(g30937), .Z(II30262) ) ;
OR4     gate19154  (.A(g29385), .B(g31376), .C(g30735), .D(g30825), .Z(II30330) ) ;
OR4     gate19155  (.A(g31672), .B(g31710), .C(g31021), .D(g30937), .Z(II30331) ) ;
OR4     gate19156  (.A(g29385), .B(g31376), .C(g30735), .D(g30825), .Z(II30399) ) ;
OR4     gate19157  (.A(g31021), .B(g30937), .C(g31327), .D(g30614), .Z(II30400) ) ;
OR4     gate19158  (.A(g29385), .B(g31376), .C(g30735), .D(g30825), .Z(II30468) ) ;
OR4     gate19159  (.A(g31672), .B(g31710), .C(g31021), .D(g30937), .Z(II30469) ) ;
OR4     gate19160  (.A(g31787), .B(g32200), .C(g31940), .D(g31949), .Z(II30717) ) ;
OR4     gate19161  (.A(g32348), .B(g32356), .C(g32097), .D(g32020), .Z(II30718) ) ;
OR4     gate19162  (.A(g31759), .B(g32196), .C(g31933), .D(g31941), .Z(II30727) ) ;
OR4     gate19163  (.A(g32345), .B(g32350), .C(g32056), .D(g32018), .Z(II30728) ) ;
OR4     gate19164  (.A(g31790), .B(g32191), .C(g32086), .D(g32095), .Z(II30734) ) ;
OR4     gate19165  (.A(g32369), .B(g32376), .C(g32089), .D(g32035), .Z(II30735) ) ;
OR4     gate19166  (.A(g31776), .B(g32188), .C(g32083), .D(g32087), .Z(II30740) ) ;
OR4     gate19167  (.A(g32085), .B(g32030), .C(g32224), .D(g32013), .Z(II30741) ) ;
OR4     gate19168  (.A(g31777), .B(g32321), .C(g32069), .D(g32084), .Z(II30745) ) ;
OR4     gate19169  (.A(g32047), .B(g31985), .C(g31991), .D(g32309), .Z(II30746) ) ;
OR4     gate19170  (.A(g31788), .B(g32310), .C(g32054), .D(g32070), .Z(II30750) ) ;
OR4     gate19171  (.A(g32042), .B(g32161), .C(g31943), .D(g31959), .Z(II30751) ) ;
OR4     gate19172  (.A(g30564), .B(g32303), .C(g32049), .D(g32055), .Z(II30755) ) ;
OR4     gate19173  (.A(g32088), .B(g32163), .C(g32098), .D(g32105), .Z(II30756) ) ;
OR4     gate19174  (.A(g31778), .B(g32295), .C(g32046), .D(g32050), .Z(II30760) ) ;
OR4     gate19175  (.A(g32071), .B(g32167), .C(g32067), .D(g32082), .Z(II30761) ) ;
OR4     gate19176  (.A(g33461), .B(g33462), .C(g33463), .D(g33464), .Z(II31838) ) ;
OR4     gate19177  (.A(g33465), .B(g33466), .C(g33467), .D(g33468), .Z(II31839) ) ;
OR3     gate19178  (.A(g33469), .B(II31838), .C(II31839), .Z(g33951) ) ;
OR4     gate19179  (.A(g33470), .B(g33471), .C(g33472), .D(g33473), .Z(II31843) ) ;
OR4     gate19180  (.A(g33474), .B(g33475), .C(g33476), .D(g33477), .Z(II31844) ) ;
OR3     gate19181  (.A(g33478), .B(II31843), .C(II31844), .Z(g33952) ) ;
OR4     gate19182  (.A(g33479), .B(g33480), .C(g33481), .D(g33482), .Z(II31848) ) ;
OR4     gate19183  (.A(g33483), .B(g33484), .C(g33485), .D(g33486), .Z(II31849) ) ;
OR3     gate19184  (.A(g33487), .B(II31848), .C(II31849), .Z(g33953) ) ;
OR4     gate19185  (.A(g33488), .B(g33489), .C(g33490), .D(g33491), .Z(II31853) ) ;
OR4     gate19186  (.A(g33492), .B(g33493), .C(g33494), .D(g33495), .Z(II31854) ) ;
OR3     gate19187  (.A(g33496), .B(II31853), .C(II31854), .Z(g33954) ) ;
OR4     gate19188  (.A(g33497), .B(g33498), .C(g33499), .D(g33500), .Z(II31858) ) ;
OR4     gate19189  (.A(g33501), .B(g33502), .C(g33503), .D(g33504), .Z(II31859) ) ;
OR3     gate19190  (.A(g33505), .B(II31858), .C(II31859), .Z(g33955) ) ;
OR4     gate19191  (.A(g33506), .B(g33507), .C(g33508), .D(g33509), .Z(II31863) ) ;
OR4     gate19192  (.A(g33510), .B(g33511), .C(g33512), .D(g33513), .Z(II31864) ) ;
OR3     gate19193  (.A(g33514), .B(II31863), .C(II31864), .Z(g33956) ) ;
OR4     gate19194  (.A(g33515), .B(g33516), .C(g33517), .D(g33518), .Z(II31868) ) ;
OR4     gate19195  (.A(g33519), .B(g33520), .C(g33521), .D(g33522), .Z(II31869) ) ;
OR3     gate19196  (.A(g33523), .B(II31868), .C(II31869), .Z(g33957) ) ;
OR4     gate19197  (.A(g33524), .B(g33525), .C(g33526), .D(g33527), .Z(II31873) ) ;
OR4     gate19198  (.A(g33528), .B(g33529), .C(g33530), .D(g33531), .Z(II31874) ) ;
OR3     gate19199  (.A(g33532), .B(II31873), .C(II31874), .Z(g33958) ) ;
NOR3    gate19200  (.A(g31566), .B(II29985), .C(II29986), .Z(g32455) ) ;
NOR3    gate19201  (.A(g31554), .B(II30054), .C(II30055), .Z(g32520) ) ;
NOR3    gate19202  (.A(g31542), .B(II30123), .C(II30124), .Z(g32585) ) ;
NOR3    gate19203  (.A(g31579), .B(II30192), .C(II30193), .Z(g32650) ) ;
NOR3    gate19204  (.A(g31327), .B(II30261), .C(II30262), .Z(g32715) ) ;
NOR3    gate19205  (.A(g31327), .B(II30330), .C(II30331), .Z(g32780) ) ;
NOR3    gate19206  (.A(g30673), .B(II30399), .C(II30400), .Z(g32845) ) ;
NOR3    gate19207  (.A(g31327), .B(II30468), .C(II30469), .Z(g32910) ) ;
NOR4    gate19208  (.A(g34883), .B(g20277), .C(g20242), .D(g21370), .Z(g34912) ) ;
NAND2   gate19209  (.A(g4593), .B(g4601), .Z(II11824) ) ;
NAND2   gate19210  (.A(g4593), .B(II11824), .Z(II11825) ) ;
NAND2   gate19211  (.A(g4601), .B(II11824), .Z(II11826) ) ;
NAND2   gate19212  (.A(II11825), .B(II11826), .Z(g7133) ) ;
NAND2   gate19213  (.A(g5016), .B(g5062), .Z(g7150) ) ;
NAND2   gate19214  (.A(g5360), .B(g5406), .Z(g7167) ) ;
NAND2   gate19215  (.A(g5706), .B(g5752), .Z(g7184) ) ;
NAND2   gate19216  (.A(g4434), .B(g4401), .Z(II11864) ) ;
NAND2   gate19217  (.A(g4434), .B(II11864), .Z(II11865) ) ;
NAND2   gate19218  (.A(g4401), .B(II11864), .Z(II11866) ) ;
NAND2   gate19219  (.A(g6052), .B(g6098), .Z(g7209) ) ;
NAND2   gate19220  (.A(g4388), .B(g4430), .Z(II11877) ) ;
NAND2   gate19221  (.A(g4388), .B(II11877), .Z(II11878) ) ;
NAND2   gate19222  (.A(g4430), .B(II11877), .Z(II11879) ) ;
NAND2   gate19223  (.A(g4584), .B(g4593), .Z(g7227) ) ;
NAND2   gate19224  (.A(g6398), .B(g6444), .Z(g7228) ) ;
NAND2   gate19225  (.A(g896), .B(g890), .Z(g7442) ) ;
NAND2   gate19226  (.A(g996), .B(g979), .Z(II12074) ) ;
NAND2   gate19227  (.A(g996), .B(II12074), .Z(II12075) ) ;
NAND2   gate19228  (.A(g979), .B(II12074), .Z(II12076) ) ;
NAND2   gate19229  (.A(g1339), .B(g1322), .Z(II12096) ) ;
NAND2   gate19230  (.A(g1339), .B(II12096), .Z(II12097) ) ;
NAND2   gate19231  (.A(g1322), .B(II12096), .Z(II12098) ) ;
NAND2   gate19232  (.A(g1094), .B(g1135), .Z(II12203) ) ;
NAND2   gate19233  (.A(g1094), .B(II12203), .Z(II12204) ) ;
NAND2   gate19234  (.A(g1135), .B(II12203), .Z(II12205) ) ;
NAND2   gate19235  (.A(g1437), .B(g1478), .Z(II12217) ) ;
NAND2   gate19236  (.A(g1437), .B(II12217), .Z(II12218) ) ;
NAND2   gate19237  (.A(g1478), .B(II12217), .Z(II12219) ) ;
NAND2   gate19238  (.A(g1111), .B(g1105), .Z(II12240) ) ;
NAND2   gate19239  (.A(g1111), .B(II12240), .Z(II12241) ) ;
NAND2   gate19240  (.A(g1105), .B(II12240), .Z(II12242) ) ;
NAND2   gate19241  (.A(g1124), .B(g1129), .Z(II12251) ) ;
NAND2   gate19242  (.A(g1124), .B(II12251), .Z(II12252) ) ;
NAND2   gate19243  (.A(g1129), .B(II12251), .Z(II12253) ) ;
NAND2   gate19244  (.A(g1454), .B(g1448), .Z(II12261) ) ;
NAND2   gate19245  (.A(g1454), .B(II12261), .Z(II12262) ) ;
NAND2   gate19246  (.A(g1448), .B(II12261), .Z(II12263) ) ;
NAND2   gate19247  (.A(g1141), .B(g956), .Z(II12269) ) ;
NAND2   gate19248  (.A(g1141), .B(II12269), .Z(II12270) ) ;
NAND2   gate19249  (.A(g956), .B(II12269), .Z(II12271) ) ;
NAND2   gate19250  (.A(g1467), .B(g1472), .Z(II12277) ) ;
NAND2   gate19251  (.A(g1467), .B(II12277), .Z(II12278) ) ;
NAND2   gate19252  (.A(g1472), .B(II12277), .Z(II12279) ) ;
NAND2   gate19253  (.A(g1484), .B(g1300), .Z(II12287) ) ;
NAND2   gate19254  (.A(g1484), .B(II12287), .Z(II12288) ) ;
NAND2   gate19255  (.A(g1300), .B(II12287), .Z(II12289) ) ;
NAND2   gate19256  (.A(g3106), .B(g3111), .Z(II12344) ) ;
NAND2   gate19257  (.A(g3106), .B(II12344), .Z(II12345) ) ;
NAND2   gate19258  (.A(g3111), .B(II12344), .Z(II12346) ) ;
NAND2   gate19259  (.A(g3457), .B(g3462), .Z(II12372) ) ;
NAND2   gate19260  (.A(g3457), .B(II12372), .Z(II12373) ) ;
NAND2   gate19261  (.A(g3462), .B(II12372), .Z(II12374) ) ;
NAND2   gate19262  (.A(g3068), .B(g3072), .Z(g8105) ) ;
NAND2   gate19263  (.A(g3808), .B(g3813), .Z(II12401) ) ;
NAND2   gate19264  (.A(g3808), .B(II12401), .Z(II12402) ) ;
NAND2   gate19265  (.A(g3813), .B(II12401), .Z(II12403) ) ;
NAND2   gate19266  (.A(g3419), .B(g3423), .Z(g8163) ) ;
NAND2   gate19267  (.A(g3770), .B(g3774), .Z(g8227) ) ;
NAND2   gate19268  (.A(g405), .B(g392), .Z(II12468) ) ;
NAND2   gate19269  (.A(g405), .B(II12468), .Z(II12469) ) ;
NAND2   gate19270  (.A(g392), .B(II12468), .Z(II12470) ) ;
NAND3   gate19271  (.A(g4358), .B(g4349), .C(g4340), .Z(g8347) ) ;
NAND2   gate19272  (.A(g191), .B(g194), .Z(II12544) ) ;
NAND2   gate19273  (.A(g191), .B(II12544), .Z(II12545) ) ;
NAND2   gate19274  (.A(g194), .B(II12544), .Z(II12546) ) ;
NAND2   gate19275  (.A(g376), .B(g358), .Z(g8678) ) ;
NAND2   gate19276  (.A(g4291), .B(g4287), .Z(II12728) ) ;
NAND2   gate19277  (.A(g4291), .B(II12728), .Z(II12729) ) ;
NAND2   gate19278  (.A(g4287), .B(II12728), .Z(II12730) ) ;
NAND2   gate19279  (.A(g128), .B(g4646), .Z(g8803) ) ;
NAND2   gate19280  (.A(g5011), .B(g4836), .Z(g8829) ) ;
NAND2   gate19281  (.A(g4831), .B(g4681), .Z(g8847) ) ;
NAND2   gate19282  (.A(g4222), .B(g4235), .Z(II12840) ) ;
NAND2   gate19283  (.A(g4222), .B(II12840), .Z(II12841) ) ;
NAND2   gate19284  (.A(g4235), .B(II12840), .Z(II12842) ) ;
NAND2   gate19285  (.A(g4281), .B(g4277), .Z(II12848) ) ;
NAND2   gate19286  (.A(g4281), .B(II12848), .Z(II12849) ) ;
NAND2   gate19287  (.A(g4277), .B(II12848), .Z(II12850) ) ;
NAND2   gate19288  (.A(g3684), .B(g4871), .Z(g8889) ) ;
NAND2   gate19289  (.A(g4200), .B(g4180), .Z(II12876) ) ;
NAND2   gate19290  (.A(g4200), .B(II12876), .Z(II12877) ) ;
NAND2   gate19291  (.A(g4180), .B(II12876), .Z(II12878) ) ;
NAND2   gate19292  (.A(g3004), .B(g3050), .Z(g9092) ) ;
NAND2   gate19293  (.A(g3355), .B(g3401), .Z(g9177) ) ;
NAND2   gate19294  (.A(g3706), .B(g3752), .Z(g9203) ) ;
NAND2   gate19295  (.A(g847), .B(g812), .Z(g9246) ) ;
NAND2   gate19296  (.A(g5115), .B(g5120), .Z(II13043) ) ;
NAND2   gate19297  (.A(g5115), .B(II13043), .Z(II13044) ) ;
NAND2   gate19298  (.A(g5120), .B(II13043), .Z(II13045) ) ;
NAND2   gate19299  (.A(g4308), .B(g4304), .Z(II13065) ) ;
NAND2   gate19300  (.A(g4308), .B(II13065), .Z(II13066) ) ;
NAND2   gate19301  (.A(g4304), .B(II13065), .Z(II13067) ) ;
NAND2   gate19302  (.A(g5462), .B(g5467), .Z(II13077) ) ;
NAND2   gate19303  (.A(g5462), .B(II13077), .Z(II13078) ) ;
NAND2   gate19304  (.A(g5467), .B(II13077), .Z(II13079) ) ;
NAND2   gate19305  (.A(g827), .B(g832), .Z(g9334) ) ;
NAND2   gate19306  (.A(g5080), .B(g5084), .Z(g9372) ) ;
NAND2   gate19307  (.A(g5808), .B(g5813), .Z(II13109) ) ;
NAND2   gate19308  (.A(g5808), .B(II13109), .Z(II13110) ) ;
NAND2   gate19309  (.A(g5813), .B(II13109), .Z(II13111) ) ;
NAND2   gate19310  (.A(g5424), .B(g5428), .Z(g9442) ) ;
NAND2   gate19311  (.A(g6154), .B(g6159), .Z(II13139) ) ;
NAND2   gate19312  (.A(g6154), .B(II13139), .Z(II13140) ) ;
NAND2   gate19313  (.A(g6159), .B(II13139), .Z(II13141) ) ;
NAND2   gate19314  (.A(g5770), .B(g5774), .Z(g9509) ) ;
NAND2   gate19315  (.A(g6500), .B(g6505), .Z(II13182) ) ;
NAND2   gate19316  (.A(g6500), .B(II13182), .Z(II13183) ) ;
NAND2   gate19317  (.A(g6505), .B(II13182), .Z(II13184) ) ;
NAND2   gate19318  (.A(g6116), .B(g6120), .Z(g9567) ) ;
NAND2   gate19319  (.A(g6462), .B(g6466), .Z(g9629) ) ;
NAND2   gate19320  (.A(g128), .B(g4646), .Z(g9663) ) ;
NAND2   gate19321  (.A(g5011), .B(g4836), .Z(g9715) ) ;
NAND2   gate19322  (.A(g1687), .B(g1691), .Z(II13334) ) ;
NAND2   gate19323  (.A(g1687), .B(II13334), .Z(II13335) ) ;
NAND2   gate19324  (.A(g1691), .B(II13334), .Z(II13336) ) ;
NAND2   gate19325  (.A(g4831), .B(g4681), .Z(g9775) ) ;
NAND2   gate19326  (.A(g269), .B(g246), .Z(II13382) ) ;
NAND2   gate19327  (.A(g269), .B(II13382), .Z(II13383) ) ;
NAND2   gate19328  (.A(g246), .B(II13382), .Z(II13384) ) ;
NAND2   gate19329  (.A(II13383), .B(II13384), .Z(g9823) ) ;
NAND2   gate19330  (.A(g1821), .B(g1825), .Z(II13390) ) ;
NAND2   gate19331  (.A(g1821), .B(II13390), .Z(II13391) ) ;
NAND2   gate19332  (.A(g1825), .B(II13390), .Z(II13392) ) ;
NAND2   gate19333  (.A(g2246), .B(g2250), .Z(II13401) ) ;
NAND2   gate19334  (.A(g2246), .B(II13401), .Z(II13402) ) ;
NAND2   gate19335  (.A(g2250), .B(II13401), .Z(II13403) ) ;
NAND2   gate19336  (.A(g3684), .B(g4871), .Z(g9852) ) ;
NAND2   gate19337  (.A(g262), .B(g239), .Z(II13442) ) ;
NAND2   gate19338  (.A(g262), .B(II13442), .Z(II13443) ) ;
NAND2   gate19339  (.A(g239), .B(II13442), .Z(II13444) ) ;
NAND2   gate19340  (.A(II13443), .B(II13444), .Z(g9904) ) ;
NAND2   gate19341  (.A(g1955), .B(g1959), .Z(II13452) ) ;
NAND2   gate19342  (.A(g1955), .B(II13452), .Z(II13453) ) ;
NAND2   gate19343  (.A(g1959), .B(II13452), .Z(II13454) ) ;
NAND2   gate19344  (.A(g2380), .B(g2384), .Z(II13462) ) ;
NAND2   gate19345  (.A(g2380), .B(II13462), .Z(II13463) ) ;
NAND2   gate19346  (.A(g2384), .B(II13462), .Z(II13464) ) ;
NAND2   gate19347  (.A(g255), .B(g232), .Z(II13497) ) ;
NAND2   gate19348  (.A(g255), .B(II13497), .Z(II13498) ) ;
NAND2   gate19349  (.A(g232), .B(II13497), .Z(II13499) ) ;
NAND2   gate19350  (.A(II13498), .B(II13499), .Z(g9966) ) ;
NAND2   gate19351  (.A(g2089), .B(g2093), .Z(II13509) ) ;
NAND2   gate19352  (.A(g2089), .B(II13509), .Z(II13510) ) ;
NAND2   gate19353  (.A(g2093), .B(II13509), .Z(II13511) ) ;
NAND2   gate19354  (.A(g2514), .B(g2518), .Z(II13518) ) ;
NAND2   gate19355  (.A(g2514), .B(II13518), .Z(II13519) ) ;
NAND2   gate19356  (.A(g2518), .B(II13518), .Z(II13520) ) ;
NAND2   gate19357  (.A(g2648), .B(g2652), .Z(II13564) ) ;
NAND2   gate19358  (.A(g2648), .B(II13564), .Z(II13565) ) ;
NAND2   gate19359  (.A(g2652), .B(II13564), .Z(II13566) ) ;
NAND2   gate19360  (.A(g4534), .B(g4537), .Z(II13729) ) ;
NAND2   gate19361  (.A(g4534), .B(II13729), .Z(II13730) ) ;
NAND2   gate19362  (.A(g4537), .B(II13729), .Z(II13731) ) ;
NAND2   gate19363  (.A(g4608), .B(g4584), .Z(II13749) ) ;
NAND2   gate19364  (.A(g4608), .B(II13749), .Z(II13750) ) ;
NAND2   gate19365  (.A(g4584), .B(II13749), .Z(II13751) ) ;
NAND2   gate19366  (.A(II13750), .B(II13751), .Z(g10336) ) ;
NAND2   gate19367  (.A(g862), .B(g7397), .Z(II13850) ) ;
NAND2   gate19368  (.A(g862), .B(II13850), .Z(II13851) ) ;
NAND2   gate19369  (.A(g7397), .B(II13850), .Z(II13852) ) ;
NAND2   gate19370  (.A(g10337), .B(g5022), .Z(g10515) ) ;
NAND2   gate19371  (.A(g7138), .B(g5366), .Z(g10537) ) ;
NAND2   gate19372  (.A(g7157), .B(g5712), .Z(g10561) ) ;
NAND2   gate19373  (.A(g7174), .B(g6058), .Z(g10578) ) ;
NAND2   gate19374  (.A(g7475), .B(g862), .Z(g10583) ) ;
NAND2   gate19375  (.A(g7191), .B(g6404), .Z(g10598) ) ;
NAND2   gate19376  (.A(g896), .B(g7397), .Z(g10601) ) ;
NAND2   gate19377  (.A(g10077), .B(g9751), .Z(g10603) ) ;
NAND2   gate19378  (.A(g10111), .B(g9826), .Z(g10609) ) ;
NAND2   gate19379  (.A(g10115), .B(g9831), .Z(g10611) ) ;
NAND3   gate19380  (.A(g9024), .B(g8977), .C(g8928), .Z(g10614) ) ;
NAND2   gate19381  (.A(g10151), .B(g9909), .Z(g10617) ) ;
NAND2   gate19382  (.A(g10153), .B(g9913), .Z(g10618) ) ;
NAND2   gate19383  (.A(g10178), .B(g9973), .Z(g10622) ) ;
NAND2   gate19384  (.A(g10181), .B(g9976), .Z(g10623) ) ;
NAND2   gate19385  (.A(g10204), .B(g10042), .Z(g10653) ) ;
NOR2    gate19386  (.A(g1183), .B(g1171), .Z(g7304) ) ;
NOR4    gate19387  (.A(g1211), .B(g1216), .C(g1221), .D(g1205), .Z(g7661) ) ;
NAND2   gate19388  (.A(g6961), .B(g9848), .Z(g10737) ) ;
NAND3   gate19389  (.A(g7936), .B(g7913), .C(g8411), .Z(g10754) ) ;
NOR2    gate19390  (.A(g1526), .B(g1514), .Z(g7352) ) ;
NOR4    gate19391  (.A(g1554), .B(g1559), .C(g1564), .D(g1548), .Z(g7675) ) ;
NAND2   gate19392  (.A(g7537), .B(g324), .Z(g10759) ) ;
NAND3   gate19393  (.A(g7960), .B(g7943), .C(g8470), .Z(g10775) ) ;
NAND2   gate19394  (.A(g1146), .B(g7854), .Z(g10916) ) ;
NAND3   gate19395  (.A(g8181), .B(g8137), .C(g417), .Z(g10928) ) ;
NAND2   gate19396  (.A(g1099), .B(g7854), .Z(g10929) ) ;
NAND2   gate19397  (.A(g1489), .B(g7876), .Z(g10946) ) ;
NAND2   gate19398  (.A(g1442), .B(g7876), .Z(g10961) ) ;
NAND2   gate19399  (.A(g7475), .B(g862), .Z(g11002) ) ;
NAND2   gate19400  (.A(g9187), .B(g9040), .Z(g11020) ) ;
NAND3   gate19401  (.A(g8087), .B(g8186), .C(g8239), .Z(g11117) ) ;
NAND2   gate19402  (.A(g8389), .B(g3119), .Z(II14169) ) ;
NAND2   gate19403  (.A(g8389), .B(II14169), .Z(II14170) ) ;
NAND2   gate19404  (.A(g3119), .B(II14169), .Z(II14171) ) ;
NAND3   gate19405  (.A(g8138), .B(g8240), .C(g8301), .Z(g11134) ) ;
NAND2   gate19406  (.A(g8442), .B(g3470), .Z(II14185) ) ;
NAND2   gate19407  (.A(g8442), .B(II14185), .Z(II14186) ) ;
NAND2   gate19408  (.A(g3470), .B(II14185), .Z(II14187) ) ;
NAND2   gate19409  (.A(g8508), .B(g3821), .Z(II14204) ) ;
NAND2   gate19410  (.A(g8508), .B(II14204), .Z(II14205) ) ;
NAND2   gate19411  (.A(g3821), .B(II14204), .Z(II14206) ) ;
NAND2   gate19412  (.A(g9252), .B(g9295), .Z(II14211) ) ;
NAND2   gate19413  (.A(g9252), .B(II14211), .Z(II14212) ) ;
NAND2   gate19414  (.A(g9295), .B(II14211), .Z(II14213) ) ;
NAND3   gate19415  (.A(g4776), .B(g7892), .C(g9030), .Z(g11155) ) ;
NAND2   gate19416  (.A(g979), .B(g8055), .Z(II14228) ) ;
NAND2   gate19417  (.A(g979), .B(II14228), .Z(II14229) ) ;
NAND2   gate19418  (.A(g8055), .B(II14228), .Z(II14230) ) ;
NAND2   gate19419  (.A(II14229), .B(II14230), .Z(g11169) ) ;
NAND2   gate19420  (.A(g8478), .B(g3096), .Z(g11172) ) ;
NAND3   gate19421  (.A(g4966), .B(g7898), .C(g9064), .Z(g11173) ) ;
NAND2   gate19422  (.A(g1322), .B(g8091), .Z(II14247) ) ;
NAND2   gate19423  (.A(g1322), .B(II14247), .Z(II14248) ) ;
NAND2   gate19424  (.A(g8091), .B(II14247), .Z(II14249) ) ;
NAND2   gate19425  (.A(II14248), .B(II14249), .Z(g11189) ) ;
NAND2   gate19426  (.A(g8539), .B(g3447), .Z(g11190) ) ;
NAND2   gate19427  (.A(g8154), .B(g3133), .Z(II14257) ) ;
NAND2   gate19428  (.A(g8154), .B(II14257), .Z(II14258) ) ;
NAND2   gate19429  (.A(g3133), .B(II14257), .Z(II14259) ) ;
NAND2   gate19430  (.A(g8592), .B(g3798), .Z(g11200) ) ;
NAND2   gate19431  (.A(g8218), .B(g3484), .Z(II14275) ) ;
NAND2   gate19432  (.A(g8218), .B(II14275), .Z(II14276) ) ;
NAND2   gate19433  (.A(g3484), .B(II14275), .Z(II14277) ) ;
NAND2   gate19434  (.A(g8282), .B(g3835), .Z(II14289) ) ;
NAND2   gate19435  (.A(g8282), .B(II14289), .Z(II14290) ) ;
NAND2   gate19436  (.A(g3835), .B(II14289), .Z(II14291) ) ;
NAND3   gate19437  (.A(g7636), .B(g7733), .C(g7697), .Z(g11245) ) ;
NAND2   gate19438  (.A(g8438), .B(g3092), .Z(g11251) ) ;
NAND2   gate19439  (.A(g8504), .B(g3443), .Z(g11279) ) ;
NAND2   gate19440  (.A(g225), .B(g9966), .Z(II14330) ) ;
NAND2   gate19441  (.A(g225), .B(II14330), .Z(II14331) ) ;
NAND2   gate19442  (.A(g9966), .B(II14330), .Z(II14332) ) ;
NAND2   gate19443  (.A(II14331), .B(II14332), .Z(g11292) ) ;
NAND2   gate19444  (.A(g8565), .B(g3794), .Z(g11312) ) ;
NAND3   gate19445  (.A(g4633), .B(g4621), .C(g7202), .Z(g11320) ) ;
NAND2   gate19446  (.A(g8890), .B(g8848), .Z(II14350) ) ;
NAND2   gate19447  (.A(g8890), .B(II14350), .Z(II14351) ) ;
NAND2   gate19448  (.A(g8848), .B(II14350), .Z(II14352) ) ;
NAND2   gate19449  (.A(g8481), .B(g3303), .Z(II14368) ) ;
NAND2   gate19450  (.A(g8481), .B(II14368), .Z(II14369) ) ;
NAND2   gate19451  (.A(g3303), .B(II14368), .Z(II14370) ) ;
NAND3   gate19452  (.A(g8644), .B(g6895), .C(g8663), .Z(g11382) ) ;
NAND2   gate19453  (.A(g8542), .B(g3654), .Z(II14398) ) ;
NAND2   gate19454  (.A(g8542), .B(II14398), .Z(II14399) ) ;
NAND2   gate19455  (.A(g3654), .B(II14398), .Z(II14400) ) ;
NAND2   gate19456  (.A(g8713), .B(g4688), .Z(g11396) ) ;
NAND3   gate19457  (.A(g6875), .B(g6895), .C(g8696), .Z(g11410) ) ;
NAND3   gate19458  (.A(g8666), .B(g6918), .C(g8697), .Z(g11412) ) ;
NAND2   gate19459  (.A(g8595), .B(g4005), .Z(II14427) ) ;
NAND2   gate19460  (.A(g8595), .B(II14427), .Z(II14428) ) ;
NAND2   gate19461  (.A(g4005), .B(II14427), .Z(II14429) ) ;
NAND2   gate19462  (.A(g8742), .B(g4878), .Z(g11426) ) ;
NOR2    gate19463  (.A(g3179), .B(g3171), .Z(g8864) ) ;
NAND3   gate19464  (.A(g8644), .B(g3288), .C(g3343), .Z(g11442) ) ;
NAND3   gate19465  (.A(g6905), .B(g6918), .C(g8733), .Z(g11444) ) ;
NAND3   gate19466  (.A(g8700), .B(g6941), .C(g8734), .Z(g11446) ) ;
NAND3   gate19467  (.A(g6875), .B(g3288), .C(g3347), .Z(g11479) ) ;
NOR2    gate19468  (.A(g3530), .B(g3522), .Z(g8906) ) ;
NAND3   gate19469  (.A(g8666), .B(g3639), .C(g3694), .Z(g11490) ) ;
NAND3   gate19470  (.A(g6928), .B(g6941), .C(g8756), .Z(g11492) ) ;
NAND2   gate19471  (.A(g10074), .B(g655), .Z(II14480) ) ;
NAND2   gate19472  (.A(g10074), .B(II14480), .Z(II14481) ) ;
NAND2   gate19473  (.A(g655), .B(II14480), .Z(II14482) ) ;
NAND3   gate19474  (.A(g6905), .B(g3639), .C(g3698), .Z(g11533) ) ;
NOR2    gate19475  (.A(g3881), .B(g3873), .Z(g8958) ) ;
NAND3   gate19476  (.A(g8700), .B(g3990), .C(g4045), .Z(g11544) ) ;
NAND2   gate19477  (.A(g9020), .B(g8737), .Z(II14497) ) ;
NAND2   gate19478  (.A(g9020), .B(II14497), .Z(II14498) ) ;
NAND2   gate19479  (.A(g8737), .B(II14497), .Z(II14499) ) ;
NAND2   gate19480  (.A(g370), .B(g8721), .Z(II14508) ) ;
NAND2   gate19481  (.A(g370), .B(II14508), .Z(II14509) ) ;
NAND2   gate19482  (.A(g8721), .B(II14508), .Z(II14510) ) ;
NAND2   gate19483  (.A(g10147), .B(g661), .Z(II14516) ) ;
NAND2   gate19484  (.A(g10147), .B(II14516), .Z(II14517) ) ;
NAND2   gate19485  (.A(g661), .B(II14516), .Z(II14518) ) ;
NAND3   gate19486  (.A(g6928), .B(g3990), .C(g4049), .Z(g11590) ) ;
NAND2   gate19487  (.A(g8840), .B(g8873), .Z(II14530) ) ;
NAND2   gate19488  (.A(g8840), .B(II14530), .Z(II14531) ) ;
NAND2   gate19489  (.A(g8873), .B(II14530), .Z(II14532) ) ;
NAND2   gate19490  (.A(g8933), .B(g4722), .Z(g11639) ) ;
NAND2   gate19491  (.A(g8676), .B(g4674), .Z(g11674) ) ;
NAND2   gate19492  (.A(g8984), .B(g4912), .Z(g11675) ) ;
NAND2   gate19493  (.A(g8836), .B(g802), .Z(g11679) ) ;
NAND2   gate19494  (.A(g8718), .B(g4864), .Z(g11707) ) ;
NAND2   gate19495  (.A(g8993), .B(g8678), .Z(II14609) ) ;
NAND2   gate19496  (.A(g8993), .B(II14609), .Z(II14610) ) ;
NAND2   gate19497  (.A(g8678), .B(II14609), .Z(II14611) ) ;
NAND2   gate19498  (.A(g9014), .B(g3010), .Z(g11858) ) ;
NAND2   gate19499  (.A(g9060), .B(g3361), .Z(g11881) ) ;
NAND2   gate19500  (.A(g7777), .B(g9086), .Z(g11892) ) ;
NAND2   gate19501  (.A(g9099), .B(g3712), .Z(g11903) ) ;
NAND2   gate19502  (.A(g9671), .B(g5128), .Z(II14712) ) ;
NAND2   gate19503  (.A(g9671), .B(II14712), .Z(II14713) ) ;
NAND2   gate19504  (.A(g5128), .B(II14712), .Z(II14714) ) ;
NAND2   gate19505  (.A(g8187), .B(g1648), .Z(g11914) ) ;
NAND2   gate19506  (.A(g9732), .B(g5475), .Z(II14733) ) ;
NAND2   gate19507  (.A(g9732), .B(II14733), .Z(II14734) ) ;
NAND2   gate19508  (.A(g5475), .B(II14733), .Z(II14735) ) ;
NAND3   gate19509  (.A(g837), .B(g9334), .C(g7197), .Z(g11933) ) ;
NAND2   gate19510  (.A(g8241), .B(g1783), .Z(g11936) ) ;
NAND2   gate19511  (.A(g8259), .B(g2208), .Z(g11938) ) ;
NAND2   gate19512  (.A(g9808), .B(g5821), .Z(II14764) ) ;
NAND2   gate19513  (.A(g9808), .B(II14764), .Z(II14765) ) ;
NAND2   gate19514  (.A(g5821), .B(II14764), .Z(II14766) ) ;
NAND3   gate19515  (.A(g9166), .B(g847), .C(g703), .Z(g11951) ) ;
NAND2   gate19516  (.A(g8302), .B(g1917), .Z(g11955) ) ;
NAND2   gate19517  (.A(g8316), .B(g2342), .Z(g11959) ) ;
NAND2   gate19518  (.A(g9777), .B(g5105), .Z(g11961) ) ;
NAND2   gate19519  (.A(g9891), .B(g6167), .Z(II14788) ) ;
NAND2   gate19520  (.A(g9891), .B(II14788), .Z(II14789) ) ;
NAND2   gate19521  (.A(g6167), .B(II14788), .Z(II14790) ) ;
NAND3   gate19522  (.A(g837), .B(g9334), .C(g9086), .Z(g11968) ) ;
NAND2   gate19523  (.A(g8365), .B(g2051), .Z(g11973) ) ;
NAND2   gate19524  (.A(g8373), .B(g2476), .Z(g11977) ) ;
NAND2   gate19525  (.A(g9861), .B(g5452), .Z(g11979) ) ;
NAND2   gate19526  (.A(g9962), .B(g6513), .Z(II14816) ) ;
NAND2   gate19527  (.A(g9962), .B(II14816), .Z(II14817) ) ;
NAND2   gate19528  (.A(g6513), .B(II14816), .Z(II14818) ) ;
NAND2   gate19529  (.A(g9166), .B(g703), .Z(g11990) ) ;
NAND2   gate19530  (.A(g8418), .B(g2610), .Z(g12000) ) ;
NAND2   gate19531  (.A(g9433), .B(g5142), .Z(II14853) ) ;
NAND2   gate19532  (.A(g9433), .B(II14853), .Z(II14854) ) ;
NAND2   gate19533  (.A(g5142), .B(II14853), .Z(II14855) ) ;
NAND2   gate19534  (.A(g9932), .B(g5798), .Z(g12008) ) ;
NAND2   gate19535  (.A(g7197), .B(g703), .Z(g12014) ) ;
NAND2   gate19536  (.A(g1648), .B(g8093), .Z(g12016) ) ;
NAND2   gate19537  (.A(g9500), .B(g5489), .Z(II14883) ) ;
NAND2   gate19538  (.A(g9500), .B(II14883), .Z(II14884) ) ;
NAND2   gate19539  (.A(g5489), .B(II14883), .Z(II14885) ) ;
NAND2   gate19540  (.A(g10000), .B(g6144), .Z(g12035) ) ;
NAND2   gate19541  (.A(g9086), .B(g703), .Z(g12042) ) ;
NAND2   gate19542  (.A(g1657), .B(g8139), .Z(g12044) ) ;
NAND2   gate19543  (.A(g1783), .B(g8146), .Z(g12045) ) ;
NAND2   gate19544  (.A(g2208), .B(g8150), .Z(g12049) ) ;
NAND2   gate19545  (.A(g9558), .B(g5835), .Z(II14923) ) ;
NAND2   gate19546  (.A(g9558), .B(II14923), .Z(II14924) ) ;
NAND2   gate19547  (.A(g5835), .B(II14923), .Z(II14925) ) ;
NAND2   gate19548  (.A(g10058), .B(g6490), .Z(g12073) ) ;
NAND2   gate19549  (.A(g8187), .B(g8093), .Z(g12078) ) ;
NAND2   gate19550  (.A(g1792), .B(g8195), .Z(g12079) ) ;
NAND2   gate19551  (.A(g1917), .B(g8201), .Z(g12080) ) ;
NAND2   gate19552  (.A(g2217), .B(g8205), .Z(g12083) ) ;
NAND2   gate19553  (.A(g2342), .B(g8211), .Z(g12084) ) ;
NAND2   gate19554  (.A(g9620), .B(g6181), .Z(II14955) ) ;
NAND2   gate19555  (.A(g9620), .B(II14955), .Z(II14956) ) ;
NAND2   gate19556  (.A(g6181), .B(II14955), .Z(II14957) ) ;
NAND2   gate19557  (.A(g847), .B(g9166), .Z(g12111) ) ;
NAND2   gate19558  (.A(g8139), .B(g1624), .Z(g12112) ) ;
NAND2   gate19559  (.A(g8241), .B(g8146), .Z(g12114) ) ;
NAND2   gate19560  (.A(g1926), .B(g8249), .Z(g12115) ) ;
NAND2   gate19561  (.A(g2051), .B(g8255), .Z(g12116) ) ;
NAND2   gate19562  (.A(g8259), .B(g8150), .Z(g12118) ) ;
NAND2   gate19563  (.A(g2351), .B(g8267), .Z(g12119) ) ;
NAND2   gate19564  (.A(g2476), .B(g8273), .Z(g12120) ) ;
NAND2   gate19565  (.A(g8741), .B(g4674), .Z(g12124) ) ;
NAND2   gate19566  (.A(g9728), .B(g5101), .Z(g12125) ) ;
NAND2   gate19567  (.A(g9685), .B(g6527), .Z(II14991) ) ;
NAND2   gate19568  (.A(g9685), .B(II14991), .Z(II14992) ) ;
NAND2   gate19569  (.A(g6527), .B(II14991), .Z(II14993) ) ;
NAND2   gate19570  (.A(g9691), .B(g1700), .Z(II15002) ) ;
NAND2   gate19571  (.A(g9691), .B(II15002), .Z(II15003) ) ;
NAND2   gate19572  (.A(g1700), .B(II15002), .Z(II15004) ) ;
NAND2   gate19573  (.A(g8195), .B(g1760), .Z(g12145) ) ;
NAND2   gate19574  (.A(g8302), .B(g8201), .Z(g12147) ) ;
NAND2   gate19575  (.A(g2060), .B(g8310), .Z(g12148) ) ;
NAND2   gate19576  (.A(g8205), .B(g2185), .Z(g12149) ) ;
NAND2   gate19577  (.A(g8316), .B(g8211), .Z(g12151) ) ;
NAND2   gate19578  (.A(g2485), .B(g8324), .Z(g12152) ) ;
NAND2   gate19579  (.A(g2610), .B(g8330), .Z(g12153) ) ;
NAND2   gate19580  (.A(g8765), .B(g4864), .Z(g12159) ) ;
NAND2   gate19581  (.A(g9804), .B(g5448), .Z(g12169) ) ;
NAND2   gate19582  (.A(g9905), .B(g799), .Z(g12185) ) ;
NAND2   gate19583  (.A(g9752), .B(g1834), .Z(II15041) ) ;
NAND2   gate19584  (.A(g9752), .B(II15041), .Z(II15042) ) ;
NAND2   gate19585  (.A(g1834), .B(II15041), .Z(II15043) ) ;
NAND2   gate19586  (.A(g8249), .B(g1894), .Z(g12188) ) ;
NAND2   gate19587  (.A(g8365), .B(g8255), .Z(g12190) ) ;
NAND2   gate19588  (.A(g9759), .B(g2259), .Z(II15051) ) ;
NAND2   gate19589  (.A(g9759), .B(II15051), .Z(II15052) ) ;
NAND2   gate19590  (.A(g2259), .B(II15051), .Z(II15053) ) ;
NAND2   gate19591  (.A(g8267), .B(g2319), .Z(g12192) ) ;
NAND2   gate19592  (.A(g8373), .B(g8273), .Z(g12194) ) ;
NAND2   gate19593  (.A(g2619), .B(g8381), .Z(g12195) ) ;
NAND2   gate19594  (.A(g8764), .B(g4688), .Z(g12196) ) ;
NAND2   gate19595  (.A(g9887), .B(g5794), .Z(g12207) ) ;
NAND2   gate19596  (.A(g9827), .B(g1968), .Z(II15078) ) ;
NAND2   gate19597  (.A(g9827), .B(II15078), .Z(II15079) ) ;
NAND2   gate19598  (.A(g1968), .B(II15078), .Z(II15080) ) ;
NAND2   gate19599  (.A(g8310), .B(g2028), .Z(g12222) ) ;
NAND2   gate19600  (.A(g9832), .B(g2393), .Z(II15087) ) ;
NAND2   gate19601  (.A(g9832), .B(II15087), .Z(II15088) ) ;
NAND2   gate19602  (.A(g2393), .B(II15087), .Z(II15089) ) ;
NAND2   gate19603  (.A(g8324), .B(g2453), .Z(g12225) ) ;
NAND2   gate19604  (.A(g8418), .B(g8330), .Z(g12227) ) ;
NAND2   gate19605  (.A(g8804), .B(g4878), .Z(g12232) ) ;
NAND2   gate19606  (.A(g9780), .B(g5313), .Z(II15105) ) ;
NAND2   gate19607  (.A(g9780), .B(II15105), .Z(II15106) ) ;
NAND2   gate19608  (.A(g5313), .B(II15105), .Z(II15107) ) ;
NAND2   gate19609  (.A(g9958), .B(g6140), .Z(g12255) ) ;
NAND2   gate19610  (.A(g9910), .B(g2102), .Z(II15121) ) ;
NAND2   gate19611  (.A(g9910), .B(II15121), .Z(II15122) ) ;
NAND2   gate19612  (.A(g2102), .B(II15121), .Z(II15123) ) ;
NAND2   gate19613  (.A(g9914), .B(g2527), .Z(II15128) ) ;
NAND2   gate19614  (.A(g9914), .B(II15128), .Z(II15129) ) ;
NAND2   gate19615  (.A(g2527), .B(II15128), .Z(II15130) ) ;
NAND2   gate19616  (.A(g8381), .B(g2587), .Z(g12287) ) ;
NAND3   gate19617  (.A(g9978), .B(g9766), .C(g9708), .Z(g12289) ) ;
NAND2   gate19618  (.A(g4698), .B(g8933), .Z(g12292) ) ;
NAND3   gate19619  (.A(g10044), .B(g7018), .C(g10090), .Z(g12294) ) ;
NAND2   gate19620  (.A(g9864), .B(g5659), .Z(II15147) ) ;
NAND2   gate19621  (.A(g9864), .B(II15147), .Z(II15148) ) ;
NAND2   gate19622  (.A(g5659), .B(II15147), .Z(II15149) ) ;
NAND2   gate19623  (.A(g10026), .B(g6486), .Z(g12317) ) ;
NAND2   gate19624  (.A(g9480), .B(g640), .Z(g12323) ) ;
NAND2   gate19625  (.A(g9904), .B(g9823), .Z(II15166) ) ;
NAND2   gate19626  (.A(g9904), .B(II15166), .Z(II15167) ) ;
NAND2   gate19627  (.A(g9823), .B(II15166), .Z(II15168) ) ;
NAND2   gate19628  (.A(II15167), .B(II15168), .Z(g12332) ) ;
NAND2   gate19629  (.A(g9977), .B(g2661), .Z(II15174) ) ;
NAND2   gate19630  (.A(g9977), .B(II15174), .Z(II15175) ) ;
NAND2   gate19631  (.A(g2661), .B(II15174), .Z(II15176) ) ;
NAND2   gate19632  (.A(g4888), .B(g8984), .Z(g12340) ) ;
NAND3   gate19633  (.A(g7004), .B(g7018), .C(g10129), .Z(g12342) ) ;
NAND3   gate19634  (.A(g10093), .B(g7041), .C(g10130), .Z(g12344) ) ;
NAND2   gate19635  (.A(g9935), .B(g6005), .Z(II15193) ) ;
NAND2   gate19636  (.A(g9935), .B(II15193), .Z(II15194) ) ;
NAND2   gate19637  (.A(g6005), .B(II15193), .Z(II15195) ) ;
NAND2   gate19638  (.A(g10035), .B(g1714), .Z(II15212) ) ;
NAND2   gate19639  (.A(g10035), .B(II15212), .Z(II15213) ) ;
NAND2   gate19640  (.A(g1714), .B(II15212), .Z(II15214) ) ;
NOR2    gate19641  (.A(g5188), .B(g5180), .Z(g10266) ) ;
NAND3   gate19642  (.A(g10044), .B(g5297), .C(g5348), .Z(g12412) ) ;
NAND3   gate19643  (.A(g7028), .B(g7041), .C(g10165), .Z(g12414) ) ;
NAND3   gate19644  (.A(g10133), .B(g7064), .C(g10166), .Z(g12416) ) ;
NAND2   gate19645  (.A(g10003), .B(g6351), .Z(II15241) ) ;
NAND2   gate19646  (.A(g10003), .B(II15241), .Z(II15242) ) ;
NAND2   gate19647  (.A(g6351), .B(II15241), .Z(II15243) ) ;
NAND2   gate19648  (.A(g10078), .B(g1848), .Z(II15253) ) ;
NAND2   gate19649  (.A(g10078), .B(II15253), .Z(II15254) ) ;
NAND2   gate19650  (.A(g1848), .B(II15253), .Z(II15255) ) ;
NAND2   gate19651  (.A(g10081), .B(g2273), .Z(II15262) ) ;
NAND2   gate19652  (.A(g10081), .B(II15262), .Z(II15263) ) ;
NAND2   gate19653  (.A(g2273), .B(II15262), .Z(II15264) ) ;
NAND3   gate19654  (.A(g7004), .B(g5297), .C(g5352), .Z(g12449) ) ;
NOR2    gate19655  (.A(g5535), .B(g5527), .Z(g10281) ) ;
NAND3   gate19656  (.A(g10093), .B(g5644), .C(g5694), .Z(g12460) ) ;
NAND3   gate19657  (.A(g7051), .B(g7064), .C(g10190), .Z(g12462) ) ;
NAND3   gate19658  (.A(g10169), .B(g7087), .C(g10191), .Z(g12464) ) ;
NAND2   gate19659  (.A(g10061), .B(g6697), .Z(II15287) ) ;
NAND2   gate19660  (.A(g10061), .B(II15287), .Z(II15288) ) ;
NAND2   gate19661  (.A(g6697), .B(II15287), .Z(II15289) ) ;
NAND2   gate19662  (.A(g10112), .B(g1982), .Z(II15298) ) ;
NAND2   gate19663  (.A(g10112), .B(II15298), .Z(II15299) ) ;
NAND2   gate19664  (.A(g1982), .B(II15298), .Z(II15300) ) ;
NAND2   gate19665  (.A(g10116), .B(g2407), .Z(II15306) ) ;
NAND2   gate19666  (.A(g10116), .B(II15306), .Z(II15307) ) ;
NAND2   gate19667  (.A(g2407), .B(II15306), .Z(II15308) ) ;
NAND3   gate19668  (.A(g7285), .B(g4462), .C(g6961), .Z(g12491) ) ;
NAND3   gate19669  (.A(g7028), .B(g5644), .C(g5698), .Z(g12511) ) ;
NOR2    gate19670  (.A(g5881), .B(g5873), .Z(g10312) ) ;
NAND3   gate19671  (.A(g10133), .B(g5990), .C(g6040), .Z(g12522) ) ;
NAND3   gate19672  (.A(g7074), .B(g7087), .C(g10212), .Z(g12524) ) ;
NAND3   gate19673  (.A(g10194), .B(g7110), .C(g10213), .Z(g12526) ) ;
NAND2   gate19674  (.A(g10152), .B(g2116), .Z(II15333) ) ;
NAND2   gate19675  (.A(g10152), .B(II15333), .Z(II15334) ) ;
NAND2   gate19676  (.A(g2116), .B(II15333), .Z(II15335) ) ;
NAND2   gate19677  (.A(g10154), .B(g2541), .Z(II15340) ) ;
NAND2   gate19678  (.A(g10154), .B(II15340), .Z(II15341) ) ;
NAND2   gate19679  (.A(g2541), .B(II15340), .Z(II15342) ) ;
NAND3   gate19680  (.A(g7051), .B(g5990), .C(g6044), .Z(g12577) ) ;
NOR2    gate19681  (.A(g6227), .B(g6219), .Z(g10341) ) ;
NAND3   gate19682  (.A(g10169), .B(g6336), .C(g6386), .Z(g12588) ) ;
NAND3   gate19683  (.A(g7097), .B(g7110), .C(g10229), .Z(g12590) ) ;
NAND2   gate19684  (.A(g10182), .B(g2675), .Z(II15363) ) ;
NAND2   gate19685  (.A(g10182), .B(II15363), .Z(II15364) ) ;
NAND2   gate19686  (.A(g2675), .B(II15363), .Z(II15365) ) ;
NAND3   gate19687  (.A(g7074), .B(g6336), .C(g6390), .Z(g12628) ) ;
NOR2    gate19688  (.A(g6573), .B(g6565), .Z(g7142) ) ;
NAND3   gate19689  (.A(g10194), .B(g6682), .C(g6732), .Z(g12639) ) ;
NAND3   gate19690  (.A(g7097), .B(g6682), .C(g6736), .Z(g12686) ) ;
NAND2   gate19691  (.A(g4467), .B(g6961), .Z(g12767) ) ;
NAND2   gate19692  (.A(g4467), .B(g6961), .Z(g12796) ) ;
NAND4   gate19693  (.A(g10275), .B(g7655), .C(g7643), .D(g7627), .Z(g12797) ) ;
NAND2   gate19694  (.A(g9848), .B(g6961), .Z(g12819) ) ;
NAND4   gate19695  (.A(g6978), .B(g7236), .C(g7224), .D(g7163), .Z(g12822) ) ;
NOR2    gate19696  (.A(g9472), .B(g9407), .Z(g12806) ) ;
NOR2    gate19697  (.A(g9631), .B(g6565), .Z(g12632) ) ;
NAND3   gate19698  (.A(g4388), .B(g7178), .C(g10476), .Z(g12969) ) ;
NAND3   gate19699  (.A(g9024), .B(g8977), .C(g10664), .Z(g12971) ) ;
NAND3   gate19700  (.A(g4392), .B(g10476), .C(g4401), .Z(g12999) ) ;
NOR2    gate19701  (.A(g5297), .B(g7004), .Z(g12002) ) ;
NAND4   gate19702  (.A(g5196), .B(g12002), .C(g5308), .D(g9780), .Z(g13040) ) ;
NAND2   gate19703  (.A(g10521), .B(g969), .Z(g13043) ) ;
NOR2    gate19704  (.A(g5644), .B(g7028), .Z(g12029) ) ;
NAND4   gate19705  (.A(g5543), .B(g12029), .C(g5654), .D(g9864), .Z(g13050) ) ;
NAND2   gate19706  (.A(g969), .B(g11294), .Z(g13057) ) ;
NAND2   gate19707  (.A(g10544), .B(g1312), .Z(g13058) ) ;
NAND3   gate19708  (.A(g4430), .B(g7178), .C(g10590), .Z(g13066) ) ;
NOR2    gate19709  (.A(g9853), .B(g7004), .Z(g12059) ) ;
NAND4   gate19710  (.A(g5240), .B(g12059), .C(g5331), .D(g9780), .Z(g13067) ) ;
NOR2    gate19711  (.A(g5990), .B(g7051), .Z(g12067) ) ;
NAND4   gate19712  (.A(g5889), .B(g12067), .C(g6000), .D(g9935), .Z(g13069) ) ;
NAND2   gate19713  (.A(g1312), .B(g11336), .Z(g13079) ) ;
NAND3   gate19714  (.A(g4392), .B(g10590), .C(g4434), .Z(g13083) ) ;
NOR2    gate19715  (.A(g9924), .B(g7028), .Z(g12093) ) ;
NAND4   gate19716  (.A(g5587), .B(g12093), .C(g5677), .D(g9864), .Z(g13084) ) ;
NOR2    gate19717  (.A(g6336), .B(g7074), .Z(g12101) ) ;
NAND4   gate19718  (.A(g6235), .B(g12101), .C(g6346), .D(g10003), .Z(g13086) ) ;
NAND2   gate19719  (.A(g1061), .B(g10761), .Z(g13092) ) ;
NOR2    gate19720  (.A(g1183), .B(g8407), .Z(g10649) ) ;
NAND4   gate19721  (.A(g5204), .B(g12002), .C(g5339), .D(g9780), .Z(g13097) ) ;
NOR2    gate19722  (.A(g9992), .B(g7051), .Z(g12129) ) ;
NAND4   gate19723  (.A(g5933), .B(g12129), .C(g6023), .D(g9935), .Z(g13098) ) ;
NOR2    gate19724  (.A(g6682), .B(g7097), .Z(g12137) ) ;
NAND4   gate19725  (.A(g6581), .B(g12137), .C(g6692), .D(g10061), .Z(g13100) ) ;
NAND2   gate19726  (.A(g1404), .B(g10794), .Z(g13104) ) ;
NOR2    gate19727  (.A(g1526), .B(g8466), .Z(g10671) ) ;
NAND4   gate19728  (.A(g5551), .B(g12029), .C(g5685), .D(g9864), .Z(g13108) ) ;
NOR2    gate19729  (.A(g10050), .B(g7074), .Z(g12173) ) ;
NAND4   gate19730  (.A(g6279), .B(g12173), .C(g6369), .D(g10003), .Z(g13109) ) ;
NAND3   gate19731  (.A(g1008), .B(g11786), .C(g11294), .Z(g13115) ) ;
NAND4   gate19732  (.A(g5897), .B(g12067), .C(g6031), .D(g9935), .Z(g13118) ) ;
NOR2    gate19733  (.A(g10099), .B(g7097), .Z(g12211) ) ;
NAND4   gate19734  (.A(g6625), .B(g12211), .C(g6715), .D(g10061), .Z(g13119) ) ;
NAND3   gate19735  (.A(g1351), .B(g11815), .C(g11336), .Z(g13130) ) ;
NAND4   gate19736  (.A(g6243), .B(g12101), .C(g6377), .D(g10003), .Z(g13131) ) ;
NAND4   gate19737  (.A(g6589), .B(g12137), .C(g6723), .D(g10061), .Z(g13139) ) ;
NOR2    gate19738  (.A(g8462), .B(g8407), .Z(g10695) ) ;
NOR2    gate19739  (.A(g8526), .B(g8466), .Z(g10715) ) ;
NAND2   gate19740  (.A(g7479), .B(g10521), .Z(g13210) ) ;
NAND2   gate19741  (.A(g1046), .B(g10521), .Z(g13240) ) ;
NAND2   gate19742  (.A(g7503), .B(g10544), .Z(g13241) ) ;
NOR3    gate19743  (.A(g7635), .B(g7518), .C(g7548), .Z(g11846) ) ;
NAND3   gate19744  (.A(g11846), .B(g11294), .C(g11812), .Z(g13256) ) ;
NAND2   gate19745  (.A(g1389), .B(g10544), .Z(g13257) ) ;
NOR3    gate19746  (.A(g7649), .B(g7534), .C(g7581), .Z(g11869) ) ;
NAND3   gate19747  (.A(g11869), .B(g11336), .C(g11849), .Z(g13264) ) ;
NAND3   gate19748  (.A(g7479), .B(g11294), .C(g11846), .Z(g13459) ) ;
NAND4   gate19749  (.A(g12449), .B(g12412), .C(g12342), .D(g12294), .Z(g13462) ) ;
NAND3   gate19750  (.A(g1008), .B(g11294), .C(g11786), .Z(g13475) ) ;
NAND3   gate19751  (.A(g7503), .B(g11336), .C(g11869), .Z(g13476) ) ;
NAND4   gate19752  (.A(g12511), .B(g12460), .C(g12414), .D(g12344), .Z(g13478) ) ;
NAND4   gate19753  (.A(g12686), .B(g12639), .C(g12590), .D(g12526), .Z(g13479) ) ;
NAND3   gate19754  (.A(g1008), .B(g11786), .C(g7972), .Z(g13495) ) ;
NAND3   gate19755  (.A(g1351), .B(g11336), .C(g11815), .Z(g13496) ) ;
NAND4   gate19756  (.A(g12577), .B(g12522), .C(g12462), .D(g12416), .Z(g13498) ) ;
NAND4   gate19757  (.A(g11479), .B(g11442), .C(g11410), .D(g11382), .Z(g13499) ) ;
NAND4   gate19758  (.A(g182), .B(g174), .C(g203), .D(g12812), .Z(g13511) ) ;
NAND3   gate19759  (.A(g1351), .B(g11815), .C(g8002), .Z(g13513) ) ;
NAND4   gate19760  (.A(g12628), .B(g12588), .C(g12524), .D(g12464), .Z(g13515) ) ;
NAND4   gate19761  (.A(g11533), .B(g11490), .C(g11444), .D(g11412), .Z(g13516) ) ;
NAND4   gate19762  (.A(g182), .B(g168), .C(g203), .D(g12812), .Z(g13527) ) ;
NAND3   gate19763  (.A(g11294), .B(g7549), .C(g1008), .Z(g13528) ) ;
NAND4   gate19764  (.A(g11590), .B(g11544), .C(g11492), .D(g11446), .Z(g13529) ) ;
NAND4   gate19765  (.A(g7972), .B(g10521), .C(g7549), .D(g1008), .Z(g13544) ) ;
NAND4   gate19766  (.A(g11812), .B(g7479), .C(g7903), .D(g10521), .Z(g13551) ) ;
NAND3   gate19767  (.A(g11336), .B(g7582), .C(g1351), .Z(g13554) ) ;
NAND4   gate19768  (.A(g8002), .B(g10544), .C(g7582), .D(g1351), .Z(g13573) ) ;
NAND4   gate19769  (.A(g11849), .B(g7503), .C(g7922), .D(g10544), .Z(g13580) ) ;
NOR2    gate19770  (.A(g9056), .B(g9092), .Z(g11039) ) ;
NAND2   gate19771  (.A(g3021), .B(g11039), .Z(g13600) ) ;
NOR2    gate19772  (.A(g9095), .B(g9177), .Z(g11107) ) ;
NAND2   gate19773  (.A(g3372), .B(g11107), .Z(g13628) ) ;
NAND2   gate19774  (.A(g11797), .B(g11261), .Z(g13634) ) ;
NOR2    gate19775  (.A(g9180), .B(g9203), .Z(g11119) ) ;
NAND2   gate19776  (.A(g3723), .B(g11119), .Z(g13667) ) ;
NAND2   gate19777  (.A(g8933), .B(g11261), .Z(g13672) ) ;
NAND2   gate19778  (.A(g11834), .B(g11283), .Z(g13676) ) ;
NAND2   gate19779  (.A(g11755), .B(g11261), .Z(g13709) ) ;
NAND2   gate19780  (.A(g8984), .B(g11283), .Z(g13712) ) ;
NAND4   gate19781  (.A(g174), .B(g203), .C(g168), .D(g12812), .Z(g13727) ) ;
NAND2   gate19782  (.A(g11773), .B(g11261), .Z(g13739) ) ;
NAND2   gate19783  (.A(g11780), .B(g11283), .Z(g13742) ) ;
NAND2   gate19784  (.A(g11252), .B(g3072), .Z(g13764) ) ;
NAND2   gate19785  (.A(g11804), .B(g11283), .Z(g13779) ) ;
NOR2    gate19786  (.A(g7998), .B(g8037), .Z(g11216) ) ;
NAND2   gate19787  (.A(g11216), .B(g401), .Z(g13795) ) ;
NAND2   gate19788  (.A(g8102), .B(g11273), .Z(g13797) ) ;
NAND2   gate19789  (.A(g11280), .B(g3423), .Z(g13798) ) ;
NAND2   gate19790  (.A(g8160), .B(g11306), .Z(g13822) ) ;
NAND2   gate19791  (.A(g11313), .B(g3774), .Z(g13823) ) ;
NAND2   gate19792  (.A(g4754), .B(g11773), .Z(g13834) ) ;
NAND2   gate19793  (.A(g8224), .B(g11360), .Z(g13851) ) ;
NAND2   gate19794  (.A(g4765), .B(g11797), .Z(g13854) ) ;
NAND2   gate19795  (.A(g4944), .B(g11804), .Z(g13855) ) ;
NOR2    gate19796  (.A(g3288), .B(g6875), .Z(g11194) ) ;
NAND4   gate19797  (.A(g3239), .B(g11194), .C(g3321), .D(g11519), .Z(g13866) ) ;
NAND2   gate19798  (.A(g11773), .B(g4732), .Z(g13870) ) ;
NAND2   gate19799  (.A(g4955), .B(g11834), .Z(g13871) ) ;
NOR2    gate19800  (.A(g3161), .B(g7964), .Z(g11566) ) ;
NOR2    gate19801  (.A(g3179), .B(g8059), .Z(g11729) ) ;
NOR2    gate19802  (.A(g3639), .B(g6905), .Z(g11207) ) ;
NAND4   gate19803  (.A(g3590), .B(g11207), .C(g3672), .D(g11576), .Z(g13882) ) ;
NAND2   gate19804  (.A(g11797), .B(g4727), .Z(g13884) ) ;
NAND2   gate19805  (.A(g11804), .B(g4922), .Z(g13886) ) ;
NOR2    gate19806  (.A(g8107), .B(g3171), .Z(g11435) ) ;
NOR2    gate19807  (.A(g7980), .B(g7964), .Z(g11653) ) ;
NOR2    gate19808  (.A(g8107), .B(g8059), .Z(g11473) ) ;
NAND4   gate19809  (.A(g3227), .B(g11194), .C(g3281), .D(g11350), .Z(g13896) ) ;
NOR2    gate19810  (.A(g8531), .B(g6875), .Z(g11217) ) ;
NAND4   gate19811  (.A(g3211), .B(g11217), .C(g3329), .D(g11519), .Z(g13897) ) ;
NOR2    gate19812  (.A(g3512), .B(g7985), .Z(g11621) ) ;
NOR2    gate19813  (.A(g3530), .B(g8114), .Z(g11747) ) ;
NOR2    gate19814  (.A(g3990), .B(g6928), .Z(g11225) ) ;
NAND4   gate19815  (.A(g3941), .B(g11225), .C(g4023), .D(g11631), .Z(g13907) ) ;
NAND2   gate19816  (.A(g11834), .B(g4917), .Z(g13911) ) ;
NAND4   gate19817  (.A(g3259), .B(g11217), .C(g3267), .D(g11350), .Z(g13918) ) ;
NOR2    gate19818  (.A(g8165), .B(g3522), .Z(g11483) ) ;
NOR2    gate19819  (.A(g8021), .B(g7985), .Z(g11692) ) ;
NOR2    gate19820  (.A(g8165), .B(g8114), .Z(g11527) ) ;
NAND4   gate19821  (.A(g3578), .B(g11207), .C(g3632), .D(g11389), .Z(g13927) ) ;
NOR2    gate19822  (.A(g8584), .B(g6905), .Z(g11238) ) ;
NAND4   gate19823  (.A(g3562), .B(g11238), .C(g3680), .D(g11576), .Z(g13928) ) ;
NOR2    gate19824  (.A(g3863), .B(g8026), .Z(g11669) ) ;
NOR2    gate19825  (.A(g3881), .B(g8172), .Z(g11763) ) ;
NAND2   gate19826  (.A(g691), .B(g11740), .Z(g13945) ) ;
NOR2    gate19827  (.A(g7980), .B(g3155), .Z(g11610) ) ;
NAND4   gate19828  (.A(g3610), .B(g11238), .C(g3618), .D(g11389), .Z(g13958) ) ;
NOR2    gate19829  (.A(g8229), .B(g3873), .Z(g11537) ) ;
NOR2    gate19830  (.A(g8080), .B(g8026), .Z(g11715) ) ;
NOR2    gate19831  (.A(g8229), .B(g8172), .Z(g11584) ) ;
NAND4   gate19832  (.A(g3929), .B(g11225), .C(g3983), .D(g11419), .Z(g13967) ) ;
NOR2    gate19833  (.A(g8623), .B(g6928), .Z(g11255) ) ;
NAND4   gate19834  (.A(g3913), .B(g11255), .C(g4031), .D(g11631), .Z(g13968) ) ;
NOR2    gate19835  (.A(g8021), .B(g3506), .Z(g11658) ) ;
NAND4   gate19836  (.A(g3961), .B(g11255), .C(g3969), .D(g11419), .Z(g13993) ) ;
NOR3    gate19837  (.A(g10295), .B(g3161), .C(g3155), .Z(g11514) ) ;
NAND4   gate19838  (.A(g3199), .B(g11217), .C(g3298), .D(g11519), .Z(g14014) ) ;
NOR2    gate19839  (.A(g8080), .B(g3857), .Z(g11697) ) ;
NOR3    gate19840  (.A(g10323), .B(g3512), .C(g3506), .Z(g11571) ) ;
NAND4   gate19841  (.A(g3550), .B(g11238), .C(g3649), .D(g11576), .Z(g14054) ) ;
NOR3    gate19842  (.A(g7121), .B(g3863), .C(g3857), .Z(g11626) ) ;
NAND4   gate19843  (.A(g3901), .B(g11255), .C(g4000), .D(g11631), .Z(g14088) ) ;
NAND2   gate19844  (.A(g11755), .B(g4717), .Z(g14089) ) ;
NAND2   gate19845  (.A(g11780), .B(g4907), .Z(g14120) ) ;
NAND2   gate19846  (.A(g10685), .B(g10928), .Z(g14123) ) ;
NAND2   gate19847  (.A(g11020), .B(g691), .Z(g14146) ) ;
NAND2   gate19848  (.A(g12111), .B(g9246), .Z(g14279) ) ;
NOR2    gate19849  (.A(g7134), .B(g7150), .Z(g11862) ) ;
NAND2   gate19850  (.A(g5033), .B(g11862), .Z(g14317) ) ;
NOR2    gate19851  (.A(g7153), .B(g7167), .Z(g11885) ) ;
NAND2   gate19852  (.A(g5377), .B(g11885), .Z(g14344) ) ;
NOR2    gate19853  (.A(g7170), .B(g7184), .Z(g11907) ) ;
NAND2   gate19854  (.A(g5723), .B(g11907), .Z(g14379) ) ;
NOR2    gate19855  (.A(g7187), .B(g7209), .Z(g11924) ) ;
NAND2   gate19856  (.A(g6069), .B(g11924), .Z(g14408) ) ;
NAND4   gate19857  (.A(g3187), .B(g11194), .C(g3298), .D(g8481), .Z(g14422) ) ;
NOR2    gate19858  (.A(g7212), .B(g7228), .Z(g11945) ) ;
NAND2   gate19859  (.A(g6415), .B(g11945), .Z(g14434) ) ;
NAND4   gate19860  (.A(g3538), .B(g11207), .C(g3649), .D(g8542), .Z(g14452) ) ;
NAND2   gate19861  (.A(g12126), .B(g5084), .Z(g14489) ) ;
NAND4   gate19862  (.A(g3231), .B(g11217), .C(g3321), .D(g8481), .Z(g14517) ) ;
NAND4   gate19863  (.A(g3889), .B(g11225), .C(g4000), .D(g8595), .Z(g14519) ) ;
NAND2   gate19864  (.A(g9369), .B(g12163), .Z(g14520) ) ;
NAND2   gate19865  (.A(g12170), .B(g5428), .Z(g14521) ) ;
NAND4   gate19866  (.A(g3582), .B(g11238), .C(g3672), .D(g8542), .Z(g14542) ) ;
NAND2   gate19867  (.A(g9439), .B(g12201), .Z(g14547) ) ;
NAND2   gate19868  (.A(g12208), .B(g5774), .Z(g14548) ) ;
NAND4   gate19869  (.A(g3195), .B(g11194), .C(g3329), .D(g8481), .Z(g14569) ) ;
NAND4   gate19870  (.A(g3933), .B(g11255), .C(g4023), .D(g8595), .Z(g14570) ) ;
NAND2   gate19871  (.A(g9506), .B(g12249), .Z(g14573) ) ;
NAND2   gate19872  (.A(g12256), .B(g6120), .Z(g14574) ) ;
NAND4   gate19873  (.A(g3546), .B(g11207), .C(g3680), .D(g8542), .Z(g14590) ) ;
NAND4   gate19874  (.A(g5248), .B(g12002), .C(g5331), .D(g12497), .Z(g14598) ) ;
NAND2   gate19875  (.A(g9564), .B(g12311), .Z(g14600) ) ;
NAND2   gate19876  (.A(g12318), .B(g6466), .Z(g14601) ) ;
NAND4   gate19877  (.A(g3897), .B(g11225), .C(g4031), .D(g8595), .Z(g14625) ) ;
NOR2    gate19878  (.A(g5170), .B(g9206), .Z(g12553) ) ;
NOR2    gate19879  (.A(g5188), .B(g9300), .Z(g12772) ) ;
NAND4   gate19880  (.A(g5595), .B(g12029), .C(g5677), .D(g12563), .Z(g14636) ) ;
NAND2   gate19881  (.A(g9626), .B(g12361), .Z(g14638) ) ;
NAND2   gate19882  (.A(g4743), .B(g11755), .Z(g14655) ) ;
NOR2    gate19883  (.A(g9374), .B(g5180), .Z(g12405) ) ;
NOR2    gate19884  (.A(g9234), .B(g9206), .Z(g12646) ) ;
NOR2    gate19885  (.A(g9374), .B(g9300), .Z(g12443) ) ;
NAND4   gate19886  (.A(g5236), .B(g12002), .C(g5290), .D(g12239), .Z(g14663) ) ;
NAND4   gate19887  (.A(g5220), .B(g12059), .C(g5339), .D(g12497), .Z(g14664) ) ;
NOR2    gate19888  (.A(g5517), .B(g9239), .Z(g12604) ) ;
NOR2    gate19889  (.A(g5535), .B(g9381), .Z(g12798) ) ;
NAND4   gate19890  (.A(g5941), .B(g12067), .C(g6023), .D(g12614), .Z(g14674) ) ;
NAND2   gate19891  (.A(g11292), .B(g12332), .Z(II16778) ) ;
NAND2   gate19892  (.A(g11292), .B(II16778), .Z(II16779) ) ;
NAND2   gate19893  (.A(g12332), .B(II16778), .Z(II16780) ) ;
NAND2   gate19894  (.A(II16779), .B(II16780), .Z(g14677) ) ;
NAND2   gate19895  (.A(g4933), .B(g11780), .Z(g14682) ) ;
NAND4   gate19896  (.A(g5268), .B(g12059), .C(g5276), .D(g12239), .Z(g14686) ) ;
NOR2    gate19897  (.A(g9444), .B(g5527), .Z(g12453) ) ;
NOR2    gate19898  (.A(g9269), .B(g9239), .Z(g12695) ) ;
NOR2    gate19899  (.A(g9444), .B(g9381), .Z(g12505) ) ;
NAND4   gate19900  (.A(g5583), .B(g12029), .C(g5637), .D(g12301), .Z(g14695) ) ;
NAND4   gate19901  (.A(g5567), .B(g12093), .C(g5685), .D(g12563), .Z(g14696) ) ;
NOR2    gate19902  (.A(g5863), .B(g9274), .Z(g12662) ) ;
NOR2    gate19903  (.A(g5881), .B(g9451), .Z(g12824) ) ;
NAND4   gate19904  (.A(g6287), .B(g12101), .C(g6369), .D(g12672), .Z(g14706) ) ;
NOR2    gate19905  (.A(g9234), .B(g5164), .Z(g12593) ) ;
NAND4   gate19906  (.A(g5615), .B(g12093), .C(g5623), .D(g12301), .Z(g14730) ) ;
NOR2    gate19907  (.A(g9511), .B(g5873), .Z(g12515) ) ;
NOR2    gate19908  (.A(g9321), .B(g9274), .Z(g12739) ) ;
NOR2    gate19909  (.A(g9511), .B(g9451), .Z(g12571) ) ;
NAND4   gate19910  (.A(g5929), .B(g12067), .C(g5983), .D(g12351), .Z(g14739) ) ;
NAND4   gate19911  (.A(g5913), .B(g12129), .C(g6031), .D(g12614), .Z(g14740) ) ;
NOR2    gate19912  (.A(g6209), .B(g9326), .Z(g12711) ) ;
NOR2    gate19913  (.A(g6227), .B(g9518), .Z(g10421) ) ;
NAND4   gate19914  (.A(g6633), .B(g12137), .C(g6715), .D(g12721), .Z(g14750) ) ;
NOR2    gate19915  (.A(g9269), .B(g5511), .Z(g12651) ) ;
NAND4   gate19916  (.A(g5961), .B(g12129), .C(g5969), .D(g12351), .Z(g14771) ) ;
NOR2    gate19917  (.A(g9569), .B(g6219), .Z(g12581) ) ;
NOR2    gate19918  (.A(g9402), .B(g9326), .Z(g12780) ) ;
NOR2    gate19919  (.A(g9569), .B(g9518), .Z(g12622) ) ;
NAND4   gate19920  (.A(g6275), .B(g12101), .C(g6329), .D(g12423), .Z(g14780) ) ;
NAND4   gate19921  (.A(g6259), .B(g12173), .C(g6377), .D(g12672), .Z(g14781) ) ;
NOR2    gate19922  (.A(g6555), .B(g9407), .Z(g12755) ) ;
NOR2    gate19923  (.A(g6573), .B(g9576), .Z(g10491) ) ;
NOR3    gate19924  (.A(g7704), .B(g5170), .C(g5164), .Z(g12492) ) ;
NAND4   gate19925  (.A(g5208), .B(g12059), .C(g5308), .D(g12497), .Z(g14803) ) ;
NOR2    gate19926  (.A(g9321), .B(g5857), .Z(g12700) ) ;
NAND4   gate19927  (.A(g6307), .B(g12173), .C(g6315), .D(g12423), .Z(g14820) ) ;
NOR2    gate19928  (.A(g9631), .B(g9576), .Z(g12680) ) ;
NAND4   gate19929  (.A(g6621), .B(g12137), .C(g6675), .D(g12471), .Z(g14829) ) ;
NAND4   gate19930  (.A(g6605), .B(g12211), .C(g6723), .D(g12721), .Z(g14830) ) ;
NOR3    gate19931  (.A(g7738), .B(g5517), .C(g5511), .Z(g12558) ) ;
NAND4   gate19932  (.A(g5555), .B(g12093), .C(g5654), .D(g12563), .Z(g14854) ) ;
NOR2    gate19933  (.A(g9402), .B(g6203), .Z(g12744) ) ;
NAND4   gate19934  (.A(g6653), .B(g12211), .C(g6661), .D(g12471), .Z(g14871) ) ;
NOR3    gate19935  (.A(g7766), .B(g5863), .C(g5857), .Z(g12609) ) ;
NAND4   gate19936  (.A(g5901), .B(g12129), .C(g6000), .D(g12614), .Z(g14898) ) ;
NOR2    gate19937  (.A(g9472), .B(g6549), .Z(g12785) ) ;
NOR3    gate19938  (.A(g7791), .B(g6209), .C(g6203), .Z(g12667) ) ;
NAND4   gate19939  (.A(g6247), .B(g12173), .C(g6346), .D(g12672), .Z(g14946) ) ;
NOR3    gate19940  (.A(g7812), .B(g6555), .C(g6549), .Z(g12716) ) ;
NAND4   gate19941  (.A(g6593), .B(g12211), .C(g6692), .D(g12721), .Z(g14987) ) ;
NOR2    gate19942  (.A(g5297), .B(g12598), .Z(g14399) ) ;
NAND4   gate19943  (.A(g5224), .B(g14399), .C(g5327), .D(g9780), .Z(g15709) ) ;
NAND2   gate19944  (.A(g319), .B(g13385), .Z(g15710) ) ;
NOR2    gate19945  (.A(g5644), .B(g12656), .Z(g14425) ) ;
NAND4   gate19946  (.A(g5571), .B(g14425), .C(g5673), .D(g9864), .Z(g15713) ) ;
NAND3   gate19947  (.A(g336), .B(g305), .C(g13385), .Z(g15715) ) ;
NAND2   gate19948  (.A(g10754), .B(g13092), .Z(g15717) ) ;
NOR2    gate19949  (.A(g9853), .B(g12598), .Z(g14490) ) ;
NAND4   gate19950  (.A(g5256), .B(g14490), .C(g5335), .D(g9780), .Z(g15719) ) ;
NOR2    gate19951  (.A(g5990), .B(g12705), .Z(g14497) ) ;
NAND4   gate19952  (.A(g5917), .B(g14497), .C(g6019), .D(g9935), .Z(g15720) ) ;
NAND3   gate19953  (.A(g7564), .B(g311), .C(g13385), .Z(g15721) ) ;
NAND2   gate19954  (.A(g10775), .B(g13104), .Z(g15723) ) ;
NOR2    gate19955  (.A(g9924), .B(g12656), .Z(g14522) ) ;
NAND4   gate19956  (.A(g5603), .B(g14522), .C(g5681), .D(g9864), .Z(g15725) ) ;
NOR2    gate19957  (.A(g6336), .B(g12749), .Z(g14529) ) ;
NAND4   gate19958  (.A(g6263), .B(g14529), .C(g6365), .D(g10003), .Z(g15726) ) ;
NAND4   gate19959  (.A(g5200), .B(g14399), .C(g5313), .D(g9780), .Z(g15728) ) ;
NOR2    gate19960  (.A(g9992), .B(g12705), .Z(g14549) ) ;
NAND4   gate19961  (.A(g5949), .B(g14549), .C(g6027), .D(g9935), .Z(g15729) ) ;
NOR2    gate19962  (.A(g6682), .B(g12790), .Z(g14556) ) ;
NAND4   gate19963  (.A(g6609), .B(g14556), .C(g6711), .D(g10061), .Z(g15730) ) ;
NAND4   gate19964  (.A(g5228), .B(g12059), .C(g5290), .D(g14631), .Z(g15734) ) ;
NAND4   gate19965  (.A(g5547), .B(g14425), .C(g5659), .D(g9864), .Z(g15735) ) ;
NOR2    gate19966  (.A(g10050), .B(g12749), .Z(g14575) ) ;
NAND4   gate19967  (.A(g6295), .B(g14575), .C(g6373), .D(g10003), .Z(g15736) ) ;
NAND4   gate19968  (.A(g5244), .B(g14490), .C(g5320), .D(g14631), .Z(g15741) ) ;
NAND4   gate19969  (.A(g5575), .B(g12093), .C(g5637), .D(g14669), .Z(g15742) ) ;
NAND4   gate19970  (.A(g5893), .B(g14497), .C(g6005), .D(g9935), .Z(g15743) ) ;
NOR2    gate19971  (.A(g10099), .B(g12790), .Z(g14602) ) ;
NAND4   gate19972  (.A(g6641), .B(g14602), .C(g6719), .D(g10061), .Z(g15744) ) ;
NAND4   gate19973  (.A(g5591), .B(g14522), .C(g5666), .D(g14669), .Z(g15751) ) ;
NAND4   gate19974  (.A(g5921), .B(g12129), .C(g5983), .D(g14701), .Z(g15752) ) ;
NAND4   gate19975  (.A(g6239), .B(g14529), .C(g6351), .D(g10003), .Z(g15753) ) ;
NAND4   gate19976  (.A(g5937), .B(g14549), .C(g6012), .D(g14701), .Z(g15780) ) ;
NAND4   gate19977  (.A(g6267), .B(g12173), .C(g6329), .D(g14745), .Z(g15781) ) ;
NAND4   gate19978  (.A(g6585), .B(g14556), .C(g6697), .D(g10061), .Z(g15782) ) ;
NAND4   gate19979  (.A(g6283), .B(g14575), .C(g6358), .D(g14745), .Z(g15787) ) ;
NAND4   gate19980  (.A(g6613), .B(g12211), .C(g6675), .D(g14786), .Z(g15788) ) ;
NAND4   gate19981  (.A(g6629), .B(g14602), .C(g6704), .D(g14786), .Z(g15798) ) ;
NOR2    gate19982  (.A(g11245), .B(g7666), .Z(g13831) ) ;
NAND2   gate19983  (.A(g4112), .B(g13831), .Z(g15829) ) ;
NOR2    gate19984  (.A(g11330), .B(g11011), .Z(g13336) ) ;
NAND2   gate19985  (.A(g13336), .B(g1129), .Z(II17379) ) ;
NAND2   gate19986  (.A(g13336), .B(II17379), .Z(II17380) ) ;
NAND2   gate19987  (.A(g1129), .B(II17379), .Z(II17381) ) ;
NOR2    gate19988  (.A(g11374), .B(g11017), .Z(g13378) ) ;
NAND2   gate19989  (.A(g13378), .B(g1472), .Z(II17404) ) ;
NAND2   gate19990  (.A(g13378), .B(II17404), .Z(II17405) ) ;
NAND2   gate19991  (.A(g1472), .B(II17404), .Z(II17406) ) ;
NAND2   gate19992  (.A(g13336), .B(g956), .Z(II17446) ) ;
NAND2   gate19993  (.A(g13336), .B(II17446), .Z(II17447) ) ;
NAND2   gate19994  (.A(g956), .B(II17446), .Z(II17448) ) ;
NAND2   gate19995  (.A(g13378), .B(g1300), .Z(II17460) ) ;
NAND2   gate19996  (.A(g13378), .B(II17460), .Z(II17461) ) ;
NAND2   gate19997  (.A(g1300), .B(II17460), .Z(II17462) ) ;
NAND2   gate19998  (.A(g13336), .B(g1105), .Z(II17474) ) ;
NAND2   gate19999  (.A(g13336), .B(II17474), .Z(II17475) ) ;
NAND2   gate20000  (.A(g1105), .B(II17474), .Z(II17476) ) ;
NAND2   gate20001  (.A(g13378), .B(g1448), .Z(II17494) ) ;
NAND2   gate20002  (.A(g13378), .B(II17494), .Z(II17495) ) ;
NAND2   gate20003  (.A(g1448), .B(II17494), .Z(II17496) ) ;
NOR3    gate20004  (.A(g4709), .B(g4785), .C(g11155), .Z(g13883) ) ;
NOR3    gate20005  (.A(g4709), .B(g8796), .C(g11155), .Z(g13908) ) ;
NOR3    gate20006  (.A(g4899), .B(g4975), .C(g11173), .Z(g13910) ) ;
NOR2    gate20007  (.A(g3017), .B(g11858), .Z(g13480) ) ;
NAND2   gate20008  (.A(g9291), .B(g13480), .Z(g16275) ) ;
NAND3   gate20009  (.A(g8102), .B(g8057), .C(g13664), .Z(g16278) ) ;
NOR3    gate20010  (.A(g8883), .B(g4785), .C(g11155), .Z(g13937) ) ;
NOR3    gate20011  (.A(g4899), .B(g8822), .C(g11173), .Z(g13939) ) ;
NOR2    gate20012  (.A(g3368), .B(g11881), .Z(g13501) ) ;
NAND2   gate20013  (.A(g9360), .B(g13501), .Z(g16296) ) ;
NAND3   gate20014  (.A(g8160), .B(g8112), .C(g13706), .Z(g16299) ) ;
NOR3    gate20015  (.A(g8883), .B(g8796), .C(g11155), .Z(g13970) ) ;
NOR3    gate20016  (.A(g8938), .B(g4975), .C(g11173), .Z(g13971) ) ;
NOR2    gate20017  (.A(g3719), .B(g11903), .Z(g13518) ) ;
NAND2   gate20018  (.A(g9429), .B(g13518), .Z(g16316) ) ;
NAND3   gate20019  (.A(g8224), .B(g8170), .C(g13736), .Z(g16319) ) ;
NOR3    gate20020  (.A(g8938), .B(g8822), .C(g11173), .Z(g13996) ) ;
NAND4   gate20021  (.A(g3251), .B(g11194), .C(g3267), .D(g13877), .Z(g16604) ) ;
NOR2    gate20022  (.A(g3288), .B(g11615), .Z(g13700) ) ;
NAND4   gate20023  (.A(g3203), .B(g13700), .C(g3274), .D(g11519), .Z(g16625) ) ;
NAND4   gate20024  (.A(g3602), .B(g11207), .C(g3618), .D(g13902), .Z(g16628) ) ;
NOR2    gate20025  (.A(g3639), .B(g11663), .Z(g13730) ) ;
NAND4   gate20026  (.A(g3554), .B(g13730), .C(g3625), .D(g11576), .Z(g16657) ) ;
NAND4   gate20027  (.A(g3953), .B(g11225), .C(g3969), .D(g13933), .Z(g16660) ) ;
NAND4   gate20028  (.A(g13854), .B(g13834), .C(g14655), .D(g12292), .Z(g16663) ) ;
NAND2   gate20029  (.A(g13336), .B(g1135), .Z(II17883) ) ;
NAND2   gate20030  (.A(g13336), .B(II17883), .Z(II17884) ) ;
NAND2   gate20031  (.A(g1135), .B(II17883), .Z(II17885) ) ;
NAND4   gate20032  (.A(g3255), .B(g13700), .C(g3325), .D(g11519), .Z(g16687) ) ;
NOR2    gate20033  (.A(g3990), .B(g11702), .Z(g13772) ) ;
NAND4   gate20034  (.A(g3905), .B(g13772), .C(g3976), .D(g11631), .Z(g16694) ) ;
NAND4   gate20035  (.A(g13871), .B(g13855), .C(g14682), .D(g12340), .Z(g16696) ) ;
NAND2   gate20036  (.A(g13378), .B(g1478), .Z(II17923) ) ;
NAND2   gate20037  (.A(g13378), .B(II17923), .Z(II17924) ) ;
NAND2   gate20038  (.A(g1478), .B(II17923), .Z(II17925) ) ;
NAND4   gate20039  (.A(g3243), .B(g13700), .C(g3310), .D(g11350), .Z(g16719) ) ;
NAND4   gate20040  (.A(g3606), .B(g13730), .C(g3676), .D(g11576), .Z(g16723) ) ;
NAND4   gate20041  (.A(g13884), .B(g13870), .C(g14089), .D(g11639), .Z(g16728) ) ;
NOR2    gate20042  (.A(g8531), .B(g11615), .Z(g13765) ) ;
NAND4   gate20043  (.A(g3207), .B(g13765), .C(g3303), .D(g11519), .Z(g16741) ) ;
NAND4   gate20044  (.A(g3594), .B(g13730), .C(g3661), .D(g11389), .Z(g16745) ) ;
NAND4   gate20045  (.A(g3957), .B(g13772), .C(g4027), .D(g11631), .Z(g16749) ) ;
NAND4   gate20046  (.A(g13911), .B(g13886), .C(g14120), .D(g11675), .Z(g16757) ) ;
NAND4   gate20047  (.A(g3263), .B(g13765), .C(g3274), .D(g8481), .Z(g16770) ) ;
NOR2    gate20048  (.A(g8584), .B(g11663), .Z(g13799) ) ;
NAND4   gate20049  (.A(g3558), .B(g13799), .C(g3654), .D(g11576), .Z(g16772) ) ;
NAND4   gate20050  (.A(g3945), .B(g13772), .C(g4012), .D(g11419), .Z(g16776) ) ;
NAND4   gate20051  (.A(g3614), .B(g13799), .C(g3625), .D(g8542), .Z(g16813) ) ;
NOR2    gate20052  (.A(g8623), .B(g11702), .Z(g13824) ) ;
NAND4   gate20053  (.A(g3909), .B(g13824), .C(g4005), .D(g11631), .Z(g16815) ) ;
NAND4   gate20054  (.A(g3965), .B(g13824), .C(g3976), .D(g8595), .Z(g16854) ) ;
NAND4   gate20055  (.A(g3223), .B(g13765), .C(g3317), .D(g11519), .Z(g16875) ) ;
NAND4   gate20056  (.A(g3574), .B(g13799), .C(g3668), .D(g11576), .Z(g16925) ) ;
NAND4   gate20057  (.A(g3925), .B(g13824), .C(g4019), .D(g11631), .Z(g16956) ) ;
NOR2    gate20058  (.A(g5029), .B(g10515), .Z(g14194) ) ;
NAND2   gate20059  (.A(g7239), .B(g14194), .Z(g17217) ) ;
NAND3   gate20060  (.A(g9369), .B(g9298), .C(g14376), .Z(g17220) ) ;
NOR2    gate20061  (.A(g9547), .B(g12289), .Z(g14367) ) ;
NAND2   gate20062  (.A(g8612), .B(g14367), .Z(g17225) ) ;
NOR2    gate20063  (.A(g5373), .B(g10537), .Z(g14212) ) ;
NAND2   gate20064  (.A(g7247), .B(g14212), .Z(g17243) ) ;
NAND3   gate20065  (.A(g9439), .B(g9379), .C(g14405), .Z(g17246) ) ;
NOR2    gate20066  (.A(g5719), .B(g10561), .Z(g14228) ) ;
NAND2   gate20067  (.A(g7262), .B(g14228), .Z(g17287) ) ;
NAND3   gate20068  (.A(g9506), .B(g9449), .C(g14431), .Z(g17290) ) ;
NOR2    gate20069  (.A(g6065), .B(g10578), .Z(g14248) ) ;
NAND2   gate20070  (.A(g7297), .B(g14248), .Z(g17312) ) ;
NAND3   gate20071  (.A(g9564), .B(g9516), .C(g14503), .Z(g17315) ) ;
NAND2   gate20072  (.A(g8635), .B(g14367), .Z(g17363) ) ;
NAND2   gate20073  (.A(g8639), .B(g14367), .Z(g17364) ) ;
NOR2    gate20074  (.A(g6411), .B(g10598), .Z(g14272) ) ;
NAND2   gate20075  (.A(g7345), .B(g14272), .Z(g17396) ) ;
NAND3   gate20076  (.A(g9626), .B(g9574), .C(g14535), .Z(g17399) ) ;
NAND4   gate20077  (.A(g3215), .B(g13700), .C(g3317), .D(g8481), .Z(g17468) ) ;
NAND2   gate20078  (.A(g8655), .B(g14367), .Z(g17492) ) ;
NAND2   gate20079  (.A(g8659), .B(g14367), .Z(g17493) ) ;
NAND4   gate20080  (.A(g3566), .B(g13730), .C(g3668), .D(g8542), .Z(g17495) ) ;
NAND4   gate20081  (.A(g3247), .B(g13765), .C(g3325), .D(g8481), .Z(g17513) ) ;
NAND4   gate20082  (.A(g3917), .B(g13772), .C(g4019), .D(g8595), .Z(g17514) ) ;
NAND4   gate20083  (.A(g5260), .B(g12002), .C(g5276), .D(g14631), .Z(g17520) ) ;
NOR2    gate20084  (.A(g12333), .B(g9749), .Z(g14611) ) ;
NAND2   gate20085  (.A(g1677), .B(g14611), .Z(II18485) ) ;
NAND2   gate20086  (.A(g1677), .B(II18485), .Z(II18486) ) ;
NAND2   gate20087  (.A(g14611), .B(II18485), .Z(II18487) ) ;
NAND2   gate20088  (.A(g8579), .B(g14367), .Z(g17571) ) ;
NAND4   gate20089  (.A(g3598), .B(g13799), .C(g3676), .D(g8542), .Z(g17572) ) ;
NAND4   gate20090  (.A(g5212), .B(g14399), .C(g5283), .D(g12497), .Z(g17578) ) ;
NAND4   gate20091  (.A(g5607), .B(g12029), .C(g5623), .D(g14669), .Z(g17581) ) ;
NOR2    gate20092  (.A(g12371), .B(g9824), .Z(g14640) ) ;
NAND2   gate20093  (.A(g1811), .B(g14640), .Z(II18529) ) ;
NAND2   gate20094  (.A(g1811), .B(II18529), .Z(II18530) ) ;
NAND2   gate20095  (.A(g14640), .B(II18529), .Z(II18531) ) ;
NOR2    gate20096  (.A(g12374), .B(g9829), .Z(g14642) ) ;
NAND2   gate20097  (.A(g2236), .B(g14642), .Z(II18536) ) ;
NAND2   gate20098  (.A(g2236), .B(II18536), .Z(II18537) ) ;
NAND2   gate20099  (.A(g14642), .B(II18536), .Z(II18538) ) ;
NAND2   gate20100  (.A(g8616), .B(g14367), .Z(g17595) ) ;
NAND2   gate20101  (.A(g8686), .B(g14367), .Z(g17596) ) ;
NAND4   gate20102  (.A(g3191), .B(g13700), .C(g3303), .D(g8481), .Z(g17597) ) ;
NAND4   gate20103  (.A(g3949), .B(g13824), .C(g4027), .D(g8595), .Z(g17598) ) ;
NAND4   gate20104  (.A(g5559), .B(g14425), .C(g5630), .D(g12563), .Z(g17605) ) ;
NAND4   gate20105  (.A(g5953), .B(g12067), .C(g5969), .D(g14701), .Z(g17608) ) ;
NOR2    gate20106  (.A(g12432), .B(g9907), .Z(g14678) ) ;
NAND2   gate20107  (.A(g1945), .B(g14678), .Z(II18579) ) ;
NAND2   gate20108  (.A(g1945), .B(II18579), .Z(II18580) ) ;
NAND2   gate20109  (.A(g14678), .B(II18579), .Z(II18581) ) ;
NOR2    gate20110  (.A(g12437), .B(g9911), .Z(g14679) ) ;
NAND2   gate20111  (.A(g2370), .B(g14679), .Z(II18587) ) ;
NAND2   gate20112  (.A(g2370), .B(II18587), .Z(II18588) ) ;
NAND2   gate20113  (.A(g14679), .B(II18587), .Z(II18589) ) ;
NAND4   gate20114  (.A(g3219), .B(g11217), .C(g3281), .D(g13877), .Z(g17634) ) ;
NAND4   gate20115  (.A(g3542), .B(g13730), .C(g3654), .D(g8542), .Z(g17635) ) ;
NAND4   gate20116  (.A(g5264), .B(g14399), .C(g5335), .D(g12497), .Z(g17640) ) ;
NAND4   gate20117  (.A(g5905), .B(g14497), .C(g5976), .D(g12614), .Z(g17647) ) ;
NAND4   gate20118  (.A(g6299), .B(g12101), .C(g6315), .D(g14745), .Z(g17650) ) ;
NOR2    gate20119  (.A(g12479), .B(g9971), .Z(g14712) ) ;
NAND2   gate20120  (.A(g2079), .B(g14712), .Z(II18625) ) ;
NAND2   gate20121  (.A(g2079), .B(II18625), .Z(II18626) ) ;
NAND2   gate20122  (.A(g14712), .B(II18625), .Z(II18627) ) ;
NOR2    gate20123  (.A(g12483), .B(g9974), .Z(g14713) ) ;
NAND2   gate20124  (.A(g2504), .B(g14713), .Z(II18633) ) ;
NAND2   gate20125  (.A(g2504), .B(II18633), .Z(II18634) ) ;
NAND2   gate20126  (.A(g14713), .B(II18633), .Z(II18635) ) ;
NAND4   gate20127  (.A(g3235), .B(g13765), .C(g3310), .D(g13877), .Z(g17668) ) ;
NAND4   gate20128  (.A(g3570), .B(g11238), .C(g3632), .D(g13902), .Z(g17669) ) ;
NAND4   gate20129  (.A(g3893), .B(g13772), .C(g4005), .D(g8595), .Z(g17670) ) ;
NAND4   gate20130  (.A(g5252), .B(g14399), .C(g5320), .D(g12239), .Z(g17675) ) ;
NAND4   gate20131  (.A(g5611), .B(g14425), .C(g5681), .D(g12563), .Z(g17679) ) ;
NAND4   gate20132  (.A(g6251), .B(g14529), .C(g6322), .D(g12672), .Z(g17686) ) ;
NAND4   gate20133  (.A(g6645), .B(g12137), .C(g6661), .D(g14786), .Z(g17689) ) ;
NOR2    gate20134  (.A(g12540), .B(g10040), .Z(g14752) ) ;
NAND2   gate20135  (.A(g2638), .B(g14752), .Z(II18680) ) ;
NAND2   gate20136  (.A(g2638), .B(II18680), .Z(II18681) ) ;
NAND2   gate20137  (.A(g14752), .B(II18680), .Z(II18682) ) ;
NAND4   gate20138  (.A(g3586), .B(g13799), .C(g3661), .D(g13902), .Z(g17705) ) ;
NAND4   gate20139  (.A(g3921), .B(g11255), .C(g3983), .D(g13933), .Z(g17706) ) ;
NAND4   gate20140  (.A(g5216), .B(g14490), .C(g5313), .D(g12497), .Z(g17708) ) ;
NAND4   gate20141  (.A(g5599), .B(g14425), .C(g5666), .D(g12301), .Z(g17712) ) ;
NAND4   gate20142  (.A(g5957), .B(g14497), .C(g6027), .D(g12614), .Z(g17716) ) ;
NAND4   gate20143  (.A(g6597), .B(g14556), .C(g6668), .D(g12721), .Z(g17723) ) ;
NAND4   gate20144  (.A(g3937), .B(g13824), .C(g4012), .D(g13933), .Z(g17732) ) ;
NAND4   gate20145  (.A(g5272), .B(g14490), .C(g5283), .D(g9780), .Z(g17734) ) ;
NAND4   gate20146  (.A(g5563), .B(g14522), .C(g5659), .D(g12563), .Z(g17736) ) ;
NAND4   gate20147  (.A(g5945), .B(g14497), .C(g6012), .D(g12351), .Z(g17740) ) ;
NAND4   gate20148  (.A(g6303), .B(g14529), .C(g6373), .D(g12672), .Z(g17744) ) ;
NAND4   gate20149  (.A(g5619), .B(g14522), .C(g5630), .D(g9864), .Z(g17755) ) ;
NAND4   gate20150  (.A(g5909), .B(g14549), .C(g6005), .D(g12614), .Z(g17757) ) ;
NAND4   gate20151  (.A(g6291), .B(g14529), .C(g6358), .D(g12423), .Z(g17761) ) ;
NAND4   gate20152  (.A(g6649), .B(g14556), .C(g6719), .D(g12721), .Z(g17765) ) ;
NAND4   gate20153  (.A(g5965), .B(g14549), .C(g5976), .D(g9935), .Z(g17773) ) ;
NAND4   gate20154  (.A(g6255), .B(g14575), .C(g6351), .D(g12672), .Z(g17775) ) ;
NAND4   gate20155  (.A(g6637), .B(g14556), .C(g6704), .D(g12471), .Z(g17779) ) ;
NAND4   gate20156  (.A(g5232), .B(g14490), .C(g5327), .D(g12497), .Z(g17788) ) ;
NAND4   gate20157  (.A(g6311), .B(g14575), .C(g6322), .D(g10003), .Z(g17790) ) ;
NAND4   gate20158  (.A(g6601), .B(g14602), .C(g6697), .D(g12721), .Z(g17792) ) ;
NAND4   gate20159  (.A(g5579), .B(g14522), .C(g5673), .D(g12563), .Z(g17814) ) ;
NAND4   gate20160  (.A(g6657), .B(g14602), .C(g6668), .D(g10061), .Z(g17816) ) ;
NAND4   gate20161  (.A(g5925), .B(g14549), .C(g6019), .D(g12614), .Z(g17820) ) ;
NAND4   gate20162  (.A(g6271), .B(g14575), .C(g6365), .D(g12672), .Z(g17846) ) ;
NAND4   gate20163  (.A(g6617), .B(g14602), .C(g6711), .D(g12721), .Z(g17872) ) ;
NAND2   gate20164  (.A(g11431), .B(g17794), .Z(g19442) ) ;
NAND2   gate20165  (.A(g11471), .B(g17794), .Z(g19450) ) ;
NAND2   gate20166  (.A(g11562), .B(g17794), .Z(g19466) ) ;
NAND2   gate20167  (.A(g11609), .B(g17794), .Z(g19474) ) ;
NOR2    gate20168  (.A(g7650), .B(g4057), .Z(g10922) ) ;
NOR2    gate20169  (.A(g4064), .B(g8451), .Z(g10899) ) ;
NOR2    gate20170  (.A(g7650), .B(g8451), .Z(g10884) ) ;
NAND3   gate20171  (.A(g1070), .B(g1199), .C(g15995), .Z(g19611) ) ;
NAND3   gate20172  (.A(g1413), .B(g1542), .C(g16047), .Z(g19632) ) ;
NOR2    gate20173  (.A(g13551), .B(g11169), .Z(g16246) ) ;
NAND2   gate20174  (.A(g16246), .B(g990), .Z(II20165) ) ;
NAND2   gate20175  (.A(g16246), .B(II20165), .Z(II20166) ) ;
NAND2   gate20176  (.A(g990), .B(II20165), .Z(II20167) ) ;
NOR2    gate20177  (.A(g13580), .B(g11189), .Z(g16272) ) ;
NAND2   gate20178  (.A(g16272), .B(g1333), .Z(II20187) ) ;
NAND2   gate20179  (.A(g16272), .B(II20187), .Z(II20188) ) ;
NAND2   gate20180  (.A(g1333), .B(II20187), .Z(II20189) ) ;
NAND2   gate20181  (.A(g16246), .B(g11147), .Z(II20203) ) ;
NAND2   gate20182  (.A(g16246), .B(II20203), .Z(II20204) ) ;
NAND2   gate20183  (.A(g11147), .B(II20203), .Z(II20205) ) ;
NAND2   gate20184  (.A(g16272), .B(g11170), .Z(II20221) ) ;
NAND2   gate20185  (.A(g16272), .B(II20221), .Z(II20222) ) ;
NAND2   gate20186  (.A(g11170), .B(II20221), .Z(II20223) ) ;
NAND2   gate20187  (.A(g11403), .B(g17794), .Z(g19886) ) ;
NAND2   gate20188  (.A(g11430), .B(g17794), .Z(g19913) ) ;
NOR2    gate20189  (.A(g8005), .B(g13600), .Z(g16313) ) ;
NAND2   gate20190  (.A(g3029), .B(g16313), .Z(g19916) ) ;
NAND2   gate20191  (.A(g11470), .B(g17794), .Z(g19962) ) ;
NOR2    gate20192  (.A(g8064), .B(g13628), .Z(g16424) ) ;
NAND2   gate20193  (.A(g3380), .B(g16424), .Z(g19965) ) ;
NAND2   gate20194  (.A(g11512), .B(g17794), .Z(g20007) ) ;
NOR2    gate20195  (.A(g8119), .B(g13667), .Z(g16476) ) ;
NAND2   gate20196  (.A(g3731), .B(g16476), .Z(g20011) ) ;
NAND2   gate20197  (.A(g11250), .B(g17794), .Z(g20039) ) ;
NAND2   gate20198  (.A(g11269), .B(g17794), .Z(g20055) ) ;
NAND2   gate20199  (.A(g11293), .B(g17794), .Z(g20068) ) ;
NAND2   gate20200  (.A(g13795), .B(g16521), .Z(g20076) ) ;
NAND2   gate20201  (.A(g11325), .B(g17794), .Z(g20081) ) ;
NAND2   gate20202  (.A(g11373), .B(g17794), .Z(g20092) ) ;
NAND2   gate20203  (.A(g11404), .B(g17794), .Z(g20107) ) ;
NAND2   gate20204  (.A(g16663), .B(g13938), .Z(g20163) ) ;
NOR3    gate20205  (.A(g4776), .B(g4801), .C(g4793), .Z(g8131) ) ;
NAND2   gate20206  (.A(g16876), .B(g8131), .Z(g20172) ) ;
NAND2   gate20207  (.A(g16696), .B(g13972), .Z(g20173) ) ;
NAND2   gate20208  (.A(g13252), .B(g16846), .Z(g20181) ) ;
NOR3    gate20209  (.A(g4966), .B(g4991), .C(g4983), .Z(g8177) ) ;
NAND2   gate20210  (.A(g16926), .B(g8177), .Z(g20186) ) ;
NAND2   gate20211  (.A(g17515), .B(g14187), .Z(II20460) ) ;
NAND2   gate20212  (.A(g17515), .B(II20460), .Z(II20461) ) ;
NAND2   gate20213  (.A(g14187), .B(II20460), .Z(II20462) ) ;
NAND2   gate20214  (.A(g16663), .B(g16728), .Z(II20467) ) ;
NAND2   gate20215  (.A(g16663), .B(II20467), .Z(II20468) ) ;
NAND2   gate20216  (.A(g16728), .B(II20467), .Z(II20469) ) ;
NAND2   gate20217  (.A(II20468), .B(II20469), .Z(g20201) ) ;
NAND2   gate20218  (.A(g16696), .B(g16757), .Z(II20486) ) ;
NAND2   gate20219  (.A(g16696), .B(II20486), .Z(II20487) ) ;
NAND2   gate20220  (.A(g16757), .B(II20486), .Z(II20488) ) ;
NAND2   gate20221  (.A(II20487), .B(II20488), .Z(g20216) ) ;
NOR2    gate20222  (.A(g9253), .B(g14317), .Z(g17284) ) ;
NAND2   gate20223  (.A(g5041), .B(g17284), .Z(g20838) ) ;
NOR2    gate20224  (.A(g9305), .B(g14344), .Z(g17309) ) ;
NAND2   gate20225  (.A(g5385), .B(g17309), .Z(g20979) ) ;
NOR2    gate20226  (.A(g9386), .B(g14379), .Z(g17393) ) ;
NAND2   gate20227  (.A(g5731), .B(g17393), .Z(g21124) ) ;
NOR2    gate20228  (.A(g9456), .B(g14408), .Z(g17420) ) ;
NAND2   gate20229  (.A(g6077), .B(g17420), .Z(g21190) ) ;
NOR2    gate20230  (.A(g9523), .B(g14434), .Z(g17482) ) ;
NAND2   gate20231  (.A(g6423), .B(g17482), .Z(g21253) ) ;
NAND2   gate20232  (.A(g11268), .B(g17157), .Z(g21272) ) ;
NAND2   gate20233  (.A(g11291), .B(g17157), .Z(g21283) ) ;
NAND2   gate20234  (.A(g11324), .B(g17157), .Z(g21294) ) ;
NAND2   gate20235  (.A(g11371), .B(g17157), .Z(g21301) ) ;
NAND2   gate20236  (.A(g11401), .B(g17157), .Z(g21330) ) ;
NAND2   gate20237  (.A(g11402), .B(g17157), .Z(g21331) ) ;
NAND2   gate20238  (.A(g11428), .B(g17157), .Z(g21344) ) ;
NAND2   gate20239  (.A(g11429), .B(g17157), .Z(g21345) ) ;
NAND2   gate20240  (.A(g11467), .B(g17157), .Z(g21353) ) ;
NAND2   gate20241  (.A(g11468), .B(g17157), .Z(g21354) ) ;
NAND2   gate20242  (.A(g11509), .B(g17157), .Z(g21359) ) ;
NAND2   gate20243  (.A(g11510), .B(g17157), .Z(g21360) ) ;
NAND2   gate20244  (.A(g11560), .B(g17157), .Z(g21377) ) ;
NAND2   gate20245  (.A(g11608), .B(g17157), .Z(g21388) ) ;
NAND2   gate20246  (.A(g11652), .B(g17157), .Z(g21403) ) ;
NAND2   gate20247  (.A(g11677), .B(g17157), .Z(g21417) ) ;
NAND4   gate20248  (.A(g4584), .B(g4616), .C(g13202), .D(g19071), .Z(g22306) ) ;
NAND2   gate20249  (.A(g18957), .B(g2886), .Z(g22638) ) ;
NAND2   gate20250  (.A(g7870), .B(g19560), .Z(g22642) ) ;
NAND2   gate20251  (.A(g20136), .B(g18954), .Z(g22643) ) ;
NAND2   gate20252  (.A(g7888), .B(g19581), .Z(g22650) ) ;
NAND2   gate20253  (.A(g20114), .B(g2873), .Z(g22651) ) ;
NAND2   gate20254  (.A(g20136), .B(g94), .Z(g22661) ) ;
NAND2   gate20255  (.A(g7680), .B(g19620), .Z(II21976) ) ;
NAND2   gate20256  (.A(g7680), .B(II21976), .Z(II21977) ) ;
NAND2   gate20257  (.A(g19620), .B(II21976), .Z(II21978) ) ;
NAND2   gate20258  (.A(g18957), .B(g2878), .Z(g22666) ) ;
NAND2   gate20259  (.A(g20219), .B(g2912), .Z(g22668) ) ;
NAND2   gate20260  (.A(g7670), .B(g19638), .Z(II21992) ) ;
NAND2   gate20261  (.A(g7670), .B(II21992), .Z(II21993) ) ;
NAND2   gate20262  (.A(g19638), .B(II21992), .Z(II21994) ) ;
NAND2   gate20263  (.A(g19560), .B(g7870), .Z(g22687) ) ;
NAND2   gate20264  (.A(g20219), .B(g2936), .Z(g22688) ) ;
NAND2   gate20265  (.A(g1193), .B(g19611), .Z(g22709) ) ;
NAND2   gate20266  (.A(g19581), .B(g7888), .Z(g22711) ) ;
NAND2   gate20267  (.A(g18957), .B(g2864), .Z(g22712) ) ;
NAND2   gate20268  (.A(g20114), .B(g2890), .Z(g22713) ) ;
NAND2   gate20269  (.A(g20114), .B(g2999), .Z(g22715) ) ;
NAND2   gate20270  (.A(g1536), .B(g19632), .Z(g22753) ) ;
NAND2   gate20271  (.A(g20114), .B(g19376), .Z(g22754) ) ;
NAND2   gate20272  (.A(g20136), .B(g18984), .Z(g22755) ) ;
NAND2   gate20273  (.A(g20114), .B(g7891), .Z(g22757) ) ;
NAND3   gate20274  (.A(g1193), .B(g19560), .C(g10666), .Z(g22833) ) ;
NAND2   gate20275  (.A(g18918), .B(g2852), .Z(g22836) ) ;
NAND2   gate20276  (.A(g20219), .B(g2907), .Z(g22837) ) ;
NAND2   gate20277  (.A(g20219), .B(g2960), .Z(g22838) ) ;
NAND2   gate20278  (.A(g20114), .B(g2988), .Z(g22839) ) ;
NAND3   gate20279  (.A(g1536), .B(g19581), .C(g10699), .Z(g22850) ) ;
NAND2   gate20280  (.A(g18957), .B(g2856), .Z(g22852) ) ;
NAND2   gate20281  (.A(g20219), .B(g2922), .Z(g22853) ) ;
NAND2   gate20282  (.A(g18918), .B(g2844), .Z(g22874) ) ;
NAND2   gate20283  (.A(g20516), .B(g2980), .Z(g22875) ) ;
NAND2   gate20284  (.A(g18957), .B(g2848), .Z(g22902) ) ;
NAND2   gate20285  (.A(g20219), .B(g2950), .Z(g22921) ) ;
NAND2   gate20286  (.A(g18918), .B(g2860), .Z(g22940) ) ;
NAND2   gate20287  (.A(g20219), .B(g2970), .Z(g22941) ) ;
NAND2   gate20288  (.A(g20114), .B(g2868), .Z(g22984) ) ;
NAND2   gate20289  (.A(g20516), .B(g2984), .Z(g23010) ) ;
NOR2    gate20290  (.A(g3025), .B(g16275), .Z(g19887) ) ;
NAND2   gate20291  (.A(g8097), .B(g19887), .Z(g23105) ) ;
NOR2    gate20292  (.A(g3376), .B(g16296), .Z(g19932) ) ;
NAND2   gate20293  (.A(g8155), .B(g19932), .Z(g23132) ) ;
NOR2    gate20294  (.A(g3727), .B(g16316), .Z(g19981) ) ;
NAND2   gate20295  (.A(g8219), .B(g19981), .Z(g23167) ) ;
NAND2   gate20296  (.A(g20136), .B(g37), .Z(g23195) ) ;
NAND2   gate20297  (.A(g18957), .B(g2882), .Z(g23210) ) ;
NAND2   gate20298  (.A(g18918), .B(g2894), .Z(g23266) ) ;
NAND2   gate20299  (.A(g18957), .B(g2898), .Z(g23281) ) ;
NAND2   gate20300  (.A(g703), .B(g20181), .Z(g23324) ) ;
NOR3    gate20301  (.A(g7928), .B(g4801), .C(g4793), .Z(g11231) ) ;
NAND2   gate20302  (.A(g20201), .B(g11231), .Z(g23357) ) ;
NOR3    gate20303  (.A(g7953), .B(g4991), .C(g4983), .Z(g11248) ) ;
NAND2   gate20304  (.A(g20216), .B(g11248), .Z(g23379) ) ;
NAND2   gate20305  (.A(g11893), .B(g21434), .Z(II22683) ) ;
NAND2   gate20306  (.A(g11893), .B(II22683), .Z(II22684) ) ;
NAND2   gate20307  (.A(g21434), .B(II22683), .Z(II22685) ) ;
NAND2   gate20308  (.A(g11915), .B(g21434), .Z(II22710) ) ;
NAND2   gate20309  (.A(g11915), .B(II22710), .Z(II22711) ) ;
NAND2   gate20310  (.A(g21434), .B(II22710), .Z(II22712) ) ;
NAND2   gate20311  (.A(g11916), .B(g21434), .Z(II22717) ) ;
NAND2   gate20312  (.A(g11916), .B(II22717), .Z(II22718) ) ;
NAND2   gate20313  (.A(g21434), .B(II22717), .Z(II22719) ) ;
NAND2   gate20314  (.A(g11937), .B(g21434), .Z(II22753) ) ;
NAND2   gate20315  (.A(g11937), .B(II22753), .Z(II22754) ) ;
NAND2   gate20316  (.A(g21434), .B(II22753), .Z(II22755) ) ;
NAND2   gate20317  (.A(g11939), .B(g21434), .Z(II22760) ) ;
NAND2   gate20318  (.A(g11939), .B(II22760), .Z(II22761) ) ;
NAND2   gate20319  (.A(g21434), .B(II22760), .Z(II22762) ) ;
NOR2    gate20320  (.A(g5037), .B(g17217), .Z(g20717) ) ;
NAND2   gate20321  (.A(g9364), .B(g20717), .Z(g23623) ) ;
NAND2   gate20322  (.A(g11956), .B(g21434), .Z(II22792) ) ;
NAND2   gate20323  (.A(g11956), .B(II22792), .Z(II22793) ) ;
NAND2   gate20324  (.A(g21434), .B(II22792), .Z(II22794) ) ;
NAND2   gate20325  (.A(g11960), .B(g21434), .Z(II22799) ) ;
NAND2   gate20326  (.A(g11960), .B(II22799), .Z(II22800) ) ;
NAND2   gate20327  (.A(g21434), .B(II22799), .Z(II22801) ) ;
NOR2    gate20328  (.A(g5381), .B(g17243), .Z(g20854) ) ;
NAND2   gate20329  (.A(g9434), .B(g20854), .Z(g23659) ) ;
NAND2   gate20330  (.A(g11978), .B(g21434), .Z(II22822) ) ;
NAND2   gate20331  (.A(g11978), .B(II22822), .Z(II22823) ) ;
NAND2   gate20332  (.A(g21434), .B(II22822), .Z(II22824) ) ;
NOR2    gate20333  (.A(g5727), .B(g17287), .Z(g20995) ) ;
NAND2   gate20334  (.A(g9501), .B(g20995), .Z(g23692) ) ;
NOR2    gate20335  (.A(g1648), .B(g8187), .Z(g12113) ) ;
NAND2   gate20336  (.A(g12113), .B(g21228), .Z(II22844) ) ;
NAND2   gate20337  (.A(g12113), .B(II22844), .Z(II22845) ) ;
NAND2   gate20338  (.A(g21228), .B(II22844), .Z(II22846) ) ;
NOR2    gate20339  (.A(g6073), .B(g17312), .Z(g21140) ) ;
NAND2   gate20340  (.A(g9559), .B(g21140), .Z(g23726) ) ;
NOR2    gate20341  (.A(g1783), .B(g8241), .Z(g12146) ) ;
NAND2   gate20342  (.A(g12146), .B(g21228), .Z(II22864) ) ;
NAND2   gate20343  (.A(g12146), .B(II22864), .Z(II22865) ) ;
NAND2   gate20344  (.A(g21228), .B(II22864), .Z(II22866) ) ;
NOR2    gate20345  (.A(g2208), .B(g8259), .Z(g12150) ) ;
NAND2   gate20346  (.A(g12150), .B(g21228), .Z(II22871) ) ;
NAND2   gate20347  (.A(g12150), .B(II22871), .Z(II22872) ) ;
NAND2   gate20348  (.A(g21228), .B(II22871), .Z(II22873) ) ;
NOR2    gate20349  (.A(g6419), .B(g17396), .Z(g21206) ) ;
NAND2   gate20350  (.A(g9621), .B(g21206), .Z(g23756) ) ;
NOR2    gate20351  (.A(g1917), .B(g8302), .Z(g12189) ) ;
NAND2   gate20352  (.A(g12189), .B(g21228), .Z(II22892) ) ;
NAND2   gate20353  (.A(g12189), .B(II22892), .Z(II22893) ) ;
NAND2   gate20354  (.A(g21228), .B(II22892), .Z(II22894) ) ;
NOR2    gate20355  (.A(g2342), .B(g8316), .Z(g12193) ) ;
NAND2   gate20356  (.A(g12193), .B(g21228), .Z(II22899) ) ;
NAND2   gate20357  (.A(g12193), .B(II22899), .Z(II22900) ) ;
NAND2   gate20358  (.A(g21228), .B(II22899), .Z(II22901) ) ;
NOR2    gate20359  (.A(g16646), .B(g9690), .Z(g21284) ) ;
NAND2   gate20360  (.A(g14677), .B(g21284), .Z(II22921) ) ;
NAND2   gate20361  (.A(g14677), .B(II22921), .Z(II22922) ) ;
NAND2   gate20362  (.A(g21284), .B(II22921), .Z(II22923) ) ;
NOR2    gate20363  (.A(g2051), .B(g8365), .Z(g12223) ) ;
NAND2   gate20364  (.A(g12223), .B(g21228), .Z(II22929) ) ;
NAND2   gate20365  (.A(g12223), .B(II22929), .Z(II22930) ) ;
NAND2   gate20366  (.A(g21228), .B(II22929), .Z(II22931) ) ;
NOR2    gate20367  (.A(g2476), .B(g8373), .Z(g12226) ) ;
NAND2   gate20368  (.A(g12226), .B(g21228), .Z(II22936) ) ;
NAND2   gate20369  (.A(g12226), .B(II22936), .Z(II22937) ) ;
NAND2   gate20370  (.A(g21228), .B(II22936), .Z(II22938) ) ;
NAND2   gate20371  (.A(g9492), .B(g19620), .Z(II22944) ) ;
NAND2   gate20372  (.A(g9492), .B(II22944), .Z(II22945) ) ;
NAND2   gate20373  (.A(g19620), .B(II22944), .Z(II22946) ) ;
NOR2    gate20374  (.A(g2610), .B(g8418), .Z(g12288) ) ;
NAND2   gate20375  (.A(g12288), .B(g21228), .Z(II22965) ) ;
NAND2   gate20376  (.A(g12288), .B(II22965), .Z(II22966) ) ;
NAND2   gate20377  (.A(g21228), .B(II22965), .Z(II22967) ) ;
NAND2   gate20378  (.A(g9657), .B(g19638), .Z(II22972) ) ;
NAND2   gate20379  (.A(g9657), .B(II22972), .Z(II22973) ) ;
NAND2   gate20380  (.A(g19638), .B(II22972), .Z(II22974) ) ;
NAND2   gate20381  (.A(g20076), .B(g417), .Z(II23118) ) ;
NAND2   gate20382  (.A(g20076), .B(II23118), .Z(II23119) ) ;
NAND2   gate20383  (.A(g417), .B(II23118), .Z(II23120) ) ;
NAND2   gate20384  (.A(II23119), .B(II23120), .Z(g23975) ) ;
NAND2   gate20385  (.A(g21370), .B(g22136), .Z(g24362) ) ;
NAND2   gate20386  (.A(g22409), .B(g4332), .Z(II23585) ) ;
NAND2   gate20387  (.A(g22409), .B(II23585), .Z(II23586) ) ;
NAND2   gate20388  (.A(g4332), .B(II23585), .Z(II23587) ) ;
NAND2   gate20389  (.A(II23586), .B(II23587), .Z(g24369) ) ;
NAND2   gate20390  (.A(g22360), .B(g4322), .Z(II23600) ) ;
NAND2   gate20391  (.A(g22360), .B(II23600), .Z(II23601) ) ;
NAND2   gate20392  (.A(g4322), .B(II23600), .Z(II23602) ) ;
NAND2   gate20393  (.A(II23601), .B(II23602), .Z(g24380) ) ;
NAND2   gate20394  (.A(g22957), .B(g2917), .Z(g24567) ) ;
NAND2   gate20395  (.A(g22957), .B(g2941), .Z(g24570) ) ;
NAND2   gate20396  (.A(g22957), .B(g2902), .Z(g24576) ) ;
NAND2   gate20397  (.A(g22957), .B(g2965), .Z(g24601) ) ;
NAND2   gate20398  (.A(g22957), .B(g2927), .Z(g24621) ) ;
NAND2   gate20399  (.A(g22957), .B(g2955), .Z(g24662) ) ;
NAND2   gate20400  (.A(g22957), .B(g2975), .Z(g24677) ) ;
NAND2   gate20401  (.A(g23975), .B(g9333), .Z(II23917) ) ;
NAND2   gate20402  (.A(g23975), .B(II23917), .Z(II23918) ) ;
NAND2   gate20403  (.A(g9333), .B(II23917), .Z(II23919) ) ;
NOR2    gate20404  (.A(g8334), .B(g19916), .Z(g23052) ) ;
NAND2   gate20405  (.A(g3040), .B(g23052), .Z(g24776) ) ;
NOR2    gate20406  (.A(g8390), .B(g19965), .Z(g23079) ) ;
NAND2   gate20407  (.A(g3391), .B(g23079), .Z(g24787) ) ;
NOR2    gate20408  (.A(g8009), .B(g10721), .Z(g13603) ) ;
NAND2   gate20409  (.A(g23162), .B(g13603), .Z(II23949) ) ;
NAND2   gate20410  (.A(g23162), .B(II23949), .Z(II23950) ) ;
NAND2   gate20411  (.A(g13603), .B(II23949), .Z(II23951) ) ;
NOR2    gate20412  (.A(g8443), .B(g20011), .Z(g23124) ) ;
NAND2   gate20413  (.A(g3742), .B(g23124), .Z(g24793) ) ;
NOR2    gate20414  (.A(g8068), .B(g10733), .Z(g13631) ) ;
NAND2   gate20415  (.A(g23184), .B(g13631), .Z(II23961) ) ;
NAND2   gate20416  (.A(g23184), .B(II23961), .Z(II23962) ) ;
NAND2   gate20417  (.A(g13631), .B(II23961), .Z(II23963) ) ;
NAND2   gate20418  (.A(g22202), .B(g490), .Z(II23969) ) ;
NAND2   gate20419  (.A(g22202), .B(II23969), .Z(II23970) ) ;
NAND2   gate20420  (.A(g490), .B(II23969), .Z(II23971) ) ;
NAND2   gate20421  (.A(II23970), .B(II23971), .Z(g24802) ) ;
NOR2    gate20422  (.A(g8123), .B(g10756), .Z(g13670) ) ;
NAND2   gate20423  (.A(g23198), .B(g13670), .Z(II23978) ) ;
NAND2   gate20424  (.A(g23198), .B(II23978), .Z(II23979) ) ;
NAND2   gate20425  (.A(g13670), .B(II23978), .Z(II23980) ) ;
NAND2   gate20426  (.A(g22182), .B(g482), .Z(II23985) ) ;
NAND2   gate20427  (.A(g22182), .B(II23985), .Z(II23986) ) ;
NAND2   gate20428  (.A(g482), .B(II23985), .Z(II23987) ) ;
NAND2   gate20429  (.A(II23986), .B(II23987), .Z(g24808) ) ;
NOR2    gate20430  (.A(g11320), .B(g8347), .Z(g13852) ) ;
NAND2   gate20431  (.A(g534), .B(g23088), .Z(g24905) ) ;
NAND2   gate20432  (.A(g8743), .B(g23088), .Z(g24906) ) ;
NAND2   gate20433  (.A(g19450), .B(g23154), .Z(g24916) ) ;
NAND2   gate20434  (.A(g19913), .B(g23172), .Z(g24917) ) ;
NAND2   gate20435  (.A(g136), .B(g23088), .Z(g24918) ) ;
NAND2   gate20436  (.A(g20007), .B(g23172), .Z(g24924) ) ;
NAND2   gate20437  (.A(g20092), .B(g23154), .Z(g24925) ) ;
NAND2   gate20438  (.A(g19886), .B(g23172), .Z(g24932) ) ;
NAND2   gate20439  (.A(g19466), .B(g23154), .Z(g24933) ) ;
NAND2   gate20440  (.A(g20039), .B(g23172), .Z(g24942) ) ;
NAND2   gate20441  (.A(g20068), .B(g23172), .Z(g24943) ) ;
NAND2   gate20442  (.A(g19442), .B(g23154), .Z(g24950) ) ;
NAND2   gate20443  (.A(g199), .B(g23088), .Z(g24951) ) ;
NAND2   gate20444  (.A(g19962), .B(g23172), .Z(g24972) ) ;
NAND2   gate20445  (.A(g546), .B(g23088), .Z(g24988) ) ;
NAND2   gate20446  (.A(g19474), .B(g23154), .Z(g25002) ) ;
NAND2   gate20447  (.A(g20107), .B(g23154), .Z(g25018) ) ;
NAND2   gate20448  (.A(g20055), .B(g23172), .Z(g25019) ) ;
NAND2   gate20449  (.A(g542), .B(g23088), .Z(g25048) ) ;
NOR2    gate20450  (.A(g9607), .B(g20838), .Z(g23560) ) ;
NAND2   gate20451  (.A(g5052), .B(g23560), .Z(g25172) ) ;
NOR2    gate20452  (.A(g9672), .B(g20979), .Z(g23602) ) ;
NAND2   gate20453  (.A(g5396), .B(g23602), .Z(g25186) ) ;
NOR2    gate20454  (.A(g9257), .B(g11111), .Z(g14320) ) ;
NAND2   gate20455  (.A(g23687), .B(g14320), .Z(II24363) ) ;
NAND2   gate20456  (.A(g23687), .B(II24363), .Z(II24364) ) ;
NAND2   gate20457  (.A(g14320), .B(II24363), .Z(II24365) ) ;
NOR2    gate20458  (.A(g9733), .B(g21124), .Z(g23642) ) ;
NAND2   gate20459  (.A(g5742), .B(g23642), .Z(g25200) ) ;
NOR2    gate20460  (.A(g9309), .B(g11123), .Z(g14347) ) ;
NAND2   gate20461  (.A(g23721), .B(g14347), .Z(II24383) ) ;
NAND2   gate20462  (.A(g23721), .B(II24383), .Z(II24384) ) ;
NAND2   gate20463  (.A(g14347), .B(II24383), .Z(II24385) ) ;
NOR2    gate20464  (.A(g9809), .B(g21190), .Z(g23678) ) ;
NAND2   gate20465  (.A(g6088), .B(g23678), .Z(g25216) ) ;
NOR2    gate20466  (.A(g9390), .B(g11139), .Z(g14382) ) ;
NAND2   gate20467  (.A(g23751), .B(g14382), .Z(II24414) ) ;
NAND2   gate20468  (.A(g23751), .B(II24414), .Z(II24415) ) ;
NAND2   gate20469  (.A(g14382), .B(II24414), .Z(II24416) ) ;
NOR2    gate20470  (.A(g9892), .B(g21253), .Z(g23711) ) ;
NAND2   gate20471  (.A(g6434), .B(g23711), .Z(g25237) ) ;
NOR2    gate20472  (.A(g9460), .B(g11160), .Z(g14411) ) ;
NAND2   gate20473  (.A(g23771), .B(g14411), .Z(II24438) ) ;
NAND2   gate20474  (.A(g23771), .B(II24438), .Z(II24439) ) ;
NAND2   gate20475  (.A(g14411), .B(II24438), .Z(II24440) ) ;
NOR2    gate20476  (.A(g9527), .B(g11178), .Z(g14437) ) ;
NAND2   gate20477  (.A(g23796), .B(g14437), .Z(II24461) ) ;
NAND2   gate20478  (.A(g23796), .B(II24461), .Z(II24462) ) ;
NAND2   gate20479  (.A(g14437), .B(II24461), .Z(II24463) ) ;
NAND2   gate20480  (.A(g538), .B(g23088), .Z(g25381) ) ;
NOR2    gate20481  (.A(g1624), .B(g8139), .Z(g12333) ) ;
NAND2   gate20482  (.A(g20081), .B(g23172), .Z(g25425) ) ;
NOR2    gate20483  (.A(g1760), .B(g8195), .Z(g12371) ) ;
NOR2    gate20484  (.A(g2185), .B(g8205), .Z(g12374) ) ;
NOR2    gate20485  (.A(g1894), .B(g8249), .Z(g12432) ) ;
NOR2    gate20486  (.A(g2319), .B(g8267), .Z(g12437) ) ;
NOR2    gate20487  (.A(g2028), .B(g8310), .Z(g12479) ) ;
NOR2    gate20488  (.A(g2453), .B(g8324), .Z(g12483) ) ;
NOR2    gate20489  (.A(g2587), .B(g8381), .Z(g12540) ) ;
NAND2   gate20490  (.A(g19694), .B(g24362), .Z(g25779) ) ;
NOR4    gate20491  (.A(g20516), .B(g20436), .C(g20219), .D(g22957), .Z(g24631) ) ;
NOR4    gate20492  (.A(g18957), .B(g18918), .C(g20136), .D(g20114), .Z(g23956) ) ;
NOR3    gate20493  (.A(g18957), .B(g20136), .C(g20114), .Z(g22405) ) ;
NOR2    gate20494  (.A(g3034), .B(g23105), .Z(g24751) ) ;
NAND2   gate20495  (.A(g7975), .B(g24751), .Z(g26208) ) ;
NOR2    gate20496  (.A(g3385), .B(g23132), .Z(g24766) ) ;
NAND2   gate20497  (.A(g8016), .B(g24766), .Z(g26235) ) ;
NAND2   gate20498  (.A(g482), .B(g24718), .Z(II25219) ) ;
NAND2   gate20499  (.A(g482), .B(II25219), .Z(II25220) ) ;
NAND2   gate20500  (.A(g24718), .B(II25219), .Z(II25221) ) ;
NAND2   gate20501  (.A(II25220), .B(II25221), .Z(g26248) ) ;
NOR2    gate20502  (.A(g3736), .B(g23167), .Z(g24779) ) ;
NAND2   gate20503  (.A(g8075), .B(g24779), .Z(g26255) ) ;
NAND2   gate20504  (.A(g490), .B(g24744), .Z(II25242) ) ;
NAND2   gate20505  (.A(g490), .B(II25242), .Z(II25243) ) ;
NAND2   gate20506  (.A(g24744), .B(II25242), .Z(II25244) ) ;
NAND2   gate20507  (.A(II25243), .B(II25244), .Z(g26269) ) ;
NOR2    gate20508  (.A(g5046), .B(g23623), .Z(g25144) ) ;
NAND2   gate20509  (.A(g9229), .B(g25144), .Z(g26666) ) ;
NOR2    gate20510  (.A(g5390), .B(g23659), .Z(g25160) ) ;
NAND2   gate20511  (.A(g9264), .B(g25160), .Z(g26685) ) ;
NOR2    gate20512  (.A(g5736), .B(g23692), .Z(g25175) ) ;
NAND2   gate20513  (.A(g9316), .B(g25175), .Z(g26714) ) ;
NOR2    gate20514  (.A(g6082), .B(g23726), .Z(g25189) ) ;
NAND2   gate20515  (.A(g9397), .B(g25189), .Z(g26752) ) ;
NOR2    gate20516  (.A(g6428), .B(g23756), .Z(g25203) ) ;
NAND2   gate20517  (.A(g9467), .B(g25203), .Z(g26782) ) ;
NOR2    gate20518  (.A(g23837), .B(g25408), .Z(g26212) ) ;
NAND2   gate20519  (.A(g26212), .B(g24799), .Z(II25845) ) ;
NAND2   gate20520  (.A(g26212), .B(II25845), .Z(II25846) ) ;
NAND2   gate20521  (.A(g24799), .B(II25845), .Z(II25847) ) ;
NOR2    gate20522  (.A(g23873), .B(g25479), .Z(g26256) ) ;
NAND2   gate20523  (.A(g26256), .B(g24782), .Z(II25907) ) ;
NAND2   gate20524  (.A(g26256), .B(II25907), .Z(II25908) ) ;
NAND2   gate20525  (.A(g24782), .B(II25907), .Z(II25909) ) ;
NOR2    gate20526  (.A(g8480), .B(g12641), .Z(g13500) ) ;
NAND2   gate20527  (.A(g25997), .B(g13500), .Z(II26049) ) ;
NAND2   gate20528  (.A(g25997), .B(II26049), .Z(II26050) ) ;
NAND2   gate20529  (.A(g13500), .B(II26049), .Z(II26051) ) ;
NAND2   gate20530  (.A(g10685), .B(g25930), .Z(g27377) ) ;
NOR2    gate20531  (.A(g8541), .B(g12692), .Z(g13517) ) ;
NAND2   gate20532  (.A(g26026), .B(g13517), .Z(II26070) ) ;
NAND2   gate20533  (.A(g26026), .B(II26070), .Z(II26071) ) ;
NAND2   gate20534  (.A(g13517), .B(II26070), .Z(II26072) ) ;
NOR2    gate20535  (.A(g8594), .B(g12735), .Z(g13539) ) ;
NAND2   gate20536  (.A(g26055), .B(g13539), .Z(II26093) ) ;
NAND2   gate20537  (.A(g26055), .B(II26093), .Z(II26094) ) ;
NAND2   gate20538  (.A(g13539), .B(II26093), .Z(II26095) ) ;
NAND4   gate20539  (.A(g21228), .B(g25243), .C(g26424), .D(g26148), .Z(g27738) ) ;
NOR2    gate20540  (.A(g9779), .B(g10823), .Z(g14211) ) ;
NAND2   gate20541  (.A(g26400), .B(g14211), .Z(II26366) ) ;
NAND2   gate20542  (.A(g26400), .B(II26366), .Z(II26367) ) ;
NAND2   gate20543  (.A(g14211), .B(II26366), .Z(II26368) ) ;
NAND4   gate20544  (.A(g21228), .B(g25262), .C(g26424), .D(g26166), .Z(g27775) ) ;
NAND4   gate20545  (.A(g21228), .B(g25263), .C(g26424), .D(g26171), .Z(g27796) ) ;
NOR2    gate20546  (.A(g9863), .B(g10838), .Z(g14227) ) ;
NAND2   gate20547  (.A(g26488), .B(g14227), .Z(II26393) ) ;
NAND2   gate20548  (.A(g26488), .B(II26393), .Z(II26394) ) ;
NAND2   gate20549  (.A(g14227), .B(II26393), .Z(II26395) ) ;
NAND4   gate20550  (.A(g21228), .B(g25282), .C(g26424), .D(g26190), .Z(g27833) ) ;
NAND4   gate20551  (.A(g21228), .B(g25283), .C(g26424), .D(g26195), .Z(g27854) ) ;
NOR2    gate20552  (.A(g9934), .B(g10869), .Z(g14247) ) ;
NAND2   gate20553  (.A(g26519), .B(g14247), .Z(II26417) ) ;
NAND2   gate20554  (.A(g26519), .B(II26417), .Z(II26418) ) ;
NAND2   gate20555  (.A(g14247), .B(II26417), .Z(II26419) ) ;
NAND4   gate20556  (.A(g21228), .B(g25307), .C(g26424), .D(g26213), .Z(g27882) ) ;
NAND4   gate20557  (.A(g21228), .B(g25316), .C(g26424), .D(g26218), .Z(g27903) ) ;
NOR2    gate20558  (.A(g10002), .B(g10874), .Z(g14271) ) ;
NAND2   gate20559  (.A(g26549), .B(g14271), .Z(II26438) ) ;
NAND2   gate20560  (.A(g26549), .B(II26438), .Z(II26439) ) ;
NAND2   gate20561  (.A(g14271), .B(II26438), .Z(II26440) ) ;
NAND4   gate20562  (.A(g21228), .B(g25356), .C(g26424), .D(g26236), .Z(g27933) ) ;
NOR2    gate20563  (.A(g10060), .B(g10887), .Z(g14306) ) ;
NAND2   gate20564  (.A(g26576), .B(g14306), .Z(II26459) ) ;
NAND2   gate20565  (.A(g26576), .B(II26459), .Z(II26460) ) ;
NAND2   gate20566  (.A(g14306), .B(II26459), .Z(II26461) ) ;
NAND2   gate20567  (.A(g27051), .B(g25783), .Z(g28109) ) ;
NAND2   gate20568  (.A(g27051), .B(g25838), .Z(g28131) ) ;
NOR2    gate20569  (.A(g1668), .B(g1592), .Z(g9586) ) ;
NOR2    gate20570  (.A(g1802), .B(g1728), .Z(g9640) ) ;
NOR2    gate20571  (.A(g2227), .B(g2153), .Z(g9649) ) ;
NOR2    gate20572  (.A(g1936), .B(g1862), .Z(g9694) ) ;
NOR2    gate20573  (.A(g2361), .B(g2287), .Z(g9700) ) ;
NOR2    gate20574  (.A(g2070), .B(g1996), .Z(g9755) ) ;
NOR2    gate20575  (.A(g2495), .B(g2421), .Z(g9762) ) ;
NOR2    gate20576  (.A(g2629), .B(g2555), .Z(g9835) ) ;
NOR2    gate20577  (.A(g22409), .B(g22360), .Z(g25540) ) ;
NAND2   gate20578  (.A(g25540), .B(g28131), .Z(g29335) ) ;
NOR2    gate20579  (.A(g22409), .B(g22360), .Z(g24383) ) ;
NAND2   gate20580  (.A(g28336), .B(g13464), .Z(g29540) ) ;
NAND2   gate20581  (.A(g28349), .B(g13486), .Z(g29556) ) ;
NAND2   gate20582  (.A(g28448), .B(g9582), .Z(g29660) ) ;
NAND2   gate20583  (.A(g29355), .B(g19666), .Z(g30573) ) ;
NAND2   gate20584  (.A(g29335), .B(g19666), .Z(g30580) ) ;
NOR2    gate20585  (.A(g22763), .B(g28241), .Z(g29497) ) ;
NOR2    gate20586  (.A(g22763), .B(g28250), .Z(g29503) ) ;
NOR2    gate20587  (.A(g9969), .B(g9586), .Z(g12017) ) ;
NAND2   gate20588  (.A(g29482), .B(g12017), .Z(II29253) ) ;
NAND2   gate20589  (.A(g29482), .B(II29253), .Z(II29254) ) ;
NAND2   gate20590  (.A(g12017), .B(II29253), .Z(II29255) ) ;
NOR2    gate20591  (.A(g10036), .B(g9640), .Z(g12046) ) ;
NAND2   gate20592  (.A(g29485), .B(g12046), .Z(II29261) ) ;
NAND2   gate20593  (.A(g29485), .B(II29261), .Z(II29262) ) ;
NAND2   gate20594  (.A(g12046), .B(II29261), .Z(II29263) ) ;
NOR2    gate20595  (.A(g10038), .B(g9649), .Z(g12050) ) ;
NAND2   gate20596  (.A(g29486), .B(g12050), .Z(II29269) ) ;
NAND2   gate20597  (.A(g29486), .B(II29269), .Z(II29270) ) ;
NAND2   gate20598  (.A(g12050), .B(II29269), .Z(II29271) ) ;
NOR2    gate20599  (.A(g10079), .B(g9694), .Z(g12081) ) ;
NAND2   gate20600  (.A(g29488), .B(g12081), .Z(II29277) ) ;
NAND2   gate20601  (.A(g29488), .B(II29277), .Z(II29278) ) ;
NAND2   gate20602  (.A(g12081), .B(II29277), .Z(II29279) ) ;
NOR2    gate20603  (.A(g10082), .B(g9700), .Z(g12085) ) ;
NAND2   gate20604  (.A(g29489), .B(g12085), .Z(II29284) ) ;
NAND2   gate20605  (.A(g29489), .B(II29284), .Z(II29285) ) ;
NAND2   gate20606  (.A(g12085), .B(II29284), .Z(II29286) ) ;
NOR2    gate20607  (.A(g10113), .B(g9755), .Z(g12117) ) ;
NAND2   gate20608  (.A(g29495), .B(g12117), .Z(II29295) ) ;
NAND2   gate20609  (.A(g29495), .B(II29295), .Z(II29296) ) ;
NAND2   gate20610  (.A(g12117), .B(II29295), .Z(II29297) ) ;
NOR2    gate20611  (.A(g10117), .B(g9762), .Z(g12121) ) ;
NAND2   gate20612  (.A(g29496), .B(g12121), .Z(II29302) ) ;
NAND2   gate20613  (.A(g29496), .B(II29302), .Z(II29303) ) ;
NAND2   gate20614  (.A(g12121), .B(II29302), .Z(II29304) ) ;
NOR2    gate20615  (.A(g10155), .B(g9835), .Z(g12154) ) ;
NAND2   gate20616  (.A(g29501), .B(g12154), .Z(II29313) ) ;
NAND2   gate20617  (.A(g29501), .B(II29313), .Z(II29314) ) ;
NAND2   gate20618  (.A(g12154), .B(II29313), .Z(II29315) ) ;
NAND2   gate20619  (.A(g30580), .B(g15591), .Z(g31978) ) ;
NAND2   gate20620  (.A(g22306), .B(g30580), .Z(g31997) ) ;
NAND2   gate20621  (.A(g7805), .B(g32118), .Z(g33083) ) ;
NAND3   gate20622  (.A(g10159), .B(g4474), .C(g32426), .Z(g33394) ) ;
NAND2   gate20623  (.A(g33378), .B(g862), .Z(g33669) ) ;
NAND2   gate20624  (.A(g33641), .B(g33631), .Z(II31972) ) ;
NAND2   gate20625  (.A(g33641), .B(II31972), .Z(II31973) ) ;
NAND2   gate20626  (.A(g33631), .B(II31972), .Z(II31974) ) ;
NAND2   gate20627  (.A(II31973), .B(II31974), .Z(g34051) ) ;
NAND2   gate20628  (.A(g33653), .B(g33648), .Z(II31983) ) ;
NAND2   gate20629  (.A(g33653), .B(II31983), .Z(II31984) ) ;
NAND2   gate20630  (.A(g33648), .B(II31983), .Z(II31985) ) ;
NAND2   gate20631  (.A(II31984), .B(II31985), .Z(g34056) ) ;
NAND2   gate20632  (.A(g33665), .B(g33661), .Z(II32185) ) ;
NAND2   gate20633  (.A(g33665), .B(II32185), .Z(II32186) ) ;
NAND2   gate20634  (.A(g33661), .B(II32185), .Z(II32187) ) ;
NAND2   gate20635  (.A(II32186), .B(II32187), .Z(g34220) ) ;
NAND2   gate20636  (.A(g33937), .B(g33670), .Z(II32202) ) ;
NAND2   gate20637  (.A(g33937), .B(II32202), .Z(II32203) ) ;
NAND2   gate20638  (.A(g33670), .B(II32202), .Z(II32204) ) ;
NAND2   gate20639  (.A(II32203), .B(II32204), .Z(g34227) ) ;
NAND2   gate20640  (.A(g34056), .B(g34051), .Z(II32431) ) ;
NAND2   gate20641  (.A(g34056), .B(II32431), .Z(II32432) ) ;
NAND2   gate20642  (.A(g34051), .B(II32431), .Z(II32433) ) ;
NAND2   gate20643  (.A(II32432), .B(II32433), .Z(g34422) ) ;
NAND2   gate20644  (.A(g34227), .B(g34220), .Z(II32439) ) ;
NAND2   gate20645  (.A(g34227), .B(II32439), .Z(II32440) ) ;
NAND2   gate20646  (.A(g34220), .B(II32439), .Z(II32441) ) ;
NAND2   gate20647  (.A(II32440), .B(II32441), .Z(g34424) ) ;
NAND2   gate20648  (.A(g34424), .B(g34422), .Z(II32516) ) ;
NAND2   gate20649  (.A(g34424), .B(II32516), .Z(II32517) ) ;
NAND2   gate20650  (.A(g34422), .B(II32516), .Z(II32518) ) ;
NAND2   gate20651  (.A(II32517), .B(II32518), .Z(g34469) ) ;
NAND2   gate20652  (.A(g34469), .B(g25779), .Z(II32756) ) ;
NAND2   gate20653  (.A(g34469), .B(II32756), .Z(II32757) ) ;
NAND2   gate20654  (.A(g25779), .B(II32756), .Z(II32758) ) ;
NOR3    gate20655  (.A(g168), .B(g174), .C(g182), .Z(g8086) ) ;
NOR4    gate20656  (.A(g2098), .B(g1964), .C(g1830), .D(g1696), .Z(g10179) ) ;
NOR4    gate20657  (.A(g2657), .B(g2523), .C(g2389), .D(g2255), .Z(g10205) ) ;
NOR3    gate20658  (.A(g4616), .B(g7133), .C(g10336), .Z(g10488) ) ;
NOR3    gate20659  (.A(g7183), .B(g4593), .C(g4584), .Z(g10510) ) ;
NOR3    gate20660  (.A(g7227), .B(g4601), .C(g4608), .Z(g10555) ) ;
NOR2    gate20661  (.A(g8534), .B(g8691), .Z(g11276) ) ;
NOR2    gate20662  (.A(g8587), .B(g8728), .Z(g11309) ) ;
NOR2    gate20663  (.A(g8626), .B(g8751), .Z(g11363) ) ;
NOR2    gate20664  (.A(g6856), .B(g2748), .Z(g12123) ) ;
NOR2    gate20665  (.A(g9856), .B(g10124), .Z(g12166) ) ;
NOR2    gate20666  (.A(g9927), .B(g10160), .Z(g12204) ) ;
NOR2    gate20667  (.A(g9995), .B(g10185), .Z(g12252) ) ;
NOR2    gate20668  (.A(g10053), .B(g10207), .Z(g12314) ) ;
NOR2    gate20669  (.A(g10102), .B(g10224), .Z(g12364) ) ;
NOR4    gate20670  (.A(g9012), .B(g8956), .C(g8904), .D(g8863), .Z(g12435) ) ;
NOR4    gate20671  (.A(g9055), .B(g9013), .C(g8957), .D(g8905), .Z(g12486) ) ;
NOR4    gate20672  (.A(g7132), .B(g10223), .C(g7149), .D(g10261), .Z(g12821) ) ;
NOR3    gate20673  (.A(g10555), .B(g10510), .C(g10488), .Z(g12970) ) ;
NOR2    gate20674  (.A(g278), .B(g11166), .Z(g13622) ) ;
NOR2    gate20675  (.A(g528), .B(g11185), .Z(g13661) ) ;
NOR4    gate20676  (.A(g10622), .B(g10617), .C(g10609), .D(g10603), .Z(g14751) ) ;
NOR4    gate20677  (.A(g10653), .B(g10623), .C(g10618), .D(g10611), .Z(g14792) ) ;
NOR2    gate20678  (.A(g13858), .B(g11330), .Z(g15718) ) ;
NOR2    gate20679  (.A(g13858), .B(g11374), .Z(g15724) ) ;
NOR2    gate20680  (.A(g13462), .B(g4704), .Z(g16201) ) ;
NOR2    gate20681  (.A(g13478), .B(g4749), .Z(g16209) ) ;
NOR2    gate20682  (.A(g13479), .B(g4894), .Z(g16210) ) ;
NOR2    gate20683  (.A(g13498), .B(g4760), .Z(g16219) ) ;
NOR2    gate20684  (.A(g13499), .B(g4939), .Z(g16220) ) ;
NOR2    gate20685  (.A(g13515), .B(g4771), .Z(g16231) ) ;
NOR2    gate20686  (.A(g13516), .B(g4950), .Z(g16232) ) ;
NOR2    gate20687  (.A(g13529), .B(g4961), .Z(g16242) ) ;
NOR2    gate20688  (.A(g13697), .B(g13656), .Z(g16488) ) ;
NOR2    gate20689  (.A(g13756), .B(g8086), .Z(g16581) ) ;
NOR2    gate20690  (.A(g16268), .B(g1061), .Z(g19778) ) ;
NOR2    gate20691  (.A(g16292), .B(g1404), .Z(g19793) ) ;
NOR2    gate20692  (.A(g15746), .B(g1052), .Z(g19853) ) ;
NOR2    gate20693  (.A(g15755), .B(g1395), .Z(g19873) ) ;
NOR2    gate20694  (.A(g2827), .B(g18949), .Z(g22190) ) ;
NOR2    gate20695  (.A(g7936), .B(g19407), .Z(g23024) ) ;
NOR2    gate20696  (.A(g7960), .B(g19427), .Z(g23051) ) ;
NOR2    gate20697  (.A(g2767), .B(g21066), .Z(g23686) ) ;
NOR2    gate20698  (.A(g2795), .B(g21276), .Z(g23763) ) ;
NOR2    gate20699  (.A(g2791), .B(g21303), .Z(g23835) ) ;
NOR2    gate20700  (.A(g2811), .B(g21348), .Z(g23871) ) ;
NOR2    gate20701  (.A(g2779), .B(g21067), .Z(g23883) ) ;
NOR2    gate20702  (.A(g2799), .B(g21382), .Z(g23918) ) ;
NOR2    gate20703  (.A(g2823), .B(g18890), .Z(g23955) ) ;
NOR2    gate20704  (.A(g11326), .B(g29660), .Z(g31294) ) ;

endmodule
